
module SubBytes_0 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;

  XNOR U2962 ( .A(n886), .B(n930), .Z(n905) );
  XNOR U2963 ( .A(n775), .B(n1434), .Z(n794) );
  XNOR U2964 ( .A(n1144), .B(n1188), .Z(n1163) );
  XOR U2965 ( .A(n1814), .B(n1777), .Z(n1784) );
  XNOR U2966 ( .A(n1390), .B(n1449), .Z(n1409) );
  XOR U2967 ( .A(n1048), .B(n1011), .Z(n1018) );
  XOR U2968 ( .A(n1690), .B(n1653), .Z(n1660) );
  XOR U2969 ( .A(n467), .B(n430), .Z(n437) );
  XNOR U2970 ( .A(n1900), .B(n1946), .Z(n1919) );
  XNOR U2971 ( .A(n1267), .B(n1311), .Z(n1286) );
  XOR U2972 ( .A(n622), .B(n585), .Z(n592) );
  XNOR U2973 ( .A(n1528), .B(n1572), .Z(n1547) );
  XNOR U2974 ( .A(n253), .B(n297), .Z(n272) );
  XOR U2975 ( .A(n800), .B(n738), .Z(n745) );
  XOR U2976 ( .A(n923), .B(n886), .Z(n893) );
  XOR U2977 ( .A(n1427), .B(n775), .Z(n782) );
  XNOR U2978 ( .A(n1777), .B(n1821), .Z(n1796) );
  XOR U2979 ( .A(n1181), .B(n1144), .Z(n1151) );
  XOR U2980 ( .A(n1442), .B(n1390), .Z(n1397) );
  XNOR U2981 ( .A(n1011), .B(n1055), .Z(n1030) );
  XNOR U2982 ( .A(n430), .B(n474), .Z(n449) );
  XNOR U2983 ( .A(n1653), .B(n1697), .Z(n1672) );
  XOR U2984 ( .A(n1304), .B(n1267), .Z(n1274) );
  XOR U2985 ( .A(n1939), .B(n1900), .Z(n1907) );
  XNOR U2986 ( .A(n585), .B(n629), .Z(n604) );
  NOR U2987 ( .A(n654), .B(x[9]), .Z(n1) );
  XNOR U2988 ( .A(n329), .B(n328), .Z(n2) );
  XNOR U2989 ( .A(n1), .B(n2), .Z(n3) );
  XNOR U2990 ( .A(n312), .B(n3), .Z(n345) );
  XOR U2991 ( .A(n290), .B(n253), .Z(n260) );
  XOR U2992 ( .A(n1565), .B(n1528), .Z(n1535) );
  XNOR U2993 ( .A(n738), .B(n807), .Z(n757) );
  XOR U2994 ( .A(n163), .B(n134), .Z(n157) );
  XOR U2995 ( .A(n77), .B(n78), .Z(n129) );
  XNOR U2996 ( .A(x[9]), .B(n323), .Z(n318) );
  XOR U2997 ( .A(n604), .B(n588), .Z(n590) );
  XOR U2998 ( .A(n905), .B(n889), .Z(n891) );
  XOR U2999 ( .A(n794), .B(n778), .Z(n780) );
  XOR U3000 ( .A(n1409), .B(n1393), .Z(n1395) );
  XOR U3001 ( .A(n1030), .B(n1014), .Z(n1016) );
  XOR U3002 ( .A(n1163), .B(n1147), .Z(n1149) );
  XOR U3003 ( .A(n1286), .B(n1270), .Z(n1272) );
  XOR U3004 ( .A(n1919), .B(n1903), .Z(n1905) );
  XOR U3005 ( .A(n1796), .B(n1780), .Z(n1782) );
  XOR U3006 ( .A(n1547), .B(n1531), .Z(n1533) );
  XOR U3007 ( .A(n1672), .B(n1656), .Z(n1658) );
  XOR U3008 ( .A(n272), .B(n256), .Z(n258) );
  XOR U3009 ( .A(n449), .B(n433), .Z(n435) );
  NANDN U3010 ( .A(n116), .B(n121), .Z(n4) );
  XOR U3011 ( .A(n116), .B(n119), .Z(n5) );
  OR U3012 ( .A(n121), .B(n5), .Z(n6) );
  NANDN U3013 ( .A(n117), .B(n6), .Z(n7) );
  NAND U3014 ( .A(n4), .B(n7), .Z(n169) );
  XOR U3015 ( .A(n643), .B(n508), .Z(n511) );
  XOR U3016 ( .A(n757), .B(n741), .Z(n743) );
  XOR U3017 ( .A(x[3]), .B(x[1]), .Z(n10) );
  XNOR U3018 ( .A(x[0]), .B(x[6]), .Z(n9) );
  XOR U3019 ( .A(n9), .B(x[2]), .Z(n8) );
  XNOR U3020 ( .A(n10), .B(n8), .Z(n45) );
  XNOR U3021 ( .A(x[5]), .B(n9), .Z(n1432) );
  XOR U3022 ( .A(n1432), .B(x[4]), .Z(n787) );
  IV U3023 ( .A(n787), .Z(n19) );
  XNOR U3024 ( .A(x[7]), .B(x[4]), .Z(n13) );
  XNOR U3025 ( .A(n10), .B(n13), .Z(n73) );
  NOR U3026 ( .A(n19), .B(n73), .Z(n12) );
  XNOR U3027 ( .A(n1432), .B(x[7]), .Z(n1067) );
  XNOR U3028 ( .A(x[2]), .B(n1067), .Z(n28) );
  XNOR U3029 ( .A(x[1]), .B(n28), .Z(n23) );
  AND U3030 ( .A(x[0]), .B(n23), .Z(n11) );
  XNOR U3031 ( .A(n12), .B(n11), .Z(n16) );
  XNOR U3032 ( .A(n45), .B(n1067), .Z(n35) );
  IV U3033 ( .A(n45), .Z(n30) );
  XNOR U3034 ( .A(x[0]), .B(n30), .Z(n50) );
  IV U3035 ( .A(n13), .Z(n777) );
  AND U3036 ( .A(n50), .B(n777), .Z(n18) );
  IV U3037 ( .A(n1432), .Z(n37) );
  XNOR U3038 ( .A(n45), .B(n37), .Z(n67) );
  XOR U3039 ( .A(n67), .B(n73), .Z(n70) );
  XOR U3040 ( .A(x[2]), .B(x[4]), .Z(n779) );
  NAND U3041 ( .A(n70), .B(n779), .Z(n14) );
  XNOR U3042 ( .A(n18), .B(n14), .Z(n39) );
  XNOR U3043 ( .A(n35), .B(n39), .Z(n15) );
  XNOR U3044 ( .A(n16), .B(n15), .Z(n62) );
  XOR U3045 ( .A(x[2]), .B(x[7]), .Z(n793) );
  XNOR U3046 ( .A(x[0]), .B(n73), .Z(n74) );
  XNOR U3047 ( .A(n1432), .B(n74), .Z(n65) );
  NAND U3048 ( .A(n793), .B(n65), .Z(n17) );
  XNOR U3049 ( .A(n18), .B(n17), .Z(n31) );
  IV U3050 ( .A(n23), .Z(n776) );
  XNOR U3051 ( .A(n776), .B(n19), .Z(n783) );
  AND U3052 ( .A(n73), .B(n783), .Z(n21) );
  AND U3053 ( .A(x[0]), .B(n787), .Z(n20) );
  XNOR U3054 ( .A(n21), .B(n20), .Z(n22) );
  NANDN U3055 ( .A(n74), .B(n22), .Z(n26) );
  NAND U3056 ( .A(x[0]), .B(n73), .Z(n24) );
  OR U3057 ( .A(n24), .B(n23), .Z(n25) );
  NAND U3058 ( .A(n26), .B(n25), .Z(n27) );
  XNOR U3059 ( .A(n28), .B(n27), .Z(n29) );
  XNOR U3060 ( .A(n31), .B(n29), .Z(n51) );
  IV U3061 ( .A(n51), .Z(n58) );
  AND U3062 ( .A(n1067), .B(n30), .Z(n33) );
  XOR U3063 ( .A(x[1]), .B(x[7]), .Z(n1069) );
  AND U3064 ( .A(n67), .B(n1069), .Z(n36) );
  XNOR U3065 ( .A(n36), .B(n31), .Z(n32) );
  XNOR U3066 ( .A(n33), .B(n32), .Z(n57) );
  NANDN U3067 ( .A(n58), .B(n57), .Z(n34) );
  NAND U3068 ( .A(n62), .B(n34), .Z(n44) );
  XNOR U3069 ( .A(n36), .B(n35), .Z(n41) );
  ANDN U3070 ( .B(n37), .A(x[1]), .Z(n38) );
  XNOR U3071 ( .A(n39), .B(n38), .Z(n40) );
  XNOR U3072 ( .A(n41), .B(n40), .Z(n54) );
  XOR U3073 ( .A(n57), .B(n54), .Z(n42) );
  NAND U3074 ( .A(n58), .B(n42), .Z(n43) );
  NAND U3075 ( .A(n44), .B(n43), .Z(n1066) );
  ANDN U3076 ( .B(n45), .A(n1066), .Z(n69) );
  IV U3077 ( .A(n54), .Z(n60) );
  XOR U3078 ( .A(n62), .B(n58), .Z(n46) );
  NANDN U3079 ( .A(n60), .B(n46), .Z(n49) );
  NANDN U3080 ( .A(n58), .B(n60), .Z(n47) );
  NANDN U3081 ( .A(n57), .B(n47), .Z(n48) );
  NAND U3082 ( .A(n49), .B(n48), .Z(n1427) );
  XNOR U3083 ( .A(n1066), .B(n1427), .Z(n778) );
  AND U3084 ( .A(n50), .B(n778), .Z(n72) );
  OR U3085 ( .A(n57), .B(n54), .Z(n56) );
  ANDN U3086 ( .B(n57), .A(n51), .Z(n52) );
  XNOR U3087 ( .A(n52), .B(n62), .Z(n53) );
  NAND U3088 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3089 ( .A(n56), .B(n55), .Z(n775) );
  NAND U3090 ( .A(n58), .B(n62), .Z(n64) );
  NAND U3091 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U3092 ( .A(n60), .B(n59), .Z(n61) );
  NANDN U3093 ( .A(n62), .B(n61), .Z(n63) );
  NAND U3094 ( .A(n64), .B(n63), .Z(n1434) );
  NAND U3095 ( .A(n794), .B(n65), .Z(n66) );
  XNOR U3096 ( .A(n72), .B(n66), .Z(n1429) );
  XOR U3097 ( .A(n1066), .B(n1434), .Z(n1068) );
  AND U3098 ( .A(n67), .B(n1068), .Z(n789) );
  XNOR U3099 ( .A(n1429), .B(n789), .Z(n68) );
  XNOR U3100 ( .A(n69), .B(n68), .Z(n1437) );
  NAND U3101 ( .A(n780), .B(n70), .Z(n71) );
  XNOR U3102 ( .A(n72), .B(n71), .Z(n797) );
  AND U3103 ( .A(n73), .B(n782), .Z(n1428) );
  NANDN U3104 ( .A(n74), .B(n775), .Z(n75) );
  XNOR U3105 ( .A(n1428), .B(n75), .Z(n939) );
  XNOR U3106 ( .A(n797), .B(n939), .Z(n786) );
  XOR U3107 ( .A(n1437), .B(n786), .Z(z[0]) );
  XOR U3108 ( .A(x[99]), .B(x[97]), .Z(n76) );
  XNOR U3109 ( .A(n76), .B(x[98]), .Z(n77) );
  XNOR U3110 ( .A(x[101]), .B(n77), .Z(n114) );
  XOR U3111 ( .A(x[98]), .B(x[100]), .Z(n135) );
  XNOR U3112 ( .A(x[102]), .B(n77), .Z(n128) );
  XOR U3113 ( .A(x[103]), .B(x[100]), .Z(n133) );
  XOR U3114 ( .A(n76), .B(n133), .Z(n124) );
  XNOR U3115 ( .A(x[96]), .B(n124), .Z(n93) );
  IV U3116 ( .A(n93), .Z(n125) );
  XNOR U3117 ( .A(x[102]), .B(x[96]), .Z(n78) );
  XNOR U3118 ( .A(x[101]), .B(n78), .Z(n139) );
  XOR U3119 ( .A(n125), .B(n139), .Z(n127) );
  XOR U3120 ( .A(n128), .B(n127), .Z(n156) );
  AND U3121 ( .A(n135), .B(n156), .Z(n80) );
  AND U3122 ( .A(n128), .B(n133), .Z(n86) );
  IV U3123 ( .A(n139), .Z(n102) );
  XNOR U3124 ( .A(x[103]), .B(n102), .Z(n161) );
  XOR U3125 ( .A(n129), .B(n161), .Z(n84) );
  XNOR U3126 ( .A(n86), .B(n84), .Z(n79) );
  XNOR U3127 ( .A(n80), .B(n79), .Z(n103) );
  XOR U3128 ( .A(x[98]), .B(n161), .Z(n98) );
  XOR U3129 ( .A(x[97]), .B(n98), .Z(n150) );
  ANDN U3130 ( .B(x[96]), .A(n150), .Z(n82) );
  XNOR U3131 ( .A(x[100]), .B(n102), .Z(n170) );
  NANDN U3132 ( .A(n124), .B(n170), .Z(n81) );
  XNOR U3133 ( .A(n82), .B(n81), .Z(n83) );
  XOR U3134 ( .A(n103), .B(n83), .Z(n119) );
  XOR U3135 ( .A(x[97]), .B(x[103]), .Z(n138) );
  AND U3136 ( .A(n138), .B(n114), .Z(n104) );
  XOR U3137 ( .A(n84), .B(n104), .Z(n89) );
  XOR U3138 ( .A(x[98]), .B(x[103]), .Z(n162) );
  NAND U3139 ( .A(n162), .B(n127), .Z(n85) );
  XOR U3140 ( .A(n86), .B(n85), .Z(n99) );
  AND U3141 ( .A(n129), .B(n161), .Z(n87) );
  XOR U3142 ( .A(n99), .B(n87), .Z(n88) );
  XNOR U3143 ( .A(n89), .B(n88), .Z(n117) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n152) );
  AND U3145 ( .A(n124), .B(n152), .Z(n91) );
  AND U3146 ( .A(x[96]), .B(n170), .Z(n90) );
  XNOR U3147 ( .A(n91), .B(n90), .Z(n92) );
  NANDN U3148 ( .A(n93), .B(n92), .Z(n96) );
  NAND U3149 ( .A(n124), .B(x[96]), .Z(n94) );
  NANDN U3150 ( .A(n94), .B(n150), .Z(n95) );
  NAND U3151 ( .A(n96), .B(n95), .Z(n97) );
  XNOR U3152 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U3153 ( .A(n100), .B(n99), .Z(n116) );
  OR U3154 ( .A(n117), .B(n116), .Z(n101) );
  NANDN U3155 ( .A(n119), .B(n101), .Z(n109) );
  ANDN U3156 ( .B(n102), .A(x[97]), .Z(n106) );
  XNOR U3157 ( .A(n104), .B(n103), .Z(n105) );
  XNOR U3158 ( .A(n106), .B(n105), .Z(n121) );
  XOR U3159 ( .A(n117), .B(n121), .Z(n107) );
  NAND U3160 ( .A(n116), .B(n107), .Z(n108) );
  NAND U3161 ( .A(n109), .B(n108), .Z(n160) );
  OR U3162 ( .A(n119), .B(n116), .Z(n113) );
  ANDN U3163 ( .B(n116), .A(n117), .Z(n110) );
  XNOR U3164 ( .A(n110), .B(n121), .Z(n111) );
  NAND U3165 ( .A(n119), .B(n111), .Z(n112) );
  NAND U3166 ( .A(n113), .B(n112), .Z(n141) );
  XNOR U3167 ( .A(n160), .B(n141), .Z(n137) );
  AND U3168 ( .A(n114), .B(n137), .Z(n131) );
  NAND U3169 ( .A(n139), .B(n141), .Z(n115) );
  XNOR U3170 ( .A(n131), .B(n115), .Z(n172) );
  NANDN U3171 ( .A(n117), .B(n121), .Z(n123) );
  NANDN U3172 ( .A(n117), .B(n116), .Z(n118) );
  XOR U3173 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U3174 ( .A(n121), .B(n120), .Z(n122) );
  NAND U3175 ( .A(n123), .B(n122), .Z(n149) );
  XOR U3176 ( .A(n169), .B(n149), .Z(n151) );
  AND U3177 ( .A(n124), .B(n151), .Z(n144) );
  NANDN U3178 ( .A(n149), .B(n125), .Z(n126) );
  XNOR U3179 ( .A(n144), .B(n126), .Z(n159) );
  XNOR U3180 ( .A(n172), .B(n159), .Z(z[98]) );
  XNOR U3181 ( .A(n149), .B(n141), .Z(n163) );
  AND U3182 ( .A(n127), .B(n163), .Z(n183) );
  XOR U3183 ( .A(n169), .B(n160), .Z(n134) );
  AND U3184 ( .A(n128), .B(n134), .Z(n181) );
  NANDN U3185 ( .A(n160), .B(n129), .Z(n130) );
  XNOR U3186 ( .A(n131), .B(n130), .Z(n145) );
  XNOR U3187 ( .A(n181), .B(n145), .Z(n132) );
  XNOR U3188 ( .A(n183), .B(n132), .Z(n1958) );
  XOR U3189 ( .A(n1958), .B(z[98]), .Z(z[100]) );
  AND U3190 ( .A(n133), .B(n134), .Z(n165) );
  NAND U3191 ( .A(n157), .B(n135), .Z(n136) );
  XNOR U3192 ( .A(n165), .B(n136), .Z(n153) );
  AND U3193 ( .A(n138), .B(n137), .Z(n166) );
  XOR U3194 ( .A(x[97]), .B(n139), .Z(n140) );
  NAND U3195 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U3196 ( .A(n166), .B(n142), .Z(n147) );
  NANDN U3197 ( .A(n169), .B(x[96]), .Z(n143) );
  XNOR U3198 ( .A(n144), .B(n143), .Z(n180) );
  XNOR U3199 ( .A(n180), .B(n145), .Z(n146) );
  XNOR U3200 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U3201 ( .A(n153), .B(n148), .Z(z[101]) );
  ANDN U3202 ( .B(n150), .A(n149), .Z(n155) );
  AND U3203 ( .A(n152), .B(n151), .Z(n171) );
  XNOR U3204 ( .A(n171), .B(n153), .Z(n154) );
  XNOR U3205 ( .A(n155), .B(n154), .Z(n1959) );
  NAND U3206 ( .A(n157), .B(n156), .Z(n158) );
  XNOR U3207 ( .A(n181), .B(n158), .Z(n175) );
  XNOR U3208 ( .A(n175), .B(n159), .Z(n1957) );
  XNOR U3209 ( .A(n1959), .B(n1957), .Z(n179) );
  ANDN U3210 ( .B(n161), .A(n160), .Z(n168) );
  NAND U3211 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U3212 ( .A(n165), .B(n164), .Z(n176) );
  XNOR U3213 ( .A(n176), .B(n166), .Z(n167) );
  XNOR U3214 ( .A(n168), .B(n167), .Z(n1962) );
  XNOR U3215 ( .A(n179), .B(n1962), .Z(z[102]) );
  ANDN U3216 ( .B(n170), .A(n169), .Z(n174) );
  XNOR U3217 ( .A(n172), .B(n171), .Z(n173) );
  XNOR U3218 ( .A(n174), .B(n173), .Z(n178) );
  XNOR U3219 ( .A(n176), .B(n175), .Z(n177) );
  XNOR U3220 ( .A(n178), .B(n177), .Z(n1960) );
  XNOR U3221 ( .A(n1960), .B(n179), .Z(z[97]) );
  XNOR U3222 ( .A(n181), .B(n180), .Z(n182) );
  XNOR U3223 ( .A(n183), .B(n182), .Z(n184) );
  XOR U3224 ( .A(n184), .B(z[97]), .Z(z[103]) );
  XOR U3225 ( .A(x[107]), .B(x[105]), .Z(n187) );
  XNOR U3226 ( .A(x[104]), .B(x[110]), .Z(n186) );
  XOR U3227 ( .A(n186), .B(x[106]), .Z(n185) );
  XNOR U3228 ( .A(n187), .B(n185), .Z(n222) );
  XNOR U3229 ( .A(x[109]), .B(n186), .Z(n295) );
  XOR U3230 ( .A(n295), .B(x[108]), .Z(n265) );
  IV U3231 ( .A(n265), .Z(n196) );
  XNOR U3232 ( .A(x[111]), .B(x[108]), .Z(n190) );
  XNOR U3233 ( .A(n187), .B(n190), .Z(n250) );
  NOR U3234 ( .A(n196), .B(n250), .Z(n189) );
  XNOR U3235 ( .A(n295), .B(x[111]), .Z(n281) );
  XNOR U3236 ( .A(x[106]), .B(n281), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n205), .Z(n200) );
  AND U3238 ( .A(x[104]), .B(n200), .Z(n188) );
  XNOR U3239 ( .A(n189), .B(n188), .Z(n193) );
  XNOR U3240 ( .A(n222), .B(n281), .Z(n212) );
  IV U3241 ( .A(n222), .Z(n207) );
  XNOR U3242 ( .A(x[104]), .B(n207), .Z(n227) );
  IV U3243 ( .A(n190), .Z(n255) );
  AND U3244 ( .A(n227), .B(n255), .Z(n195) );
  IV U3245 ( .A(n295), .Z(n214) );
  XNOR U3246 ( .A(n222), .B(n214), .Z(n244) );
  XOR U3247 ( .A(n244), .B(n250), .Z(n247) );
  XOR U3248 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NAND U3249 ( .A(n247), .B(n257), .Z(n191) );
  XNOR U3250 ( .A(n195), .B(n191), .Z(n216) );
  XNOR U3251 ( .A(n212), .B(n216), .Z(n192) );
  XNOR U3252 ( .A(n193), .B(n192), .Z(n239) );
  XOR U3253 ( .A(x[106]), .B(x[111]), .Z(n271) );
  XNOR U3254 ( .A(x[104]), .B(n250), .Z(n251) );
  XNOR U3255 ( .A(n295), .B(n251), .Z(n242) );
  NAND U3256 ( .A(n271), .B(n242), .Z(n194) );
  XNOR U3257 ( .A(n195), .B(n194), .Z(n208) );
  IV U3258 ( .A(n200), .Z(n254) );
  XNOR U3259 ( .A(n254), .B(n196), .Z(n261) );
  AND U3260 ( .A(n250), .B(n261), .Z(n198) );
  AND U3261 ( .A(x[104]), .B(n265), .Z(n197) );
  XNOR U3262 ( .A(n198), .B(n197), .Z(n199) );
  NANDN U3263 ( .A(n251), .B(n199), .Z(n203) );
  NAND U3264 ( .A(x[104]), .B(n250), .Z(n201) );
  OR U3265 ( .A(n201), .B(n200), .Z(n202) );
  NAND U3266 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U3267 ( .A(n205), .B(n204), .Z(n206) );
  XNOR U3268 ( .A(n208), .B(n206), .Z(n228) );
  IV U3269 ( .A(n228), .Z(n235) );
  AND U3270 ( .A(n281), .B(n207), .Z(n210) );
  XOR U3271 ( .A(x[105]), .B(x[111]), .Z(n283) );
  AND U3272 ( .A(n244), .B(n283), .Z(n213) );
  XNOR U3273 ( .A(n213), .B(n208), .Z(n209) );
  XNOR U3274 ( .A(n210), .B(n209), .Z(n234) );
  NANDN U3275 ( .A(n235), .B(n234), .Z(n211) );
  NAND U3276 ( .A(n239), .B(n211), .Z(n221) );
  XNOR U3277 ( .A(n213), .B(n212), .Z(n218) );
  ANDN U3278 ( .B(n214), .A(x[105]), .Z(n215) );
  XNOR U3279 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3280 ( .A(n218), .B(n217), .Z(n231) );
  XOR U3281 ( .A(n234), .B(n231), .Z(n219) );
  NAND U3282 ( .A(n235), .B(n219), .Z(n220) );
  NAND U3283 ( .A(n221), .B(n220), .Z(n280) );
  ANDN U3284 ( .B(n222), .A(n280), .Z(n246) );
  IV U3285 ( .A(n231), .Z(n237) );
  XOR U3286 ( .A(n239), .B(n235), .Z(n223) );
  NANDN U3287 ( .A(n237), .B(n223), .Z(n226) );
  NANDN U3288 ( .A(n235), .B(n237), .Z(n224) );
  NANDN U3289 ( .A(n234), .B(n224), .Z(n225) );
  NAND U3290 ( .A(n226), .B(n225), .Z(n290) );
  XNOR U3291 ( .A(n280), .B(n290), .Z(n256) );
  AND U3292 ( .A(n227), .B(n256), .Z(n249) );
  OR U3293 ( .A(n234), .B(n231), .Z(n233) );
  ANDN U3294 ( .B(n234), .A(n228), .Z(n229) );
  XNOR U3295 ( .A(n229), .B(n239), .Z(n230) );
  NAND U3296 ( .A(n231), .B(n230), .Z(n232) );
  NAND U3297 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3298 ( .A(n235), .B(n239), .Z(n241) );
  NAND U3299 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U3300 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U3301 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3302 ( .A(n241), .B(n240), .Z(n297) );
  NAND U3303 ( .A(n272), .B(n242), .Z(n243) );
  XNOR U3304 ( .A(n249), .B(n243), .Z(n292) );
  XOR U3305 ( .A(n280), .B(n297), .Z(n282) );
  AND U3306 ( .A(n244), .B(n282), .Z(n267) );
  XNOR U3307 ( .A(n292), .B(n267), .Z(n245) );
  XNOR U3308 ( .A(n246), .B(n245), .Z(n300) );
  NAND U3309 ( .A(n258), .B(n247), .Z(n248) );
  XNOR U3310 ( .A(n249), .B(n248), .Z(n275) );
  AND U3311 ( .A(n250), .B(n260), .Z(n291) );
  NANDN U3312 ( .A(n251), .B(n253), .Z(n252) );
  XNOR U3313 ( .A(n291), .B(n252), .Z(n279) );
  XNOR U3314 ( .A(n275), .B(n279), .Z(n264) );
  XOR U3315 ( .A(n300), .B(n264), .Z(z[104]) );
  AND U3316 ( .A(n254), .B(n253), .Z(n263) );
  AND U3317 ( .A(n256), .B(n255), .Z(n274) );
  NAND U3318 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3319 ( .A(n274), .B(n259), .Z(n301) );
  AND U3320 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3321 ( .A(n301), .B(n268), .Z(n262) );
  XNOR U3322 ( .A(n263), .B(n262), .Z(n288) );
  XNOR U3323 ( .A(n288), .B(n264), .Z(n360) );
  AND U3324 ( .A(n265), .B(n290), .Z(n270) );
  NANDN U3325 ( .A(n297), .B(n295), .Z(n266) );
  XNOR U3326 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3327 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3328 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3329 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3330 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3331 ( .A(n275), .B(n284), .Z(n276) );
  XNOR U3332 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3333 ( .A(n360), .B(n287), .Z(z[105]) );
  XNOR U3334 ( .A(n279), .B(n278), .Z(z[106]) );
  NOR U3335 ( .A(n281), .B(n280), .Z(n286) );
  AND U3336 ( .A(n283), .B(n282), .Z(n299) );
  XNOR U3337 ( .A(n284), .B(n299), .Z(n285) );
  XNOR U3338 ( .A(n286), .B(n285), .Z(n359) );
  XOR U3339 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U3340 ( .A(n359), .B(n289), .Z(z[107]) );
  XOR U3341 ( .A(n300), .B(z[106]), .Z(z[108]) );
  AND U3342 ( .A(x[104]), .B(n290), .Z(n294) );
  XNOR U3343 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U3344 ( .A(n294), .B(n293), .Z(n361) );
  XOR U3345 ( .A(n295), .B(x[105]), .Z(n296) );
  NANDN U3346 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U3347 ( .A(n299), .B(n298), .Z(n303) );
  XNOR U3348 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U3349 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U3350 ( .A(n361), .B(n304), .Z(z[109]) );
  XOR U3351 ( .A(x[9]), .B(x[11]), .Z(n305) );
  XOR U3352 ( .A(x[15]), .B(x[12]), .Z(n486) );
  XOR U3353 ( .A(n305), .B(n486), .Z(n341) );
  XNOR U3354 ( .A(x[8]), .B(x[14]), .Z(n307) );
  XNOR U3355 ( .A(x[13]), .B(n307), .Z(n654) );
  XNOR U3356 ( .A(x[15]), .B(n654), .Z(n485) );
  XNOR U3357 ( .A(n305), .B(x[10]), .Z(n306) );
  XNOR U3358 ( .A(n307), .B(n306), .Z(n308) );
  AND U3359 ( .A(n485), .B(n308), .Z(n311) );
  IV U3360 ( .A(n308), .Z(n641) );
  XOR U3361 ( .A(n641), .B(n654), .Z(n357) );
  XOR U3362 ( .A(x[9]), .B(x[15]), .Z(n491) );
  AND U3363 ( .A(n357), .B(n491), .Z(n312) );
  XNOR U3364 ( .A(x[8]), .B(n308), .Z(n509) );
  AND U3365 ( .A(n486), .B(n509), .Z(n314) );
  XOR U3366 ( .A(x[15]), .B(x[10]), .Z(n488) );
  XNOR U3367 ( .A(n341), .B(x[8]), .Z(n342) );
  XNOR U3368 ( .A(n654), .B(n342), .Z(n642) );
  NAND U3369 ( .A(n488), .B(n642), .Z(n309) );
  XNOR U3370 ( .A(n314), .B(n309), .Z(n325) );
  XNOR U3371 ( .A(n312), .B(n325), .Z(n310) );
  XNOR U3372 ( .A(n311), .B(n310), .Z(n349) );
  XNOR U3373 ( .A(n641), .B(n485), .Z(n329) );
  XOR U3374 ( .A(x[12]), .B(x[10]), .Z(n496) );
  XOR U3375 ( .A(n341), .B(n357), .Z(n510) );
  NAND U3376 ( .A(n496), .B(n510), .Z(n313) );
  XNOR U3377 ( .A(n314), .B(n313), .Z(n328) );
  OR U3378 ( .A(n349), .B(n345), .Z(n335) );
  XNOR U3379 ( .A(x[10]), .B(n485), .Z(n323) );
  IV U3380 ( .A(n318), .Z(n495) );
  XNOR U3381 ( .A(x[12]), .B(n654), .Z(n503) );
  XNOR U3382 ( .A(n495), .B(n503), .Z(n500) );
  AND U3383 ( .A(n341), .B(n500), .Z(n316) );
  ANDN U3384 ( .B(x[8]), .A(n503), .Z(n315) );
  XNOR U3385 ( .A(n316), .B(n315), .Z(n317) );
  NANDN U3386 ( .A(n342), .B(n317), .Z(n321) );
  NAND U3387 ( .A(n341), .B(x[8]), .Z(n319) );
  OR U3388 ( .A(n319), .B(n318), .Z(n320) );
  NAND U3389 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U3390 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U3391 ( .A(n325), .B(n324), .Z(n336) );
  ANDN U3392 ( .B(n349), .A(n336), .Z(n332) );
  NOR U3393 ( .A(n503), .B(n341), .Z(n327) );
  ANDN U3394 ( .B(x[8]), .A(n495), .Z(n326) );
  XNOR U3395 ( .A(n327), .B(n326), .Z(n331) );
  XNOR U3396 ( .A(n329), .B(n328), .Z(n330) );
  XNOR U3397 ( .A(n331), .B(n330), .Z(n354) );
  XNOR U3398 ( .A(n332), .B(n354), .Z(n333) );
  NAND U3399 ( .A(n345), .B(n333), .Z(n334) );
  NAND U3400 ( .A(n335), .B(n334), .Z(n494) );
  IV U3401 ( .A(n494), .Z(n487) );
  IV U3402 ( .A(n345), .Z(n352) );
  IV U3403 ( .A(n336), .Z(n350) );
  XOR U3404 ( .A(n354), .B(n350), .Z(n337) );
  NANDN U3405 ( .A(n352), .B(n337), .Z(n340) );
  NANDN U3406 ( .A(n350), .B(n352), .Z(n338) );
  NANDN U3407 ( .A(n349), .B(n338), .Z(n339) );
  NAND U3408 ( .A(n340), .B(n339), .Z(n649) );
  XNOR U3409 ( .A(n487), .B(n649), .Z(n499) );
  AND U3410 ( .A(n341), .B(n499), .Z(n651) );
  NANDN U3411 ( .A(n342), .B(n494), .Z(n343) );
  XNOR U3412 ( .A(n651), .B(n343), .Z(n663) );
  NANDN U3413 ( .A(n350), .B(n349), .Z(n344) );
  NAND U3414 ( .A(n354), .B(n344), .Z(n348) );
  XOR U3415 ( .A(n349), .B(n345), .Z(n346) );
  NAND U3416 ( .A(n350), .B(n346), .Z(n347) );
  NAND U3417 ( .A(n348), .B(n347), .Z(n640) );
  NAND U3418 ( .A(n350), .B(n354), .Z(n356) );
  NAND U3419 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U3420 ( .A(n352), .B(n351), .Z(n353) );
  NANDN U3421 ( .A(n354), .B(n353), .Z(n355) );
  NAND U3422 ( .A(n356), .B(n355), .Z(n656) );
  XOR U3423 ( .A(n640), .B(n656), .Z(n490) );
  AND U3424 ( .A(n357), .B(n490), .Z(n646) );
  NANDN U3425 ( .A(n656), .B(n654), .Z(n358) );
  XNOR U3426 ( .A(n646), .B(n358), .Z(n513) );
  XNOR U3427 ( .A(n663), .B(n513), .Z(z[10]) );
  XNOR U3428 ( .A(n360), .B(n359), .Z(z[110]) );
  XOR U3429 ( .A(n361), .B(z[105]), .Z(z[111]) );
  XOR U3430 ( .A(x[115]), .B(x[113]), .Z(n364) );
  XNOR U3431 ( .A(x[112]), .B(x[118]), .Z(n363) );
  XOR U3432 ( .A(n363), .B(x[114]), .Z(n362) );
  XNOR U3433 ( .A(n364), .B(n362), .Z(n399) );
  XNOR U3434 ( .A(x[117]), .B(n363), .Z(n472) );
  XOR U3435 ( .A(n472), .B(x[116]), .Z(n442) );
  IV U3436 ( .A(n442), .Z(n373) );
  XNOR U3437 ( .A(x[119]), .B(x[116]), .Z(n367) );
  XNOR U3438 ( .A(n364), .B(n367), .Z(n427) );
  NOR U3439 ( .A(n373), .B(n427), .Z(n366) );
  XNOR U3440 ( .A(n472), .B(x[119]), .Z(n458) );
  XNOR U3441 ( .A(x[114]), .B(n458), .Z(n382) );
  XNOR U3442 ( .A(x[113]), .B(n382), .Z(n377) );
  AND U3443 ( .A(x[112]), .B(n377), .Z(n365) );
  XNOR U3444 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U3445 ( .A(n399), .B(n458), .Z(n389) );
  IV U3446 ( .A(n399), .Z(n384) );
  XNOR U3447 ( .A(x[112]), .B(n384), .Z(n404) );
  IV U3448 ( .A(n367), .Z(n432) );
  AND U3449 ( .A(n404), .B(n432), .Z(n372) );
  IV U3450 ( .A(n472), .Z(n391) );
  XNOR U3451 ( .A(n399), .B(n391), .Z(n421) );
  XOR U3452 ( .A(n421), .B(n427), .Z(n424) );
  XOR U3453 ( .A(x[114]), .B(x[116]), .Z(n434) );
  NAND U3454 ( .A(n424), .B(n434), .Z(n368) );
  XNOR U3455 ( .A(n372), .B(n368), .Z(n393) );
  XNOR U3456 ( .A(n389), .B(n393), .Z(n369) );
  XNOR U3457 ( .A(n370), .B(n369), .Z(n416) );
  XOR U3458 ( .A(x[114]), .B(x[119]), .Z(n448) );
  XNOR U3459 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3460 ( .A(n472), .B(n428), .Z(n419) );
  NAND U3461 ( .A(n448), .B(n419), .Z(n371) );
  XNOR U3462 ( .A(n372), .B(n371), .Z(n385) );
  IV U3463 ( .A(n377), .Z(n431) );
  XNOR U3464 ( .A(n431), .B(n373), .Z(n438) );
  AND U3465 ( .A(n427), .B(n438), .Z(n375) );
  AND U3466 ( .A(x[112]), .B(n442), .Z(n374) );
  XNOR U3467 ( .A(n375), .B(n374), .Z(n376) );
  NANDN U3468 ( .A(n428), .B(n376), .Z(n380) );
  NAND U3469 ( .A(x[112]), .B(n427), .Z(n378) );
  OR U3470 ( .A(n378), .B(n377), .Z(n379) );
  NAND U3471 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U3472 ( .A(n382), .B(n381), .Z(n383) );
  XNOR U3473 ( .A(n385), .B(n383), .Z(n405) );
  IV U3474 ( .A(n405), .Z(n412) );
  AND U3475 ( .A(n458), .B(n384), .Z(n387) );
  XOR U3476 ( .A(x[113]), .B(x[119]), .Z(n460) );
  AND U3477 ( .A(n421), .B(n460), .Z(n390) );
  XNOR U3478 ( .A(n390), .B(n385), .Z(n386) );
  XNOR U3479 ( .A(n387), .B(n386), .Z(n411) );
  NANDN U3480 ( .A(n412), .B(n411), .Z(n388) );
  NAND U3481 ( .A(n416), .B(n388), .Z(n398) );
  XNOR U3482 ( .A(n390), .B(n389), .Z(n395) );
  ANDN U3483 ( .B(n391), .A(x[113]), .Z(n392) );
  XNOR U3484 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U3485 ( .A(n395), .B(n394), .Z(n408) );
  XOR U3486 ( .A(n411), .B(n408), .Z(n396) );
  NAND U3487 ( .A(n412), .B(n396), .Z(n397) );
  NAND U3488 ( .A(n398), .B(n397), .Z(n457) );
  ANDN U3489 ( .B(n399), .A(n457), .Z(n423) );
  IV U3490 ( .A(n408), .Z(n414) );
  XOR U3491 ( .A(n416), .B(n412), .Z(n400) );
  NANDN U3492 ( .A(n414), .B(n400), .Z(n403) );
  NANDN U3493 ( .A(n412), .B(n414), .Z(n401) );
  NANDN U3494 ( .A(n411), .B(n401), .Z(n402) );
  NAND U3495 ( .A(n403), .B(n402), .Z(n467) );
  XNOR U3496 ( .A(n457), .B(n467), .Z(n433) );
  AND U3497 ( .A(n404), .B(n433), .Z(n426) );
  OR U3498 ( .A(n411), .B(n408), .Z(n410) );
  ANDN U3499 ( .B(n411), .A(n405), .Z(n406) );
  XNOR U3500 ( .A(n406), .B(n416), .Z(n407) );
  NAND U3501 ( .A(n408), .B(n407), .Z(n409) );
  NAND U3502 ( .A(n410), .B(n409), .Z(n430) );
  NAND U3503 ( .A(n412), .B(n416), .Z(n418) );
  NAND U3504 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U3505 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U3506 ( .A(n416), .B(n415), .Z(n417) );
  NAND U3507 ( .A(n418), .B(n417), .Z(n474) );
  NAND U3508 ( .A(n449), .B(n419), .Z(n420) );
  XNOR U3509 ( .A(n426), .B(n420), .Z(n469) );
  XOR U3510 ( .A(n457), .B(n474), .Z(n459) );
  AND U3511 ( .A(n421), .B(n459), .Z(n444) );
  XNOR U3512 ( .A(n469), .B(n444), .Z(n422) );
  XNOR U3513 ( .A(n423), .B(n422), .Z(n477) );
  NAND U3514 ( .A(n435), .B(n424), .Z(n425) );
  XNOR U3515 ( .A(n426), .B(n425), .Z(n452) );
  AND U3516 ( .A(n427), .B(n437), .Z(n468) );
  NANDN U3517 ( .A(n428), .B(n430), .Z(n429) );
  XNOR U3518 ( .A(n468), .B(n429), .Z(n456) );
  XNOR U3519 ( .A(n452), .B(n456), .Z(n441) );
  XOR U3520 ( .A(n477), .B(n441), .Z(z[112]) );
  AND U3521 ( .A(n431), .B(n430), .Z(n440) );
  AND U3522 ( .A(n433), .B(n432), .Z(n451) );
  NAND U3523 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U3524 ( .A(n451), .B(n436), .Z(n478) );
  AND U3525 ( .A(n438), .B(n437), .Z(n445) );
  XNOR U3526 ( .A(n478), .B(n445), .Z(n439) );
  XNOR U3527 ( .A(n440), .B(n439), .Z(n465) );
  XNOR U3528 ( .A(n465), .B(n441), .Z(n483) );
  AND U3529 ( .A(n442), .B(n467), .Z(n447) );
  NANDN U3530 ( .A(n474), .B(n472), .Z(n443) );
  XNOR U3531 ( .A(n444), .B(n443), .Z(n455) );
  XNOR U3532 ( .A(n445), .B(n455), .Z(n446) );
  XNOR U3533 ( .A(n447), .B(n446), .Z(n454) );
  NAND U3534 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U3535 ( .A(n451), .B(n450), .Z(n461) );
  XNOR U3536 ( .A(n452), .B(n461), .Z(n453) );
  XNOR U3537 ( .A(n454), .B(n453), .Z(n464) );
  XNOR U3538 ( .A(n483), .B(n464), .Z(z[113]) );
  XNOR U3539 ( .A(n456), .B(n455), .Z(z[114]) );
  NOR U3540 ( .A(n458), .B(n457), .Z(n463) );
  AND U3541 ( .A(n460), .B(n459), .Z(n476) );
  XNOR U3542 ( .A(n461), .B(n476), .Z(n462) );
  XNOR U3543 ( .A(n463), .B(n462), .Z(n482) );
  XOR U3544 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U3545 ( .A(n482), .B(n466), .Z(z[115]) );
  XOR U3546 ( .A(n477), .B(z[114]), .Z(z[116]) );
  AND U3547 ( .A(x[112]), .B(n467), .Z(n471) );
  XNOR U3548 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U3549 ( .A(n471), .B(n470), .Z(n484) );
  XOR U3550 ( .A(n472), .B(x[113]), .Z(n473) );
  NANDN U3551 ( .A(n474), .B(n473), .Z(n475) );
  XNOR U3552 ( .A(n476), .B(n475), .Z(n480) );
  XNOR U3553 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U3554 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U3555 ( .A(n484), .B(n481), .Z(z[117]) );
  XNOR U3556 ( .A(n483), .B(n482), .Z(z[118]) );
  XOR U3557 ( .A(n484), .B(z[113]), .Z(z[119]) );
  NOR U3558 ( .A(n485), .B(n640), .Z(n493) );
  XNOR U3559 ( .A(n640), .B(n649), .Z(n508) );
  AND U3560 ( .A(n486), .B(n508), .Z(n498) );
  XOR U3561 ( .A(n487), .B(n656), .Z(n643) );
  NAND U3562 ( .A(n643), .B(n488), .Z(n489) );
  XNOR U3563 ( .A(n498), .B(n489), .Z(n504) );
  AND U3564 ( .A(n491), .B(n490), .Z(n658) );
  XNOR U3565 ( .A(n504), .B(n658), .Z(n492) );
  XNOR U3566 ( .A(n493), .B(n492), .Z(n666) );
  AND U3567 ( .A(n495), .B(n494), .Z(n502) );
  NAND U3568 ( .A(n511), .B(n496), .Z(n497) );
  XNOR U3569 ( .A(n498), .B(n497), .Z(n659) );
  AND U3570 ( .A(n500), .B(n499), .Z(n505) );
  XNOR U3571 ( .A(n659), .B(n505), .Z(n501) );
  XNOR U3572 ( .A(n502), .B(n501), .Z(n665) );
  ANDN U3573 ( .B(n649), .A(n503), .Z(n507) );
  XNOR U3574 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U3575 ( .A(n507), .B(n506), .Z(n515) );
  AND U3576 ( .A(n509), .B(n508), .Z(n645) );
  NAND U3577 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U3578 ( .A(n645), .B(n512), .Z(n664) );
  XNOR U3579 ( .A(n664), .B(n513), .Z(n514) );
  XNOR U3580 ( .A(n515), .B(n514), .Z(n667) );
  XOR U3581 ( .A(n665), .B(n667), .Z(n516) );
  XNOR U3582 ( .A(n666), .B(n516), .Z(z[11]) );
  XOR U3583 ( .A(x[123]), .B(x[121]), .Z(n519) );
  XNOR U3584 ( .A(x[120]), .B(x[126]), .Z(n518) );
  XOR U3585 ( .A(n518), .B(x[122]), .Z(n517) );
  XNOR U3586 ( .A(n519), .B(n517), .Z(n554) );
  XNOR U3587 ( .A(x[125]), .B(n518), .Z(n627) );
  XOR U3588 ( .A(n627), .B(x[124]), .Z(n597) );
  IV U3589 ( .A(n597), .Z(n528) );
  XNOR U3590 ( .A(x[127]), .B(x[124]), .Z(n522) );
  XNOR U3591 ( .A(n519), .B(n522), .Z(n582) );
  NOR U3592 ( .A(n528), .B(n582), .Z(n521) );
  XNOR U3593 ( .A(n627), .B(x[127]), .Z(n613) );
  XNOR U3594 ( .A(x[122]), .B(n613), .Z(n537) );
  XNOR U3595 ( .A(x[121]), .B(n537), .Z(n532) );
  AND U3596 ( .A(x[120]), .B(n532), .Z(n520) );
  XNOR U3597 ( .A(n521), .B(n520), .Z(n525) );
  XNOR U3598 ( .A(n554), .B(n613), .Z(n544) );
  IV U3599 ( .A(n554), .Z(n539) );
  XNOR U3600 ( .A(x[120]), .B(n539), .Z(n559) );
  IV U3601 ( .A(n522), .Z(n587) );
  AND U3602 ( .A(n559), .B(n587), .Z(n527) );
  IV U3603 ( .A(n627), .Z(n546) );
  XNOR U3604 ( .A(n554), .B(n546), .Z(n576) );
  XOR U3605 ( .A(n576), .B(n582), .Z(n579) );
  XOR U3606 ( .A(x[122]), .B(x[124]), .Z(n589) );
  NAND U3607 ( .A(n579), .B(n589), .Z(n523) );
  XNOR U3608 ( .A(n527), .B(n523), .Z(n548) );
  XNOR U3609 ( .A(n544), .B(n548), .Z(n524) );
  XNOR U3610 ( .A(n525), .B(n524), .Z(n571) );
  XOR U3611 ( .A(x[122]), .B(x[127]), .Z(n603) );
  XNOR U3612 ( .A(x[120]), .B(n582), .Z(n583) );
  XNOR U3613 ( .A(n627), .B(n583), .Z(n574) );
  NAND U3614 ( .A(n603), .B(n574), .Z(n526) );
  XNOR U3615 ( .A(n527), .B(n526), .Z(n540) );
  IV U3616 ( .A(n532), .Z(n586) );
  XNOR U3617 ( .A(n586), .B(n528), .Z(n593) );
  AND U3618 ( .A(n582), .B(n593), .Z(n530) );
  AND U3619 ( .A(x[120]), .B(n597), .Z(n529) );
  XNOR U3620 ( .A(n530), .B(n529), .Z(n531) );
  NANDN U3621 ( .A(n583), .B(n531), .Z(n535) );
  NAND U3622 ( .A(x[120]), .B(n582), .Z(n533) );
  OR U3623 ( .A(n533), .B(n532), .Z(n534) );
  NAND U3624 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U3625 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U3626 ( .A(n540), .B(n538), .Z(n560) );
  IV U3627 ( .A(n560), .Z(n567) );
  AND U3628 ( .A(n613), .B(n539), .Z(n542) );
  XOR U3629 ( .A(x[121]), .B(x[127]), .Z(n615) );
  AND U3630 ( .A(n576), .B(n615), .Z(n545) );
  XNOR U3631 ( .A(n545), .B(n540), .Z(n541) );
  XNOR U3632 ( .A(n542), .B(n541), .Z(n566) );
  NANDN U3633 ( .A(n567), .B(n566), .Z(n543) );
  NAND U3634 ( .A(n571), .B(n543), .Z(n553) );
  XNOR U3635 ( .A(n545), .B(n544), .Z(n550) );
  ANDN U3636 ( .B(n546), .A(x[121]), .Z(n547) );
  XNOR U3637 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U3638 ( .A(n550), .B(n549), .Z(n563) );
  XOR U3639 ( .A(n566), .B(n563), .Z(n551) );
  NAND U3640 ( .A(n567), .B(n551), .Z(n552) );
  NAND U3641 ( .A(n553), .B(n552), .Z(n612) );
  ANDN U3642 ( .B(n554), .A(n612), .Z(n578) );
  IV U3643 ( .A(n563), .Z(n569) );
  XOR U3644 ( .A(n571), .B(n567), .Z(n555) );
  NANDN U3645 ( .A(n569), .B(n555), .Z(n558) );
  NANDN U3646 ( .A(n567), .B(n569), .Z(n556) );
  NANDN U3647 ( .A(n566), .B(n556), .Z(n557) );
  NAND U3648 ( .A(n558), .B(n557), .Z(n622) );
  XNOR U3649 ( .A(n612), .B(n622), .Z(n588) );
  AND U3650 ( .A(n559), .B(n588), .Z(n581) );
  OR U3651 ( .A(n566), .B(n563), .Z(n565) );
  ANDN U3652 ( .B(n566), .A(n560), .Z(n561) );
  XNOR U3653 ( .A(n561), .B(n571), .Z(n562) );
  NAND U3654 ( .A(n563), .B(n562), .Z(n564) );
  NAND U3655 ( .A(n565), .B(n564), .Z(n585) );
  NAND U3656 ( .A(n567), .B(n571), .Z(n573) );
  NAND U3657 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U3658 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U3659 ( .A(n571), .B(n570), .Z(n572) );
  NAND U3660 ( .A(n573), .B(n572), .Z(n629) );
  NAND U3661 ( .A(n604), .B(n574), .Z(n575) );
  XNOR U3662 ( .A(n581), .B(n575), .Z(n624) );
  XOR U3663 ( .A(n612), .B(n629), .Z(n614) );
  AND U3664 ( .A(n576), .B(n614), .Z(n599) );
  XNOR U3665 ( .A(n624), .B(n599), .Z(n577) );
  XNOR U3666 ( .A(n578), .B(n577), .Z(n632) );
  NAND U3667 ( .A(n590), .B(n579), .Z(n580) );
  XNOR U3668 ( .A(n581), .B(n580), .Z(n607) );
  AND U3669 ( .A(n582), .B(n592), .Z(n623) );
  NANDN U3670 ( .A(n583), .B(n585), .Z(n584) );
  XNOR U3671 ( .A(n623), .B(n584), .Z(n611) );
  XNOR U3672 ( .A(n607), .B(n611), .Z(n596) );
  XOR U3673 ( .A(n632), .B(n596), .Z(z[120]) );
  AND U3674 ( .A(n586), .B(n585), .Z(n595) );
  AND U3675 ( .A(n588), .B(n587), .Z(n606) );
  NAND U3676 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U3677 ( .A(n606), .B(n591), .Z(n633) );
  AND U3678 ( .A(n593), .B(n592), .Z(n600) );
  XNOR U3679 ( .A(n633), .B(n600), .Z(n594) );
  XNOR U3680 ( .A(n595), .B(n594), .Z(n620) );
  XNOR U3681 ( .A(n620), .B(n596), .Z(n638) );
  AND U3682 ( .A(n597), .B(n622), .Z(n602) );
  NANDN U3683 ( .A(n629), .B(n627), .Z(n598) );
  XNOR U3684 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U3685 ( .A(n600), .B(n610), .Z(n601) );
  XNOR U3686 ( .A(n602), .B(n601), .Z(n609) );
  NAND U3687 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U3688 ( .A(n606), .B(n605), .Z(n616) );
  XNOR U3689 ( .A(n607), .B(n616), .Z(n608) );
  XNOR U3690 ( .A(n609), .B(n608), .Z(n619) );
  XNOR U3691 ( .A(n638), .B(n619), .Z(z[121]) );
  XNOR U3692 ( .A(n611), .B(n610), .Z(z[122]) );
  NOR U3693 ( .A(n613), .B(n612), .Z(n618) );
  AND U3694 ( .A(n615), .B(n614), .Z(n631) );
  XNOR U3695 ( .A(n616), .B(n631), .Z(n617) );
  XNOR U3696 ( .A(n618), .B(n617), .Z(n637) );
  XOR U3697 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U3698 ( .A(n637), .B(n621), .Z(z[123]) );
  XOR U3699 ( .A(n632), .B(z[122]), .Z(z[124]) );
  AND U3700 ( .A(x[120]), .B(n622), .Z(n626) );
  XNOR U3701 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U3702 ( .A(n626), .B(n625), .Z(n639) );
  XOR U3703 ( .A(n627), .B(x[121]), .Z(n628) );
  NANDN U3704 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U3705 ( .A(n631), .B(n630), .Z(n635) );
  XNOR U3706 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U3707 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U3708 ( .A(n639), .B(n636), .Z(z[125]) );
  XNOR U3709 ( .A(n638), .B(n637), .Z(z[126]) );
  XOR U3710 ( .A(n639), .B(z[121]), .Z(z[127]) );
  ANDN U3711 ( .B(n641), .A(n640), .Z(n648) );
  NAND U3712 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U3713 ( .A(n645), .B(n644), .Z(n650) );
  XNOR U3714 ( .A(n650), .B(n646), .Z(n647) );
  XNOR U3715 ( .A(n648), .B(n647), .Z(n1926) );
  XOR U3716 ( .A(n1926), .B(z[10]), .Z(z[12]) );
  AND U3717 ( .A(x[8]), .B(n649), .Z(n653) );
  XNOR U3718 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U3719 ( .A(n653), .B(n652), .Z(n669) );
  XOR U3720 ( .A(n654), .B(x[9]), .Z(n655) );
  NANDN U3721 ( .A(n656), .B(n655), .Z(n657) );
  XNOR U3722 ( .A(n658), .B(n657), .Z(n661) );
  XNOR U3723 ( .A(n659), .B(n1926), .Z(n660) );
  XNOR U3724 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U3725 ( .A(n669), .B(n662), .Z(z[13]) );
  XNOR U3726 ( .A(n664), .B(n663), .Z(n1925) );
  XNOR U3727 ( .A(n665), .B(n1925), .Z(n668) );
  XNOR U3728 ( .A(n668), .B(n666), .Z(z[14]) );
  XNOR U3729 ( .A(n668), .B(n667), .Z(z[9]) );
  XOR U3730 ( .A(n669), .B(z[9]), .Z(z[15]) );
  XOR U3731 ( .A(x[19]), .B(x[17]), .Z(n672) );
  XNOR U3732 ( .A(x[16]), .B(x[22]), .Z(n671) );
  XOR U3733 ( .A(n671), .B(x[18]), .Z(n670) );
  XNOR U3734 ( .A(n672), .B(n670), .Z(n707) );
  XNOR U3735 ( .A(x[21]), .B(n671), .Z(n805) );
  XOR U3736 ( .A(n805), .B(x[20]), .Z(n750) );
  IV U3737 ( .A(n750), .Z(n681) );
  XNOR U3738 ( .A(x[23]), .B(x[20]), .Z(n675) );
  XNOR U3739 ( .A(n672), .B(n675), .Z(n735) );
  NOR U3740 ( .A(n681), .B(n735), .Z(n674) );
  XNOR U3741 ( .A(n805), .B(x[23]), .Z(n766) );
  XNOR U3742 ( .A(x[18]), .B(n766), .Z(n690) );
  XNOR U3743 ( .A(x[17]), .B(n690), .Z(n685) );
  AND U3744 ( .A(x[16]), .B(n685), .Z(n673) );
  XNOR U3745 ( .A(n674), .B(n673), .Z(n678) );
  XNOR U3746 ( .A(n707), .B(n766), .Z(n697) );
  IV U3747 ( .A(n707), .Z(n692) );
  XNOR U3748 ( .A(x[16]), .B(n692), .Z(n712) );
  IV U3749 ( .A(n675), .Z(n740) );
  AND U3750 ( .A(n712), .B(n740), .Z(n680) );
  IV U3751 ( .A(n805), .Z(n699) );
  XNOR U3752 ( .A(n707), .B(n699), .Z(n729) );
  XOR U3753 ( .A(n729), .B(n735), .Z(n732) );
  XOR U3754 ( .A(x[18]), .B(x[20]), .Z(n742) );
  NAND U3755 ( .A(n732), .B(n742), .Z(n676) );
  XNOR U3756 ( .A(n680), .B(n676), .Z(n701) );
  XNOR U3757 ( .A(n697), .B(n701), .Z(n677) );
  XNOR U3758 ( .A(n678), .B(n677), .Z(n724) );
  XOR U3759 ( .A(x[18]), .B(x[23]), .Z(n756) );
  XNOR U3760 ( .A(x[16]), .B(n735), .Z(n736) );
  XNOR U3761 ( .A(n805), .B(n736), .Z(n727) );
  NAND U3762 ( .A(n756), .B(n727), .Z(n679) );
  XNOR U3763 ( .A(n680), .B(n679), .Z(n693) );
  IV U3764 ( .A(n685), .Z(n739) );
  XNOR U3765 ( .A(n739), .B(n681), .Z(n746) );
  AND U3766 ( .A(n735), .B(n746), .Z(n683) );
  AND U3767 ( .A(x[16]), .B(n750), .Z(n682) );
  XNOR U3768 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U3769 ( .A(n736), .B(n684), .Z(n688) );
  NAND U3770 ( .A(x[16]), .B(n735), .Z(n686) );
  OR U3771 ( .A(n686), .B(n685), .Z(n687) );
  NAND U3772 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U3773 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U3774 ( .A(n693), .B(n691), .Z(n713) );
  IV U3775 ( .A(n713), .Z(n720) );
  AND U3776 ( .A(n766), .B(n692), .Z(n695) );
  XOR U3777 ( .A(x[17]), .B(x[23]), .Z(n768) );
  AND U3778 ( .A(n729), .B(n768), .Z(n698) );
  XNOR U3779 ( .A(n698), .B(n693), .Z(n694) );
  XNOR U3780 ( .A(n695), .B(n694), .Z(n719) );
  NANDN U3781 ( .A(n720), .B(n719), .Z(n696) );
  NAND U3782 ( .A(n724), .B(n696), .Z(n706) );
  XNOR U3783 ( .A(n698), .B(n697), .Z(n703) );
  ANDN U3784 ( .B(n699), .A(x[17]), .Z(n700) );
  XNOR U3785 ( .A(n701), .B(n700), .Z(n702) );
  XNOR U3786 ( .A(n703), .B(n702), .Z(n716) );
  XOR U3787 ( .A(n719), .B(n716), .Z(n704) );
  NAND U3788 ( .A(n720), .B(n704), .Z(n705) );
  NAND U3789 ( .A(n706), .B(n705), .Z(n765) );
  ANDN U3790 ( .B(n707), .A(n765), .Z(n731) );
  IV U3791 ( .A(n716), .Z(n722) );
  XOR U3792 ( .A(n724), .B(n720), .Z(n708) );
  NANDN U3793 ( .A(n722), .B(n708), .Z(n711) );
  NANDN U3794 ( .A(n720), .B(n722), .Z(n709) );
  NANDN U3795 ( .A(n719), .B(n709), .Z(n710) );
  NAND U3796 ( .A(n711), .B(n710), .Z(n800) );
  XNOR U3797 ( .A(n765), .B(n800), .Z(n741) );
  AND U3798 ( .A(n712), .B(n741), .Z(n734) );
  OR U3799 ( .A(n719), .B(n716), .Z(n718) );
  ANDN U3800 ( .B(n719), .A(n713), .Z(n714) );
  XNOR U3801 ( .A(n714), .B(n724), .Z(n715) );
  NAND U3802 ( .A(n716), .B(n715), .Z(n717) );
  NAND U3803 ( .A(n718), .B(n717), .Z(n738) );
  NAND U3804 ( .A(n720), .B(n724), .Z(n726) );
  NAND U3805 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U3806 ( .A(n722), .B(n721), .Z(n723) );
  NANDN U3807 ( .A(n724), .B(n723), .Z(n725) );
  NAND U3808 ( .A(n726), .B(n725), .Z(n807) );
  NAND U3809 ( .A(n757), .B(n727), .Z(n728) );
  XNOR U3810 ( .A(n734), .B(n728), .Z(n802) );
  XOR U3811 ( .A(n765), .B(n807), .Z(n767) );
  AND U3812 ( .A(n729), .B(n767), .Z(n752) );
  XNOR U3813 ( .A(n802), .B(n752), .Z(n730) );
  XNOR U3814 ( .A(n731), .B(n730), .Z(n810) );
  NAND U3815 ( .A(n743), .B(n732), .Z(n733) );
  XNOR U3816 ( .A(n734), .B(n733), .Z(n760) );
  AND U3817 ( .A(n735), .B(n745), .Z(n801) );
  NANDN U3818 ( .A(n736), .B(n738), .Z(n737) );
  XNOR U3819 ( .A(n801), .B(n737), .Z(n764) );
  XNOR U3820 ( .A(n760), .B(n764), .Z(n749) );
  XOR U3821 ( .A(n810), .B(n749), .Z(z[16]) );
  AND U3822 ( .A(n739), .B(n738), .Z(n748) );
  AND U3823 ( .A(n741), .B(n740), .Z(n759) );
  NAND U3824 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U3825 ( .A(n759), .B(n744), .Z(n811) );
  AND U3826 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U3827 ( .A(n811), .B(n753), .Z(n747) );
  XNOR U3828 ( .A(n748), .B(n747), .Z(n773) );
  XNOR U3829 ( .A(n773), .B(n749), .Z(n816) );
  AND U3830 ( .A(n750), .B(n800), .Z(n755) );
  NANDN U3831 ( .A(n807), .B(n805), .Z(n751) );
  XNOR U3832 ( .A(n752), .B(n751), .Z(n763) );
  XNOR U3833 ( .A(n753), .B(n763), .Z(n754) );
  XNOR U3834 ( .A(n755), .B(n754), .Z(n762) );
  NAND U3835 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U3836 ( .A(n759), .B(n758), .Z(n769) );
  XNOR U3837 ( .A(n760), .B(n769), .Z(n761) );
  XNOR U3838 ( .A(n762), .B(n761), .Z(n772) );
  XNOR U3839 ( .A(n816), .B(n772), .Z(z[17]) );
  XNOR U3840 ( .A(n764), .B(n763), .Z(z[18]) );
  NOR U3841 ( .A(n766), .B(n765), .Z(n771) );
  AND U3842 ( .A(n768), .B(n767), .Z(n809) );
  XNOR U3843 ( .A(n769), .B(n809), .Z(n770) );
  XNOR U3844 ( .A(n771), .B(n770), .Z(n815) );
  XOR U3845 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U3846 ( .A(n815), .B(n774), .Z(z[19]) );
  AND U3847 ( .A(n776), .B(n775), .Z(n785) );
  AND U3848 ( .A(n778), .B(n777), .Z(n796) );
  NAND U3849 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U3850 ( .A(n796), .B(n781), .Z(n1438) );
  AND U3851 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U3852 ( .A(n1438), .B(n790), .Z(n784) );
  XNOR U3853 ( .A(n785), .B(n784), .Z(n1074) );
  XNOR U3854 ( .A(n1074), .B(n786), .Z(n1581) );
  AND U3855 ( .A(n787), .B(n1427), .Z(n792) );
  NANDN U3856 ( .A(n1434), .B(n1432), .Z(n788) );
  XNOR U3857 ( .A(n789), .B(n788), .Z(n938) );
  XNOR U3858 ( .A(n790), .B(n938), .Z(n791) );
  XNOR U3859 ( .A(n792), .B(n791), .Z(n799) );
  NAND U3860 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U3861 ( .A(n796), .B(n795), .Z(n1070) );
  XNOR U3862 ( .A(n797), .B(n1070), .Z(n798) );
  XNOR U3863 ( .A(n799), .B(n798), .Z(n1073) );
  XNOR U3864 ( .A(n1581), .B(n1073), .Z(z[1]) );
  XOR U3865 ( .A(n810), .B(z[18]), .Z(z[20]) );
  AND U3866 ( .A(x[16]), .B(n800), .Z(n804) );
  XNOR U3867 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U3868 ( .A(n804), .B(n803), .Z(n817) );
  XOR U3869 ( .A(n805), .B(x[17]), .Z(n806) );
  NANDN U3870 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3871 ( .A(n809), .B(n808), .Z(n813) );
  XNOR U3872 ( .A(n811), .B(n810), .Z(n812) );
  XNOR U3873 ( .A(n813), .B(n812), .Z(n814) );
  XNOR U3874 ( .A(n817), .B(n814), .Z(z[21]) );
  XNOR U3875 ( .A(n816), .B(n815), .Z(z[22]) );
  XOR U3876 ( .A(n817), .B(z[17]), .Z(z[23]) );
  XOR U3877 ( .A(x[27]), .B(x[25]), .Z(n820) );
  XNOR U3878 ( .A(x[24]), .B(x[30]), .Z(n819) );
  XOR U3879 ( .A(n819), .B(x[26]), .Z(n818) );
  XNOR U3880 ( .A(n820), .B(n818), .Z(n855) );
  XNOR U3881 ( .A(x[29]), .B(n819), .Z(n928) );
  XOR U3882 ( .A(n928), .B(x[28]), .Z(n898) );
  IV U3883 ( .A(n898), .Z(n829) );
  XNOR U3884 ( .A(x[31]), .B(x[28]), .Z(n823) );
  XNOR U3885 ( .A(n820), .B(n823), .Z(n883) );
  NOR U3886 ( .A(n829), .B(n883), .Z(n822) );
  XNOR U3887 ( .A(n928), .B(x[31]), .Z(n914) );
  XNOR U3888 ( .A(x[26]), .B(n914), .Z(n838) );
  XNOR U3889 ( .A(x[25]), .B(n838), .Z(n833) );
  AND U3890 ( .A(x[24]), .B(n833), .Z(n821) );
  XNOR U3891 ( .A(n822), .B(n821), .Z(n826) );
  XNOR U3892 ( .A(n855), .B(n914), .Z(n845) );
  IV U3893 ( .A(n855), .Z(n840) );
  XNOR U3894 ( .A(x[24]), .B(n840), .Z(n860) );
  IV U3895 ( .A(n823), .Z(n888) );
  AND U3896 ( .A(n860), .B(n888), .Z(n828) );
  IV U3897 ( .A(n928), .Z(n847) );
  XNOR U3898 ( .A(n855), .B(n847), .Z(n877) );
  XOR U3899 ( .A(n877), .B(n883), .Z(n880) );
  XOR U3900 ( .A(x[26]), .B(x[28]), .Z(n890) );
  NAND U3901 ( .A(n880), .B(n890), .Z(n824) );
  XNOR U3902 ( .A(n828), .B(n824), .Z(n849) );
  XNOR U3903 ( .A(n845), .B(n849), .Z(n825) );
  XNOR U3904 ( .A(n826), .B(n825), .Z(n872) );
  XOR U3905 ( .A(x[26]), .B(x[31]), .Z(n904) );
  XNOR U3906 ( .A(x[24]), .B(n883), .Z(n884) );
  XNOR U3907 ( .A(n928), .B(n884), .Z(n875) );
  NAND U3908 ( .A(n904), .B(n875), .Z(n827) );
  XNOR U3909 ( .A(n828), .B(n827), .Z(n841) );
  IV U3910 ( .A(n833), .Z(n887) );
  XNOR U3911 ( .A(n887), .B(n829), .Z(n894) );
  AND U3912 ( .A(n883), .B(n894), .Z(n831) );
  AND U3913 ( .A(x[24]), .B(n898), .Z(n830) );
  XNOR U3914 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U3915 ( .A(n884), .B(n832), .Z(n836) );
  NAND U3916 ( .A(x[24]), .B(n883), .Z(n834) );
  OR U3917 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3918 ( .A(n836), .B(n835), .Z(n837) );
  XNOR U3919 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U3920 ( .A(n841), .B(n839), .Z(n861) );
  IV U3921 ( .A(n861), .Z(n868) );
  AND U3922 ( .A(n914), .B(n840), .Z(n843) );
  XOR U3923 ( .A(x[25]), .B(x[31]), .Z(n916) );
  AND U3924 ( .A(n877), .B(n916), .Z(n846) );
  XNOR U3925 ( .A(n846), .B(n841), .Z(n842) );
  XNOR U3926 ( .A(n843), .B(n842), .Z(n867) );
  NANDN U3927 ( .A(n868), .B(n867), .Z(n844) );
  NAND U3928 ( .A(n872), .B(n844), .Z(n854) );
  XNOR U3929 ( .A(n846), .B(n845), .Z(n851) );
  ANDN U3930 ( .B(n847), .A(x[25]), .Z(n848) );
  XNOR U3931 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U3932 ( .A(n851), .B(n850), .Z(n864) );
  XOR U3933 ( .A(n867), .B(n864), .Z(n852) );
  NAND U3934 ( .A(n868), .B(n852), .Z(n853) );
  NAND U3935 ( .A(n854), .B(n853), .Z(n913) );
  ANDN U3936 ( .B(n855), .A(n913), .Z(n879) );
  IV U3937 ( .A(n864), .Z(n870) );
  XOR U3938 ( .A(n872), .B(n868), .Z(n856) );
  NANDN U3939 ( .A(n870), .B(n856), .Z(n859) );
  NANDN U3940 ( .A(n868), .B(n870), .Z(n857) );
  NANDN U3941 ( .A(n867), .B(n857), .Z(n858) );
  NAND U3942 ( .A(n859), .B(n858), .Z(n923) );
  XNOR U3943 ( .A(n913), .B(n923), .Z(n889) );
  AND U3944 ( .A(n860), .B(n889), .Z(n882) );
  OR U3945 ( .A(n867), .B(n864), .Z(n866) );
  ANDN U3946 ( .B(n867), .A(n861), .Z(n862) );
  XNOR U3947 ( .A(n862), .B(n872), .Z(n863) );
  NAND U3948 ( .A(n864), .B(n863), .Z(n865) );
  NAND U3949 ( .A(n866), .B(n865), .Z(n886) );
  NAND U3950 ( .A(n868), .B(n872), .Z(n874) );
  NAND U3951 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U3952 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U3953 ( .A(n872), .B(n871), .Z(n873) );
  NAND U3954 ( .A(n874), .B(n873), .Z(n930) );
  NAND U3955 ( .A(n905), .B(n875), .Z(n876) );
  XNOR U3956 ( .A(n882), .B(n876), .Z(n925) );
  XOR U3957 ( .A(n913), .B(n930), .Z(n915) );
  AND U3958 ( .A(n877), .B(n915), .Z(n900) );
  XNOR U3959 ( .A(n925), .B(n900), .Z(n878) );
  XNOR U3960 ( .A(n879), .B(n878), .Z(n933) );
  NAND U3961 ( .A(n891), .B(n880), .Z(n881) );
  XNOR U3962 ( .A(n882), .B(n881), .Z(n908) );
  AND U3963 ( .A(n883), .B(n893), .Z(n924) );
  NANDN U3964 ( .A(n884), .B(n886), .Z(n885) );
  XNOR U3965 ( .A(n924), .B(n885), .Z(n912) );
  XNOR U3966 ( .A(n908), .B(n912), .Z(n897) );
  XOR U3967 ( .A(n933), .B(n897), .Z(z[24]) );
  AND U3968 ( .A(n887), .B(n886), .Z(n896) );
  AND U3969 ( .A(n889), .B(n888), .Z(n907) );
  NAND U3970 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U3971 ( .A(n907), .B(n892), .Z(n934) );
  AND U3972 ( .A(n894), .B(n893), .Z(n901) );
  XNOR U3973 ( .A(n934), .B(n901), .Z(n895) );
  XNOR U3974 ( .A(n896), .B(n895), .Z(n921) );
  XNOR U3975 ( .A(n921), .B(n897), .Z(n941) );
  AND U3976 ( .A(n898), .B(n923), .Z(n903) );
  NANDN U3977 ( .A(n930), .B(n928), .Z(n899) );
  XNOR U3978 ( .A(n900), .B(n899), .Z(n911) );
  XNOR U3979 ( .A(n901), .B(n911), .Z(n902) );
  XNOR U3980 ( .A(n903), .B(n902), .Z(n910) );
  NAND U3981 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3982 ( .A(n907), .B(n906), .Z(n917) );
  XNOR U3983 ( .A(n908), .B(n917), .Z(n909) );
  XNOR U3984 ( .A(n910), .B(n909), .Z(n920) );
  XNOR U3985 ( .A(n941), .B(n920), .Z(z[25]) );
  XNOR U3986 ( .A(n912), .B(n911), .Z(z[26]) );
  NOR U3987 ( .A(n914), .B(n913), .Z(n919) );
  AND U3988 ( .A(n916), .B(n915), .Z(n932) );
  XNOR U3989 ( .A(n917), .B(n932), .Z(n918) );
  XNOR U3990 ( .A(n919), .B(n918), .Z(n940) );
  XOR U3991 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U3992 ( .A(n940), .B(n922), .Z(z[27]) );
  XOR U3993 ( .A(n933), .B(z[26]), .Z(z[28]) );
  AND U3994 ( .A(x[24]), .B(n923), .Z(n927) );
  XNOR U3995 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U3996 ( .A(n927), .B(n926), .Z(n942) );
  XOR U3997 ( .A(n928), .B(x[25]), .Z(n929) );
  NANDN U3998 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U3999 ( .A(n932), .B(n931), .Z(n936) );
  XNOR U4000 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U4001 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U4002 ( .A(n942), .B(n937), .Z(z[29]) );
  XNOR U4003 ( .A(n939), .B(n938), .Z(z[2]) );
  XNOR U4004 ( .A(n941), .B(n940), .Z(z[30]) );
  XOR U4005 ( .A(n942), .B(z[25]), .Z(z[31]) );
  XOR U4006 ( .A(x[35]), .B(x[33]), .Z(n945) );
  XNOR U4007 ( .A(x[32]), .B(x[38]), .Z(n944) );
  XOR U4008 ( .A(n944), .B(x[34]), .Z(n943) );
  XNOR U4009 ( .A(n945), .B(n943), .Z(n980) );
  XNOR U4010 ( .A(x[37]), .B(n944), .Z(n1053) );
  XOR U4011 ( .A(n1053), .B(x[36]), .Z(n1023) );
  IV U4012 ( .A(n1023), .Z(n954) );
  XNOR U4013 ( .A(x[39]), .B(x[36]), .Z(n948) );
  XNOR U4014 ( .A(n945), .B(n948), .Z(n1008) );
  NOR U4015 ( .A(n954), .B(n1008), .Z(n947) );
  XNOR U4016 ( .A(n1053), .B(x[39]), .Z(n1039) );
  XNOR U4017 ( .A(x[34]), .B(n1039), .Z(n963) );
  XNOR U4018 ( .A(x[33]), .B(n963), .Z(n958) );
  AND U4019 ( .A(x[32]), .B(n958), .Z(n946) );
  XNOR U4020 ( .A(n947), .B(n946), .Z(n951) );
  XNOR U4021 ( .A(n980), .B(n1039), .Z(n970) );
  IV U4022 ( .A(n980), .Z(n965) );
  XNOR U4023 ( .A(x[32]), .B(n965), .Z(n985) );
  IV U4024 ( .A(n948), .Z(n1013) );
  AND U4025 ( .A(n985), .B(n1013), .Z(n953) );
  IV U4026 ( .A(n1053), .Z(n972) );
  XNOR U4027 ( .A(n980), .B(n972), .Z(n1002) );
  XOR U4028 ( .A(n1002), .B(n1008), .Z(n1005) );
  XOR U4029 ( .A(x[34]), .B(x[36]), .Z(n1015) );
  NAND U4030 ( .A(n1005), .B(n1015), .Z(n949) );
  XNOR U4031 ( .A(n953), .B(n949), .Z(n974) );
  XNOR U4032 ( .A(n970), .B(n974), .Z(n950) );
  XNOR U4033 ( .A(n951), .B(n950), .Z(n997) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1029) );
  XNOR U4035 ( .A(x[32]), .B(n1008), .Z(n1009) );
  XNOR U4036 ( .A(n1053), .B(n1009), .Z(n1000) );
  NAND U4037 ( .A(n1029), .B(n1000), .Z(n952) );
  XNOR U4038 ( .A(n953), .B(n952), .Z(n966) );
  IV U4039 ( .A(n958), .Z(n1012) );
  XNOR U4040 ( .A(n1012), .B(n954), .Z(n1019) );
  AND U4041 ( .A(n1008), .B(n1019), .Z(n956) );
  AND U4042 ( .A(x[32]), .B(n1023), .Z(n955) );
  XNOR U4043 ( .A(n956), .B(n955), .Z(n957) );
  NANDN U4044 ( .A(n1009), .B(n957), .Z(n961) );
  NAND U4045 ( .A(x[32]), .B(n1008), .Z(n959) );
  OR U4046 ( .A(n959), .B(n958), .Z(n960) );
  NAND U4047 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U4048 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U4049 ( .A(n966), .B(n964), .Z(n986) );
  IV U4050 ( .A(n986), .Z(n993) );
  AND U4051 ( .A(n1039), .B(n965), .Z(n968) );
  XOR U4052 ( .A(x[33]), .B(x[39]), .Z(n1041) );
  AND U4053 ( .A(n1002), .B(n1041), .Z(n971) );
  XNOR U4054 ( .A(n971), .B(n966), .Z(n967) );
  XNOR U4055 ( .A(n968), .B(n967), .Z(n992) );
  NANDN U4056 ( .A(n993), .B(n992), .Z(n969) );
  NAND U4057 ( .A(n997), .B(n969), .Z(n979) );
  XNOR U4058 ( .A(n971), .B(n970), .Z(n976) );
  ANDN U4059 ( .B(n972), .A(x[33]), .Z(n973) );
  XNOR U4060 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U4061 ( .A(n976), .B(n975), .Z(n989) );
  XOR U4062 ( .A(n992), .B(n989), .Z(n977) );
  NAND U4063 ( .A(n993), .B(n977), .Z(n978) );
  NAND U4064 ( .A(n979), .B(n978), .Z(n1038) );
  ANDN U4065 ( .B(n980), .A(n1038), .Z(n1004) );
  IV U4066 ( .A(n989), .Z(n995) );
  XOR U4067 ( .A(n997), .B(n993), .Z(n981) );
  NANDN U4068 ( .A(n995), .B(n981), .Z(n984) );
  NANDN U4069 ( .A(n993), .B(n995), .Z(n982) );
  NANDN U4070 ( .A(n992), .B(n982), .Z(n983) );
  NAND U4071 ( .A(n984), .B(n983), .Z(n1048) );
  XNOR U4072 ( .A(n1038), .B(n1048), .Z(n1014) );
  AND U4073 ( .A(n985), .B(n1014), .Z(n1007) );
  OR U4074 ( .A(n992), .B(n989), .Z(n991) );
  ANDN U4075 ( .B(n992), .A(n986), .Z(n987) );
  XNOR U4076 ( .A(n987), .B(n997), .Z(n988) );
  NAND U4077 ( .A(n989), .B(n988), .Z(n990) );
  NAND U4078 ( .A(n991), .B(n990), .Z(n1011) );
  NAND U4079 ( .A(n993), .B(n997), .Z(n999) );
  NAND U4080 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U4081 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U4082 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4083 ( .A(n999), .B(n998), .Z(n1055) );
  NAND U4084 ( .A(n1030), .B(n1000), .Z(n1001) );
  XNOR U4085 ( .A(n1007), .B(n1001), .Z(n1050) );
  XOR U4086 ( .A(n1038), .B(n1055), .Z(n1040) );
  AND U4087 ( .A(n1002), .B(n1040), .Z(n1025) );
  XNOR U4088 ( .A(n1050), .B(n1025), .Z(n1003) );
  XNOR U4089 ( .A(n1004), .B(n1003), .Z(n1058) );
  NAND U4090 ( .A(n1016), .B(n1005), .Z(n1006) );
  XNOR U4091 ( .A(n1007), .B(n1006), .Z(n1033) );
  AND U4092 ( .A(n1008), .B(n1018), .Z(n1049) );
  NANDN U4093 ( .A(n1009), .B(n1011), .Z(n1010) );
  XNOR U4094 ( .A(n1049), .B(n1010), .Z(n1037) );
  XNOR U4095 ( .A(n1033), .B(n1037), .Z(n1022) );
  XOR U4096 ( .A(n1058), .B(n1022), .Z(z[32]) );
  AND U4097 ( .A(n1012), .B(n1011), .Z(n1021) );
  AND U4098 ( .A(n1014), .B(n1013), .Z(n1032) );
  NAND U4099 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U4100 ( .A(n1032), .B(n1017), .Z(n1059) );
  AND U4101 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U4102 ( .A(n1059), .B(n1026), .Z(n1020) );
  XNOR U4103 ( .A(n1021), .B(n1020), .Z(n1046) );
  XNOR U4104 ( .A(n1046), .B(n1022), .Z(n1064) );
  AND U4105 ( .A(n1023), .B(n1048), .Z(n1028) );
  NANDN U4106 ( .A(n1055), .B(n1053), .Z(n1024) );
  XNOR U4107 ( .A(n1025), .B(n1024), .Z(n1036) );
  XNOR U4108 ( .A(n1026), .B(n1036), .Z(n1027) );
  XNOR U4109 ( .A(n1028), .B(n1027), .Z(n1035) );
  NAND U4110 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U4111 ( .A(n1032), .B(n1031), .Z(n1042) );
  XNOR U4112 ( .A(n1033), .B(n1042), .Z(n1034) );
  XNOR U4113 ( .A(n1035), .B(n1034), .Z(n1045) );
  XNOR U4114 ( .A(n1064), .B(n1045), .Z(z[33]) );
  XNOR U4115 ( .A(n1037), .B(n1036), .Z(z[34]) );
  NOR U4116 ( .A(n1039), .B(n1038), .Z(n1044) );
  AND U4117 ( .A(n1041), .B(n1040), .Z(n1057) );
  XNOR U4118 ( .A(n1042), .B(n1057), .Z(n1043) );
  XNOR U4119 ( .A(n1044), .B(n1043), .Z(n1063) );
  XOR U4120 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U4121 ( .A(n1063), .B(n1047), .Z(z[35]) );
  XOR U4122 ( .A(n1058), .B(z[34]), .Z(z[36]) );
  AND U4123 ( .A(x[32]), .B(n1048), .Z(n1052) );
  XNOR U4124 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U4125 ( .A(n1052), .B(n1051), .Z(n1065) );
  XOR U4126 ( .A(n1053), .B(x[33]), .Z(n1054) );
  NANDN U4127 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U4128 ( .A(n1057), .B(n1056), .Z(n1061) );
  XNOR U4129 ( .A(n1059), .B(n1058), .Z(n1060) );
  XNOR U4130 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U4131 ( .A(n1065), .B(n1062), .Z(z[37]) );
  XNOR U4132 ( .A(n1064), .B(n1063), .Z(z[38]) );
  XOR U4133 ( .A(n1065), .B(z[33]), .Z(z[39]) );
  NOR U4134 ( .A(n1067), .B(n1066), .Z(n1072) );
  AND U4135 ( .A(n1069), .B(n1068), .Z(n1436) );
  XNOR U4136 ( .A(n1070), .B(n1436), .Z(n1071) );
  XNOR U4137 ( .A(n1072), .B(n1071), .Z(n1580) );
  XOR U4138 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U4139 ( .A(n1580), .B(n1075), .Z(z[3]) );
  XOR U4140 ( .A(x[43]), .B(x[41]), .Z(n1078) );
  XNOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1077) );
  XOR U4142 ( .A(n1077), .B(x[42]), .Z(n1076) );
  XNOR U4143 ( .A(n1078), .B(n1076), .Z(n1113) );
  XNOR U4144 ( .A(x[45]), .B(n1077), .Z(n1186) );
  XOR U4145 ( .A(n1186), .B(x[44]), .Z(n1156) );
  IV U4146 ( .A(n1156), .Z(n1087) );
  XNOR U4147 ( .A(x[47]), .B(x[44]), .Z(n1081) );
  XNOR U4148 ( .A(n1078), .B(n1081), .Z(n1141) );
  NOR U4149 ( .A(n1087), .B(n1141), .Z(n1080) );
  XNOR U4150 ( .A(n1186), .B(x[47]), .Z(n1172) );
  XNOR U4151 ( .A(x[42]), .B(n1172), .Z(n1096) );
  XNOR U4152 ( .A(x[41]), .B(n1096), .Z(n1091) );
  AND U4153 ( .A(x[40]), .B(n1091), .Z(n1079) );
  XNOR U4154 ( .A(n1080), .B(n1079), .Z(n1084) );
  XNOR U4155 ( .A(n1113), .B(n1172), .Z(n1103) );
  IV U4156 ( .A(n1113), .Z(n1098) );
  XNOR U4157 ( .A(x[40]), .B(n1098), .Z(n1118) );
  IV U4158 ( .A(n1081), .Z(n1146) );
  AND U4159 ( .A(n1118), .B(n1146), .Z(n1086) );
  IV U4160 ( .A(n1186), .Z(n1105) );
  XNOR U4161 ( .A(n1113), .B(n1105), .Z(n1135) );
  XOR U4162 ( .A(n1135), .B(n1141), .Z(n1138) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1148) );
  NAND U4164 ( .A(n1138), .B(n1148), .Z(n1082) );
  XNOR U4165 ( .A(n1086), .B(n1082), .Z(n1107) );
  XNOR U4166 ( .A(n1103), .B(n1107), .Z(n1083) );
  XNOR U4167 ( .A(n1084), .B(n1083), .Z(n1130) );
  XOR U4168 ( .A(x[42]), .B(x[47]), .Z(n1162) );
  XNOR U4169 ( .A(x[40]), .B(n1141), .Z(n1142) );
  XNOR U4170 ( .A(n1186), .B(n1142), .Z(n1133) );
  NAND U4171 ( .A(n1162), .B(n1133), .Z(n1085) );
  XNOR U4172 ( .A(n1086), .B(n1085), .Z(n1099) );
  IV U4173 ( .A(n1091), .Z(n1145) );
  XNOR U4174 ( .A(n1145), .B(n1087), .Z(n1152) );
  AND U4175 ( .A(n1141), .B(n1152), .Z(n1089) );
  AND U4176 ( .A(x[40]), .B(n1156), .Z(n1088) );
  XNOR U4177 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U4178 ( .A(n1142), .B(n1090), .Z(n1094) );
  NAND U4179 ( .A(x[40]), .B(n1141), .Z(n1092) );
  OR U4180 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U4181 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U4182 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U4183 ( .A(n1099), .B(n1097), .Z(n1119) );
  IV U4184 ( .A(n1119), .Z(n1126) );
  AND U4185 ( .A(n1172), .B(n1098), .Z(n1101) );
  XOR U4186 ( .A(x[41]), .B(x[47]), .Z(n1174) );
  AND U4187 ( .A(n1135), .B(n1174), .Z(n1104) );
  XNOR U4188 ( .A(n1104), .B(n1099), .Z(n1100) );
  XNOR U4189 ( .A(n1101), .B(n1100), .Z(n1125) );
  NANDN U4190 ( .A(n1126), .B(n1125), .Z(n1102) );
  NAND U4191 ( .A(n1130), .B(n1102), .Z(n1112) );
  XNOR U4192 ( .A(n1104), .B(n1103), .Z(n1109) );
  ANDN U4193 ( .B(n1105), .A(x[41]), .Z(n1106) );
  XNOR U4194 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U4195 ( .A(n1109), .B(n1108), .Z(n1122) );
  XOR U4196 ( .A(n1125), .B(n1122), .Z(n1110) );
  NAND U4197 ( .A(n1126), .B(n1110), .Z(n1111) );
  NAND U4198 ( .A(n1112), .B(n1111), .Z(n1171) );
  ANDN U4199 ( .B(n1113), .A(n1171), .Z(n1137) );
  IV U4200 ( .A(n1122), .Z(n1128) );
  XOR U4201 ( .A(n1130), .B(n1126), .Z(n1114) );
  NANDN U4202 ( .A(n1128), .B(n1114), .Z(n1117) );
  NANDN U4203 ( .A(n1126), .B(n1128), .Z(n1115) );
  NANDN U4204 ( .A(n1125), .B(n1115), .Z(n1116) );
  NAND U4205 ( .A(n1117), .B(n1116), .Z(n1181) );
  XNOR U4206 ( .A(n1171), .B(n1181), .Z(n1147) );
  AND U4207 ( .A(n1118), .B(n1147), .Z(n1140) );
  OR U4208 ( .A(n1125), .B(n1122), .Z(n1124) );
  ANDN U4209 ( .B(n1125), .A(n1119), .Z(n1120) );
  XNOR U4210 ( .A(n1120), .B(n1130), .Z(n1121) );
  NAND U4211 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U4212 ( .A(n1124), .B(n1123), .Z(n1144) );
  NAND U4213 ( .A(n1126), .B(n1130), .Z(n1132) );
  NAND U4214 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U4215 ( .A(n1128), .B(n1127), .Z(n1129) );
  NANDN U4216 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U4217 ( .A(n1132), .B(n1131), .Z(n1188) );
  NAND U4218 ( .A(n1163), .B(n1133), .Z(n1134) );
  XNOR U4219 ( .A(n1140), .B(n1134), .Z(n1183) );
  XOR U4220 ( .A(n1171), .B(n1188), .Z(n1173) );
  AND U4221 ( .A(n1135), .B(n1173), .Z(n1158) );
  XNOR U4222 ( .A(n1183), .B(n1158), .Z(n1136) );
  XNOR U4223 ( .A(n1137), .B(n1136), .Z(n1191) );
  NAND U4224 ( .A(n1149), .B(n1138), .Z(n1139) );
  XNOR U4225 ( .A(n1140), .B(n1139), .Z(n1166) );
  AND U4226 ( .A(n1141), .B(n1151), .Z(n1182) );
  NANDN U4227 ( .A(n1142), .B(n1144), .Z(n1143) );
  XNOR U4228 ( .A(n1182), .B(n1143), .Z(n1170) );
  XNOR U4229 ( .A(n1166), .B(n1170), .Z(n1155) );
  XOR U4230 ( .A(n1191), .B(n1155), .Z(z[40]) );
  AND U4231 ( .A(n1145), .B(n1144), .Z(n1154) );
  AND U4232 ( .A(n1147), .B(n1146), .Z(n1165) );
  NAND U4233 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U4234 ( .A(n1165), .B(n1150), .Z(n1192) );
  AND U4235 ( .A(n1152), .B(n1151), .Z(n1159) );
  XNOR U4236 ( .A(n1192), .B(n1159), .Z(n1153) );
  XNOR U4237 ( .A(n1154), .B(n1153), .Z(n1179) );
  XNOR U4238 ( .A(n1179), .B(n1155), .Z(n1197) );
  AND U4239 ( .A(n1156), .B(n1181), .Z(n1161) );
  NANDN U4240 ( .A(n1188), .B(n1186), .Z(n1157) );
  XNOR U4241 ( .A(n1158), .B(n1157), .Z(n1169) );
  XNOR U4242 ( .A(n1159), .B(n1169), .Z(n1160) );
  XNOR U4243 ( .A(n1161), .B(n1160), .Z(n1168) );
  NAND U4244 ( .A(n1163), .B(n1162), .Z(n1164) );
  XNOR U4245 ( .A(n1165), .B(n1164), .Z(n1175) );
  XNOR U4246 ( .A(n1166), .B(n1175), .Z(n1167) );
  XNOR U4247 ( .A(n1168), .B(n1167), .Z(n1178) );
  XNOR U4248 ( .A(n1197), .B(n1178), .Z(z[41]) );
  XNOR U4249 ( .A(n1170), .B(n1169), .Z(z[42]) );
  NOR U4250 ( .A(n1172), .B(n1171), .Z(n1177) );
  AND U4251 ( .A(n1174), .B(n1173), .Z(n1190) );
  XNOR U4252 ( .A(n1175), .B(n1190), .Z(n1176) );
  XNOR U4253 ( .A(n1177), .B(n1176), .Z(n1196) );
  XOR U4254 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4255 ( .A(n1196), .B(n1180), .Z(z[43]) );
  XOR U4256 ( .A(n1191), .B(z[42]), .Z(z[44]) );
  AND U4257 ( .A(x[40]), .B(n1181), .Z(n1185) );
  XNOR U4258 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U4259 ( .A(n1185), .B(n1184), .Z(n1198) );
  XOR U4260 ( .A(n1186), .B(x[41]), .Z(n1187) );
  NANDN U4261 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U4262 ( .A(n1190), .B(n1189), .Z(n1194) );
  XNOR U4263 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U4264 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U4265 ( .A(n1198), .B(n1195), .Z(z[45]) );
  XNOR U4266 ( .A(n1197), .B(n1196), .Z(z[46]) );
  XOR U4267 ( .A(n1198), .B(z[41]), .Z(z[47]) );
  XOR U4268 ( .A(x[51]), .B(x[49]), .Z(n1201) );
  XNOR U4269 ( .A(x[48]), .B(x[54]), .Z(n1200) );
  XOR U4270 ( .A(n1200), .B(x[50]), .Z(n1199) );
  XNOR U4271 ( .A(n1201), .B(n1199), .Z(n1236) );
  XNOR U4272 ( .A(x[53]), .B(n1200), .Z(n1309) );
  XOR U4273 ( .A(n1309), .B(x[52]), .Z(n1279) );
  IV U4274 ( .A(n1279), .Z(n1210) );
  XNOR U4275 ( .A(x[55]), .B(x[52]), .Z(n1204) );
  XNOR U4276 ( .A(n1201), .B(n1204), .Z(n1264) );
  NOR U4277 ( .A(n1210), .B(n1264), .Z(n1203) );
  XNOR U4278 ( .A(n1309), .B(x[55]), .Z(n1295) );
  XNOR U4279 ( .A(x[50]), .B(n1295), .Z(n1219) );
  XNOR U4280 ( .A(x[49]), .B(n1219), .Z(n1214) );
  AND U4281 ( .A(x[48]), .B(n1214), .Z(n1202) );
  XNOR U4282 ( .A(n1203), .B(n1202), .Z(n1207) );
  XNOR U4283 ( .A(n1236), .B(n1295), .Z(n1226) );
  IV U4284 ( .A(n1236), .Z(n1221) );
  XNOR U4285 ( .A(x[48]), .B(n1221), .Z(n1241) );
  IV U4286 ( .A(n1204), .Z(n1269) );
  AND U4287 ( .A(n1241), .B(n1269), .Z(n1209) );
  IV U4288 ( .A(n1309), .Z(n1228) );
  XNOR U4289 ( .A(n1236), .B(n1228), .Z(n1258) );
  XOR U4290 ( .A(n1258), .B(n1264), .Z(n1261) );
  XOR U4291 ( .A(x[50]), .B(x[52]), .Z(n1271) );
  NAND U4292 ( .A(n1261), .B(n1271), .Z(n1205) );
  XNOR U4293 ( .A(n1209), .B(n1205), .Z(n1230) );
  XNOR U4294 ( .A(n1226), .B(n1230), .Z(n1206) );
  XNOR U4295 ( .A(n1207), .B(n1206), .Z(n1253) );
  XOR U4296 ( .A(x[50]), .B(x[55]), .Z(n1285) );
  XNOR U4297 ( .A(x[48]), .B(n1264), .Z(n1265) );
  XNOR U4298 ( .A(n1309), .B(n1265), .Z(n1256) );
  NAND U4299 ( .A(n1285), .B(n1256), .Z(n1208) );
  XNOR U4300 ( .A(n1209), .B(n1208), .Z(n1222) );
  IV U4301 ( .A(n1214), .Z(n1268) );
  XNOR U4302 ( .A(n1268), .B(n1210), .Z(n1275) );
  AND U4303 ( .A(n1264), .B(n1275), .Z(n1212) );
  AND U4304 ( .A(x[48]), .B(n1279), .Z(n1211) );
  XNOR U4305 ( .A(n1212), .B(n1211), .Z(n1213) );
  NANDN U4306 ( .A(n1265), .B(n1213), .Z(n1217) );
  NAND U4307 ( .A(x[48]), .B(n1264), .Z(n1215) );
  OR U4308 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4309 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U4310 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U4311 ( .A(n1222), .B(n1220), .Z(n1242) );
  IV U4312 ( .A(n1242), .Z(n1249) );
  AND U4313 ( .A(n1295), .B(n1221), .Z(n1224) );
  XOR U4314 ( .A(x[49]), .B(x[55]), .Z(n1297) );
  AND U4315 ( .A(n1258), .B(n1297), .Z(n1227) );
  XNOR U4316 ( .A(n1227), .B(n1222), .Z(n1223) );
  XNOR U4317 ( .A(n1224), .B(n1223), .Z(n1248) );
  NANDN U4318 ( .A(n1249), .B(n1248), .Z(n1225) );
  NAND U4319 ( .A(n1253), .B(n1225), .Z(n1235) );
  XNOR U4320 ( .A(n1227), .B(n1226), .Z(n1232) );
  ANDN U4321 ( .B(n1228), .A(x[49]), .Z(n1229) );
  XNOR U4322 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U4323 ( .A(n1232), .B(n1231), .Z(n1245) );
  XOR U4324 ( .A(n1248), .B(n1245), .Z(n1233) );
  NAND U4325 ( .A(n1249), .B(n1233), .Z(n1234) );
  NAND U4326 ( .A(n1235), .B(n1234), .Z(n1294) );
  ANDN U4327 ( .B(n1236), .A(n1294), .Z(n1260) );
  IV U4328 ( .A(n1245), .Z(n1251) );
  XOR U4329 ( .A(n1253), .B(n1249), .Z(n1237) );
  NANDN U4330 ( .A(n1251), .B(n1237), .Z(n1240) );
  NANDN U4331 ( .A(n1249), .B(n1251), .Z(n1238) );
  NANDN U4332 ( .A(n1248), .B(n1238), .Z(n1239) );
  NAND U4333 ( .A(n1240), .B(n1239), .Z(n1304) );
  XNOR U4334 ( .A(n1294), .B(n1304), .Z(n1270) );
  AND U4335 ( .A(n1241), .B(n1270), .Z(n1263) );
  OR U4336 ( .A(n1248), .B(n1245), .Z(n1247) );
  ANDN U4337 ( .B(n1248), .A(n1242), .Z(n1243) );
  XNOR U4338 ( .A(n1243), .B(n1253), .Z(n1244) );
  NAND U4339 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U4340 ( .A(n1247), .B(n1246), .Z(n1267) );
  NAND U4341 ( .A(n1249), .B(n1253), .Z(n1255) );
  NAND U4342 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U4343 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U4344 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U4345 ( .A(n1255), .B(n1254), .Z(n1311) );
  NAND U4346 ( .A(n1286), .B(n1256), .Z(n1257) );
  XNOR U4347 ( .A(n1263), .B(n1257), .Z(n1306) );
  XOR U4348 ( .A(n1294), .B(n1311), .Z(n1296) );
  AND U4349 ( .A(n1258), .B(n1296), .Z(n1281) );
  XNOR U4350 ( .A(n1306), .B(n1281), .Z(n1259) );
  XNOR U4351 ( .A(n1260), .B(n1259), .Z(n1314) );
  NAND U4352 ( .A(n1272), .B(n1261), .Z(n1262) );
  XNOR U4353 ( .A(n1263), .B(n1262), .Z(n1289) );
  AND U4354 ( .A(n1264), .B(n1274), .Z(n1305) );
  NANDN U4355 ( .A(n1265), .B(n1267), .Z(n1266) );
  XNOR U4356 ( .A(n1305), .B(n1266), .Z(n1293) );
  XNOR U4357 ( .A(n1289), .B(n1293), .Z(n1278) );
  XOR U4358 ( .A(n1314), .B(n1278), .Z(z[48]) );
  AND U4359 ( .A(n1268), .B(n1267), .Z(n1277) );
  AND U4360 ( .A(n1270), .B(n1269), .Z(n1288) );
  NAND U4361 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U4362 ( .A(n1288), .B(n1273), .Z(n1315) );
  AND U4363 ( .A(n1275), .B(n1274), .Z(n1282) );
  XNOR U4364 ( .A(n1315), .B(n1282), .Z(n1276) );
  XNOR U4365 ( .A(n1277), .B(n1276), .Z(n1302) );
  XNOR U4366 ( .A(n1302), .B(n1278), .Z(n1320) );
  AND U4367 ( .A(n1279), .B(n1304), .Z(n1284) );
  NANDN U4368 ( .A(n1311), .B(n1309), .Z(n1280) );
  XNOR U4369 ( .A(n1281), .B(n1280), .Z(n1292) );
  XNOR U4370 ( .A(n1282), .B(n1292), .Z(n1283) );
  XNOR U4371 ( .A(n1284), .B(n1283), .Z(n1291) );
  NAND U4372 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U4373 ( .A(n1288), .B(n1287), .Z(n1298) );
  XNOR U4374 ( .A(n1289), .B(n1298), .Z(n1290) );
  XNOR U4375 ( .A(n1291), .B(n1290), .Z(n1301) );
  XNOR U4376 ( .A(n1320), .B(n1301), .Z(z[49]) );
  XOR U4377 ( .A(n1437), .B(z[2]), .Z(z[4]) );
  XNOR U4378 ( .A(n1293), .B(n1292), .Z(z[50]) );
  NOR U4379 ( .A(n1295), .B(n1294), .Z(n1300) );
  AND U4380 ( .A(n1297), .B(n1296), .Z(n1313) );
  XNOR U4381 ( .A(n1298), .B(n1313), .Z(n1299) );
  XNOR U4382 ( .A(n1300), .B(n1299), .Z(n1319) );
  XOR U4383 ( .A(n1302), .B(n1301), .Z(n1303) );
  XNOR U4384 ( .A(n1319), .B(n1303), .Z(z[51]) );
  XOR U4385 ( .A(n1314), .B(z[50]), .Z(z[52]) );
  AND U4386 ( .A(x[48]), .B(n1304), .Z(n1308) );
  XNOR U4387 ( .A(n1306), .B(n1305), .Z(n1307) );
  XNOR U4388 ( .A(n1308), .B(n1307), .Z(n1321) );
  XOR U4389 ( .A(n1309), .B(x[49]), .Z(n1310) );
  NANDN U4390 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U4391 ( .A(n1313), .B(n1312), .Z(n1317) );
  XNOR U4392 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U4393 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U4394 ( .A(n1321), .B(n1318), .Z(z[53]) );
  XNOR U4395 ( .A(n1320), .B(n1319), .Z(z[54]) );
  XOR U4396 ( .A(n1321), .B(z[49]), .Z(z[55]) );
  XOR U4397 ( .A(x[59]), .B(x[57]), .Z(n1324) );
  XNOR U4398 ( .A(x[56]), .B(x[62]), .Z(n1323) );
  XOR U4399 ( .A(n1323), .B(x[58]), .Z(n1322) );
  XNOR U4400 ( .A(n1324), .B(n1322), .Z(n1359) );
  XNOR U4401 ( .A(x[61]), .B(n1323), .Z(n1447) );
  XOR U4402 ( .A(n1447), .B(x[60]), .Z(n1402) );
  IV U4403 ( .A(n1402), .Z(n1333) );
  XNOR U4404 ( .A(x[63]), .B(x[60]), .Z(n1327) );
  XNOR U4405 ( .A(n1324), .B(n1327), .Z(n1387) );
  NOR U4406 ( .A(n1333), .B(n1387), .Z(n1326) );
  XNOR U4407 ( .A(n1447), .B(x[63]), .Z(n1418) );
  XNOR U4408 ( .A(x[58]), .B(n1418), .Z(n1342) );
  XNOR U4409 ( .A(x[57]), .B(n1342), .Z(n1337) );
  AND U4410 ( .A(x[56]), .B(n1337), .Z(n1325) );
  XNOR U4411 ( .A(n1326), .B(n1325), .Z(n1330) );
  XNOR U4412 ( .A(n1359), .B(n1418), .Z(n1349) );
  IV U4413 ( .A(n1359), .Z(n1344) );
  XNOR U4414 ( .A(x[56]), .B(n1344), .Z(n1364) );
  IV U4415 ( .A(n1327), .Z(n1392) );
  AND U4416 ( .A(n1364), .B(n1392), .Z(n1332) );
  IV U4417 ( .A(n1447), .Z(n1351) );
  XNOR U4418 ( .A(n1359), .B(n1351), .Z(n1381) );
  XOR U4419 ( .A(n1381), .B(n1387), .Z(n1384) );
  XOR U4420 ( .A(x[58]), .B(x[60]), .Z(n1394) );
  NAND U4421 ( .A(n1384), .B(n1394), .Z(n1328) );
  XNOR U4422 ( .A(n1332), .B(n1328), .Z(n1353) );
  XNOR U4423 ( .A(n1349), .B(n1353), .Z(n1329) );
  XNOR U4424 ( .A(n1330), .B(n1329), .Z(n1376) );
  XOR U4425 ( .A(x[58]), .B(x[63]), .Z(n1408) );
  XNOR U4426 ( .A(x[56]), .B(n1387), .Z(n1388) );
  XNOR U4427 ( .A(n1447), .B(n1388), .Z(n1379) );
  NAND U4428 ( .A(n1408), .B(n1379), .Z(n1331) );
  XNOR U4429 ( .A(n1332), .B(n1331), .Z(n1345) );
  IV U4430 ( .A(n1337), .Z(n1391) );
  XNOR U4431 ( .A(n1391), .B(n1333), .Z(n1398) );
  AND U4432 ( .A(n1387), .B(n1398), .Z(n1335) );
  AND U4433 ( .A(x[56]), .B(n1402), .Z(n1334) );
  XNOR U4434 ( .A(n1335), .B(n1334), .Z(n1336) );
  NANDN U4435 ( .A(n1388), .B(n1336), .Z(n1340) );
  NAND U4436 ( .A(x[56]), .B(n1387), .Z(n1338) );
  OR U4437 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U4438 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4439 ( .A(n1342), .B(n1341), .Z(n1343) );
  XNOR U4440 ( .A(n1345), .B(n1343), .Z(n1365) );
  IV U4441 ( .A(n1365), .Z(n1372) );
  AND U4442 ( .A(n1418), .B(n1344), .Z(n1347) );
  XOR U4443 ( .A(x[57]), .B(x[63]), .Z(n1420) );
  AND U4444 ( .A(n1381), .B(n1420), .Z(n1350) );
  XNOR U4445 ( .A(n1350), .B(n1345), .Z(n1346) );
  XNOR U4446 ( .A(n1347), .B(n1346), .Z(n1371) );
  NANDN U4447 ( .A(n1372), .B(n1371), .Z(n1348) );
  NAND U4448 ( .A(n1376), .B(n1348), .Z(n1358) );
  XNOR U4449 ( .A(n1350), .B(n1349), .Z(n1355) );
  ANDN U4450 ( .B(n1351), .A(x[57]), .Z(n1352) );
  XNOR U4451 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U4452 ( .A(n1355), .B(n1354), .Z(n1368) );
  XOR U4453 ( .A(n1371), .B(n1368), .Z(n1356) );
  NAND U4454 ( .A(n1372), .B(n1356), .Z(n1357) );
  NAND U4455 ( .A(n1358), .B(n1357), .Z(n1417) );
  ANDN U4456 ( .B(n1359), .A(n1417), .Z(n1383) );
  IV U4457 ( .A(n1368), .Z(n1374) );
  XOR U4458 ( .A(n1376), .B(n1372), .Z(n1360) );
  NANDN U4459 ( .A(n1374), .B(n1360), .Z(n1363) );
  NANDN U4460 ( .A(n1372), .B(n1374), .Z(n1361) );
  NANDN U4461 ( .A(n1371), .B(n1361), .Z(n1362) );
  NAND U4462 ( .A(n1363), .B(n1362), .Z(n1442) );
  XNOR U4463 ( .A(n1417), .B(n1442), .Z(n1393) );
  AND U4464 ( .A(n1364), .B(n1393), .Z(n1386) );
  OR U4465 ( .A(n1371), .B(n1368), .Z(n1370) );
  ANDN U4466 ( .B(n1371), .A(n1365), .Z(n1366) );
  XNOR U4467 ( .A(n1366), .B(n1376), .Z(n1367) );
  NAND U4468 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U4469 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U4470 ( .A(n1372), .B(n1376), .Z(n1378) );
  NAND U4471 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4472 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U4473 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U4474 ( .A(n1378), .B(n1377), .Z(n1449) );
  NAND U4475 ( .A(n1409), .B(n1379), .Z(n1380) );
  XNOR U4476 ( .A(n1386), .B(n1380), .Z(n1444) );
  XOR U4477 ( .A(n1417), .B(n1449), .Z(n1419) );
  AND U4478 ( .A(n1381), .B(n1419), .Z(n1404) );
  XNOR U4479 ( .A(n1444), .B(n1404), .Z(n1382) );
  XNOR U4480 ( .A(n1383), .B(n1382), .Z(n1452) );
  NAND U4481 ( .A(n1395), .B(n1384), .Z(n1385) );
  XNOR U4482 ( .A(n1386), .B(n1385), .Z(n1412) );
  AND U4483 ( .A(n1387), .B(n1397), .Z(n1443) );
  NANDN U4484 ( .A(n1388), .B(n1390), .Z(n1389) );
  XNOR U4485 ( .A(n1443), .B(n1389), .Z(n1416) );
  XNOR U4486 ( .A(n1412), .B(n1416), .Z(n1401) );
  XOR U4487 ( .A(n1452), .B(n1401), .Z(z[56]) );
  AND U4488 ( .A(n1391), .B(n1390), .Z(n1400) );
  AND U4489 ( .A(n1393), .B(n1392), .Z(n1411) );
  NAND U4490 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U4491 ( .A(n1411), .B(n1396), .Z(n1453) );
  AND U4492 ( .A(n1398), .B(n1397), .Z(n1405) );
  XNOR U4493 ( .A(n1453), .B(n1405), .Z(n1399) );
  XNOR U4494 ( .A(n1400), .B(n1399), .Z(n1425) );
  XNOR U4495 ( .A(n1425), .B(n1401), .Z(n1458) );
  AND U4496 ( .A(n1402), .B(n1442), .Z(n1407) );
  NANDN U4497 ( .A(n1449), .B(n1447), .Z(n1403) );
  XNOR U4498 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U4499 ( .A(n1405), .B(n1415), .Z(n1406) );
  XNOR U4500 ( .A(n1407), .B(n1406), .Z(n1414) );
  NAND U4501 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U4502 ( .A(n1411), .B(n1410), .Z(n1421) );
  XNOR U4503 ( .A(n1412), .B(n1421), .Z(n1413) );
  XNOR U4504 ( .A(n1414), .B(n1413), .Z(n1424) );
  XNOR U4505 ( .A(n1458), .B(n1424), .Z(z[57]) );
  XNOR U4506 ( .A(n1416), .B(n1415), .Z(z[58]) );
  NOR U4507 ( .A(n1418), .B(n1417), .Z(n1423) );
  AND U4508 ( .A(n1420), .B(n1419), .Z(n1451) );
  XNOR U4509 ( .A(n1421), .B(n1451), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1457) );
  XOR U4511 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U4512 ( .A(n1457), .B(n1426), .Z(z[59]) );
  AND U4513 ( .A(x[0]), .B(n1427), .Z(n1431) );
  XNOR U4514 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U4515 ( .A(n1431), .B(n1430), .Z(n1708) );
  XOR U4516 ( .A(n1432), .B(x[1]), .Z(n1433) );
  NANDN U4517 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U4518 ( .A(n1436), .B(n1435), .Z(n1440) );
  XNOR U4519 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U4520 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U4521 ( .A(n1708), .B(n1441), .Z(z[5]) );
  XOR U4522 ( .A(n1452), .B(z[58]), .Z(z[60]) );
  AND U4523 ( .A(x[56]), .B(n1442), .Z(n1446) );
  XNOR U4524 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U4525 ( .A(n1446), .B(n1445), .Z(n1459) );
  XOR U4526 ( .A(n1447), .B(x[57]), .Z(n1448) );
  NANDN U4527 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U4528 ( .A(n1451), .B(n1450), .Z(n1455) );
  XNOR U4529 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U4530 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U4531 ( .A(n1459), .B(n1456), .Z(z[61]) );
  XNOR U4532 ( .A(n1458), .B(n1457), .Z(z[62]) );
  XOR U4533 ( .A(n1459), .B(z[57]), .Z(z[63]) );
  XOR U4534 ( .A(x[67]), .B(x[65]), .Z(n1462) );
  XNOR U4535 ( .A(x[64]), .B(x[70]), .Z(n1461) );
  XOR U4536 ( .A(n1461), .B(x[66]), .Z(n1460) );
  XNOR U4537 ( .A(n1462), .B(n1460), .Z(n1497) );
  XNOR U4538 ( .A(x[69]), .B(n1461), .Z(n1570) );
  XOR U4539 ( .A(n1570), .B(x[68]), .Z(n1540) );
  IV U4540 ( .A(n1540), .Z(n1471) );
  XNOR U4541 ( .A(x[71]), .B(x[68]), .Z(n1465) );
  XNOR U4542 ( .A(n1462), .B(n1465), .Z(n1525) );
  NOR U4543 ( .A(n1471), .B(n1525), .Z(n1464) );
  XNOR U4544 ( .A(n1570), .B(x[71]), .Z(n1556) );
  XNOR U4545 ( .A(x[66]), .B(n1556), .Z(n1480) );
  XNOR U4546 ( .A(x[65]), .B(n1480), .Z(n1475) );
  AND U4547 ( .A(x[64]), .B(n1475), .Z(n1463) );
  XNOR U4548 ( .A(n1464), .B(n1463), .Z(n1468) );
  XNOR U4549 ( .A(n1497), .B(n1556), .Z(n1487) );
  IV U4550 ( .A(n1497), .Z(n1482) );
  XNOR U4551 ( .A(x[64]), .B(n1482), .Z(n1502) );
  IV U4552 ( .A(n1465), .Z(n1530) );
  AND U4553 ( .A(n1502), .B(n1530), .Z(n1470) );
  IV U4554 ( .A(n1570), .Z(n1489) );
  XNOR U4555 ( .A(n1497), .B(n1489), .Z(n1519) );
  XOR U4556 ( .A(n1519), .B(n1525), .Z(n1522) );
  XOR U4557 ( .A(x[66]), .B(x[68]), .Z(n1532) );
  NAND U4558 ( .A(n1522), .B(n1532), .Z(n1466) );
  XNOR U4559 ( .A(n1470), .B(n1466), .Z(n1491) );
  XNOR U4560 ( .A(n1487), .B(n1491), .Z(n1467) );
  XNOR U4561 ( .A(n1468), .B(n1467), .Z(n1514) );
  XOR U4562 ( .A(x[66]), .B(x[71]), .Z(n1546) );
  XNOR U4563 ( .A(x[64]), .B(n1525), .Z(n1526) );
  XNOR U4564 ( .A(n1570), .B(n1526), .Z(n1517) );
  NAND U4565 ( .A(n1546), .B(n1517), .Z(n1469) );
  XNOR U4566 ( .A(n1470), .B(n1469), .Z(n1483) );
  IV U4567 ( .A(n1475), .Z(n1529) );
  XNOR U4568 ( .A(n1529), .B(n1471), .Z(n1536) );
  AND U4569 ( .A(n1525), .B(n1536), .Z(n1473) );
  AND U4570 ( .A(x[64]), .B(n1540), .Z(n1472) );
  XNOR U4571 ( .A(n1473), .B(n1472), .Z(n1474) );
  NANDN U4572 ( .A(n1526), .B(n1474), .Z(n1478) );
  NAND U4573 ( .A(x[64]), .B(n1525), .Z(n1476) );
  OR U4574 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U4575 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4576 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR U4577 ( .A(n1483), .B(n1481), .Z(n1503) );
  IV U4578 ( .A(n1503), .Z(n1510) );
  AND U4579 ( .A(n1556), .B(n1482), .Z(n1485) );
  XOR U4580 ( .A(x[65]), .B(x[71]), .Z(n1558) );
  AND U4581 ( .A(n1519), .B(n1558), .Z(n1488) );
  XNOR U4582 ( .A(n1488), .B(n1483), .Z(n1484) );
  XNOR U4583 ( .A(n1485), .B(n1484), .Z(n1509) );
  NANDN U4584 ( .A(n1510), .B(n1509), .Z(n1486) );
  NAND U4585 ( .A(n1514), .B(n1486), .Z(n1496) );
  XNOR U4586 ( .A(n1488), .B(n1487), .Z(n1493) );
  ANDN U4587 ( .B(n1489), .A(x[65]), .Z(n1490) );
  XNOR U4588 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U4589 ( .A(n1493), .B(n1492), .Z(n1506) );
  XOR U4590 ( .A(n1509), .B(n1506), .Z(n1494) );
  NAND U4591 ( .A(n1510), .B(n1494), .Z(n1495) );
  NAND U4592 ( .A(n1496), .B(n1495), .Z(n1555) );
  ANDN U4593 ( .B(n1497), .A(n1555), .Z(n1521) );
  IV U4594 ( .A(n1506), .Z(n1512) );
  XOR U4595 ( .A(n1514), .B(n1510), .Z(n1498) );
  NANDN U4596 ( .A(n1512), .B(n1498), .Z(n1501) );
  NANDN U4597 ( .A(n1510), .B(n1512), .Z(n1499) );
  NANDN U4598 ( .A(n1509), .B(n1499), .Z(n1500) );
  NAND U4599 ( .A(n1501), .B(n1500), .Z(n1565) );
  XNOR U4600 ( .A(n1555), .B(n1565), .Z(n1531) );
  AND U4601 ( .A(n1502), .B(n1531), .Z(n1524) );
  OR U4602 ( .A(n1509), .B(n1506), .Z(n1508) );
  ANDN U4603 ( .B(n1509), .A(n1503), .Z(n1504) );
  XNOR U4604 ( .A(n1504), .B(n1514), .Z(n1505) );
  NAND U4605 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U4606 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U4607 ( .A(n1510), .B(n1514), .Z(n1516) );
  NAND U4608 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4609 ( .A(n1512), .B(n1511), .Z(n1513) );
  NANDN U4610 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U4611 ( .A(n1516), .B(n1515), .Z(n1572) );
  NAND U4612 ( .A(n1547), .B(n1517), .Z(n1518) );
  XNOR U4613 ( .A(n1524), .B(n1518), .Z(n1567) );
  XOR U4614 ( .A(n1555), .B(n1572), .Z(n1557) );
  AND U4615 ( .A(n1519), .B(n1557), .Z(n1542) );
  XNOR U4616 ( .A(n1567), .B(n1542), .Z(n1520) );
  XNOR U4617 ( .A(n1521), .B(n1520), .Z(n1575) );
  NAND U4618 ( .A(n1533), .B(n1522), .Z(n1523) );
  XNOR U4619 ( .A(n1524), .B(n1523), .Z(n1550) );
  AND U4620 ( .A(n1525), .B(n1535), .Z(n1566) );
  NANDN U4621 ( .A(n1526), .B(n1528), .Z(n1527) );
  XNOR U4622 ( .A(n1566), .B(n1527), .Z(n1554) );
  XNOR U4623 ( .A(n1550), .B(n1554), .Z(n1539) );
  XOR U4624 ( .A(n1575), .B(n1539), .Z(z[64]) );
  AND U4625 ( .A(n1529), .B(n1528), .Z(n1538) );
  AND U4626 ( .A(n1531), .B(n1530), .Z(n1549) );
  NAND U4627 ( .A(n1533), .B(n1532), .Z(n1534) );
  XNOR U4628 ( .A(n1549), .B(n1534), .Z(n1576) );
  AND U4629 ( .A(n1536), .B(n1535), .Z(n1543) );
  XNOR U4630 ( .A(n1576), .B(n1543), .Z(n1537) );
  XNOR U4631 ( .A(n1538), .B(n1537), .Z(n1563) );
  XNOR U4632 ( .A(n1563), .B(n1539), .Z(n1583) );
  AND U4633 ( .A(n1540), .B(n1565), .Z(n1545) );
  NANDN U4634 ( .A(n1572), .B(n1570), .Z(n1541) );
  XNOR U4635 ( .A(n1542), .B(n1541), .Z(n1553) );
  XNOR U4636 ( .A(n1543), .B(n1553), .Z(n1544) );
  XNOR U4637 ( .A(n1545), .B(n1544), .Z(n1552) );
  NAND U4638 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U4639 ( .A(n1549), .B(n1548), .Z(n1559) );
  XNOR U4640 ( .A(n1550), .B(n1559), .Z(n1551) );
  XNOR U4641 ( .A(n1552), .B(n1551), .Z(n1562) );
  XNOR U4642 ( .A(n1583), .B(n1562), .Z(z[65]) );
  XNOR U4643 ( .A(n1554), .B(n1553), .Z(z[66]) );
  NOR U4644 ( .A(n1556), .B(n1555), .Z(n1561) );
  AND U4645 ( .A(n1558), .B(n1557), .Z(n1574) );
  XNOR U4646 ( .A(n1559), .B(n1574), .Z(n1560) );
  XNOR U4647 ( .A(n1561), .B(n1560), .Z(n1582) );
  XOR U4648 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U4649 ( .A(n1582), .B(n1564), .Z(z[67]) );
  XOR U4650 ( .A(n1575), .B(z[66]), .Z(z[68]) );
  AND U4651 ( .A(x[64]), .B(n1565), .Z(n1569) );
  XNOR U4652 ( .A(n1567), .B(n1566), .Z(n1568) );
  XNOR U4653 ( .A(n1569), .B(n1568), .Z(n1584) );
  XOR U4654 ( .A(n1570), .B(x[65]), .Z(n1571) );
  NANDN U4655 ( .A(n1572), .B(n1571), .Z(n1573) );
  XNOR U4656 ( .A(n1574), .B(n1573), .Z(n1578) );
  XNOR U4657 ( .A(n1576), .B(n1575), .Z(n1577) );
  XNOR U4658 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U4659 ( .A(n1584), .B(n1579), .Z(z[69]) );
  XNOR U4660 ( .A(n1581), .B(n1580), .Z(z[6]) );
  XNOR U4661 ( .A(n1583), .B(n1582), .Z(z[70]) );
  XOR U4662 ( .A(n1584), .B(z[65]), .Z(z[71]) );
  XOR U4663 ( .A(x[75]), .B(x[73]), .Z(n1587) );
  XNOR U4664 ( .A(x[72]), .B(x[78]), .Z(n1586) );
  XOR U4665 ( .A(n1586), .B(x[74]), .Z(n1585) );
  XNOR U4666 ( .A(n1587), .B(n1585), .Z(n1622) );
  XNOR U4667 ( .A(x[77]), .B(n1586), .Z(n1695) );
  XOR U4668 ( .A(n1695), .B(x[76]), .Z(n1665) );
  IV U4669 ( .A(n1665), .Z(n1596) );
  XNOR U4670 ( .A(x[79]), .B(x[76]), .Z(n1590) );
  XNOR U4671 ( .A(n1587), .B(n1590), .Z(n1650) );
  NOR U4672 ( .A(n1596), .B(n1650), .Z(n1589) );
  XNOR U4673 ( .A(n1695), .B(x[79]), .Z(n1681) );
  XNOR U4674 ( .A(x[74]), .B(n1681), .Z(n1605) );
  XNOR U4675 ( .A(x[73]), .B(n1605), .Z(n1600) );
  AND U4676 ( .A(x[72]), .B(n1600), .Z(n1588) );
  XNOR U4677 ( .A(n1589), .B(n1588), .Z(n1593) );
  XNOR U4678 ( .A(n1622), .B(n1681), .Z(n1612) );
  IV U4679 ( .A(n1622), .Z(n1607) );
  XNOR U4680 ( .A(x[72]), .B(n1607), .Z(n1627) );
  IV U4681 ( .A(n1590), .Z(n1655) );
  AND U4682 ( .A(n1627), .B(n1655), .Z(n1595) );
  IV U4683 ( .A(n1695), .Z(n1614) );
  XNOR U4684 ( .A(n1622), .B(n1614), .Z(n1644) );
  XOR U4685 ( .A(n1644), .B(n1650), .Z(n1647) );
  XOR U4686 ( .A(x[74]), .B(x[76]), .Z(n1657) );
  NAND U4687 ( .A(n1647), .B(n1657), .Z(n1591) );
  XNOR U4688 ( .A(n1595), .B(n1591), .Z(n1616) );
  XNOR U4689 ( .A(n1612), .B(n1616), .Z(n1592) );
  XNOR U4690 ( .A(n1593), .B(n1592), .Z(n1639) );
  XOR U4691 ( .A(x[74]), .B(x[79]), .Z(n1671) );
  XNOR U4692 ( .A(x[72]), .B(n1650), .Z(n1651) );
  XNOR U4693 ( .A(n1695), .B(n1651), .Z(n1642) );
  NAND U4694 ( .A(n1671), .B(n1642), .Z(n1594) );
  XNOR U4695 ( .A(n1595), .B(n1594), .Z(n1608) );
  IV U4696 ( .A(n1600), .Z(n1654) );
  XNOR U4697 ( .A(n1654), .B(n1596), .Z(n1661) );
  AND U4698 ( .A(n1650), .B(n1661), .Z(n1598) );
  AND U4699 ( .A(x[72]), .B(n1665), .Z(n1597) );
  XNOR U4700 ( .A(n1598), .B(n1597), .Z(n1599) );
  NANDN U4701 ( .A(n1651), .B(n1599), .Z(n1603) );
  NAND U4702 ( .A(x[72]), .B(n1650), .Z(n1601) );
  OR U4703 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U4704 ( .A(n1603), .B(n1602), .Z(n1604) );
  XNOR U4705 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U4706 ( .A(n1608), .B(n1606), .Z(n1628) );
  IV U4707 ( .A(n1628), .Z(n1635) );
  AND U4708 ( .A(n1681), .B(n1607), .Z(n1610) );
  XOR U4709 ( .A(x[73]), .B(x[79]), .Z(n1683) );
  AND U4710 ( .A(n1644), .B(n1683), .Z(n1613) );
  XNOR U4711 ( .A(n1613), .B(n1608), .Z(n1609) );
  XNOR U4712 ( .A(n1610), .B(n1609), .Z(n1634) );
  NANDN U4713 ( .A(n1635), .B(n1634), .Z(n1611) );
  NAND U4714 ( .A(n1639), .B(n1611), .Z(n1621) );
  XNOR U4715 ( .A(n1613), .B(n1612), .Z(n1618) );
  ANDN U4716 ( .B(n1614), .A(x[73]), .Z(n1615) );
  XNOR U4717 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4718 ( .A(n1618), .B(n1617), .Z(n1631) );
  XOR U4719 ( .A(n1634), .B(n1631), .Z(n1619) );
  NAND U4720 ( .A(n1635), .B(n1619), .Z(n1620) );
  NAND U4721 ( .A(n1621), .B(n1620), .Z(n1680) );
  ANDN U4722 ( .B(n1622), .A(n1680), .Z(n1646) );
  IV U4723 ( .A(n1631), .Z(n1637) );
  XOR U4724 ( .A(n1639), .B(n1635), .Z(n1623) );
  NANDN U4725 ( .A(n1637), .B(n1623), .Z(n1626) );
  NANDN U4726 ( .A(n1635), .B(n1637), .Z(n1624) );
  NANDN U4727 ( .A(n1634), .B(n1624), .Z(n1625) );
  NAND U4728 ( .A(n1626), .B(n1625), .Z(n1690) );
  XNOR U4729 ( .A(n1680), .B(n1690), .Z(n1656) );
  AND U4730 ( .A(n1627), .B(n1656), .Z(n1649) );
  OR U4731 ( .A(n1634), .B(n1631), .Z(n1633) );
  ANDN U4732 ( .B(n1634), .A(n1628), .Z(n1629) );
  XNOR U4733 ( .A(n1629), .B(n1639), .Z(n1630) );
  NAND U4734 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U4735 ( .A(n1633), .B(n1632), .Z(n1653) );
  NAND U4736 ( .A(n1635), .B(n1639), .Z(n1641) );
  NAND U4737 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U4738 ( .A(n1637), .B(n1636), .Z(n1638) );
  NANDN U4739 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U4740 ( .A(n1641), .B(n1640), .Z(n1697) );
  NAND U4741 ( .A(n1672), .B(n1642), .Z(n1643) );
  XNOR U4742 ( .A(n1649), .B(n1643), .Z(n1692) );
  XOR U4743 ( .A(n1680), .B(n1697), .Z(n1682) );
  AND U4744 ( .A(n1644), .B(n1682), .Z(n1667) );
  XNOR U4745 ( .A(n1692), .B(n1667), .Z(n1645) );
  XNOR U4746 ( .A(n1646), .B(n1645), .Z(n1700) );
  NAND U4747 ( .A(n1658), .B(n1647), .Z(n1648) );
  XNOR U4748 ( .A(n1649), .B(n1648), .Z(n1675) );
  AND U4749 ( .A(n1650), .B(n1660), .Z(n1691) );
  NANDN U4750 ( .A(n1651), .B(n1653), .Z(n1652) );
  XNOR U4751 ( .A(n1691), .B(n1652), .Z(n1679) );
  XNOR U4752 ( .A(n1675), .B(n1679), .Z(n1664) );
  XOR U4753 ( .A(n1700), .B(n1664), .Z(z[72]) );
  AND U4754 ( .A(n1654), .B(n1653), .Z(n1663) );
  AND U4755 ( .A(n1656), .B(n1655), .Z(n1674) );
  NAND U4756 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U4757 ( .A(n1674), .B(n1659), .Z(n1701) );
  AND U4758 ( .A(n1661), .B(n1660), .Z(n1668) );
  XNOR U4759 ( .A(n1701), .B(n1668), .Z(n1662) );
  XNOR U4760 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U4761 ( .A(n1688), .B(n1664), .Z(n1706) );
  AND U4762 ( .A(n1665), .B(n1690), .Z(n1670) );
  NANDN U4763 ( .A(n1697), .B(n1695), .Z(n1666) );
  XNOR U4764 ( .A(n1667), .B(n1666), .Z(n1678) );
  XNOR U4765 ( .A(n1668), .B(n1678), .Z(n1669) );
  XNOR U4766 ( .A(n1670), .B(n1669), .Z(n1677) );
  NAND U4767 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR U4768 ( .A(n1674), .B(n1673), .Z(n1684) );
  XNOR U4769 ( .A(n1675), .B(n1684), .Z(n1676) );
  XNOR U4770 ( .A(n1677), .B(n1676), .Z(n1687) );
  XNOR U4771 ( .A(n1706), .B(n1687), .Z(z[73]) );
  XNOR U4772 ( .A(n1679), .B(n1678), .Z(z[74]) );
  NOR U4773 ( .A(n1681), .B(n1680), .Z(n1686) );
  AND U4774 ( .A(n1683), .B(n1682), .Z(n1699) );
  XNOR U4775 ( .A(n1684), .B(n1699), .Z(n1685) );
  XNOR U4776 ( .A(n1686), .B(n1685), .Z(n1705) );
  XOR U4777 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4778 ( .A(n1705), .B(n1689), .Z(z[75]) );
  XOR U4779 ( .A(n1700), .B(z[74]), .Z(z[76]) );
  AND U4780 ( .A(x[72]), .B(n1690), .Z(n1694) );
  XNOR U4781 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4782 ( .A(n1694), .B(n1693), .Z(n1707) );
  XOR U4783 ( .A(n1695), .B(x[73]), .Z(n1696) );
  NANDN U4784 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U4785 ( .A(n1699), .B(n1698), .Z(n1703) );
  XNOR U4786 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U4787 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U4788 ( .A(n1707), .B(n1704), .Z(z[77]) );
  XNOR U4789 ( .A(n1706), .B(n1705), .Z(z[78]) );
  XOR U4790 ( .A(n1707), .B(z[73]), .Z(z[79]) );
  XOR U4791 ( .A(n1708), .B(z[1]), .Z(z[7]) );
  XOR U4792 ( .A(x[83]), .B(x[81]), .Z(n1711) );
  XNOR U4793 ( .A(x[80]), .B(x[86]), .Z(n1710) );
  XOR U4794 ( .A(n1710), .B(x[82]), .Z(n1709) );
  XNOR U4795 ( .A(n1711), .B(n1709), .Z(n1746) );
  XNOR U4796 ( .A(x[85]), .B(n1710), .Z(n1819) );
  XOR U4797 ( .A(n1819), .B(x[84]), .Z(n1789) );
  IV U4798 ( .A(n1789), .Z(n1720) );
  XNOR U4799 ( .A(x[87]), .B(x[84]), .Z(n1714) );
  XNOR U4800 ( .A(n1711), .B(n1714), .Z(n1774) );
  NOR U4801 ( .A(n1720), .B(n1774), .Z(n1713) );
  XNOR U4802 ( .A(n1819), .B(x[87]), .Z(n1805) );
  XNOR U4803 ( .A(x[82]), .B(n1805), .Z(n1729) );
  XNOR U4804 ( .A(x[81]), .B(n1729), .Z(n1724) );
  AND U4805 ( .A(x[80]), .B(n1724), .Z(n1712) );
  XNOR U4806 ( .A(n1713), .B(n1712), .Z(n1717) );
  XNOR U4807 ( .A(n1746), .B(n1805), .Z(n1736) );
  IV U4808 ( .A(n1746), .Z(n1731) );
  XNOR U4809 ( .A(x[80]), .B(n1731), .Z(n1751) );
  IV U4810 ( .A(n1714), .Z(n1779) );
  AND U4811 ( .A(n1751), .B(n1779), .Z(n1719) );
  IV U4812 ( .A(n1819), .Z(n1738) );
  XNOR U4813 ( .A(n1746), .B(n1738), .Z(n1768) );
  XOR U4814 ( .A(n1768), .B(n1774), .Z(n1771) );
  XOR U4815 ( .A(x[82]), .B(x[84]), .Z(n1781) );
  NAND U4816 ( .A(n1771), .B(n1781), .Z(n1715) );
  XNOR U4817 ( .A(n1719), .B(n1715), .Z(n1740) );
  XNOR U4818 ( .A(n1736), .B(n1740), .Z(n1716) );
  XNOR U4819 ( .A(n1717), .B(n1716), .Z(n1763) );
  XOR U4820 ( .A(x[82]), .B(x[87]), .Z(n1795) );
  XNOR U4821 ( .A(x[80]), .B(n1774), .Z(n1775) );
  XNOR U4822 ( .A(n1819), .B(n1775), .Z(n1766) );
  NAND U4823 ( .A(n1795), .B(n1766), .Z(n1718) );
  XNOR U4824 ( .A(n1719), .B(n1718), .Z(n1732) );
  IV U4825 ( .A(n1724), .Z(n1778) );
  XNOR U4826 ( .A(n1778), .B(n1720), .Z(n1785) );
  AND U4827 ( .A(n1774), .B(n1785), .Z(n1722) );
  AND U4828 ( .A(x[80]), .B(n1789), .Z(n1721) );
  XNOR U4829 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U4830 ( .A(n1775), .B(n1723), .Z(n1727) );
  NAND U4831 ( .A(x[80]), .B(n1774), .Z(n1725) );
  OR U4832 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U4833 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U4834 ( .A(n1729), .B(n1728), .Z(n1730) );
  XNOR U4835 ( .A(n1732), .B(n1730), .Z(n1752) );
  IV U4836 ( .A(n1752), .Z(n1759) );
  AND U4837 ( .A(n1805), .B(n1731), .Z(n1734) );
  XOR U4838 ( .A(x[81]), .B(x[87]), .Z(n1807) );
  AND U4839 ( .A(n1768), .B(n1807), .Z(n1737) );
  XNOR U4840 ( .A(n1737), .B(n1732), .Z(n1733) );
  XNOR U4841 ( .A(n1734), .B(n1733), .Z(n1758) );
  NANDN U4842 ( .A(n1759), .B(n1758), .Z(n1735) );
  NAND U4843 ( .A(n1763), .B(n1735), .Z(n1745) );
  XNOR U4844 ( .A(n1737), .B(n1736), .Z(n1742) );
  ANDN U4845 ( .B(n1738), .A(x[81]), .Z(n1739) );
  XNOR U4846 ( .A(n1740), .B(n1739), .Z(n1741) );
  XNOR U4847 ( .A(n1742), .B(n1741), .Z(n1755) );
  XOR U4848 ( .A(n1758), .B(n1755), .Z(n1743) );
  NAND U4849 ( .A(n1759), .B(n1743), .Z(n1744) );
  NAND U4850 ( .A(n1745), .B(n1744), .Z(n1804) );
  ANDN U4851 ( .B(n1746), .A(n1804), .Z(n1770) );
  IV U4852 ( .A(n1755), .Z(n1761) );
  XOR U4853 ( .A(n1763), .B(n1759), .Z(n1747) );
  NANDN U4854 ( .A(n1761), .B(n1747), .Z(n1750) );
  NANDN U4855 ( .A(n1759), .B(n1761), .Z(n1748) );
  NANDN U4856 ( .A(n1758), .B(n1748), .Z(n1749) );
  NAND U4857 ( .A(n1750), .B(n1749), .Z(n1814) );
  XNOR U4858 ( .A(n1804), .B(n1814), .Z(n1780) );
  AND U4859 ( .A(n1751), .B(n1780), .Z(n1773) );
  OR U4860 ( .A(n1758), .B(n1755), .Z(n1757) );
  ANDN U4861 ( .B(n1758), .A(n1752), .Z(n1753) );
  XNOR U4862 ( .A(n1753), .B(n1763), .Z(n1754) );
  NAND U4863 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U4864 ( .A(n1757), .B(n1756), .Z(n1777) );
  NAND U4865 ( .A(n1759), .B(n1763), .Z(n1765) );
  NAND U4866 ( .A(n1759), .B(n1758), .Z(n1760) );
  XNOR U4867 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U4868 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1821) );
  NAND U4870 ( .A(n1796), .B(n1766), .Z(n1767) );
  XNOR U4871 ( .A(n1773), .B(n1767), .Z(n1816) );
  XOR U4872 ( .A(n1804), .B(n1821), .Z(n1806) );
  AND U4873 ( .A(n1768), .B(n1806), .Z(n1791) );
  XNOR U4874 ( .A(n1816), .B(n1791), .Z(n1769) );
  XNOR U4875 ( .A(n1770), .B(n1769), .Z(n1824) );
  NAND U4876 ( .A(n1782), .B(n1771), .Z(n1772) );
  XNOR U4877 ( .A(n1773), .B(n1772), .Z(n1799) );
  AND U4878 ( .A(n1774), .B(n1784), .Z(n1815) );
  NANDN U4879 ( .A(n1775), .B(n1777), .Z(n1776) );
  XNOR U4880 ( .A(n1815), .B(n1776), .Z(n1803) );
  XNOR U4881 ( .A(n1799), .B(n1803), .Z(n1788) );
  XOR U4882 ( .A(n1824), .B(n1788), .Z(z[80]) );
  AND U4883 ( .A(n1778), .B(n1777), .Z(n1787) );
  AND U4884 ( .A(n1780), .B(n1779), .Z(n1798) );
  NAND U4885 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U4886 ( .A(n1798), .B(n1783), .Z(n1825) );
  AND U4887 ( .A(n1785), .B(n1784), .Z(n1792) );
  XNOR U4888 ( .A(n1825), .B(n1792), .Z(n1786) );
  XNOR U4889 ( .A(n1787), .B(n1786), .Z(n1812) );
  XNOR U4890 ( .A(n1812), .B(n1788), .Z(n1830) );
  AND U4891 ( .A(n1789), .B(n1814), .Z(n1794) );
  NANDN U4892 ( .A(n1821), .B(n1819), .Z(n1790) );
  XNOR U4893 ( .A(n1791), .B(n1790), .Z(n1802) );
  XNOR U4894 ( .A(n1792), .B(n1802), .Z(n1793) );
  XNOR U4895 ( .A(n1794), .B(n1793), .Z(n1801) );
  NAND U4896 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U4897 ( .A(n1798), .B(n1797), .Z(n1808) );
  XNOR U4898 ( .A(n1799), .B(n1808), .Z(n1800) );
  XNOR U4899 ( .A(n1801), .B(n1800), .Z(n1811) );
  XNOR U4900 ( .A(n1830), .B(n1811), .Z(z[81]) );
  XNOR U4901 ( .A(n1803), .B(n1802), .Z(z[82]) );
  NOR U4902 ( .A(n1805), .B(n1804), .Z(n1810) );
  AND U4903 ( .A(n1807), .B(n1806), .Z(n1823) );
  XNOR U4904 ( .A(n1808), .B(n1823), .Z(n1809) );
  XNOR U4905 ( .A(n1810), .B(n1809), .Z(n1829) );
  XOR U4906 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U4907 ( .A(n1829), .B(n1813), .Z(z[83]) );
  XOR U4908 ( .A(n1824), .B(z[82]), .Z(z[84]) );
  AND U4909 ( .A(x[80]), .B(n1814), .Z(n1818) );
  XNOR U4910 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U4911 ( .A(n1818), .B(n1817), .Z(n1831) );
  XOR U4912 ( .A(n1819), .B(x[81]), .Z(n1820) );
  NANDN U4913 ( .A(n1821), .B(n1820), .Z(n1822) );
  XNOR U4914 ( .A(n1823), .B(n1822), .Z(n1827) );
  XNOR U4915 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U4916 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U4917 ( .A(n1831), .B(n1828), .Z(z[85]) );
  XNOR U4918 ( .A(n1830), .B(n1829), .Z(z[86]) );
  XOR U4919 ( .A(n1831), .B(z[81]), .Z(z[87]) );
  XOR U4920 ( .A(x[91]), .B(x[89]), .Z(n1834) );
  XNOR U4921 ( .A(x[88]), .B(x[94]), .Z(n1833) );
  XOR U4922 ( .A(n1833), .B(x[90]), .Z(n1832) );
  XNOR U4923 ( .A(n1834), .B(n1832), .Z(n1869) );
  XNOR U4924 ( .A(x[93]), .B(n1833), .Z(n1944) );
  XOR U4925 ( .A(n1944), .B(x[92]), .Z(n1912) );
  IV U4926 ( .A(n1912), .Z(n1843) );
  XNOR U4927 ( .A(x[95]), .B(x[92]), .Z(n1837) );
  XNOR U4928 ( .A(n1834), .B(n1837), .Z(n1897) );
  NOR U4929 ( .A(n1843), .B(n1897), .Z(n1836) );
  XNOR U4930 ( .A(n1944), .B(x[95]), .Z(n1930) );
  XNOR U4931 ( .A(x[90]), .B(n1930), .Z(n1852) );
  XNOR U4932 ( .A(x[89]), .B(n1852), .Z(n1847) );
  AND U4933 ( .A(x[88]), .B(n1847), .Z(n1835) );
  XNOR U4934 ( .A(n1836), .B(n1835), .Z(n1840) );
  XNOR U4935 ( .A(n1869), .B(n1930), .Z(n1859) );
  IV U4936 ( .A(n1869), .Z(n1854) );
  XNOR U4937 ( .A(x[88]), .B(n1854), .Z(n1874) );
  IV U4938 ( .A(n1837), .Z(n1902) );
  AND U4939 ( .A(n1874), .B(n1902), .Z(n1842) );
  IV U4940 ( .A(n1944), .Z(n1861) );
  XNOR U4941 ( .A(n1869), .B(n1861), .Z(n1891) );
  XOR U4942 ( .A(n1891), .B(n1897), .Z(n1894) );
  XOR U4943 ( .A(x[90]), .B(x[92]), .Z(n1904) );
  NAND U4944 ( .A(n1894), .B(n1904), .Z(n1838) );
  XNOR U4945 ( .A(n1842), .B(n1838), .Z(n1863) );
  XNOR U4946 ( .A(n1859), .B(n1863), .Z(n1839) );
  XNOR U4947 ( .A(n1840), .B(n1839), .Z(n1886) );
  XOR U4948 ( .A(x[90]), .B(x[95]), .Z(n1918) );
  XNOR U4949 ( .A(x[88]), .B(n1897), .Z(n1898) );
  XNOR U4950 ( .A(n1944), .B(n1898), .Z(n1889) );
  NAND U4951 ( .A(n1918), .B(n1889), .Z(n1841) );
  XNOR U4952 ( .A(n1842), .B(n1841), .Z(n1855) );
  IV U4953 ( .A(n1847), .Z(n1901) );
  XNOR U4954 ( .A(n1901), .B(n1843), .Z(n1908) );
  AND U4955 ( .A(n1897), .B(n1908), .Z(n1845) );
  AND U4956 ( .A(x[88]), .B(n1912), .Z(n1844) );
  XNOR U4957 ( .A(n1845), .B(n1844), .Z(n1846) );
  NANDN U4958 ( .A(n1898), .B(n1846), .Z(n1850) );
  NAND U4959 ( .A(x[88]), .B(n1897), .Z(n1848) );
  OR U4960 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U4961 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U4962 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U4963 ( .A(n1855), .B(n1853), .Z(n1875) );
  IV U4964 ( .A(n1875), .Z(n1882) );
  AND U4965 ( .A(n1930), .B(n1854), .Z(n1857) );
  XOR U4966 ( .A(x[89]), .B(x[95]), .Z(n1932) );
  AND U4967 ( .A(n1891), .B(n1932), .Z(n1860) );
  XNOR U4968 ( .A(n1860), .B(n1855), .Z(n1856) );
  XNOR U4969 ( .A(n1857), .B(n1856), .Z(n1881) );
  NANDN U4970 ( .A(n1882), .B(n1881), .Z(n1858) );
  NAND U4971 ( .A(n1886), .B(n1858), .Z(n1868) );
  XNOR U4972 ( .A(n1860), .B(n1859), .Z(n1865) );
  ANDN U4973 ( .B(n1861), .A(x[89]), .Z(n1862) );
  XNOR U4974 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U4975 ( .A(n1865), .B(n1864), .Z(n1878) );
  XOR U4976 ( .A(n1881), .B(n1878), .Z(n1866) );
  NAND U4977 ( .A(n1882), .B(n1866), .Z(n1867) );
  NAND U4978 ( .A(n1868), .B(n1867), .Z(n1929) );
  ANDN U4979 ( .B(n1869), .A(n1929), .Z(n1893) );
  IV U4980 ( .A(n1878), .Z(n1884) );
  XOR U4981 ( .A(n1886), .B(n1882), .Z(n1870) );
  NANDN U4982 ( .A(n1884), .B(n1870), .Z(n1873) );
  NANDN U4983 ( .A(n1882), .B(n1884), .Z(n1871) );
  NANDN U4984 ( .A(n1881), .B(n1871), .Z(n1872) );
  NAND U4985 ( .A(n1873), .B(n1872), .Z(n1939) );
  XNOR U4986 ( .A(n1929), .B(n1939), .Z(n1903) );
  AND U4987 ( .A(n1874), .B(n1903), .Z(n1896) );
  OR U4988 ( .A(n1881), .B(n1878), .Z(n1880) );
  ANDN U4989 ( .B(n1881), .A(n1875), .Z(n1876) );
  XNOR U4990 ( .A(n1876), .B(n1886), .Z(n1877) );
  NAND U4991 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U4992 ( .A(n1880), .B(n1879), .Z(n1900) );
  NAND U4993 ( .A(n1882), .B(n1886), .Z(n1888) );
  NAND U4994 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U4995 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U4996 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4997 ( .A(n1888), .B(n1887), .Z(n1946) );
  NAND U4998 ( .A(n1919), .B(n1889), .Z(n1890) );
  XNOR U4999 ( .A(n1896), .B(n1890), .Z(n1941) );
  XOR U5000 ( .A(n1929), .B(n1946), .Z(n1931) );
  AND U5001 ( .A(n1891), .B(n1931), .Z(n1914) );
  XNOR U5002 ( .A(n1941), .B(n1914), .Z(n1892) );
  XNOR U5003 ( .A(n1893), .B(n1892), .Z(n1949) );
  NAND U5004 ( .A(n1905), .B(n1894), .Z(n1895) );
  XNOR U5005 ( .A(n1896), .B(n1895), .Z(n1922) );
  AND U5006 ( .A(n1897), .B(n1907), .Z(n1940) );
  NANDN U5007 ( .A(n1898), .B(n1900), .Z(n1899) );
  XNOR U5008 ( .A(n1940), .B(n1899), .Z(n1928) );
  XNOR U5009 ( .A(n1922), .B(n1928), .Z(n1911) );
  XOR U5010 ( .A(n1949), .B(n1911), .Z(z[88]) );
  AND U5011 ( .A(n1901), .B(n1900), .Z(n1910) );
  AND U5012 ( .A(n1903), .B(n1902), .Z(n1921) );
  NAND U5013 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U5014 ( .A(n1921), .B(n1906), .Z(n1950) );
  AND U5015 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U5016 ( .A(n1950), .B(n1915), .Z(n1909) );
  XNOR U5017 ( .A(n1910), .B(n1909), .Z(n1937) );
  XNOR U5018 ( .A(n1937), .B(n1911), .Z(n1955) );
  AND U5019 ( .A(n1912), .B(n1939), .Z(n1917) );
  NANDN U5020 ( .A(n1946), .B(n1944), .Z(n1913) );
  XNOR U5021 ( .A(n1914), .B(n1913), .Z(n1927) );
  XNOR U5022 ( .A(n1915), .B(n1927), .Z(n1916) );
  XNOR U5023 ( .A(n1917), .B(n1916), .Z(n1924) );
  NAND U5024 ( .A(n1919), .B(n1918), .Z(n1920) );
  XNOR U5025 ( .A(n1921), .B(n1920), .Z(n1933) );
  XNOR U5026 ( .A(n1922), .B(n1933), .Z(n1923) );
  XNOR U5027 ( .A(n1924), .B(n1923), .Z(n1936) );
  XNOR U5028 ( .A(n1955), .B(n1936), .Z(z[89]) );
  XOR U5029 ( .A(n1926), .B(n1925), .Z(z[8]) );
  XNOR U5030 ( .A(n1928), .B(n1927), .Z(z[90]) );
  NOR U5031 ( .A(n1930), .B(n1929), .Z(n1935) );
  AND U5032 ( .A(n1932), .B(n1931), .Z(n1948) );
  XNOR U5033 ( .A(n1933), .B(n1948), .Z(n1934) );
  XNOR U5034 ( .A(n1935), .B(n1934), .Z(n1954) );
  XOR U5035 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U5036 ( .A(n1954), .B(n1938), .Z(z[91]) );
  XOR U5037 ( .A(n1949), .B(z[90]), .Z(z[92]) );
  AND U5038 ( .A(x[88]), .B(n1939), .Z(n1943) );
  XNOR U5039 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5040 ( .A(n1943), .B(n1942), .Z(n1956) );
  XOR U5041 ( .A(n1944), .B(x[89]), .Z(n1945) );
  NANDN U5042 ( .A(n1946), .B(n1945), .Z(n1947) );
  XNOR U5043 ( .A(n1948), .B(n1947), .Z(n1952) );
  XNOR U5044 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U5045 ( .A(n1952), .B(n1951), .Z(n1953) );
  XNOR U5046 ( .A(n1956), .B(n1953), .Z(z[93]) );
  XNOR U5047 ( .A(n1955), .B(n1954), .Z(z[94]) );
  XOR U5048 ( .A(n1956), .B(z[89]), .Z(z[95]) );
  XOR U5049 ( .A(n1958), .B(n1957), .Z(z[96]) );
  XOR U5050 ( .A(n1960), .B(n1959), .Z(n1961) );
  XNOR U5051 ( .A(n1962), .B(n1961), .Z(z[99]) );
endmodule


module SubBytes_1 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;

  XOR U2962 ( .A(n1048), .B(n1011), .Z(n1018) );
  XOR U2963 ( .A(n1690), .B(n1653), .Z(n1660) );
  XOR U2964 ( .A(n467), .B(n430), .Z(n437) );
  XOR U2965 ( .A(n923), .B(n886), .Z(n893) );
  XOR U2966 ( .A(n1565), .B(n1528), .Z(n1535) );
  XOR U2967 ( .A(n290), .B(n253), .Z(n260) );
  XOR U2968 ( .A(n800), .B(n738), .Z(n745) );
  XOR U2969 ( .A(n1442), .B(n1390), .Z(n1397) );
  XOR U2970 ( .A(n1304), .B(n1267), .Z(n1274) );
  XOR U2971 ( .A(n1939), .B(n1900), .Z(n1907) );
  XOR U2972 ( .A(n1427), .B(n775), .Z(n782) );
  XOR U2973 ( .A(n1181), .B(n1144), .Z(n1151) );
  XOR U2974 ( .A(n1814), .B(n1777), .Z(n1784) );
  XOR U2975 ( .A(n622), .B(n585), .Z(n592) );
  XNOR U2976 ( .A(n1011), .B(n1055), .Z(n1030) );
  XNOR U2977 ( .A(n1653), .B(n1697), .Z(n1672) );
  XNOR U2978 ( .A(n430), .B(n474), .Z(n449) );
  XNOR U2979 ( .A(n886), .B(n930), .Z(n905) );
  XNOR U2980 ( .A(n1528), .B(n1572), .Z(n1547) );
  XNOR U2981 ( .A(n253), .B(n297), .Z(n272) );
  XNOR U2982 ( .A(n738), .B(n807), .Z(n757) );
  XNOR U2983 ( .A(n1390), .B(n1449), .Z(n1409) );
  NOR U2984 ( .A(n654), .B(x[9]), .Z(n1) );
  XNOR U2985 ( .A(n329), .B(n328), .Z(n2) );
  XNOR U2986 ( .A(n1), .B(n2), .Z(n3) );
  XNOR U2987 ( .A(n312), .B(n3), .Z(n345) );
  XNOR U2988 ( .A(n1267), .B(n1311), .Z(n1286) );
  XNOR U2989 ( .A(n1900), .B(n1946), .Z(n1919) );
  XNOR U2990 ( .A(n775), .B(n1434), .Z(n794) );
  XNOR U2991 ( .A(n1144), .B(n1188), .Z(n1163) );
  XNOR U2992 ( .A(n1777), .B(n1821), .Z(n1796) );
  XNOR U2993 ( .A(n585), .B(n629), .Z(n604) );
  XOR U2994 ( .A(n163), .B(n134), .Z(n157) );
  XOR U2995 ( .A(n77), .B(n78), .Z(n129) );
  XNOR U2996 ( .A(x[9]), .B(n323), .Z(n318) );
  XOR U2997 ( .A(n1030), .B(n1014), .Z(n1016) );
  XOR U2998 ( .A(n1672), .B(n1656), .Z(n1658) );
  XOR U2999 ( .A(n449), .B(n433), .Z(n435) );
  XOR U3000 ( .A(n905), .B(n889), .Z(n891) );
  XOR U3001 ( .A(n1547), .B(n1531), .Z(n1533) );
  XOR U3002 ( .A(n272), .B(n256), .Z(n258) );
  XOR U3003 ( .A(n757), .B(n741), .Z(n743) );
  XOR U3004 ( .A(n1409), .B(n1393), .Z(n1395) );
  XOR U3005 ( .A(n116), .B(n119), .Z(n4) );
  NANDN U3006 ( .A(n116), .B(n121), .Z(n5) );
  OR U3007 ( .A(n121), .B(n4), .Z(n6) );
  NANDN U3008 ( .A(n117), .B(n6), .Z(n7) );
  NAND U3009 ( .A(n5), .B(n7), .Z(n169) );
  XOR U3010 ( .A(n643), .B(n508), .Z(n511) );
  XOR U3011 ( .A(n1286), .B(n1270), .Z(n1272) );
  XOR U3012 ( .A(n1919), .B(n1903), .Z(n1905) );
  XOR U3013 ( .A(n794), .B(n778), .Z(n780) );
  XOR U3014 ( .A(n1163), .B(n1147), .Z(n1149) );
  XOR U3015 ( .A(n1796), .B(n1780), .Z(n1782) );
  XOR U3016 ( .A(n604), .B(n588), .Z(n590) );
  XOR U3017 ( .A(x[3]), .B(x[1]), .Z(n10) );
  XNOR U3018 ( .A(x[0]), .B(x[6]), .Z(n9) );
  XOR U3019 ( .A(n9), .B(x[2]), .Z(n8) );
  XNOR U3020 ( .A(n10), .B(n8), .Z(n45) );
  XNOR U3021 ( .A(x[5]), .B(n9), .Z(n1432) );
  XOR U3022 ( .A(n1432), .B(x[4]), .Z(n787) );
  IV U3023 ( .A(n787), .Z(n19) );
  XNOR U3024 ( .A(x[7]), .B(x[4]), .Z(n13) );
  XNOR U3025 ( .A(n10), .B(n13), .Z(n73) );
  NOR U3026 ( .A(n19), .B(n73), .Z(n12) );
  XNOR U3027 ( .A(n1432), .B(x[7]), .Z(n1067) );
  XNOR U3028 ( .A(x[2]), .B(n1067), .Z(n28) );
  XNOR U3029 ( .A(x[1]), .B(n28), .Z(n23) );
  AND U3030 ( .A(x[0]), .B(n23), .Z(n11) );
  XNOR U3031 ( .A(n12), .B(n11), .Z(n16) );
  XNOR U3032 ( .A(n45), .B(n1067), .Z(n35) );
  IV U3033 ( .A(n45), .Z(n30) );
  XNOR U3034 ( .A(x[0]), .B(n30), .Z(n50) );
  IV U3035 ( .A(n13), .Z(n777) );
  AND U3036 ( .A(n50), .B(n777), .Z(n18) );
  IV U3037 ( .A(n1432), .Z(n37) );
  XNOR U3038 ( .A(n45), .B(n37), .Z(n67) );
  XOR U3039 ( .A(n67), .B(n73), .Z(n70) );
  XOR U3040 ( .A(x[2]), .B(x[4]), .Z(n779) );
  NAND U3041 ( .A(n70), .B(n779), .Z(n14) );
  XNOR U3042 ( .A(n18), .B(n14), .Z(n39) );
  XNOR U3043 ( .A(n35), .B(n39), .Z(n15) );
  XNOR U3044 ( .A(n16), .B(n15), .Z(n62) );
  XOR U3045 ( .A(x[2]), .B(x[7]), .Z(n793) );
  XNOR U3046 ( .A(x[0]), .B(n73), .Z(n74) );
  XNOR U3047 ( .A(n1432), .B(n74), .Z(n65) );
  NAND U3048 ( .A(n793), .B(n65), .Z(n17) );
  XNOR U3049 ( .A(n18), .B(n17), .Z(n31) );
  IV U3050 ( .A(n23), .Z(n776) );
  XNOR U3051 ( .A(n776), .B(n19), .Z(n783) );
  AND U3052 ( .A(n73), .B(n783), .Z(n21) );
  AND U3053 ( .A(x[0]), .B(n787), .Z(n20) );
  XNOR U3054 ( .A(n21), .B(n20), .Z(n22) );
  NANDN U3055 ( .A(n74), .B(n22), .Z(n26) );
  NAND U3056 ( .A(x[0]), .B(n73), .Z(n24) );
  OR U3057 ( .A(n24), .B(n23), .Z(n25) );
  NAND U3058 ( .A(n26), .B(n25), .Z(n27) );
  XNOR U3059 ( .A(n28), .B(n27), .Z(n29) );
  XNOR U3060 ( .A(n31), .B(n29), .Z(n51) );
  IV U3061 ( .A(n51), .Z(n58) );
  AND U3062 ( .A(n1067), .B(n30), .Z(n33) );
  XOR U3063 ( .A(x[1]), .B(x[7]), .Z(n1069) );
  AND U3064 ( .A(n67), .B(n1069), .Z(n36) );
  XNOR U3065 ( .A(n36), .B(n31), .Z(n32) );
  XNOR U3066 ( .A(n33), .B(n32), .Z(n57) );
  NANDN U3067 ( .A(n58), .B(n57), .Z(n34) );
  NAND U3068 ( .A(n62), .B(n34), .Z(n44) );
  XNOR U3069 ( .A(n36), .B(n35), .Z(n41) );
  ANDN U3070 ( .B(n37), .A(x[1]), .Z(n38) );
  XNOR U3071 ( .A(n39), .B(n38), .Z(n40) );
  XNOR U3072 ( .A(n41), .B(n40), .Z(n54) );
  XOR U3073 ( .A(n57), .B(n54), .Z(n42) );
  NAND U3074 ( .A(n58), .B(n42), .Z(n43) );
  NAND U3075 ( .A(n44), .B(n43), .Z(n1066) );
  ANDN U3076 ( .B(n45), .A(n1066), .Z(n69) );
  IV U3077 ( .A(n54), .Z(n60) );
  XOR U3078 ( .A(n62), .B(n58), .Z(n46) );
  NANDN U3079 ( .A(n60), .B(n46), .Z(n49) );
  NANDN U3080 ( .A(n58), .B(n60), .Z(n47) );
  NANDN U3081 ( .A(n57), .B(n47), .Z(n48) );
  NAND U3082 ( .A(n49), .B(n48), .Z(n1427) );
  XNOR U3083 ( .A(n1066), .B(n1427), .Z(n778) );
  AND U3084 ( .A(n50), .B(n778), .Z(n72) );
  OR U3085 ( .A(n57), .B(n54), .Z(n56) );
  ANDN U3086 ( .B(n57), .A(n51), .Z(n52) );
  XNOR U3087 ( .A(n52), .B(n62), .Z(n53) );
  NAND U3088 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3089 ( .A(n56), .B(n55), .Z(n775) );
  NAND U3090 ( .A(n58), .B(n62), .Z(n64) );
  NAND U3091 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U3092 ( .A(n60), .B(n59), .Z(n61) );
  NANDN U3093 ( .A(n62), .B(n61), .Z(n63) );
  NAND U3094 ( .A(n64), .B(n63), .Z(n1434) );
  NAND U3095 ( .A(n794), .B(n65), .Z(n66) );
  XNOR U3096 ( .A(n72), .B(n66), .Z(n1429) );
  XOR U3097 ( .A(n1066), .B(n1434), .Z(n1068) );
  AND U3098 ( .A(n67), .B(n1068), .Z(n789) );
  XNOR U3099 ( .A(n1429), .B(n789), .Z(n68) );
  XNOR U3100 ( .A(n69), .B(n68), .Z(n1437) );
  NAND U3101 ( .A(n780), .B(n70), .Z(n71) );
  XNOR U3102 ( .A(n72), .B(n71), .Z(n797) );
  AND U3103 ( .A(n73), .B(n782), .Z(n1428) );
  NANDN U3104 ( .A(n74), .B(n775), .Z(n75) );
  XNOR U3105 ( .A(n1428), .B(n75), .Z(n939) );
  XNOR U3106 ( .A(n797), .B(n939), .Z(n786) );
  XOR U3107 ( .A(n1437), .B(n786), .Z(z[0]) );
  XOR U3108 ( .A(x[99]), .B(x[97]), .Z(n76) );
  XNOR U3109 ( .A(n76), .B(x[98]), .Z(n77) );
  XNOR U3110 ( .A(x[101]), .B(n77), .Z(n114) );
  XOR U3111 ( .A(x[98]), .B(x[100]), .Z(n135) );
  XNOR U3112 ( .A(x[102]), .B(n77), .Z(n128) );
  XOR U3113 ( .A(x[103]), .B(x[100]), .Z(n133) );
  XOR U3114 ( .A(n76), .B(n133), .Z(n124) );
  XNOR U3115 ( .A(x[96]), .B(n124), .Z(n93) );
  IV U3116 ( .A(n93), .Z(n125) );
  XNOR U3117 ( .A(x[102]), .B(x[96]), .Z(n78) );
  XNOR U3118 ( .A(x[101]), .B(n78), .Z(n139) );
  XOR U3119 ( .A(n125), .B(n139), .Z(n127) );
  XOR U3120 ( .A(n128), .B(n127), .Z(n156) );
  AND U3121 ( .A(n135), .B(n156), .Z(n80) );
  AND U3122 ( .A(n128), .B(n133), .Z(n86) );
  IV U3123 ( .A(n139), .Z(n102) );
  XNOR U3124 ( .A(x[103]), .B(n102), .Z(n161) );
  XOR U3125 ( .A(n129), .B(n161), .Z(n84) );
  XNOR U3126 ( .A(n86), .B(n84), .Z(n79) );
  XNOR U3127 ( .A(n80), .B(n79), .Z(n103) );
  XOR U3128 ( .A(x[98]), .B(n161), .Z(n98) );
  XOR U3129 ( .A(x[97]), .B(n98), .Z(n150) );
  ANDN U3130 ( .B(x[96]), .A(n150), .Z(n82) );
  XNOR U3131 ( .A(x[100]), .B(n102), .Z(n170) );
  NANDN U3132 ( .A(n124), .B(n170), .Z(n81) );
  XNOR U3133 ( .A(n82), .B(n81), .Z(n83) );
  XOR U3134 ( .A(n103), .B(n83), .Z(n119) );
  XOR U3135 ( .A(x[97]), .B(x[103]), .Z(n138) );
  AND U3136 ( .A(n138), .B(n114), .Z(n104) );
  XOR U3137 ( .A(n84), .B(n104), .Z(n89) );
  XOR U3138 ( .A(x[98]), .B(x[103]), .Z(n162) );
  NAND U3139 ( .A(n162), .B(n127), .Z(n85) );
  XOR U3140 ( .A(n86), .B(n85), .Z(n99) );
  AND U3141 ( .A(n129), .B(n161), .Z(n87) );
  XOR U3142 ( .A(n99), .B(n87), .Z(n88) );
  XNOR U3143 ( .A(n89), .B(n88), .Z(n117) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n152) );
  AND U3145 ( .A(n124), .B(n152), .Z(n91) );
  AND U3146 ( .A(x[96]), .B(n170), .Z(n90) );
  XNOR U3147 ( .A(n91), .B(n90), .Z(n92) );
  NANDN U3148 ( .A(n93), .B(n92), .Z(n96) );
  NAND U3149 ( .A(n124), .B(x[96]), .Z(n94) );
  NANDN U3150 ( .A(n94), .B(n150), .Z(n95) );
  NAND U3151 ( .A(n96), .B(n95), .Z(n97) );
  XNOR U3152 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U3153 ( .A(n100), .B(n99), .Z(n116) );
  OR U3154 ( .A(n117), .B(n116), .Z(n101) );
  NANDN U3155 ( .A(n119), .B(n101), .Z(n109) );
  ANDN U3156 ( .B(n102), .A(x[97]), .Z(n106) );
  XNOR U3157 ( .A(n104), .B(n103), .Z(n105) );
  XNOR U3158 ( .A(n106), .B(n105), .Z(n121) );
  XOR U3159 ( .A(n117), .B(n121), .Z(n107) );
  NAND U3160 ( .A(n116), .B(n107), .Z(n108) );
  NAND U3161 ( .A(n109), .B(n108), .Z(n160) );
  OR U3162 ( .A(n119), .B(n116), .Z(n113) );
  ANDN U3163 ( .B(n116), .A(n117), .Z(n110) );
  XNOR U3164 ( .A(n110), .B(n121), .Z(n111) );
  NAND U3165 ( .A(n119), .B(n111), .Z(n112) );
  NAND U3166 ( .A(n113), .B(n112), .Z(n141) );
  XNOR U3167 ( .A(n160), .B(n141), .Z(n137) );
  AND U3168 ( .A(n114), .B(n137), .Z(n131) );
  NAND U3169 ( .A(n139), .B(n141), .Z(n115) );
  XNOR U3170 ( .A(n131), .B(n115), .Z(n172) );
  NANDN U3171 ( .A(n117), .B(n121), .Z(n123) );
  NANDN U3172 ( .A(n117), .B(n116), .Z(n118) );
  XOR U3173 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U3174 ( .A(n121), .B(n120), .Z(n122) );
  NAND U3175 ( .A(n123), .B(n122), .Z(n149) );
  XOR U3176 ( .A(n169), .B(n149), .Z(n151) );
  AND U3177 ( .A(n124), .B(n151), .Z(n144) );
  NANDN U3178 ( .A(n149), .B(n125), .Z(n126) );
  XNOR U3179 ( .A(n144), .B(n126), .Z(n159) );
  XNOR U3180 ( .A(n172), .B(n159), .Z(z[98]) );
  XNOR U3181 ( .A(n149), .B(n141), .Z(n163) );
  AND U3182 ( .A(n127), .B(n163), .Z(n183) );
  XOR U3183 ( .A(n169), .B(n160), .Z(n134) );
  AND U3184 ( .A(n128), .B(n134), .Z(n181) );
  NANDN U3185 ( .A(n160), .B(n129), .Z(n130) );
  XNOR U3186 ( .A(n131), .B(n130), .Z(n145) );
  XNOR U3187 ( .A(n181), .B(n145), .Z(n132) );
  XNOR U3188 ( .A(n183), .B(n132), .Z(n1958) );
  XOR U3189 ( .A(n1958), .B(z[98]), .Z(z[100]) );
  AND U3190 ( .A(n133), .B(n134), .Z(n165) );
  NAND U3191 ( .A(n157), .B(n135), .Z(n136) );
  XNOR U3192 ( .A(n165), .B(n136), .Z(n153) );
  AND U3193 ( .A(n138), .B(n137), .Z(n166) );
  XOR U3194 ( .A(x[97]), .B(n139), .Z(n140) );
  NAND U3195 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U3196 ( .A(n166), .B(n142), .Z(n147) );
  NANDN U3197 ( .A(n169), .B(x[96]), .Z(n143) );
  XNOR U3198 ( .A(n144), .B(n143), .Z(n180) );
  XNOR U3199 ( .A(n180), .B(n145), .Z(n146) );
  XNOR U3200 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U3201 ( .A(n153), .B(n148), .Z(z[101]) );
  ANDN U3202 ( .B(n150), .A(n149), .Z(n155) );
  AND U3203 ( .A(n152), .B(n151), .Z(n171) );
  XNOR U3204 ( .A(n171), .B(n153), .Z(n154) );
  XNOR U3205 ( .A(n155), .B(n154), .Z(n1959) );
  NAND U3206 ( .A(n157), .B(n156), .Z(n158) );
  XNOR U3207 ( .A(n181), .B(n158), .Z(n175) );
  XNOR U3208 ( .A(n175), .B(n159), .Z(n1957) );
  XNOR U3209 ( .A(n1959), .B(n1957), .Z(n179) );
  ANDN U3210 ( .B(n161), .A(n160), .Z(n168) );
  NAND U3211 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U3212 ( .A(n165), .B(n164), .Z(n176) );
  XNOR U3213 ( .A(n176), .B(n166), .Z(n167) );
  XNOR U3214 ( .A(n168), .B(n167), .Z(n1962) );
  XNOR U3215 ( .A(n179), .B(n1962), .Z(z[102]) );
  ANDN U3216 ( .B(n170), .A(n169), .Z(n174) );
  XNOR U3217 ( .A(n172), .B(n171), .Z(n173) );
  XNOR U3218 ( .A(n174), .B(n173), .Z(n178) );
  XNOR U3219 ( .A(n176), .B(n175), .Z(n177) );
  XNOR U3220 ( .A(n178), .B(n177), .Z(n1960) );
  XNOR U3221 ( .A(n1960), .B(n179), .Z(z[97]) );
  XNOR U3222 ( .A(n181), .B(n180), .Z(n182) );
  XNOR U3223 ( .A(n183), .B(n182), .Z(n184) );
  XOR U3224 ( .A(n184), .B(z[97]), .Z(z[103]) );
  XOR U3225 ( .A(x[107]), .B(x[105]), .Z(n187) );
  XNOR U3226 ( .A(x[104]), .B(x[110]), .Z(n186) );
  XOR U3227 ( .A(n186), .B(x[106]), .Z(n185) );
  XNOR U3228 ( .A(n187), .B(n185), .Z(n222) );
  XNOR U3229 ( .A(x[109]), .B(n186), .Z(n295) );
  XOR U3230 ( .A(n295), .B(x[108]), .Z(n265) );
  IV U3231 ( .A(n265), .Z(n196) );
  XNOR U3232 ( .A(x[111]), .B(x[108]), .Z(n190) );
  XNOR U3233 ( .A(n187), .B(n190), .Z(n250) );
  NOR U3234 ( .A(n196), .B(n250), .Z(n189) );
  XNOR U3235 ( .A(n295), .B(x[111]), .Z(n281) );
  XNOR U3236 ( .A(x[106]), .B(n281), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n205), .Z(n200) );
  AND U3238 ( .A(x[104]), .B(n200), .Z(n188) );
  XNOR U3239 ( .A(n189), .B(n188), .Z(n193) );
  XNOR U3240 ( .A(n222), .B(n281), .Z(n212) );
  IV U3241 ( .A(n222), .Z(n207) );
  XNOR U3242 ( .A(x[104]), .B(n207), .Z(n227) );
  IV U3243 ( .A(n190), .Z(n255) );
  AND U3244 ( .A(n227), .B(n255), .Z(n195) );
  IV U3245 ( .A(n295), .Z(n214) );
  XNOR U3246 ( .A(n222), .B(n214), .Z(n244) );
  XOR U3247 ( .A(n244), .B(n250), .Z(n247) );
  XOR U3248 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NAND U3249 ( .A(n247), .B(n257), .Z(n191) );
  XNOR U3250 ( .A(n195), .B(n191), .Z(n216) );
  XNOR U3251 ( .A(n212), .B(n216), .Z(n192) );
  XNOR U3252 ( .A(n193), .B(n192), .Z(n239) );
  XOR U3253 ( .A(x[106]), .B(x[111]), .Z(n271) );
  XNOR U3254 ( .A(x[104]), .B(n250), .Z(n251) );
  XNOR U3255 ( .A(n295), .B(n251), .Z(n242) );
  NAND U3256 ( .A(n271), .B(n242), .Z(n194) );
  XNOR U3257 ( .A(n195), .B(n194), .Z(n208) );
  IV U3258 ( .A(n200), .Z(n254) );
  XNOR U3259 ( .A(n254), .B(n196), .Z(n261) );
  AND U3260 ( .A(n250), .B(n261), .Z(n198) );
  AND U3261 ( .A(x[104]), .B(n265), .Z(n197) );
  XNOR U3262 ( .A(n198), .B(n197), .Z(n199) );
  NANDN U3263 ( .A(n251), .B(n199), .Z(n203) );
  NAND U3264 ( .A(x[104]), .B(n250), .Z(n201) );
  OR U3265 ( .A(n201), .B(n200), .Z(n202) );
  NAND U3266 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U3267 ( .A(n205), .B(n204), .Z(n206) );
  XNOR U3268 ( .A(n208), .B(n206), .Z(n228) );
  IV U3269 ( .A(n228), .Z(n235) );
  AND U3270 ( .A(n281), .B(n207), .Z(n210) );
  XOR U3271 ( .A(x[105]), .B(x[111]), .Z(n283) );
  AND U3272 ( .A(n244), .B(n283), .Z(n213) );
  XNOR U3273 ( .A(n213), .B(n208), .Z(n209) );
  XNOR U3274 ( .A(n210), .B(n209), .Z(n234) );
  NANDN U3275 ( .A(n235), .B(n234), .Z(n211) );
  NAND U3276 ( .A(n239), .B(n211), .Z(n221) );
  XNOR U3277 ( .A(n213), .B(n212), .Z(n218) );
  ANDN U3278 ( .B(n214), .A(x[105]), .Z(n215) );
  XNOR U3279 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3280 ( .A(n218), .B(n217), .Z(n231) );
  XOR U3281 ( .A(n234), .B(n231), .Z(n219) );
  NAND U3282 ( .A(n235), .B(n219), .Z(n220) );
  NAND U3283 ( .A(n221), .B(n220), .Z(n280) );
  ANDN U3284 ( .B(n222), .A(n280), .Z(n246) );
  IV U3285 ( .A(n231), .Z(n237) );
  XOR U3286 ( .A(n239), .B(n235), .Z(n223) );
  NANDN U3287 ( .A(n237), .B(n223), .Z(n226) );
  NANDN U3288 ( .A(n235), .B(n237), .Z(n224) );
  NANDN U3289 ( .A(n234), .B(n224), .Z(n225) );
  NAND U3290 ( .A(n226), .B(n225), .Z(n290) );
  XNOR U3291 ( .A(n280), .B(n290), .Z(n256) );
  AND U3292 ( .A(n227), .B(n256), .Z(n249) );
  OR U3293 ( .A(n234), .B(n231), .Z(n233) );
  ANDN U3294 ( .B(n234), .A(n228), .Z(n229) );
  XNOR U3295 ( .A(n229), .B(n239), .Z(n230) );
  NAND U3296 ( .A(n231), .B(n230), .Z(n232) );
  NAND U3297 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3298 ( .A(n235), .B(n239), .Z(n241) );
  NAND U3299 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U3300 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U3301 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3302 ( .A(n241), .B(n240), .Z(n297) );
  NAND U3303 ( .A(n272), .B(n242), .Z(n243) );
  XNOR U3304 ( .A(n249), .B(n243), .Z(n292) );
  XOR U3305 ( .A(n280), .B(n297), .Z(n282) );
  AND U3306 ( .A(n244), .B(n282), .Z(n267) );
  XNOR U3307 ( .A(n292), .B(n267), .Z(n245) );
  XNOR U3308 ( .A(n246), .B(n245), .Z(n300) );
  NAND U3309 ( .A(n258), .B(n247), .Z(n248) );
  XNOR U3310 ( .A(n249), .B(n248), .Z(n275) );
  AND U3311 ( .A(n250), .B(n260), .Z(n291) );
  NANDN U3312 ( .A(n251), .B(n253), .Z(n252) );
  XNOR U3313 ( .A(n291), .B(n252), .Z(n279) );
  XNOR U3314 ( .A(n275), .B(n279), .Z(n264) );
  XOR U3315 ( .A(n300), .B(n264), .Z(z[104]) );
  AND U3316 ( .A(n254), .B(n253), .Z(n263) );
  AND U3317 ( .A(n256), .B(n255), .Z(n274) );
  NAND U3318 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3319 ( .A(n274), .B(n259), .Z(n301) );
  AND U3320 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3321 ( .A(n301), .B(n268), .Z(n262) );
  XNOR U3322 ( .A(n263), .B(n262), .Z(n288) );
  XNOR U3323 ( .A(n288), .B(n264), .Z(n360) );
  AND U3324 ( .A(n265), .B(n290), .Z(n270) );
  NANDN U3325 ( .A(n297), .B(n295), .Z(n266) );
  XNOR U3326 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3327 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3328 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3329 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3330 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3331 ( .A(n275), .B(n284), .Z(n276) );
  XNOR U3332 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3333 ( .A(n360), .B(n287), .Z(z[105]) );
  XNOR U3334 ( .A(n279), .B(n278), .Z(z[106]) );
  NOR U3335 ( .A(n281), .B(n280), .Z(n286) );
  AND U3336 ( .A(n283), .B(n282), .Z(n299) );
  XNOR U3337 ( .A(n284), .B(n299), .Z(n285) );
  XNOR U3338 ( .A(n286), .B(n285), .Z(n359) );
  XOR U3339 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U3340 ( .A(n359), .B(n289), .Z(z[107]) );
  XOR U3341 ( .A(n300), .B(z[106]), .Z(z[108]) );
  AND U3342 ( .A(x[104]), .B(n290), .Z(n294) );
  XNOR U3343 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U3344 ( .A(n294), .B(n293), .Z(n361) );
  XOR U3345 ( .A(n295), .B(x[105]), .Z(n296) );
  NANDN U3346 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U3347 ( .A(n299), .B(n298), .Z(n303) );
  XNOR U3348 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U3349 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U3350 ( .A(n361), .B(n304), .Z(z[109]) );
  XOR U3351 ( .A(x[9]), .B(x[11]), .Z(n305) );
  XOR U3352 ( .A(x[15]), .B(x[12]), .Z(n486) );
  XOR U3353 ( .A(n305), .B(n486), .Z(n341) );
  XNOR U3354 ( .A(x[8]), .B(x[14]), .Z(n307) );
  XNOR U3355 ( .A(x[13]), .B(n307), .Z(n654) );
  XNOR U3356 ( .A(x[15]), .B(n654), .Z(n485) );
  XNOR U3357 ( .A(n305), .B(x[10]), .Z(n306) );
  XNOR U3358 ( .A(n307), .B(n306), .Z(n308) );
  AND U3359 ( .A(n485), .B(n308), .Z(n311) );
  IV U3360 ( .A(n308), .Z(n641) );
  XOR U3361 ( .A(n641), .B(n654), .Z(n357) );
  XOR U3362 ( .A(x[9]), .B(x[15]), .Z(n491) );
  AND U3363 ( .A(n357), .B(n491), .Z(n312) );
  XNOR U3364 ( .A(x[8]), .B(n308), .Z(n509) );
  AND U3365 ( .A(n486), .B(n509), .Z(n314) );
  XOR U3366 ( .A(x[15]), .B(x[10]), .Z(n488) );
  XNOR U3367 ( .A(n341), .B(x[8]), .Z(n342) );
  XNOR U3368 ( .A(n654), .B(n342), .Z(n642) );
  NAND U3369 ( .A(n488), .B(n642), .Z(n309) );
  XNOR U3370 ( .A(n314), .B(n309), .Z(n325) );
  XNOR U3371 ( .A(n312), .B(n325), .Z(n310) );
  XNOR U3372 ( .A(n311), .B(n310), .Z(n349) );
  XNOR U3373 ( .A(n641), .B(n485), .Z(n329) );
  XOR U3374 ( .A(x[12]), .B(x[10]), .Z(n496) );
  XOR U3375 ( .A(n341), .B(n357), .Z(n510) );
  NAND U3376 ( .A(n496), .B(n510), .Z(n313) );
  XNOR U3377 ( .A(n314), .B(n313), .Z(n328) );
  OR U3378 ( .A(n349), .B(n345), .Z(n335) );
  XNOR U3379 ( .A(x[10]), .B(n485), .Z(n323) );
  IV U3380 ( .A(n318), .Z(n495) );
  XNOR U3381 ( .A(x[12]), .B(n654), .Z(n503) );
  XNOR U3382 ( .A(n495), .B(n503), .Z(n500) );
  AND U3383 ( .A(n341), .B(n500), .Z(n316) );
  ANDN U3384 ( .B(x[8]), .A(n503), .Z(n315) );
  XNOR U3385 ( .A(n316), .B(n315), .Z(n317) );
  NANDN U3386 ( .A(n342), .B(n317), .Z(n321) );
  NAND U3387 ( .A(n341), .B(x[8]), .Z(n319) );
  OR U3388 ( .A(n319), .B(n318), .Z(n320) );
  NAND U3389 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U3390 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U3391 ( .A(n325), .B(n324), .Z(n336) );
  ANDN U3392 ( .B(n349), .A(n336), .Z(n332) );
  NOR U3393 ( .A(n503), .B(n341), .Z(n327) );
  ANDN U3394 ( .B(x[8]), .A(n495), .Z(n326) );
  XNOR U3395 ( .A(n327), .B(n326), .Z(n331) );
  XNOR U3396 ( .A(n329), .B(n328), .Z(n330) );
  XNOR U3397 ( .A(n331), .B(n330), .Z(n354) );
  XNOR U3398 ( .A(n332), .B(n354), .Z(n333) );
  NAND U3399 ( .A(n345), .B(n333), .Z(n334) );
  NAND U3400 ( .A(n335), .B(n334), .Z(n494) );
  IV U3401 ( .A(n494), .Z(n487) );
  IV U3402 ( .A(n345), .Z(n352) );
  IV U3403 ( .A(n336), .Z(n350) );
  XOR U3404 ( .A(n354), .B(n350), .Z(n337) );
  NANDN U3405 ( .A(n352), .B(n337), .Z(n340) );
  NANDN U3406 ( .A(n350), .B(n352), .Z(n338) );
  NANDN U3407 ( .A(n349), .B(n338), .Z(n339) );
  NAND U3408 ( .A(n340), .B(n339), .Z(n649) );
  XNOR U3409 ( .A(n487), .B(n649), .Z(n499) );
  AND U3410 ( .A(n341), .B(n499), .Z(n651) );
  NANDN U3411 ( .A(n342), .B(n494), .Z(n343) );
  XNOR U3412 ( .A(n651), .B(n343), .Z(n663) );
  NANDN U3413 ( .A(n350), .B(n349), .Z(n344) );
  NAND U3414 ( .A(n354), .B(n344), .Z(n348) );
  XOR U3415 ( .A(n349), .B(n345), .Z(n346) );
  NAND U3416 ( .A(n350), .B(n346), .Z(n347) );
  NAND U3417 ( .A(n348), .B(n347), .Z(n640) );
  NAND U3418 ( .A(n350), .B(n354), .Z(n356) );
  NAND U3419 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U3420 ( .A(n352), .B(n351), .Z(n353) );
  NANDN U3421 ( .A(n354), .B(n353), .Z(n355) );
  NAND U3422 ( .A(n356), .B(n355), .Z(n656) );
  XOR U3423 ( .A(n640), .B(n656), .Z(n490) );
  AND U3424 ( .A(n357), .B(n490), .Z(n646) );
  NANDN U3425 ( .A(n656), .B(n654), .Z(n358) );
  XNOR U3426 ( .A(n646), .B(n358), .Z(n513) );
  XNOR U3427 ( .A(n663), .B(n513), .Z(z[10]) );
  XNOR U3428 ( .A(n360), .B(n359), .Z(z[110]) );
  XOR U3429 ( .A(n361), .B(z[105]), .Z(z[111]) );
  XOR U3430 ( .A(x[115]), .B(x[113]), .Z(n364) );
  XNOR U3431 ( .A(x[112]), .B(x[118]), .Z(n363) );
  XOR U3432 ( .A(n363), .B(x[114]), .Z(n362) );
  XNOR U3433 ( .A(n364), .B(n362), .Z(n399) );
  XNOR U3434 ( .A(x[117]), .B(n363), .Z(n472) );
  XOR U3435 ( .A(n472), .B(x[116]), .Z(n442) );
  IV U3436 ( .A(n442), .Z(n373) );
  XNOR U3437 ( .A(x[119]), .B(x[116]), .Z(n367) );
  XNOR U3438 ( .A(n364), .B(n367), .Z(n427) );
  NOR U3439 ( .A(n373), .B(n427), .Z(n366) );
  XNOR U3440 ( .A(n472), .B(x[119]), .Z(n458) );
  XNOR U3441 ( .A(x[114]), .B(n458), .Z(n382) );
  XNOR U3442 ( .A(x[113]), .B(n382), .Z(n377) );
  AND U3443 ( .A(x[112]), .B(n377), .Z(n365) );
  XNOR U3444 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U3445 ( .A(n399), .B(n458), .Z(n389) );
  IV U3446 ( .A(n399), .Z(n384) );
  XNOR U3447 ( .A(x[112]), .B(n384), .Z(n404) );
  IV U3448 ( .A(n367), .Z(n432) );
  AND U3449 ( .A(n404), .B(n432), .Z(n372) );
  IV U3450 ( .A(n472), .Z(n391) );
  XNOR U3451 ( .A(n399), .B(n391), .Z(n421) );
  XOR U3452 ( .A(n421), .B(n427), .Z(n424) );
  XOR U3453 ( .A(x[114]), .B(x[116]), .Z(n434) );
  NAND U3454 ( .A(n424), .B(n434), .Z(n368) );
  XNOR U3455 ( .A(n372), .B(n368), .Z(n393) );
  XNOR U3456 ( .A(n389), .B(n393), .Z(n369) );
  XNOR U3457 ( .A(n370), .B(n369), .Z(n416) );
  XOR U3458 ( .A(x[114]), .B(x[119]), .Z(n448) );
  XNOR U3459 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3460 ( .A(n472), .B(n428), .Z(n419) );
  NAND U3461 ( .A(n448), .B(n419), .Z(n371) );
  XNOR U3462 ( .A(n372), .B(n371), .Z(n385) );
  IV U3463 ( .A(n377), .Z(n431) );
  XNOR U3464 ( .A(n431), .B(n373), .Z(n438) );
  AND U3465 ( .A(n427), .B(n438), .Z(n375) );
  AND U3466 ( .A(x[112]), .B(n442), .Z(n374) );
  XNOR U3467 ( .A(n375), .B(n374), .Z(n376) );
  NANDN U3468 ( .A(n428), .B(n376), .Z(n380) );
  NAND U3469 ( .A(x[112]), .B(n427), .Z(n378) );
  OR U3470 ( .A(n378), .B(n377), .Z(n379) );
  NAND U3471 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U3472 ( .A(n382), .B(n381), .Z(n383) );
  XNOR U3473 ( .A(n385), .B(n383), .Z(n405) );
  IV U3474 ( .A(n405), .Z(n412) );
  AND U3475 ( .A(n458), .B(n384), .Z(n387) );
  XOR U3476 ( .A(x[113]), .B(x[119]), .Z(n460) );
  AND U3477 ( .A(n421), .B(n460), .Z(n390) );
  XNOR U3478 ( .A(n390), .B(n385), .Z(n386) );
  XNOR U3479 ( .A(n387), .B(n386), .Z(n411) );
  NANDN U3480 ( .A(n412), .B(n411), .Z(n388) );
  NAND U3481 ( .A(n416), .B(n388), .Z(n398) );
  XNOR U3482 ( .A(n390), .B(n389), .Z(n395) );
  ANDN U3483 ( .B(n391), .A(x[113]), .Z(n392) );
  XNOR U3484 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U3485 ( .A(n395), .B(n394), .Z(n408) );
  XOR U3486 ( .A(n411), .B(n408), .Z(n396) );
  NAND U3487 ( .A(n412), .B(n396), .Z(n397) );
  NAND U3488 ( .A(n398), .B(n397), .Z(n457) );
  ANDN U3489 ( .B(n399), .A(n457), .Z(n423) );
  IV U3490 ( .A(n408), .Z(n414) );
  XOR U3491 ( .A(n416), .B(n412), .Z(n400) );
  NANDN U3492 ( .A(n414), .B(n400), .Z(n403) );
  NANDN U3493 ( .A(n412), .B(n414), .Z(n401) );
  NANDN U3494 ( .A(n411), .B(n401), .Z(n402) );
  NAND U3495 ( .A(n403), .B(n402), .Z(n467) );
  XNOR U3496 ( .A(n457), .B(n467), .Z(n433) );
  AND U3497 ( .A(n404), .B(n433), .Z(n426) );
  OR U3498 ( .A(n411), .B(n408), .Z(n410) );
  ANDN U3499 ( .B(n411), .A(n405), .Z(n406) );
  XNOR U3500 ( .A(n406), .B(n416), .Z(n407) );
  NAND U3501 ( .A(n408), .B(n407), .Z(n409) );
  NAND U3502 ( .A(n410), .B(n409), .Z(n430) );
  NAND U3503 ( .A(n412), .B(n416), .Z(n418) );
  NAND U3504 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U3505 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U3506 ( .A(n416), .B(n415), .Z(n417) );
  NAND U3507 ( .A(n418), .B(n417), .Z(n474) );
  NAND U3508 ( .A(n449), .B(n419), .Z(n420) );
  XNOR U3509 ( .A(n426), .B(n420), .Z(n469) );
  XOR U3510 ( .A(n457), .B(n474), .Z(n459) );
  AND U3511 ( .A(n421), .B(n459), .Z(n444) );
  XNOR U3512 ( .A(n469), .B(n444), .Z(n422) );
  XNOR U3513 ( .A(n423), .B(n422), .Z(n477) );
  NAND U3514 ( .A(n435), .B(n424), .Z(n425) );
  XNOR U3515 ( .A(n426), .B(n425), .Z(n452) );
  AND U3516 ( .A(n427), .B(n437), .Z(n468) );
  NANDN U3517 ( .A(n428), .B(n430), .Z(n429) );
  XNOR U3518 ( .A(n468), .B(n429), .Z(n456) );
  XNOR U3519 ( .A(n452), .B(n456), .Z(n441) );
  XOR U3520 ( .A(n477), .B(n441), .Z(z[112]) );
  AND U3521 ( .A(n431), .B(n430), .Z(n440) );
  AND U3522 ( .A(n433), .B(n432), .Z(n451) );
  NAND U3523 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U3524 ( .A(n451), .B(n436), .Z(n478) );
  AND U3525 ( .A(n438), .B(n437), .Z(n445) );
  XNOR U3526 ( .A(n478), .B(n445), .Z(n439) );
  XNOR U3527 ( .A(n440), .B(n439), .Z(n465) );
  XNOR U3528 ( .A(n465), .B(n441), .Z(n483) );
  AND U3529 ( .A(n442), .B(n467), .Z(n447) );
  NANDN U3530 ( .A(n474), .B(n472), .Z(n443) );
  XNOR U3531 ( .A(n444), .B(n443), .Z(n455) );
  XNOR U3532 ( .A(n445), .B(n455), .Z(n446) );
  XNOR U3533 ( .A(n447), .B(n446), .Z(n454) );
  NAND U3534 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U3535 ( .A(n451), .B(n450), .Z(n461) );
  XNOR U3536 ( .A(n452), .B(n461), .Z(n453) );
  XNOR U3537 ( .A(n454), .B(n453), .Z(n464) );
  XNOR U3538 ( .A(n483), .B(n464), .Z(z[113]) );
  XNOR U3539 ( .A(n456), .B(n455), .Z(z[114]) );
  NOR U3540 ( .A(n458), .B(n457), .Z(n463) );
  AND U3541 ( .A(n460), .B(n459), .Z(n476) );
  XNOR U3542 ( .A(n461), .B(n476), .Z(n462) );
  XNOR U3543 ( .A(n463), .B(n462), .Z(n482) );
  XOR U3544 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U3545 ( .A(n482), .B(n466), .Z(z[115]) );
  XOR U3546 ( .A(n477), .B(z[114]), .Z(z[116]) );
  AND U3547 ( .A(x[112]), .B(n467), .Z(n471) );
  XNOR U3548 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U3549 ( .A(n471), .B(n470), .Z(n484) );
  XOR U3550 ( .A(n472), .B(x[113]), .Z(n473) );
  NANDN U3551 ( .A(n474), .B(n473), .Z(n475) );
  XNOR U3552 ( .A(n476), .B(n475), .Z(n480) );
  XNOR U3553 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U3554 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U3555 ( .A(n484), .B(n481), .Z(z[117]) );
  XNOR U3556 ( .A(n483), .B(n482), .Z(z[118]) );
  XOR U3557 ( .A(n484), .B(z[113]), .Z(z[119]) );
  NOR U3558 ( .A(n485), .B(n640), .Z(n493) );
  XNOR U3559 ( .A(n640), .B(n649), .Z(n508) );
  AND U3560 ( .A(n486), .B(n508), .Z(n498) );
  XOR U3561 ( .A(n487), .B(n656), .Z(n643) );
  NAND U3562 ( .A(n643), .B(n488), .Z(n489) );
  XNOR U3563 ( .A(n498), .B(n489), .Z(n504) );
  AND U3564 ( .A(n491), .B(n490), .Z(n658) );
  XNOR U3565 ( .A(n504), .B(n658), .Z(n492) );
  XNOR U3566 ( .A(n493), .B(n492), .Z(n666) );
  AND U3567 ( .A(n495), .B(n494), .Z(n502) );
  NAND U3568 ( .A(n511), .B(n496), .Z(n497) );
  XNOR U3569 ( .A(n498), .B(n497), .Z(n659) );
  AND U3570 ( .A(n500), .B(n499), .Z(n505) );
  XNOR U3571 ( .A(n659), .B(n505), .Z(n501) );
  XNOR U3572 ( .A(n502), .B(n501), .Z(n665) );
  ANDN U3573 ( .B(n649), .A(n503), .Z(n507) );
  XNOR U3574 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U3575 ( .A(n507), .B(n506), .Z(n515) );
  AND U3576 ( .A(n509), .B(n508), .Z(n645) );
  NAND U3577 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U3578 ( .A(n645), .B(n512), .Z(n664) );
  XNOR U3579 ( .A(n664), .B(n513), .Z(n514) );
  XNOR U3580 ( .A(n515), .B(n514), .Z(n667) );
  XOR U3581 ( .A(n665), .B(n667), .Z(n516) );
  XNOR U3582 ( .A(n666), .B(n516), .Z(z[11]) );
  XOR U3583 ( .A(x[123]), .B(x[121]), .Z(n519) );
  XNOR U3584 ( .A(x[120]), .B(x[126]), .Z(n518) );
  XOR U3585 ( .A(n518), .B(x[122]), .Z(n517) );
  XNOR U3586 ( .A(n519), .B(n517), .Z(n554) );
  XNOR U3587 ( .A(x[125]), .B(n518), .Z(n627) );
  XOR U3588 ( .A(n627), .B(x[124]), .Z(n597) );
  IV U3589 ( .A(n597), .Z(n528) );
  XNOR U3590 ( .A(x[127]), .B(x[124]), .Z(n522) );
  XNOR U3591 ( .A(n519), .B(n522), .Z(n582) );
  NOR U3592 ( .A(n528), .B(n582), .Z(n521) );
  XNOR U3593 ( .A(n627), .B(x[127]), .Z(n613) );
  XNOR U3594 ( .A(x[122]), .B(n613), .Z(n537) );
  XNOR U3595 ( .A(x[121]), .B(n537), .Z(n532) );
  AND U3596 ( .A(x[120]), .B(n532), .Z(n520) );
  XNOR U3597 ( .A(n521), .B(n520), .Z(n525) );
  XNOR U3598 ( .A(n554), .B(n613), .Z(n544) );
  IV U3599 ( .A(n554), .Z(n539) );
  XNOR U3600 ( .A(x[120]), .B(n539), .Z(n559) );
  IV U3601 ( .A(n522), .Z(n587) );
  AND U3602 ( .A(n559), .B(n587), .Z(n527) );
  IV U3603 ( .A(n627), .Z(n546) );
  XNOR U3604 ( .A(n554), .B(n546), .Z(n576) );
  XOR U3605 ( .A(n576), .B(n582), .Z(n579) );
  XOR U3606 ( .A(x[122]), .B(x[124]), .Z(n589) );
  NAND U3607 ( .A(n579), .B(n589), .Z(n523) );
  XNOR U3608 ( .A(n527), .B(n523), .Z(n548) );
  XNOR U3609 ( .A(n544), .B(n548), .Z(n524) );
  XNOR U3610 ( .A(n525), .B(n524), .Z(n571) );
  XOR U3611 ( .A(x[122]), .B(x[127]), .Z(n603) );
  XNOR U3612 ( .A(x[120]), .B(n582), .Z(n583) );
  XNOR U3613 ( .A(n627), .B(n583), .Z(n574) );
  NAND U3614 ( .A(n603), .B(n574), .Z(n526) );
  XNOR U3615 ( .A(n527), .B(n526), .Z(n540) );
  IV U3616 ( .A(n532), .Z(n586) );
  XNOR U3617 ( .A(n586), .B(n528), .Z(n593) );
  AND U3618 ( .A(n582), .B(n593), .Z(n530) );
  AND U3619 ( .A(x[120]), .B(n597), .Z(n529) );
  XNOR U3620 ( .A(n530), .B(n529), .Z(n531) );
  NANDN U3621 ( .A(n583), .B(n531), .Z(n535) );
  NAND U3622 ( .A(x[120]), .B(n582), .Z(n533) );
  OR U3623 ( .A(n533), .B(n532), .Z(n534) );
  NAND U3624 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U3625 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U3626 ( .A(n540), .B(n538), .Z(n560) );
  IV U3627 ( .A(n560), .Z(n567) );
  AND U3628 ( .A(n613), .B(n539), .Z(n542) );
  XOR U3629 ( .A(x[121]), .B(x[127]), .Z(n615) );
  AND U3630 ( .A(n576), .B(n615), .Z(n545) );
  XNOR U3631 ( .A(n545), .B(n540), .Z(n541) );
  XNOR U3632 ( .A(n542), .B(n541), .Z(n566) );
  NANDN U3633 ( .A(n567), .B(n566), .Z(n543) );
  NAND U3634 ( .A(n571), .B(n543), .Z(n553) );
  XNOR U3635 ( .A(n545), .B(n544), .Z(n550) );
  ANDN U3636 ( .B(n546), .A(x[121]), .Z(n547) );
  XNOR U3637 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U3638 ( .A(n550), .B(n549), .Z(n563) );
  XOR U3639 ( .A(n566), .B(n563), .Z(n551) );
  NAND U3640 ( .A(n567), .B(n551), .Z(n552) );
  NAND U3641 ( .A(n553), .B(n552), .Z(n612) );
  ANDN U3642 ( .B(n554), .A(n612), .Z(n578) );
  IV U3643 ( .A(n563), .Z(n569) );
  XOR U3644 ( .A(n571), .B(n567), .Z(n555) );
  NANDN U3645 ( .A(n569), .B(n555), .Z(n558) );
  NANDN U3646 ( .A(n567), .B(n569), .Z(n556) );
  NANDN U3647 ( .A(n566), .B(n556), .Z(n557) );
  NAND U3648 ( .A(n558), .B(n557), .Z(n622) );
  XNOR U3649 ( .A(n612), .B(n622), .Z(n588) );
  AND U3650 ( .A(n559), .B(n588), .Z(n581) );
  OR U3651 ( .A(n566), .B(n563), .Z(n565) );
  ANDN U3652 ( .B(n566), .A(n560), .Z(n561) );
  XNOR U3653 ( .A(n561), .B(n571), .Z(n562) );
  NAND U3654 ( .A(n563), .B(n562), .Z(n564) );
  NAND U3655 ( .A(n565), .B(n564), .Z(n585) );
  NAND U3656 ( .A(n567), .B(n571), .Z(n573) );
  NAND U3657 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U3658 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U3659 ( .A(n571), .B(n570), .Z(n572) );
  NAND U3660 ( .A(n573), .B(n572), .Z(n629) );
  NAND U3661 ( .A(n604), .B(n574), .Z(n575) );
  XNOR U3662 ( .A(n581), .B(n575), .Z(n624) );
  XOR U3663 ( .A(n612), .B(n629), .Z(n614) );
  AND U3664 ( .A(n576), .B(n614), .Z(n599) );
  XNOR U3665 ( .A(n624), .B(n599), .Z(n577) );
  XNOR U3666 ( .A(n578), .B(n577), .Z(n632) );
  NAND U3667 ( .A(n590), .B(n579), .Z(n580) );
  XNOR U3668 ( .A(n581), .B(n580), .Z(n607) );
  AND U3669 ( .A(n582), .B(n592), .Z(n623) );
  NANDN U3670 ( .A(n583), .B(n585), .Z(n584) );
  XNOR U3671 ( .A(n623), .B(n584), .Z(n611) );
  XNOR U3672 ( .A(n607), .B(n611), .Z(n596) );
  XOR U3673 ( .A(n632), .B(n596), .Z(z[120]) );
  AND U3674 ( .A(n586), .B(n585), .Z(n595) );
  AND U3675 ( .A(n588), .B(n587), .Z(n606) );
  NAND U3676 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U3677 ( .A(n606), .B(n591), .Z(n633) );
  AND U3678 ( .A(n593), .B(n592), .Z(n600) );
  XNOR U3679 ( .A(n633), .B(n600), .Z(n594) );
  XNOR U3680 ( .A(n595), .B(n594), .Z(n620) );
  XNOR U3681 ( .A(n620), .B(n596), .Z(n638) );
  AND U3682 ( .A(n597), .B(n622), .Z(n602) );
  NANDN U3683 ( .A(n629), .B(n627), .Z(n598) );
  XNOR U3684 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U3685 ( .A(n600), .B(n610), .Z(n601) );
  XNOR U3686 ( .A(n602), .B(n601), .Z(n609) );
  NAND U3687 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U3688 ( .A(n606), .B(n605), .Z(n616) );
  XNOR U3689 ( .A(n607), .B(n616), .Z(n608) );
  XNOR U3690 ( .A(n609), .B(n608), .Z(n619) );
  XNOR U3691 ( .A(n638), .B(n619), .Z(z[121]) );
  XNOR U3692 ( .A(n611), .B(n610), .Z(z[122]) );
  NOR U3693 ( .A(n613), .B(n612), .Z(n618) );
  AND U3694 ( .A(n615), .B(n614), .Z(n631) );
  XNOR U3695 ( .A(n616), .B(n631), .Z(n617) );
  XNOR U3696 ( .A(n618), .B(n617), .Z(n637) );
  XOR U3697 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U3698 ( .A(n637), .B(n621), .Z(z[123]) );
  XOR U3699 ( .A(n632), .B(z[122]), .Z(z[124]) );
  AND U3700 ( .A(x[120]), .B(n622), .Z(n626) );
  XNOR U3701 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U3702 ( .A(n626), .B(n625), .Z(n639) );
  XOR U3703 ( .A(n627), .B(x[121]), .Z(n628) );
  NANDN U3704 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U3705 ( .A(n631), .B(n630), .Z(n635) );
  XNOR U3706 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U3707 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U3708 ( .A(n639), .B(n636), .Z(z[125]) );
  XNOR U3709 ( .A(n638), .B(n637), .Z(z[126]) );
  XOR U3710 ( .A(n639), .B(z[121]), .Z(z[127]) );
  ANDN U3711 ( .B(n641), .A(n640), .Z(n648) );
  NAND U3712 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U3713 ( .A(n645), .B(n644), .Z(n650) );
  XNOR U3714 ( .A(n650), .B(n646), .Z(n647) );
  XNOR U3715 ( .A(n648), .B(n647), .Z(n1926) );
  XOR U3716 ( .A(n1926), .B(z[10]), .Z(z[12]) );
  AND U3717 ( .A(x[8]), .B(n649), .Z(n653) );
  XNOR U3718 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U3719 ( .A(n653), .B(n652), .Z(n669) );
  XOR U3720 ( .A(n654), .B(x[9]), .Z(n655) );
  NANDN U3721 ( .A(n656), .B(n655), .Z(n657) );
  XNOR U3722 ( .A(n658), .B(n657), .Z(n661) );
  XNOR U3723 ( .A(n659), .B(n1926), .Z(n660) );
  XNOR U3724 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U3725 ( .A(n669), .B(n662), .Z(z[13]) );
  XNOR U3726 ( .A(n664), .B(n663), .Z(n1925) );
  XNOR U3727 ( .A(n665), .B(n1925), .Z(n668) );
  XNOR U3728 ( .A(n668), .B(n666), .Z(z[14]) );
  XNOR U3729 ( .A(n668), .B(n667), .Z(z[9]) );
  XOR U3730 ( .A(n669), .B(z[9]), .Z(z[15]) );
  XOR U3731 ( .A(x[19]), .B(x[17]), .Z(n672) );
  XNOR U3732 ( .A(x[16]), .B(x[22]), .Z(n671) );
  XOR U3733 ( .A(n671), .B(x[18]), .Z(n670) );
  XNOR U3734 ( .A(n672), .B(n670), .Z(n707) );
  XNOR U3735 ( .A(x[21]), .B(n671), .Z(n805) );
  XOR U3736 ( .A(n805), .B(x[20]), .Z(n750) );
  IV U3737 ( .A(n750), .Z(n681) );
  XNOR U3738 ( .A(x[23]), .B(x[20]), .Z(n675) );
  XNOR U3739 ( .A(n672), .B(n675), .Z(n735) );
  NOR U3740 ( .A(n681), .B(n735), .Z(n674) );
  XNOR U3741 ( .A(n805), .B(x[23]), .Z(n766) );
  XNOR U3742 ( .A(x[18]), .B(n766), .Z(n690) );
  XNOR U3743 ( .A(x[17]), .B(n690), .Z(n685) );
  AND U3744 ( .A(x[16]), .B(n685), .Z(n673) );
  XNOR U3745 ( .A(n674), .B(n673), .Z(n678) );
  XNOR U3746 ( .A(n707), .B(n766), .Z(n697) );
  IV U3747 ( .A(n707), .Z(n692) );
  XNOR U3748 ( .A(x[16]), .B(n692), .Z(n712) );
  IV U3749 ( .A(n675), .Z(n740) );
  AND U3750 ( .A(n712), .B(n740), .Z(n680) );
  IV U3751 ( .A(n805), .Z(n699) );
  XNOR U3752 ( .A(n707), .B(n699), .Z(n729) );
  XOR U3753 ( .A(n729), .B(n735), .Z(n732) );
  XOR U3754 ( .A(x[18]), .B(x[20]), .Z(n742) );
  NAND U3755 ( .A(n732), .B(n742), .Z(n676) );
  XNOR U3756 ( .A(n680), .B(n676), .Z(n701) );
  XNOR U3757 ( .A(n697), .B(n701), .Z(n677) );
  XNOR U3758 ( .A(n678), .B(n677), .Z(n724) );
  XOR U3759 ( .A(x[18]), .B(x[23]), .Z(n756) );
  XNOR U3760 ( .A(x[16]), .B(n735), .Z(n736) );
  XNOR U3761 ( .A(n805), .B(n736), .Z(n727) );
  NAND U3762 ( .A(n756), .B(n727), .Z(n679) );
  XNOR U3763 ( .A(n680), .B(n679), .Z(n693) );
  IV U3764 ( .A(n685), .Z(n739) );
  XNOR U3765 ( .A(n739), .B(n681), .Z(n746) );
  AND U3766 ( .A(n735), .B(n746), .Z(n683) );
  AND U3767 ( .A(x[16]), .B(n750), .Z(n682) );
  XNOR U3768 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U3769 ( .A(n736), .B(n684), .Z(n688) );
  NAND U3770 ( .A(x[16]), .B(n735), .Z(n686) );
  OR U3771 ( .A(n686), .B(n685), .Z(n687) );
  NAND U3772 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U3773 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U3774 ( .A(n693), .B(n691), .Z(n713) );
  IV U3775 ( .A(n713), .Z(n720) );
  AND U3776 ( .A(n766), .B(n692), .Z(n695) );
  XOR U3777 ( .A(x[17]), .B(x[23]), .Z(n768) );
  AND U3778 ( .A(n729), .B(n768), .Z(n698) );
  XNOR U3779 ( .A(n698), .B(n693), .Z(n694) );
  XNOR U3780 ( .A(n695), .B(n694), .Z(n719) );
  NANDN U3781 ( .A(n720), .B(n719), .Z(n696) );
  NAND U3782 ( .A(n724), .B(n696), .Z(n706) );
  XNOR U3783 ( .A(n698), .B(n697), .Z(n703) );
  ANDN U3784 ( .B(n699), .A(x[17]), .Z(n700) );
  XNOR U3785 ( .A(n701), .B(n700), .Z(n702) );
  XNOR U3786 ( .A(n703), .B(n702), .Z(n716) );
  XOR U3787 ( .A(n719), .B(n716), .Z(n704) );
  NAND U3788 ( .A(n720), .B(n704), .Z(n705) );
  NAND U3789 ( .A(n706), .B(n705), .Z(n765) );
  ANDN U3790 ( .B(n707), .A(n765), .Z(n731) );
  IV U3791 ( .A(n716), .Z(n722) );
  XOR U3792 ( .A(n724), .B(n720), .Z(n708) );
  NANDN U3793 ( .A(n722), .B(n708), .Z(n711) );
  NANDN U3794 ( .A(n720), .B(n722), .Z(n709) );
  NANDN U3795 ( .A(n719), .B(n709), .Z(n710) );
  NAND U3796 ( .A(n711), .B(n710), .Z(n800) );
  XNOR U3797 ( .A(n765), .B(n800), .Z(n741) );
  AND U3798 ( .A(n712), .B(n741), .Z(n734) );
  OR U3799 ( .A(n719), .B(n716), .Z(n718) );
  ANDN U3800 ( .B(n719), .A(n713), .Z(n714) );
  XNOR U3801 ( .A(n714), .B(n724), .Z(n715) );
  NAND U3802 ( .A(n716), .B(n715), .Z(n717) );
  NAND U3803 ( .A(n718), .B(n717), .Z(n738) );
  NAND U3804 ( .A(n720), .B(n724), .Z(n726) );
  NAND U3805 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U3806 ( .A(n722), .B(n721), .Z(n723) );
  NANDN U3807 ( .A(n724), .B(n723), .Z(n725) );
  NAND U3808 ( .A(n726), .B(n725), .Z(n807) );
  NAND U3809 ( .A(n757), .B(n727), .Z(n728) );
  XNOR U3810 ( .A(n734), .B(n728), .Z(n802) );
  XOR U3811 ( .A(n765), .B(n807), .Z(n767) );
  AND U3812 ( .A(n729), .B(n767), .Z(n752) );
  XNOR U3813 ( .A(n802), .B(n752), .Z(n730) );
  XNOR U3814 ( .A(n731), .B(n730), .Z(n810) );
  NAND U3815 ( .A(n743), .B(n732), .Z(n733) );
  XNOR U3816 ( .A(n734), .B(n733), .Z(n760) );
  AND U3817 ( .A(n735), .B(n745), .Z(n801) );
  NANDN U3818 ( .A(n736), .B(n738), .Z(n737) );
  XNOR U3819 ( .A(n801), .B(n737), .Z(n764) );
  XNOR U3820 ( .A(n760), .B(n764), .Z(n749) );
  XOR U3821 ( .A(n810), .B(n749), .Z(z[16]) );
  AND U3822 ( .A(n739), .B(n738), .Z(n748) );
  AND U3823 ( .A(n741), .B(n740), .Z(n759) );
  NAND U3824 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U3825 ( .A(n759), .B(n744), .Z(n811) );
  AND U3826 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U3827 ( .A(n811), .B(n753), .Z(n747) );
  XNOR U3828 ( .A(n748), .B(n747), .Z(n773) );
  XNOR U3829 ( .A(n773), .B(n749), .Z(n816) );
  AND U3830 ( .A(n750), .B(n800), .Z(n755) );
  NANDN U3831 ( .A(n807), .B(n805), .Z(n751) );
  XNOR U3832 ( .A(n752), .B(n751), .Z(n763) );
  XNOR U3833 ( .A(n753), .B(n763), .Z(n754) );
  XNOR U3834 ( .A(n755), .B(n754), .Z(n762) );
  NAND U3835 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U3836 ( .A(n759), .B(n758), .Z(n769) );
  XNOR U3837 ( .A(n760), .B(n769), .Z(n761) );
  XNOR U3838 ( .A(n762), .B(n761), .Z(n772) );
  XNOR U3839 ( .A(n816), .B(n772), .Z(z[17]) );
  XNOR U3840 ( .A(n764), .B(n763), .Z(z[18]) );
  NOR U3841 ( .A(n766), .B(n765), .Z(n771) );
  AND U3842 ( .A(n768), .B(n767), .Z(n809) );
  XNOR U3843 ( .A(n769), .B(n809), .Z(n770) );
  XNOR U3844 ( .A(n771), .B(n770), .Z(n815) );
  XOR U3845 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U3846 ( .A(n815), .B(n774), .Z(z[19]) );
  AND U3847 ( .A(n776), .B(n775), .Z(n785) );
  AND U3848 ( .A(n778), .B(n777), .Z(n796) );
  NAND U3849 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U3850 ( .A(n796), .B(n781), .Z(n1438) );
  AND U3851 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U3852 ( .A(n1438), .B(n790), .Z(n784) );
  XNOR U3853 ( .A(n785), .B(n784), .Z(n1074) );
  XNOR U3854 ( .A(n1074), .B(n786), .Z(n1581) );
  AND U3855 ( .A(n787), .B(n1427), .Z(n792) );
  NANDN U3856 ( .A(n1434), .B(n1432), .Z(n788) );
  XNOR U3857 ( .A(n789), .B(n788), .Z(n938) );
  XNOR U3858 ( .A(n790), .B(n938), .Z(n791) );
  XNOR U3859 ( .A(n792), .B(n791), .Z(n799) );
  NAND U3860 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U3861 ( .A(n796), .B(n795), .Z(n1070) );
  XNOR U3862 ( .A(n797), .B(n1070), .Z(n798) );
  XNOR U3863 ( .A(n799), .B(n798), .Z(n1073) );
  XNOR U3864 ( .A(n1581), .B(n1073), .Z(z[1]) );
  XOR U3865 ( .A(n810), .B(z[18]), .Z(z[20]) );
  AND U3866 ( .A(x[16]), .B(n800), .Z(n804) );
  XNOR U3867 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U3868 ( .A(n804), .B(n803), .Z(n817) );
  XOR U3869 ( .A(n805), .B(x[17]), .Z(n806) );
  NANDN U3870 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3871 ( .A(n809), .B(n808), .Z(n813) );
  XNOR U3872 ( .A(n811), .B(n810), .Z(n812) );
  XNOR U3873 ( .A(n813), .B(n812), .Z(n814) );
  XNOR U3874 ( .A(n817), .B(n814), .Z(z[21]) );
  XNOR U3875 ( .A(n816), .B(n815), .Z(z[22]) );
  XOR U3876 ( .A(n817), .B(z[17]), .Z(z[23]) );
  XOR U3877 ( .A(x[27]), .B(x[25]), .Z(n820) );
  XNOR U3878 ( .A(x[24]), .B(x[30]), .Z(n819) );
  XOR U3879 ( .A(n819), .B(x[26]), .Z(n818) );
  XNOR U3880 ( .A(n820), .B(n818), .Z(n855) );
  XNOR U3881 ( .A(x[29]), .B(n819), .Z(n928) );
  XOR U3882 ( .A(n928), .B(x[28]), .Z(n898) );
  IV U3883 ( .A(n898), .Z(n829) );
  XNOR U3884 ( .A(x[31]), .B(x[28]), .Z(n823) );
  XNOR U3885 ( .A(n820), .B(n823), .Z(n883) );
  NOR U3886 ( .A(n829), .B(n883), .Z(n822) );
  XNOR U3887 ( .A(n928), .B(x[31]), .Z(n914) );
  XNOR U3888 ( .A(x[26]), .B(n914), .Z(n838) );
  XNOR U3889 ( .A(x[25]), .B(n838), .Z(n833) );
  AND U3890 ( .A(x[24]), .B(n833), .Z(n821) );
  XNOR U3891 ( .A(n822), .B(n821), .Z(n826) );
  XNOR U3892 ( .A(n855), .B(n914), .Z(n845) );
  IV U3893 ( .A(n855), .Z(n840) );
  XNOR U3894 ( .A(x[24]), .B(n840), .Z(n860) );
  IV U3895 ( .A(n823), .Z(n888) );
  AND U3896 ( .A(n860), .B(n888), .Z(n828) );
  IV U3897 ( .A(n928), .Z(n847) );
  XNOR U3898 ( .A(n855), .B(n847), .Z(n877) );
  XOR U3899 ( .A(n877), .B(n883), .Z(n880) );
  XOR U3900 ( .A(x[26]), .B(x[28]), .Z(n890) );
  NAND U3901 ( .A(n880), .B(n890), .Z(n824) );
  XNOR U3902 ( .A(n828), .B(n824), .Z(n849) );
  XNOR U3903 ( .A(n845), .B(n849), .Z(n825) );
  XNOR U3904 ( .A(n826), .B(n825), .Z(n872) );
  XOR U3905 ( .A(x[26]), .B(x[31]), .Z(n904) );
  XNOR U3906 ( .A(x[24]), .B(n883), .Z(n884) );
  XNOR U3907 ( .A(n928), .B(n884), .Z(n875) );
  NAND U3908 ( .A(n904), .B(n875), .Z(n827) );
  XNOR U3909 ( .A(n828), .B(n827), .Z(n841) );
  IV U3910 ( .A(n833), .Z(n887) );
  XNOR U3911 ( .A(n887), .B(n829), .Z(n894) );
  AND U3912 ( .A(n883), .B(n894), .Z(n831) );
  AND U3913 ( .A(x[24]), .B(n898), .Z(n830) );
  XNOR U3914 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U3915 ( .A(n884), .B(n832), .Z(n836) );
  NAND U3916 ( .A(x[24]), .B(n883), .Z(n834) );
  OR U3917 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3918 ( .A(n836), .B(n835), .Z(n837) );
  XNOR U3919 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U3920 ( .A(n841), .B(n839), .Z(n861) );
  IV U3921 ( .A(n861), .Z(n868) );
  AND U3922 ( .A(n914), .B(n840), .Z(n843) );
  XOR U3923 ( .A(x[25]), .B(x[31]), .Z(n916) );
  AND U3924 ( .A(n877), .B(n916), .Z(n846) );
  XNOR U3925 ( .A(n846), .B(n841), .Z(n842) );
  XNOR U3926 ( .A(n843), .B(n842), .Z(n867) );
  NANDN U3927 ( .A(n868), .B(n867), .Z(n844) );
  NAND U3928 ( .A(n872), .B(n844), .Z(n854) );
  XNOR U3929 ( .A(n846), .B(n845), .Z(n851) );
  ANDN U3930 ( .B(n847), .A(x[25]), .Z(n848) );
  XNOR U3931 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U3932 ( .A(n851), .B(n850), .Z(n864) );
  XOR U3933 ( .A(n867), .B(n864), .Z(n852) );
  NAND U3934 ( .A(n868), .B(n852), .Z(n853) );
  NAND U3935 ( .A(n854), .B(n853), .Z(n913) );
  ANDN U3936 ( .B(n855), .A(n913), .Z(n879) );
  IV U3937 ( .A(n864), .Z(n870) );
  XOR U3938 ( .A(n872), .B(n868), .Z(n856) );
  NANDN U3939 ( .A(n870), .B(n856), .Z(n859) );
  NANDN U3940 ( .A(n868), .B(n870), .Z(n857) );
  NANDN U3941 ( .A(n867), .B(n857), .Z(n858) );
  NAND U3942 ( .A(n859), .B(n858), .Z(n923) );
  XNOR U3943 ( .A(n913), .B(n923), .Z(n889) );
  AND U3944 ( .A(n860), .B(n889), .Z(n882) );
  OR U3945 ( .A(n867), .B(n864), .Z(n866) );
  ANDN U3946 ( .B(n867), .A(n861), .Z(n862) );
  XNOR U3947 ( .A(n862), .B(n872), .Z(n863) );
  NAND U3948 ( .A(n864), .B(n863), .Z(n865) );
  NAND U3949 ( .A(n866), .B(n865), .Z(n886) );
  NAND U3950 ( .A(n868), .B(n872), .Z(n874) );
  NAND U3951 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U3952 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U3953 ( .A(n872), .B(n871), .Z(n873) );
  NAND U3954 ( .A(n874), .B(n873), .Z(n930) );
  NAND U3955 ( .A(n905), .B(n875), .Z(n876) );
  XNOR U3956 ( .A(n882), .B(n876), .Z(n925) );
  XOR U3957 ( .A(n913), .B(n930), .Z(n915) );
  AND U3958 ( .A(n877), .B(n915), .Z(n900) );
  XNOR U3959 ( .A(n925), .B(n900), .Z(n878) );
  XNOR U3960 ( .A(n879), .B(n878), .Z(n933) );
  NAND U3961 ( .A(n891), .B(n880), .Z(n881) );
  XNOR U3962 ( .A(n882), .B(n881), .Z(n908) );
  AND U3963 ( .A(n883), .B(n893), .Z(n924) );
  NANDN U3964 ( .A(n884), .B(n886), .Z(n885) );
  XNOR U3965 ( .A(n924), .B(n885), .Z(n912) );
  XNOR U3966 ( .A(n908), .B(n912), .Z(n897) );
  XOR U3967 ( .A(n933), .B(n897), .Z(z[24]) );
  AND U3968 ( .A(n887), .B(n886), .Z(n896) );
  AND U3969 ( .A(n889), .B(n888), .Z(n907) );
  NAND U3970 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U3971 ( .A(n907), .B(n892), .Z(n934) );
  AND U3972 ( .A(n894), .B(n893), .Z(n901) );
  XNOR U3973 ( .A(n934), .B(n901), .Z(n895) );
  XNOR U3974 ( .A(n896), .B(n895), .Z(n921) );
  XNOR U3975 ( .A(n921), .B(n897), .Z(n941) );
  AND U3976 ( .A(n898), .B(n923), .Z(n903) );
  NANDN U3977 ( .A(n930), .B(n928), .Z(n899) );
  XNOR U3978 ( .A(n900), .B(n899), .Z(n911) );
  XNOR U3979 ( .A(n901), .B(n911), .Z(n902) );
  XNOR U3980 ( .A(n903), .B(n902), .Z(n910) );
  NAND U3981 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3982 ( .A(n907), .B(n906), .Z(n917) );
  XNOR U3983 ( .A(n908), .B(n917), .Z(n909) );
  XNOR U3984 ( .A(n910), .B(n909), .Z(n920) );
  XNOR U3985 ( .A(n941), .B(n920), .Z(z[25]) );
  XNOR U3986 ( .A(n912), .B(n911), .Z(z[26]) );
  NOR U3987 ( .A(n914), .B(n913), .Z(n919) );
  AND U3988 ( .A(n916), .B(n915), .Z(n932) );
  XNOR U3989 ( .A(n917), .B(n932), .Z(n918) );
  XNOR U3990 ( .A(n919), .B(n918), .Z(n940) );
  XOR U3991 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U3992 ( .A(n940), .B(n922), .Z(z[27]) );
  XOR U3993 ( .A(n933), .B(z[26]), .Z(z[28]) );
  AND U3994 ( .A(x[24]), .B(n923), .Z(n927) );
  XNOR U3995 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U3996 ( .A(n927), .B(n926), .Z(n942) );
  XOR U3997 ( .A(n928), .B(x[25]), .Z(n929) );
  NANDN U3998 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U3999 ( .A(n932), .B(n931), .Z(n936) );
  XNOR U4000 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U4001 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U4002 ( .A(n942), .B(n937), .Z(z[29]) );
  XNOR U4003 ( .A(n939), .B(n938), .Z(z[2]) );
  XNOR U4004 ( .A(n941), .B(n940), .Z(z[30]) );
  XOR U4005 ( .A(n942), .B(z[25]), .Z(z[31]) );
  XOR U4006 ( .A(x[35]), .B(x[33]), .Z(n945) );
  XNOR U4007 ( .A(x[32]), .B(x[38]), .Z(n944) );
  XOR U4008 ( .A(n944), .B(x[34]), .Z(n943) );
  XNOR U4009 ( .A(n945), .B(n943), .Z(n980) );
  XNOR U4010 ( .A(x[37]), .B(n944), .Z(n1053) );
  XOR U4011 ( .A(n1053), .B(x[36]), .Z(n1023) );
  IV U4012 ( .A(n1023), .Z(n954) );
  XNOR U4013 ( .A(x[39]), .B(x[36]), .Z(n948) );
  XNOR U4014 ( .A(n945), .B(n948), .Z(n1008) );
  NOR U4015 ( .A(n954), .B(n1008), .Z(n947) );
  XNOR U4016 ( .A(n1053), .B(x[39]), .Z(n1039) );
  XNOR U4017 ( .A(x[34]), .B(n1039), .Z(n963) );
  XNOR U4018 ( .A(x[33]), .B(n963), .Z(n958) );
  AND U4019 ( .A(x[32]), .B(n958), .Z(n946) );
  XNOR U4020 ( .A(n947), .B(n946), .Z(n951) );
  XNOR U4021 ( .A(n980), .B(n1039), .Z(n970) );
  IV U4022 ( .A(n980), .Z(n965) );
  XNOR U4023 ( .A(x[32]), .B(n965), .Z(n985) );
  IV U4024 ( .A(n948), .Z(n1013) );
  AND U4025 ( .A(n985), .B(n1013), .Z(n953) );
  IV U4026 ( .A(n1053), .Z(n972) );
  XNOR U4027 ( .A(n980), .B(n972), .Z(n1002) );
  XOR U4028 ( .A(n1002), .B(n1008), .Z(n1005) );
  XOR U4029 ( .A(x[34]), .B(x[36]), .Z(n1015) );
  NAND U4030 ( .A(n1005), .B(n1015), .Z(n949) );
  XNOR U4031 ( .A(n953), .B(n949), .Z(n974) );
  XNOR U4032 ( .A(n970), .B(n974), .Z(n950) );
  XNOR U4033 ( .A(n951), .B(n950), .Z(n997) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1029) );
  XNOR U4035 ( .A(x[32]), .B(n1008), .Z(n1009) );
  XNOR U4036 ( .A(n1053), .B(n1009), .Z(n1000) );
  NAND U4037 ( .A(n1029), .B(n1000), .Z(n952) );
  XNOR U4038 ( .A(n953), .B(n952), .Z(n966) );
  IV U4039 ( .A(n958), .Z(n1012) );
  XNOR U4040 ( .A(n1012), .B(n954), .Z(n1019) );
  AND U4041 ( .A(n1008), .B(n1019), .Z(n956) );
  AND U4042 ( .A(x[32]), .B(n1023), .Z(n955) );
  XNOR U4043 ( .A(n956), .B(n955), .Z(n957) );
  NANDN U4044 ( .A(n1009), .B(n957), .Z(n961) );
  NAND U4045 ( .A(x[32]), .B(n1008), .Z(n959) );
  OR U4046 ( .A(n959), .B(n958), .Z(n960) );
  NAND U4047 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U4048 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U4049 ( .A(n966), .B(n964), .Z(n986) );
  IV U4050 ( .A(n986), .Z(n993) );
  AND U4051 ( .A(n1039), .B(n965), .Z(n968) );
  XOR U4052 ( .A(x[33]), .B(x[39]), .Z(n1041) );
  AND U4053 ( .A(n1002), .B(n1041), .Z(n971) );
  XNOR U4054 ( .A(n971), .B(n966), .Z(n967) );
  XNOR U4055 ( .A(n968), .B(n967), .Z(n992) );
  NANDN U4056 ( .A(n993), .B(n992), .Z(n969) );
  NAND U4057 ( .A(n997), .B(n969), .Z(n979) );
  XNOR U4058 ( .A(n971), .B(n970), .Z(n976) );
  ANDN U4059 ( .B(n972), .A(x[33]), .Z(n973) );
  XNOR U4060 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U4061 ( .A(n976), .B(n975), .Z(n989) );
  XOR U4062 ( .A(n992), .B(n989), .Z(n977) );
  NAND U4063 ( .A(n993), .B(n977), .Z(n978) );
  NAND U4064 ( .A(n979), .B(n978), .Z(n1038) );
  ANDN U4065 ( .B(n980), .A(n1038), .Z(n1004) );
  IV U4066 ( .A(n989), .Z(n995) );
  XOR U4067 ( .A(n997), .B(n993), .Z(n981) );
  NANDN U4068 ( .A(n995), .B(n981), .Z(n984) );
  NANDN U4069 ( .A(n993), .B(n995), .Z(n982) );
  NANDN U4070 ( .A(n992), .B(n982), .Z(n983) );
  NAND U4071 ( .A(n984), .B(n983), .Z(n1048) );
  XNOR U4072 ( .A(n1038), .B(n1048), .Z(n1014) );
  AND U4073 ( .A(n985), .B(n1014), .Z(n1007) );
  OR U4074 ( .A(n992), .B(n989), .Z(n991) );
  ANDN U4075 ( .B(n992), .A(n986), .Z(n987) );
  XNOR U4076 ( .A(n987), .B(n997), .Z(n988) );
  NAND U4077 ( .A(n989), .B(n988), .Z(n990) );
  NAND U4078 ( .A(n991), .B(n990), .Z(n1011) );
  NAND U4079 ( .A(n993), .B(n997), .Z(n999) );
  NAND U4080 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U4081 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U4082 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4083 ( .A(n999), .B(n998), .Z(n1055) );
  NAND U4084 ( .A(n1030), .B(n1000), .Z(n1001) );
  XNOR U4085 ( .A(n1007), .B(n1001), .Z(n1050) );
  XOR U4086 ( .A(n1038), .B(n1055), .Z(n1040) );
  AND U4087 ( .A(n1002), .B(n1040), .Z(n1025) );
  XNOR U4088 ( .A(n1050), .B(n1025), .Z(n1003) );
  XNOR U4089 ( .A(n1004), .B(n1003), .Z(n1058) );
  NAND U4090 ( .A(n1016), .B(n1005), .Z(n1006) );
  XNOR U4091 ( .A(n1007), .B(n1006), .Z(n1033) );
  AND U4092 ( .A(n1008), .B(n1018), .Z(n1049) );
  NANDN U4093 ( .A(n1009), .B(n1011), .Z(n1010) );
  XNOR U4094 ( .A(n1049), .B(n1010), .Z(n1037) );
  XNOR U4095 ( .A(n1033), .B(n1037), .Z(n1022) );
  XOR U4096 ( .A(n1058), .B(n1022), .Z(z[32]) );
  AND U4097 ( .A(n1012), .B(n1011), .Z(n1021) );
  AND U4098 ( .A(n1014), .B(n1013), .Z(n1032) );
  NAND U4099 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U4100 ( .A(n1032), .B(n1017), .Z(n1059) );
  AND U4101 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U4102 ( .A(n1059), .B(n1026), .Z(n1020) );
  XNOR U4103 ( .A(n1021), .B(n1020), .Z(n1046) );
  XNOR U4104 ( .A(n1046), .B(n1022), .Z(n1064) );
  AND U4105 ( .A(n1023), .B(n1048), .Z(n1028) );
  NANDN U4106 ( .A(n1055), .B(n1053), .Z(n1024) );
  XNOR U4107 ( .A(n1025), .B(n1024), .Z(n1036) );
  XNOR U4108 ( .A(n1026), .B(n1036), .Z(n1027) );
  XNOR U4109 ( .A(n1028), .B(n1027), .Z(n1035) );
  NAND U4110 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U4111 ( .A(n1032), .B(n1031), .Z(n1042) );
  XNOR U4112 ( .A(n1033), .B(n1042), .Z(n1034) );
  XNOR U4113 ( .A(n1035), .B(n1034), .Z(n1045) );
  XNOR U4114 ( .A(n1064), .B(n1045), .Z(z[33]) );
  XNOR U4115 ( .A(n1037), .B(n1036), .Z(z[34]) );
  NOR U4116 ( .A(n1039), .B(n1038), .Z(n1044) );
  AND U4117 ( .A(n1041), .B(n1040), .Z(n1057) );
  XNOR U4118 ( .A(n1042), .B(n1057), .Z(n1043) );
  XNOR U4119 ( .A(n1044), .B(n1043), .Z(n1063) );
  XOR U4120 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U4121 ( .A(n1063), .B(n1047), .Z(z[35]) );
  XOR U4122 ( .A(n1058), .B(z[34]), .Z(z[36]) );
  AND U4123 ( .A(x[32]), .B(n1048), .Z(n1052) );
  XNOR U4124 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U4125 ( .A(n1052), .B(n1051), .Z(n1065) );
  XOR U4126 ( .A(n1053), .B(x[33]), .Z(n1054) );
  NANDN U4127 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U4128 ( .A(n1057), .B(n1056), .Z(n1061) );
  XNOR U4129 ( .A(n1059), .B(n1058), .Z(n1060) );
  XNOR U4130 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U4131 ( .A(n1065), .B(n1062), .Z(z[37]) );
  XNOR U4132 ( .A(n1064), .B(n1063), .Z(z[38]) );
  XOR U4133 ( .A(n1065), .B(z[33]), .Z(z[39]) );
  NOR U4134 ( .A(n1067), .B(n1066), .Z(n1072) );
  AND U4135 ( .A(n1069), .B(n1068), .Z(n1436) );
  XNOR U4136 ( .A(n1070), .B(n1436), .Z(n1071) );
  XNOR U4137 ( .A(n1072), .B(n1071), .Z(n1580) );
  XOR U4138 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U4139 ( .A(n1580), .B(n1075), .Z(z[3]) );
  XOR U4140 ( .A(x[43]), .B(x[41]), .Z(n1078) );
  XNOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1077) );
  XOR U4142 ( .A(n1077), .B(x[42]), .Z(n1076) );
  XNOR U4143 ( .A(n1078), .B(n1076), .Z(n1113) );
  XNOR U4144 ( .A(x[45]), .B(n1077), .Z(n1186) );
  XOR U4145 ( .A(n1186), .B(x[44]), .Z(n1156) );
  IV U4146 ( .A(n1156), .Z(n1087) );
  XNOR U4147 ( .A(x[47]), .B(x[44]), .Z(n1081) );
  XNOR U4148 ( .A(n1078), .B(n1081), .Z(n1141) );
  NOR U4149 ( .A(n1087), .B(n1141), .Z(n1080) );
  XNOR U4150 ( .A(n1186), .B(x[47]), .Z(n1172) );
  XNOR U4151 ( .A(x[42]), .B(n1172), .Z(n1096) );
  XNOR U4152 ( .A(x[41]), .B(n1096), .Z(n1091) );
  AND U4153 ( .A(x[40]), .B(n1091), .Z(n1079) );
  XNOR U4154 ( .A(n1080), .B(n1079), .Z(n1084) );
  XNOR U4155 ( .A(n1113), .B(n1172), .Z(n1103) );
  IV U4156 ( .A(n1113), .Z(n1098) );
  XNOR U4157 ( .A(x[40]), .B(n1098), .Z(n1118) );
  IV U4158 ( .A(n1081), .Z(n1146) );
  AND U4159 ( .A(n1118), .B(n1146), .Z(n1086) );
  IV U4160 ( .A(n1186), .Z(n1105) );
  XNOR U4161 ( .A(n1113), .B(n1105), .Z(n1135) );
  XOR U4162 ( .A(n1135), .B(n1141), .Z(n1138) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1148) );
  NAND U4164 ( .A(n1138), .B(n1148), .Z(n1082) );
  XNOR U4165 ( .A(n1086), .B(n1082), .Z(n1107) );
  XNOR U4166 ( .A(n1103), .B(n1107), .Z(n1083) );
  XNOR U4167 ( .A(n1084), .B(n1083), .Z(n1130) );
  XOR U4168 ( .A(x[42]), .B(x[47]), .Z(n1162) );
  XNOR U4169 ( .A(x[40]), .B(n1141), .Z(n1142) );
  XNOR U4170 ( .A(n1186), .B(n1142), .Z(n1133) );
  NAND U4171 ( .A(n1162), .B(n1133), .Z(n1085) );
  XNOR U4172 ( .A(n1086), .B(n1085), .Z(n1099) );
  IV U4173 ( .A(n1091), .Z(n1145) );
  XNOR U4174 ( .A(n1145), .B(n1087), .Z(n1152) );
  AND U4175 ( .A(n1141), .B(n1152), .Z(n1089) );
  AND U4176 ( .A(x[40]), .B(n1156), .Z(n1088) );
  XNOR U4177 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U4178 ( .A(n1142), .B(n1090), .Z(n1094) );
  NAND U4179 ( .A(x[40]), .B(n1141), .Z(n1092) );
  OR U4180 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U4181 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U4182 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U4183 ( .A(n1099), .B(n1097), .Z(n1119) );
  IV U4184 ( .A(n1119), .Z(n1126) );
  AND U4185 ( .A(n1172), .B(n1098), .Z(n1101) );
  XOR U4186 ( .A(x[41]), .B(x[47]), .Z(n1174) );
  AND U4187 ( .A(n1135), .B(n1174), .Z(n1104) );
  XNOR U4188 ( .A(n1104), .B(n1099), .Z(n1100) );
  XNOR U4189 ( .A(n1101), .B(n1100), .Z(n1125) );
  NANDN U4190 ( .A(n1126), .B(n1125), .Z(n1102) );
  NAND U4191 ( .A(n1130), .B(n1102), .Z(n1112) );
  XNOR U4192 ( .A(n1104), .B(n1103), .Z(n1109) );
  ANDN U4193 ( .B(n1105), .A(x[41]), .Z(n1106) );
  XNOR U4194 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U4195 ( .A(n1109), .B(n1108), .Z(n1122) );
  XOR U4196 ( .A(n1125), .B(n1122), .Z(n1110) );
  NAND U4197 ( .A(n1126), .B(n1110), .Z(n1111) );
  NAND U4198 ( .A(n1112), .B(n1111), .Z(n1171) );
  ANDN U4199 ( .B(n1113), .A(n1171), .Z(n1137) );
  IV U4200 ( .A(n1122), .Z(n1128) );
  XOR U4201 ( .A(n1130), .B(n1126), .Z(n1114) );
  NANDN U4202 ( .A(n1128), .B(n1114), .Z(n1117) );
  NANDN U4203 ( .A(n1126), .B(n1128), .Z(n1115) );
  NANDN U4204 ( .A(n1125), .B(n1115), .Z(n1116) );
  NAND U4205 ( .A(n1117), .B(n1116), .Z(n1181) );
  XNOR U4206 ( .A(n1171), .B(n1181), .Z(n1147) );
  AND U4207 ( .A(n1118), .B(n1147), .Z(n1140) );
  OR U4208 ( .A(n1125), .B(n1122), .Z(n1124) );
  ANDN U4209 ( .B(n1125), .A(n1119), .Z(n1120) );
  XNOR U4210 ( .A(n1120), .B(n1130), .Z(n1121) );
  NAND U4211 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U4212 ( .A(n1124), .B(n1123), .Z(n1144) );
  NAND U4213 ( .A(n1126), .B(n1130), .Z(n1132) );
  NAND U4214 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U4215 ( .A(n1128), .B(n1127), .Z(n1129) );
  NANDN U4216 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U4217 ( .A(n1132), .B(n1131), .Z(n1188) );
  NAND U4218 ( .A(n1163), .B(n1133), .Z(n1134) );
  XNOR U4219 ( .A(n1140), .B(n1134), .Z(n1183) );
  XOR U4220 ( .A(n1171), .B(n1188), .Z(n1173) );
  AND U4221 ( .A(n1135), .B(n1173), .Z(n1158) );
  XNOR U4222 ( .A(n1183), .B(n1158), .Z(n1136) );
  XNOR U4223 ( .A(n1137), .B(n1136), .Z(n1191) );
  NAND U4224 ( .A(n1149), .B(n1138), .Z(n1139) );
  XNOR U4225 ( .A(n1140), .B(n1139), .Z(n1166) );
  AND U4226 ( .A(n1141), .B(n1151), .Z(n1182) );
  NANDN U4227 ( .A(n1142), .B(n1144), .Z(n1143) );
  XNOR U4228 ( .A(n1182), .B(n1143), .Z(n1170) );
  XNOR U4229 ( .A(n1166), .B(n1170), .Z(n1155) );
  XOR U4230 ( .A(n1191), .B(n1155), .Z(z[40]) );
  AND U4231 ( .A(n1145), .B(n1144), .Z(n1154) );
  AND U4232 ( .A(n1147), .B(n1146), .Z(n1165) );
  NAND U4233 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U4234 ( .A(n1165), .B(n1150), .Z(n1192) );
  AND U4235 ( .A(n1152), .B(n1151), .Z(n1159) );
  XNOR U4236 ( .A(n1192), .B(n1159), .Z(n1153) );
  XNOR U4237 ( .A(n1154), .B(n1153), .Z(n1179) );
  XNOR U4238 ( .A(n1179), .B(n1155), .Z(n1197) );
  AND U4239 ( .A(n1156), .B(n1181), .Z(n1161) );
  NANDN U4240 ( .A(n1188), .B(n1186), .Z(n1157) );
  XNOR U4241 ( .A(n1158), .B(n1157), .Z(n1169) );
  XNOR U4242 ( .A(n1159), .B(n1169), .Z(n1160) );
  XNOR U4243 ( .A(n1161), .B(n1160), .Z(n1168) );
  NAND U4244 ( .A(n1163), .B(n1162), .Z(n1164) );
  XNOR U4245 ( .A(n1165), .B(n1164), .Z(n1175) );
  XNOR U4246 ( .A(n1166), .B(n1175), .Z(n1167) );
  XNOR U4247 ( .A(n1168), .B(n1167), .Z(n1178) );
  XNOR U4248 ( .A(n1197), .B(n1178), .Z(z[41]) );
  XNOR U4249 ( .A(n1170), .B(n1169), .Z(z[42]) );
  NOR U4250 ( .A(n1172), .B(n1171), .Z(n1177) );
  AND U4251 ( .A(n1174), .B(n1173), .Z(n1190) );
  XNOR U4252 ( .A(n1175), .B(n1190), .Z(n1176) );
  XNOR U4253 ( .A(n1177), .B(n1176), .Z(n1196) );
  XOR U4254 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4255 ( .A(n1196), .B(n1180), .Z(z[43]) );
  XOR U4256 ( .A(n1191), .B(z[42]), .Z(z[44]) );
  AND U4257 ( .A(x[40]), .B(n1181), .Z(n1185) );
  XNOR U4258 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U4259 ( .A(n1185), .B(n1184), .Z(n1198) );
  XOR U4260 ( .A(n1186), .B(x[41]), .Z(n1187) );
  NANDN U4261 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U4262 ( .A(n1190), .B(n1189), .Z(n1194) );
  XNOR U4263 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U4264 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U4265 ( .A(n1198), .B(n1195), .Z(z[45]) );
  XNOR U4266 ( .A(n1197), .B(n1196), .Z(z[46]) );
  XOR U4267 ( .A(n1198), .B(z[41]), .Z(z[47]) );
  XOR U4268 ( .A(x[51]), .B(x[49]), .Z(n1201) );
  XNOR U4269 ( .A(x[48]), .B(x[54]), .Z(n1200) );
  XOR U4270 ( .A(n1200), .B(x[50]), .Z(n1199) );
  XNOR U4271 ( .A(n1201), .B(n1199), .Z(n1236) );
  XNOR U4272 ( .A(x[53]), .B(n1200), .Z(n1309) );
  XOR U4273 ( .A(n1309), .B(x[52]), .Z(n1279) );
  IV U4274 ( .A(n1279), .Z(n1210) );
  XNOR U4275 ( .A(x[55]), .B(x[52]), .Z(n1204) );
  XNOR U4276 ( .A(n1201), .B(n1204), .Z(n1264) );
  NOR U4277 ( .A(n1210), .B(n1264), .Z(n1203) );
  XNOR U4278 ( .A(n1309), .B(x[55]), .Z(n1295) );
  XNOR U4279 ( .A(x[50]), .B(n1295), .Z(n1219) );
  XNOR U4280 ( .A(x[49]), .B(n1219), .Z(n1214) );
  AND U4281 ( .A(x[48]), .B(n1214), .Z(n1202) );
  XNOR U4282 ( .A(n1203), .B(n1202), .Z(n1207) );
  XNOR U4283 ( .A(n1236), .B(n1295), .Z(n1226) );
  IV U4284 ( .A(n1236), .Z(n1221) );
  XNOR U4285 ( .A(x[48]), .B(n1221), .Z(n1241) );
  IV U4286 ( .A(n1204), .Z(n1269) );
  AND U4287 ( .A(n1241), .B(n1269), .Z(n1209) );
  IV U4288 ( .A(n1309), .Z(n1228) );
  XNOR U4289 ( .A(n1236), .B(n1228), .Z(n1258) );
  XOR U4290 ( .A(n1258), .B(n1264), .Z(n1261) );
  XOR U4291 ( .A(x[50]), .B(x[52]), .Z(n1271) );
  NAND U4292 ( .A(n1261), .B(n1271), .Z(n1205) );
  XNOR U4293 ( .A(n1209), .B(n1205), .Z(n1230) );
  XNOR U4294 ( .A(n1226), .B(n1230), .Z(n1206) );
  XNOR U4295 ( .A(n1207), .B(n1206), .Z(n1253) );
  XOR U4296 ( .A(x[50]), .B(x[55]), .Z(n1285) );
  XNOR U4297 ( .A(x[48]), .B(n1264), .Z(n1265) );
  XNOR U4298 ( .A(n1309), .B(n1265), .Z(n1256) );
  NAND U4299 ( .A(n1285), .B(n1256), .Z(n1208) );
  XNOR U4300 ( .A(n1209), .B(n1208), .Z(n1222) );
  IV U4301 ( .A(n1214), .Z(n1268) );
  XNOR U4302 ( .A(n1268), .B(n1210), .Z(n1275) );
  AND U4303 ( .A(n1264), .B(n1275), .Z(n1212) );
  AND U4304 ( .A(x[48]), .B(n1279), .Z(n1211) );
  XNOR U4305 ( .A(n1212), .B(n1211), .Z(n1213) );
  NANDN U4306 ( .A(n1265), .B(n1213), .Z(n1217) );
  NAND U4307 ( .A(x[48]), .B(n1264), .Z(n1215) );
  OR U4308 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4309 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U4310 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U4311 ( .A(n1222), .B(n1220), .Z(n1242) );
  IV U4312 ( .A(n1242), .Z(n1249) );
  AND U4313 ( .A(n1295), .B(n1221), .Z(n1224) );
  XOR U4314 ( .A(x[49]), .B(x[55]), .Z(n1297) );
  AND U4315 ( .A(n1258), .B(n1297), .Z(n1227) );
  XNOR U4316 ( .A(n1227), .B(n1222), .Z(n1223) );
  XNOR U4317 ( .A(n1224), .B(n1223), .Z(n1248) );
  NANDN U4318 ( .A(n1249), .B(n1248), .Z(n1225) );
  NAND U4319 ( .A(n1253), .B(n1225), .Z(n1235) );
  XNOR U4320 ( .A(n1227), .B(n1226), .Z(n1232) );
  ANDN U4321 ( .B(n1228), .A(x[49]), .Z(n1229) );
  XNOR U4322 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U4323 ( .A(n1232), .B(n1231), .Z(n1245) );
  XOR U4324 ( .A(n1248), .B(n1245), .Z(n1233) );
  NAND U4325 ( .A(n1249), .B(n1233), .Z(n1234) );
  NAND U4326 ( .A(n1235), .B(n1234), .Z(n1294) );
  ANDN U4327 ( .B(n1236), .A(n1294), .Z(n1260) );
  IV U4328 ( .A(n1245), .Z(n1251) );
  XOR U4329 ( .A(n1253), .B(n1249), .Z(n1237) );
  NANDN U4330 ( .A(n1251), .B(n1237), .Z(n1240) );
  NANDN U4331 ( .A(n1249), .B(n1251), .Z(n1238) );
  NANDN U4332 ( .A(n1248), .B(n1238), .Z(n1239) );
  NAND U4333 ( .A(n1240), .B(n1239), .Z(n1304) );
  XNOR U4334 ( .A(n1294), .B(n1304), .Z(n1270) );
  AND U4335 ( .A(n1241), .B(n1270), .Z(n1263) );
  OR U4336 ( .A(n1248), .B(n1245), .Z(n1247) );
  ANDN U4337 ( .B(n1248), .A(n1242), .Z(n1243) );
  XNOR U4338 ( .A(n1243), .B(n1253), .Z(n1244) );
  NAND U4339 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U4340 ( .A(n1247), .B(n1246), .Z(n1267) );
  NAND U4341 ( .A(n1249), .B(n1253), .Z(n1255) );
  NAND U4342 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U4343 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U4344 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U4345 ( .A(n1255), .B(n1254), .Z(n1311) );
  NAND U4346 ( .A(n1286), .B(n1256), .Z(n1257) );
  XNOR U4347 ( .A(n1263), .B(n1257), .Z(n1306) );
  XOR U4348 ( .A(n1294), .B(n1311), .Z(n1296) );
  AND U4349 ( .A(n1258), .B(n1296), .Z(n1281) );
  XNOR U4350 ( .A(n1306), .B(n1281), .Z(n1259) );
  XNOR U4351 ( .A(n1260), .B(n1259), .Z(n1314) );
  NAND U4352 ( .A(n1272), .B(n1261), .Z(n1262) );
  XNOR U4353 ( .A(n1263), .B(n1262), .Z(n1289) );
  AND U4354 ( .A(n1264), .B(n1274), .Z(n1305) );
  NANDN U4355 ( .A(n1265), .B(n1267), .Z(n1266) );
  XNOR U4356 ( .A(n1305), .B(n1266), .Z(n1293) );
  XNOR U4357 ( .A(n1289), .B(n1293), .Z(n1278) );
  XOR U4358 ( .A(n1314), .B(n1278), .Z(z[48]) );
  AND U4359 ( .A(n1268), .B(n1267), .Z(n1277) );
  AND U4360 ( .A(n1270), .B(n1269), .Z(n1288) );
  NAND U4361 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U4362 ( .A(n1288), .B(n1273), .Z(n1315) );
  AND U4363 ( .A(n1275), .B(n1274), .Z(n1282) );
  XNOR U4364 ( .A(n1315), .B(n1282), .Z(n1276) );
  XNOR U4365 ( .A(n1277), .B(n1276), .Z(n1302) );
  XNOR U4366 ( .A(n1302), .B(n1278), .Z(n1320) );
  AND U4367 ( .A(n1279), .B(n1304), .Z(n1284) );
  NANDN U4368 ( .A(n1311), .B(n1309), .Z(n1280) );
  XNOR U4369 ( .A(n1281), .B(n1280), .Z(n1292) );
  XNOR U4370 ( .A(n1282), .B(n1292), .Z(n1283) );
  XNOR U4371 ( .A(n1284), .B(n1283), .Z(n1291) );
  NAND U4372 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U4373 ( .A(n1288), .B(n1287), .Z(n1298) );
  XNOR U4374 ( .A(n1289), .B(n1298), .Z(n1290) );
  XNOR U4375 ( .A(n1291), .B(n1290), .Z(n1301) );
  XNOR U4376 ( .A(n1320), .B(n1301), .Z(z[49]) );
  XOR U4377 ( .A(n1437), .B(z[2]), .Z(z[4]) );
  XNOR U4378 ( .A(n1293), .B(n1292), .Z(z[50]) );
  NOR U4379 ( .A(n1295), .B(n1294), .Z(n1300) );
  AND U4380 ( .A(n1297), .B(n1296), .Z(n1313) );
  XNOR U4381 ( .A(n1298), .B(n1313), .Z(n1299) );
  XNOR U4382 ( .A(n1300), .B(n1299), .Z(n1319) );
  XOR U4383 ( .A(n1302), .B(n1301), .Z(n1303) );
  XNOR U4384 ( .A(n1319), .B(n1303), .Z(z[51]) );
  XOR U4385 ( .A(n1314), .B(z[50]), .Z(z[52]) );
  AND U4386 ( .A(x[48]), .B(n1304), .Z(n1308) );
  XNOR U4387 ( .A(n1306), .B(n1305), .Z(n1307) );
  XNOR U4388 ( .A(n1308), .B(n1307), .Z(n1321) );
  XOR U4389 ( .A(n1309), .B(x[49]), .Z(n1310) );
  NANDN U4390 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U4391 ( .A(n1313), .B(n1312), .Z(n1317) );
  XNOR U4392 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U4393 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U4394 ( .A(n1321), .B(n1318), .Z(z[53]) );
  XNOR U4395 ( .A(n1320), .B(n1319), .Z(z[54]) );
  XOR U4396 ( .A(n1321), .B(z[49]), .Z(z[55]) );
  XOR U4397 ( .A(x[59]), .B(x[57]), .Z(n1324) );
  XNOR U4398 ( .A(x[56]), .B(x[62]), .Z(n1323) );
  XOR U4399 ( .A(n1323), .B(x[58]), .Z(n1322) );
  XNOR U4400 ( .A(n1324), .B(n1322), .Z(n1359) );
  XNOR U4401 ( .A(x[61]), .B(n1323), .Z(n1447) );
  XOR U4402 ( .A(n1447), .B(x[60]), .Z(n1402) );
  IV U4403 ( .A(n1402), .Z(n1333) );
  XNOR U4404 ( .A(x[63]), .B(x[60]), .Z(n1327) );
  XNOR U4405 ( .A(n1324), .B(n1327), .Z(n1387) );
  NOR U4406 ( .A(n1333), .B(n1387), .Z(n1326) );
  XNOR U4407 ( .A(n1447), .B(x[63]), .Z(n1418) );
  XNOR U4408 ( .A(x[58]), .B(n1418), .Z(n1342) );
  XNOR U4409 ( .A(x[57]), .B(n1342), .Z(n1337) );
  AND U4410 ( .A(x[56]), .B(n1337), .Z(n1325) );
  XNOR U4411 ( .A(n1326), .B(n1325), .Z(n1330) );
  XNOR U4412 ( .A(n1359), .B(n1418), .Z(n1349) );
  IV U4413 ( .A(n1359), .Z(n1344) );
  XNOR U4414 ( .A(x[56]), .B(n1344), .Z(n1364) );
  IV U4415 ( .A(n1327), .Z(n1392) );
  AND U4416 ( .A(n1364), .B(n1392), .Z(n1332) );
  IV U4417 ( .A(n1447), .Z(n1351) );
  XNOR U4418 ( .A(n1359), .B(n1351), .Z(n1381) );
  XOR U4419 ( .A(n1381), .B(n1387), .Z(n1384) );
  XOR U4420 ( .A(x[58]), .B(x[60]), .Z(n1394) );
  NAND U4421 ( .A(n1384), .B(n1394), .Z(n1328) );
  XNOR U4422 ( .A(n1332), .B(n1328), .Z(n1353) );
  XNOR U4423 ( .A(n1349), .B(n1353), .Z(n1329) );
  XNOR U4424 ( .A(n1330), .B(n1329), .Z(n1376) );
  XOR U4425 ( .A(x[58]), .B(x[63]), .Z(n1408) );
  XNOR U4426 ( .A(x[56]), .B(n1387), .Z(n1388) );
  XNOR U4427 ( .A(n1447), .B(n1388), .Z(n1379) );
  NAND U4428 ( .A(n1408), .B(n1379), .Z(n1331) );
  XNOR U4429 ( .A(n1332), .B(n1331), .Z(n1345) );
  IV U4430 ( .A(n1337), .Z(n1391) );
  XNOR U4431 ( .A(n1391), .B(n1333), .Z(n1398) );
  AND U4432 ( .A(n1387), .B(n1398), .Z(n1335) );
  AND U4433 ( .A(x[56]), .B(n1402), .Z(n1334) );
  XNOR U4434 ( .A(n1335), .B(n1334), .Z(n1336) );
  NANDN U4435 ( .A(n1388), .B(n1336), .Z(n1340) );
  NAND U4436 ( .A(x[56]), .B(n1387), .Z(n1338) );
  OR U4437 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U4438 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4439 ( .A(n1342), .B(n1341), .Z(n1343) );
  XNOR U4440 ( .A(n1345), .B(n1343), .Z(n1365) );
  IV U4441 ( .A(n1365), .Z(n1372) );
  AND U4442 ( .A(n1418), .B(n1344), .Z(n1347) );
  XOR U4443 ( .A(x[57]), .B(x[63]), .Z(n1420) );
  AND U4444 ( .A(n1381), .B(n1420), .Z(n1350) );
  XNOR U4445 ( .A(n1350), .B(n1345), .Z(n1346) );
  XNOR U4446 ( .A(n1347), .B(n1346), .Z(n1371) );
  NANDN U4447 ( .A(n1372), .B(n1371), .Z(n1348) );
  NAND U4448 ( .A(n1376), .B(n1348), .Z(n1358) );
  XNOR U4449 ( .A(n1350), .B(n1349), .Z(n1355) );
  ANDN U4450 ( .B(n1351), .A(x[57]), .Z(n1352) );
  XNOR U4451 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U4452 ( .A(n1355), .B(n1354), .Z(n1368) );
  XOR U4453 ( .A(n1371), .B(n1368), .Z(n1356) );
  NAND U4454 ( .A(n1372), .B(n1356), .Z(n1357) );
  NAND U4455 ( .A(n1358), .B(n1357), .Z(n1417) );
  ANDN U4456 ( .B(n1359), .A(n1417), .Z(n1383) );
  IV U4457 ( .A(n1368), .Z(n1374) );
  XOR U4458 ( .A(n1376), .B(n1372), .Z(n1360) );
  NANDN U4459 ( .A(n1374), .B(n1360), .Z(n1363) );
  NANDN U4460 ( .A(n1372), .B(n1374), .Z(n1361) );
  NANDN U4461 ( .A(n1371), .B(n1361), .Z(n1362) );
  NAND U4462 ( .A(n1363), .B(n1362), .Z(n1442) );
  XNOR U4463 ( .A(n1417), .B(n1442), .Z(n1393) );
  AND U4464 ( .A(n1364), .B(n1393), .Z(n1386) );
  OR U4465 ( .A(n1371), .B(n1368), .Z(n1370) );
  ANDN U4466 ( .B(n1371), .A(n1365), .Z(n1366) );
  XNOR U4467 ( .A(n1366), .B(n1376), .Z(n1367) );
  NAND U4468 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U4469 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U4470 ( .A(n1372), .B(n1376), .Z(n1378) );
  NAND U4471 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4472 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U4473 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U4474 ( .A(n1378), .B(n1377), .Z(n1449) );
  NAND U4475 ( .A(n1409), .B(n1379), .Z(n1380) );
  XNOR U4476 ( .A(n1386), .B(n1380), .Z(n1444) );
  XOR U4477 ( .A(n1417), .B(n1449), .Z(n1419) );
  AND U4478 ( .A(n1381), .B(n1419), .Z(n1404) );
  XNOR U4479 ( .A(n1444), .B(n1404), .Z(n1382) );
  XNOR U4480 ( .A(n1383), .B(n1382), .Z(n1452) );
  NAND U4481 ( .A(n1395), .B(n1384), .Z(n1385) );
  XNOR U4482 ( .A(n1386), .B(n1385), .Z(n1412) );
  AND U4483 ( .A(n1387), .B(n1397), .Z(n1443) );
  NANDN U4484 ( .A(n1388), .B(n1390), .Z(n1389) );
  XNOR U4485 ( .A(n1443), .B(n1389), .Z(n1416) );
  XNOR U4486 ( .A(n1412), .B(n1416), .Z(n1401) );
  XOR U4487 ( .A(n1452), .B(n1401), .Z(z[56]) );
  AND U4488 ( .A(n1391), .B(n1390), .Z(n1400) );
  AND U4489 ( .A(n1393), .B(n1392), .Z(n1411) );
  NAND U4490 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U4491 ( .A(n1411), .B(n1396), .Z(n1453) );
  AND U4492 ( .A(n1398), .B(n1397), .Z(n1405) );
  XNOR U4493 ( .A(n1453), .B(n1405), .Z(n1399) );
  XNOR U4494 ( .A(n1400), .B(n1399), .Z(n1425) );
  XNOR U4495 ( .A(n1425), .B(n1401), .Z(n1458) );
  AND U4496 ( .A(n1402), .B(n1442), .Z(n1407) );
  NANDN U4497 ( .A(n1449), .B(n1447), .Z(n1403) );
  XNOR U4498 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U4499 ( .A(n1405), .B(n1415), .Z(n1406) );
  XNOR U4500 ( .A(n1407), .B(n1406), .Z(n1414) );
  NAND U4501 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U4502 ( .A(n1411), .B(n1410), .Z(n1421) );
  XNOR U4503 ( .A(n1412), .B(n1421), .Z(n1413) );
  XNOR U4504 ( .A(n1414), .B(n1413), .Z(n1424) );
  XNOR U4505 ( .A(n1458), .B(n1424), .Z(z[57]) );
  XNOR U4506 ( .A(n1416), .B(n1415), .Z(z[58]) );
  NOR U4507 ( .A(n1418), .B(n1417), .Z(n1423) );
  AND U4508 ( .A(n1420), .B(n1419), .Z(n1451) );
  XNOR U4509 ( .A(n1421), .B(n1451), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1457) );
  XOR U4511 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U4512 ( .A(n1457), .B(n1426), .Z(z[59]) );
  AND U4513 ( .A(x[0]), .B(n1427), .Z(n1431) );
  XNOR U4514 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U4515 ( .A(n1431), .B(n1430), .Z(n1708) );
  XOR U4516 ( .A(n1432), .B(x[1]), .Z(n1433) );
  NANDN U4517 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U4518 ( .A(n1436), .B(n1435), .Z(n1440) );
  XNOR U4519 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U4520 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U4521 ( .A(n1708), .B(n1441), .Z(z[5]) );
  XOR U4522 ( .A(n1452), .B(z[58]), .Z(z[60]) );
  AND U4523 ( .A(x[56]), .B(n1442), .Z(n1446) );
  XNOR U4524 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U4525 ( .A(n1446), .B(n1445), .Z(n1459) );
  XOR U4526 ( .A(n1447), .B(x[57]), .Z(n1448) );
  NANDN U4527 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U4528 ( .A(n1451), .B(n1450), .Z(n1455) );
  XNOR U4529 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U4530 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U4531 ( .A(n1459), .B(n1456), .Z(z[61]) );
  XNOR U4532 ( .A(n1458), .B(n1457), .Z(z[62]) );
  XOR U4533 ( .A(n1459), .B(z[57]), .Z(z[63]) );
  XOR U4534 ( .A(x[67]), .B(x[65]), .Z(n1462) );
  XNOR U4535 ( .A(x[64]), .B(x[70]), .Z(n1461) );
  XOR U4536 ( .A(n1461), .B(x[66]), .Z(n1460) );
  XNOR U4537 ( .A(n1462), .B(n1460), .Z(n1497) );
  XNOR U4538 ( .A(x[69]), .B(n1461), .Z(n1570) );
  XOR U4539 ( .A(n1570), .B(x[68]), .Z(n1540) );
  IV U4540 ( .A(n1540), .Z(n1471) );
  XNOR U4541 ( .A(x[71]), .B(x[68]), .Z(n1465) );
  XNOR U4542 ( .A(n1462), .B(n1465), .Z(n1525) );
  NOR U4543 ( .A(n1471), .B(n1525), .Z(n1464) );
  XNOR U4544 ( .A(n1570), .B(x[71]), .Z(n1556) );
  XNOR U4545 ( .A(x[66]), .B(n1556), .Z(n1480) );
  XNOR U4546 ( .A(x[65]), .B(n1480), .Z(n1475) );
  AND U4547 ( .A(x[64]), .B(n1475), .Z(n1463) );
  XNOR U4548 ( .A(n1464), .B(n1463), .Z(n1468) );
  XNOR U4549 ( .A(n1497), .B(n1556), .Z(n1487) );
  IV U4550 ( .A(n1497), .Z(n1482) );
  XNOR U4551 ( .A(x[64]), .B(n1482), .Z(n1502) );
  IV U4552 ( .A(n1465), .Z(n1530) );
  AND U4553 ( .A(n1502), .B(n1530), .Z(n1470) );
  IV U4554 ( .A(n1570), .Z(n1489) );
  XNOR U4555 ( .A(n1497), .B(n1489), .Z(n1519) );
  XOR U4556 ( .A(n1519), .B(n1525), .Z(n1522) );
  XOR U4557 ( .A(x[66]), .B(x[68]), .Z(n1532) );
  NAND U4558 ( .A(n1522), .B(n1532), .Z(n1466) );
  XNOR U4559 ( .A(n1470), .B(n1466), .Z(n1491) );
  XNOR U4560 ( .A(n1487), .B(n1491), .Z(n1467) );
  XNOR U4561 ( .A(n1468), .B(n1467), .Z(n1514) );
  XOR U4562 ( .A(x[66]), .B(x[71]), .Z(n1546) );
  XNOR U4563 ( .A(x[64]), .B(n1525), .Z(n1526) );
  XNOR U4564 ( .A(n1570), .B(n1526), .Z(n1517) );
  NAND U4565 ( .A(n1546), .B(n1517), .Z(n1469) );
  XNOR U4566 ( .A(n1470), .B(n1469), .Z(n1483) );
  IV U4567 ( .A(n1475), .Z(n1529) );
  XNOR U4568 ( .A(n1529), .B(n1471), .Z(n1536) );
  AND U4569 ( .A(n1525), .B(n1536), .Z(n1473) );
  AND U4570 ( .A(x[64]), .B(n1540), .Z(n1472) );
  XNOR U4571 ( .A(n1473), .B(n1472), .Z(n1474) );
  NANDN U4572 ( .A(n1526), .B(n1474), .Z(n1478) );
  NAND U4573 ( .A(x[64]), .B(n1525), .Z(n1476) );
  OR U4574 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U4575 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4576 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR U4577 ( .A(n1483), .B(n1481), .Z(n1503) );
  IV U4578 ( .A(n1503), .Z(n1510) );
  AND U4579 ( .A(n1556), .B(n1482), .Z(n1485) );
  XOR U4580 ( .A(x[65]), .B(x[71]), .Z(n1558) );
  AND U4581 ( .A(n1519), .B(n1558), .Z(n1488) );
  XNOR U4582 ( .A(n1488), .B(n1483), .Z(n1484) );
  XNOR U4583 ( .A(n1485), .B(n1484), .Z(n1509) );
  NANDN U4584 ( .A(n1510), .B(n1509), .Z(n1486) );
  NAND U4585 ( .A(n1514), .B(n1486), .Z(n1496) );
  XNOR U4586 ( .A(n1488), .B(n1487), .Z(n1493) );
  ANDN U4587 ( .B(n1489), .A(x[65]), .Z(n1490) );
  XNOR U4588 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U4589 ( .A(n1493), .B(n1492), .Z(n1506) );
  XOR U4590 ( .A(n1509), .B(n1506), .Z(n1494) );
  NAND U4591 ( .A(n1510), .B(n1494), .Z(n1495) );
  NAND U4592 ( .A(n1496), .B(n1495), .Z(n1555) );
  ANDN U4593 ( .B(n1497), .A(n1555), .Z(n1521) );
  IV U4594 ( .A(n1506), .Z(n1512) );
  XOR U4595 ( .A(n1514), .B(n1510), .Z(n1498) );
  NANDN U4596 ( .A(n1512), .B(n1498), .Z(n1501) );
  NANDN U4597 ( .A(n1510), .B(n1512), .Z(n1499) );
  NANDN U4598 ( .A(n1509), .B(n1499), .Z(n1500) );
  NAND U4599 ( .A(n1501), .B(n1500), .Z(n1565) );
  XNOR U4600 ( .A(n1555), .B(n1565), .Z(n1531) );
  AND U4601 ( .A(n1502), .B(n1531), .Z(n1524) );
  OR U4602 ( .A(n1509), .B(n1506), .Z(n1508) );
  ANDN U4603 ( .B(n1509), .A(n1503), .Z(n1504) );
  XNOR U4604 ( .A(n1504), .B(n1514), .Z(n1505) );
  NAND U4605 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U4606 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U4607 ( .A(n1510), .B(n1514), .Z(n1516) );
  NAND U4608 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4609 ( .A(n1512), .B(n1511), .Z(n1513) );
  NANDN U4610 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U4611 ( .A(n1516), .B(n1515), .Z(n1572) );
  NAND U4612 ( .A(n1547), .B(n1517), .Z(n1518) );
  XNOR U4613 ( .A(n1524), .B(n1518), .Z(n1567) );
  XOR U4614 ( .A(n1555), .B(n1572), .Z(n1557) );
  AND U4615 ( .A(n1519), .B(n1557), .Z(n1542) );
  XNOR U4616 ( .A(n1567), .B(n1542), .Z(n1520) );
  XNOR U4617 ( .A(n1521), .B(n1520), .Z(n1575) );
  NAND U4618 ( .A(n1533), .B(n1522), .Z(n1523) );
  XNOR U4619 ( .A(n1524), .B(n1523), .Z(n1550) );
  AND U4620 ( .A(n1525), .B(n1535), .Z(n1566) );
  NANDN U4621 ( .A(n1526), .B(n1528), .Z(n1527) );
  XNOR U4622 ( .A(n1566), .B(n1527), .Z(n1554) );
  XNOR U4623 ( .A(n1550), .B(n1554), .Z(n1539) );
  XOR U4624 ( .A(n1575), .B(n1539), .Z(z[64]) );
  AND U4625 ( .A(n1529), .B(n1528), .Z(n1538) );
  AND U4626 ( .A(n1531), .B(n1530), .Z(n1549) );
  NAND U4627 ( .A(n1533), .B(n1532), .Z(n1534) );
  XNOR U4628 ( .A(n1549), .B(n1534), .Z(n1576) );
  AND U4629 ( .A(n1536), .B(n1535), .Z(n1543) );
  XNOR U4630 ( .A(n1576), .B(n1543), .Z(n1537) );
  XNOR U4631 ( .A(n1538), .B(n1537), .Z(n1563) );
  XNOR U4632 ( .A(n1563), .B(n1539), .Z(n1583) );
  AND U4633 ( .A(n1540), .B(n1565), .Z(n1545) );
  NANDN U4634 ( .A(n1572), .B(n1570), .Z(n1541) );
  XNOR U4635 ( .A(n1542), .B(n1541), .Z(n1553) );
  XNOR U4636 ( .A(n1543), .B(n1553), .Z(n1544) );
  XNOR U4637 ( .A(n1545), .B(n1544), .Z(n1552) );
  NAND U4638 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U4639 ( .A(n1549), .B(n1548), .Z(n1559) );
  XNOR U4640 ( .A(n1550), .B(n1559), .Z(n1551) );
  XNOR U4641 ( .A(n1552), .B(n1551), .Z(n1562) );
  XNOR U4642 ( .A(n1583), .B(n1562), .Z(z[65]) );
  XNOR U4643 ( .A(n1554), .B(n1553), .Z(z[66]) );
  NOR U4644 ( .A(n1556), .B(n1555), .Z(n1561) );
  AND U4645 ( .A(n1558), .B(n1557), .Z(n1574) );
  XNOR U4646 ( .A(n1559), .B(n1574), .Z(n1560) );
  XNOR U4647 ( .A(n1561), .B(n1560), .Z(n1582) );
  XOR U4648 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U4649 ( .A(n1582), .B(n1564), .Z(z[67]) );
  XOR U4650 ( .A(n1575), .B(z[66]), .Z(z[68]) );
  AND U4651 ( .A(x[64]), .B(n1565), .Z(n1569) );
  XNOR U4652 ( .A(n1567), .B(n1566), .Z(n1568) );
  XNOR U4653 ( .A(n1569), .B(n1568), .Z(n1584) );
  XOR U4654 ( .A(n1570), .B(x[65]), .Z(n1571) );
  NANDN U4655 ( .A(n1572), .B(n1571), .Z(n1573) );
  XNOR U4656 ( .A(n1574), .B(n1573), .Z(n1578) );
  XNOR U4657 ( .A(n1576), .B(n1575), .Z(n1577) );
  XNOR U4658 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U4659 ( .A(n1584), .B(n1579), .Z(z[69]) );
  XNOR U4660 ( .A(n1581), .B(n1580), .Z(z[6]) );
  XNOR U4661 ( .A(n1583), .B(n1582), .Z(z[70]) );
  XOR U4662 ( .A(n1584), .B(z[65]), .Z(z[71]) );
  XOR U4663 ( .A(x[75]), .B(x[73]), .Z(n1587) );
  XNOR U4664 ( .A(x[72]), .B(x[78]), .Z(n1586) );
  XOR U4665 ( .A(n1586), .B(x[74]), .Z(n1585) );
  XNOR U4666 ( .A(n1587), .B(n1585), .Z(n1622) );
  XNOR U4667 ( .A(x[77]), .B(n1586), .Z(n1695) );
  XOR U4668 ( .A(n1695), .B(x[76]), .Z(n1665) );
  IV U4669 ( .A(n1665), .Z(n1596) );
  XNOR U4670 ( .A(x[79]), .B(x[76]), .Z(n1590) );
  XNOR U4671 ( .A(n1587), .B(n1590), .Z(n1650) );
  NOR U4672 ( .A(n1596), .B(n1650), .Z(n1589) );
  XNOR U4673 ( .A(n1695), .B(x[79]), .Z(n1681) );
  XNOR U4674 ( .A(x[74]), .B(n1681), .Z(n1605) );
  XNOR U4675 ( .A(x[73]), .B(n1605), .Z(n1600) );
  AND U4676 ( .A(x[72]), .B(n1600), .Z(n1588) );
  XNOR U4677 ( .A(n1589), .B(n1588), .Z(n1593) );
  XNOR U4678 ( .A(n1622), .B(n1681), .Z(n1612) );
  IV U4679 ( .A(n1622), .Z(n1607) );
  XNOR U4680 ( .A(x[72]), .B(n1607), .Z(n1627) );
  IV U4681 ( .A(n1590), .Z(n1655) );
  AND U4682 ( .A(n1627), .B(n1655), .Z(n1595) );
  IV U4683 ( .A(n1695), .Z(n1614) );
  XNOR U4684 ( .A(n1622), .B(n1614), .Z(n1644) );
  XOR U4685 ( .A(n1644), .B(n1650), .Z(n1647) );
  XOR U4686 ( .A(x[74]), .B(x[76]), .Z(n1657) );
  NAND U4687 ( .A(n1647), .B(n1657), .Z(n1591) );
  XNOR U4688 ( .A(n1595), .B(n1591), .Z(n1616) );
  XNOR U4689 ( .A(n1612), .B(n1616), .Z(n1592) );
  XNOR U4690 ( .A(n1593), .B(n1592), .Z(n1639) );
  XOR U4691 ( .A(x[74]), .B(x[79]), .Z(n1671) );
  XNOR U4692 ( .A(x[72]), .B(n1650), .Z(n1651) );
  XNOR U4693 ( .A(n1695), .B(n1651), .Z(n1642) );
  NAND U4694 ( .A(n1671), .B(n1642), .Z(n1594) );
  XNOR U4695 ( .A(n1595), .B(n1594), .Z(n1608) );
  IV U4696 ( .A(n1600), .Z(n1654) );
  XNOR U4697 ( .A(n1654), .B(n1596), .Z(n1661) );
  AND U4698 ( .A(n1650), .B(n1661), .Z(n1598) );
  AND U4699 ( .A(x[72]), .B(n1665), .Z(n1597) );
  XNOR U4700 ( .A(n1598), .B(n1597), .Z(n1599) );
  NANDN U4701 ( .A(n1651), .B(n1599), .Z(n1603) );
  NAND U4702 ( .A(x[72]), .B(n1650), .Z(n1601) );
  OR U4703 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U4704 ( .A(n1603), .B(n1602), .Z(n1604) );
  XNOR U4705 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U4706 ( .A(n1608), .B(n1606), .Z(n1628) );
  IV U4707 ( .A(n1628), .Z(n1635) );
  AND U4708 ( .A(n1681), .B(n1607), .Z(n1610) );
  XOR U4709 ( .A(x[73]), .B(x[79]), .Z(n1683) );
  AND U4710 ( .A(n1644), .B(n1683), .Z(n1613) );
  XNOR U4711 ( .A(n1613), .B(n1608), .Z(n1609) );
  XNOR U4712 ( .A(n1610), .B(n1609), .Z(n1634) );
  NANDN U4713 ( .A(n1635), .B(n1634), .Z(n1611) );
  NAND U4714 ( .A(n1639), .B(n1611), .Z(n1621) );
  XNOR U4715 ( .A(n1613), .B(n1612), .Z(n1618) );
  ANDN U4716 ( .B(n1614), .A(x[73]), .Z(n1615) );
  XNOR U4717 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4718 ( .A(n1618), .B(n1617), .Z(n1631) );
  XOR U4719 ( .A(n1634), .B(n1631), .Z(n1619) );
  NAND U4720 ( .A(n1635), .B(n1619), .Z(n1620) );
  NAND U4721 ( .A(n1621), .B(n1620), .Z(n1680) );
  ANDN U4722 ( .B(n1622), .A(n1680), .Z(n1646) );
  IV U4723 ( .A(n1631), .Z(n1637) );
  XOR U4724 ( .A(n1639), .B(n1635), .Z(n1623) );
  NANDN U4725 ( .A(n1637), .B(n1623), .Z(n1626) );
  NANDN U4726 ( .A(n1635), .B(n1637), .Z(n1624) );
  NANDN U4727 ( .A(n1634), .B(n1624), .Z(n1625) );
  NAND U4728 ( .A(n1626), .B(n1625), .Z(n1690) );
  XNOR U4729 ( .A(n1680), .B(n1690), .Z(n1656) );
  AND U4730 ( .A(n1627), .B(n1656), .Z(n1649) );
  OR U4731 ( .A(n1634), .B(n1631), .Z(n1633) );
  ANDN U4732 ( .B(n1634), .A(n1628), .Z(n1629) );
  XNOR U4733 ( .A(n1629), .B(n1639), .Z(n1630) );
  NAND U4734 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U4735 ( .A(n1633), .B(n1632), .Z(n1653) );
  NAND U4736 ( .A(n1635), .B(n1639), .Z(n1641) );
  NAND U4737 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U4738 ( .A(n1637), .B(n1636), .Z(n1638) );
  NANDN U4739 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U4740 ( .A(n1641), .B(n1640), .Z(n1697) );
  NAND U4741 ( .A(n1672), .B(n1642), .Z(n1643) );
  XNOR U4742 ( .A(n1649), .B(n1643), .Z(n1692) );
  XOR U4743 ( .A(n1680), .B(n1697), .Z(n1682) );
  AND U4744 ( .A(n1644), .B(n1682), .Z(n1667) );
  XNOR U4745 ( .A(n1692), .B(n1667), .Z(n1645) );
  XNOR U4746 ( .A(n1646), .B(n1645), .Z(n1700) );
  NAND U4747 ( .A(n1658), .B(n1647), .Z(n1648) );
  XNOR U4748 ( .A(n1649), .B(n1648), .Z(n1675) );
  AND U4749 ( .A(n1650), .B(n1660), .Z(n1691) );
  NANDN U4750 ( .A(n1651), .B(n1653), .Z(n1652) );
  XNOR U4751 ( .A(n1691), .B(n1652), .Z(n1679) );
  XNOR U4752 ( .A(n1675), .B(n1679), .Z(n1664) );
  XOR U4753 ( .A(n1700), .B(n1664), .Z(z[72]) );
  AND U4754 ( .A(n1654), .B(n1653), .Z(n1663) );
  AND U4755 ( .A(n1656), .B(n1655), .Z(n1674) );
  NAND U4756 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U4757 ( .A(n1674), .B(n1659), .Z(n1701) );
  AND U4758 ( .A(n1661), .B(n1660), .Z(n1668) );
  XNOR U4759 ( .A(n1701), .B(n1668), .Z(n1662) );
  XNOR U4760 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U4761 ( .A(n1688), .B(n1664), .Z(n1706) );
  AND U4762 ( .A(n1665), .B(n1690), .Z(n1670) );
  NANDN U4763 ( .A(n1697), .B(n1695), .Z(n1666) );
  XNOR U4764 ( .A(n1667), .B(n1666), .Z(n1678) );
  XNOR U4765 ( .A(n1668), .B(n1678), .Z(n1669) );
  XNOR U4766 ( .A(n1670), .B(n1669), .Z(n1677) );
  NAND U4767 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR U4768 ( .A(n1674), .B(n1673), .Z(n1684) );
  XNOR U4769 ( .A(n1675), .B(n1684), .Z(n1676) );
  XNOR U4770 ( .A(n1677), .B(n1676), .Z(n1687) );
  XNOR U4771 ( .A(n1706), .B(n1687), .Z(z[73]) );
  XNOR U4772 ( .A(n1679), .B(n1678), .Z(z[74]) );
  NOR U4773 ( .A(n1681), .B(n1680), .Z(n1686) );
  AND U4774 ( .A(n1683), .B(n1682), .Z(n1699) );
  XNOR U4775 ( .A(n1684), .B(n1699), .Z(n1685) );
  XNOR U4776 ( .A(n1686), .B(n1685), .Z(n1705) );
  XOR U4777 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4778 ( .A(n1705), .B(n1689), .Z(z[75]) );
  XOR U4779 ( .A(n1700), .B(z[74]), .Z(z[76]) );
  AND U4780 ( .A(x[72]), .B(n1690), .Z(n1694) );
  XNOR U4781 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4782 ( .A(n1694), .B(n1693), .Z(n1707) );
  XOR U4783 ( .A(n1695), .B(x[73]), .Z(n1696) );
  NANDN U4784 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U4785 ( .A(n1699), .B(n1698), .Z(n1703) );
  XNOR U4786 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U4787 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U4788 ( .A(n1707), .B(n1704), .Z(z[77]) );
  XNOR U4789 ( .A(n1706), .B(n1705), .Z(z[78]) );
  XOR U4790 ( .A(n1707), .B(z[73]), .Z(z[79]) );
  XOR U4791 ( .A(n1708), .B(z[1]), .Z(z[7]) );
  XOR U4792 ( .A(x[83]), .B(x[81]), .Z(n1711) );
  XNOR U4793 ( .A(x[80]), .B(x[86]), .Z(n1710) );
  XOR U4794 ( .A(n1710), .B(x[82]), .Z(n1709) );
  XNOR U4795 ( .A(n1711), .B(n1709), .Z(n1746) );
  XNOR U4796 ( .A(x[85]), .B(n1710), .Z(n1819) );
  XOR U4797 ( .A(n1819), .B(x[84]), .Z(n1789) );
  IV U4798 ( .A(n1789), .Z(n1720) );
  XNOR U4799 ( .A(x[87]), .B(x[84]), .Z(n1714) );
  XNOR U4800 ( .A(n1711), .B(n1714), .Z(n1774) );
  NOR U4801 ( .A(n1720), .B(n1774), .Z(n1713) );
  XNOR U4802 ( .A(n1819), .B(x[87]), .Z(n1805) );
  XNOR U4803 ( .A(x[82]), .B(n1805), .Z(n1729) );
  XNOR U4804 ( .A(x[81]), .B(n1729), .Z(n1724) );
  AND U4805 ( .A(x[80]), .B(n1724), .Z(n1712) );
  XNOR U4806 ( .A(n1713), .B(n1712), .Z(n1717) );
  XNOR U4807 ( .A(n1746), .B(n1805), .Z(n1736) );
  IV U4808 ( .A(n1746), .Z(n1731) );
  XNOR U4809 ( .A(x[80]), .B(n1731), .Z(n1751) );
  IV U4810 ( .A(n1714), .Z(n1779) );
  AND U4811 ( .A(n1751), .B(n1779), .Z(n1719) );
  IV U4812 ( .A(n1819), .Z(n1738) );
  XNOR U4813 ( .A(n1746), .B(n1738), .Z(n1768) );
  XOR U4814 ( .A(n1768), .B(n1774), .Z(n1771) );
  XOR U4815 ( .A(x[82]), .B(x[84]), .Z(n1781) );
  NAND U4816 ( .A(n1771), .B(n1781), .Z(n1715) );
  XNOR U4817 ( .A(n1719), .B(n1715), .Z(n1740) );
  XNOR U4818 ( .A(n1736), .B(n1740), .Z(n1716) );
  XNOR U4819 ( .A(n1717), .B(n1716), .Z(n1763) );
  XOR U4820 ( .A(x[82]), .B(x[87]), .Z(n1795) );
  XNOR U4821 ( .A(x[80]), .B(n1774), .Z(n1775) );
  XNOR U4822 ( .A(n1819), .B(n1775), .Z(n1766) );
  NAND U4823 ( .A(n1795), .B(n1766), .Z(n1718) );
  XNOR U4824 ( .A(n1719), .B(n1718), .Z(n1732) );
  IV U4825 ( .A(n1724), .Z(n1778) );
  XNOR U4826 ( .A(n1778), .B(n1720), .Z(n1785) );
  AND U4827 ( .A(n1774), .B(n1785), .Z(n1722) );
  AND U4828 ( .A(x[80]), .B(n1789), .Z(n1721) );
  XNOR U4829 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U4830 ( .A(n1775), .B(n1723), .Z(n1727) );
  NAND U4831 ( .A(x[80]), .B(n1774), .Z(n1725) );
  OR U4832 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U4833 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U4834 ( .A(n1729), .B(n1728), .Z(n1730) );
  XNOR U4835 ( .A(n1732), .B(n1730), .Z(n1752) );
  IV U4836 ( .A(n1752), .Z(n1759) );
  AND U4837 ( .A(n1805), .B(n1731), .Z(n1734) );
  XOR U4838 ( .A(x[81]), .B(x[87]), .Z(n1807) );
  AND U4839 ( .A(n1768), .B(n1807), .Z(n1737) );
  XNOR U4840 ( .A(n1737), .B(n1732), .Z(n1733) );
  XNOR U4841 ( .A(n1734), .B(n1733), .Z(n1758) );
  NANDN U4842 ( .A(n1759), .B(n1758), .Z(n1735) );
  NAND U4843 ( .A(n1763), .B(n1735), .Z(n1745) );
  XNOR U4844 ( .A(n1737), .B(n1736), .Z(n1742) );
  ANDN U4845 ( .B(n1738), .A(x[81]), .Z(n1739) );
  XNOR U4846 ( .A(n1740), .B(n1739), .Z(n1741) );
  XNOR U4847 ( .A(n1742), .B(n1741), .Z(n1755) );
  XOR U4848 ( .A(n1758), .B(n1755), .Z(n1743) );
  NAND U4849 ( .A(n1759), .B(n1743), .Z(n1744) );
  NAND U4850 ( .A(n1745), .B(n1744), .Z(n1804) );
  ANDN U4851 ( .B(n1746), .A(n1804), .Z(n1770) );
  IV U4852 ( .A(n1755), .Z(n1761) );
  XOR U4853 ( .A(n1763), .B(n1759), .Z(n1747) );
  NANDN U4854 ( .A(n1761), .B(n1747), .Z(n1750) );
  NANDN U4855 ( .A(n1759), .B(n1761), .Z(n1748) );
  NANDN U4856 ( .A(n1758), .B(n1748), .Z(n1749) );
  NAND U4857 ( .A(n1750), .B(n1749), .Z(n1814) );
  XNOR U4858 ( .A(n1804), .B(n1814), .Z(n1780) );
  AND U4859 ( .A(n1751), .B(n1780), .Z(n1773) );
  OR U4860 ( .A(n1758), .B(n1755), .Z(n1757) );
  ANDN U4861 ( .B(n1758), .A(n1752), .Z(n1753) );
  XNOR U4862 ( .A(n1753), .B(n1763), .Z(n1754) );
  NAND U4863 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U4864 ( .A(n1757), .B(n1756), .Z(n1777) );
  NAND U4865 ( .A(n1759), .B(n1763), .Z(n1765) );
  NAND U4866 ( .A(n1759), .B(n1758), .Z(n1760) );
  XNOR U4867 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U4868 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1821) );
  NAND U4870 ( .A(n1796), .B(n1766), .Z(n1767) );
  XNOR U4871 ( .A(n1773), .B(n1767), .Z(n1816) );
  XOR U4872 ( .A(n1804), .B(n1821), .Z(n1806) );
  AND U4873 ( .A(n1768), .B(n1806), .Z(n1791) );
  XNOR U4874 ( .A(n1816), .B(n1791), .Z(n1769) );
  XNOR U4875 ( .A(n1770), .B(n1769), .Z(n1824) );
  NAND U4876 ( .A(n1782), .B(n1771), .Z(n1772) );
  XNOR U4877 ( .A(n1773), .B(n1772), .Z(n1799) );
  AND U4878 ( .A(n1774), .B(n1784), .Z(n1815) );
  NANDN U4879 ( .A(n1775), .B(n1777), .Z(n1776) );
  XNOR U4880 ( .A(n1815), .B(n1776), .Z(n1803) );
  XNOR U4881 ( .A(n1799), .B(n1803), .Z(n1788) );
  XOR U4882 ( .A(n1824), .B(n1788), .Z(z[80]) );
  AND U4883 ( .A(n1778), .B(n1777), .Z(n1787) );
  AND U4884 ( .A(n1780), .B(n1779), .Z(n1798) );
  NAND U4885 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U4886 ( .A(n1798), .B(n1783), .Z(n1825) );
  AND U4887 ( .A(n1785), .B(n1784), .Z(n1792) );
  XNOR U4888 ( .A(n1825), .B(n1792), .Z(n1786) );
  XNOR U4889 ( .A(n1787), .B(n1786), .Z(n1812) );
  XNOR U4890 ( .A(n1812), .B(n1788), .Z(n1830) );
  AND U4891 ( .A(n1789), .B(n1814), .Z(n1794) );
  NANDN U4892 ( .A(n1821), .B(n1819), .Z(n1790) );
  XNOR U4893 ( .A(n1791), .B(n1790), .Z(n1802) );
  XNOR U4894 ( .A(n1792), .B(n1802), .Z(n1793) );
  XNOR U4895 ( .A(n1794), .B(n1793), .Z(n1801) );
  NAND U4896 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U4897 ( .A(n1798), .B(n1797), .Z(n1808) );
  XNOR U4898 ( .A(n1799), .B(n1808), .Z(n1800) );
  XNOR U4899 ( .A(n1801), .B(n1800), .Z(n1811) );
  XNOR U4900 ( .A(n1830), .B(n1811), .Z(z[81]) );
  XNOR U4901 ( .A(n1803), .B(n1802), .Z(z[82]) );
  NOR U4902 ( .A(n1805), .B(n1804), .Z(n1810) );
  AND U4903 ( .A(n1807), .B(n1806), .Z(n1823) );
  XNOR U4904 ( .A(n1808), .B(n1823), .Z(n1809) );
  XNOR U4905 ( .A(n1810), .B(n1809), .Z(n1829) );
  XOR U4906 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U4907 ( .A(n1829), .B(n1813), .Z(z[83]) );
  XOR U4908 ( .A(n1824), .B(z[82]), .Z(z[84]) );
  AND U4909 ( .A(x[80]), .B(n1814), .Z(n1818) );
  XNOR U4910 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U4911 ( .A(n1818), .B(n1817), .Z(n1831) );
  XOR U4912 ( .A(n1819), .B(x[81]), .Z(n1820) );
  NANDN U4913 ( .A(n1821), .B(n1820), .Z(n1822) );
  XNOR U4914 ( .A(n1823), .B(n1822), .Z(n1827) );
  XNOR U4915 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U4916 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U4917 ( .A(n1831), .B(n1828), .Z(z[85]) );
  XNOR U4918 ( .A(n1830), .B(n1829), .Z(z[86]) );
  XOR U4919 ( .A(n1831), .B(z[81]), .Z(z[87]) );
  XOR U4920 ( .A(x[91]), .B(x[89]), .Z(n1834) );
  XNOR U4921 ( .A(x[88]), .B(x[94]), .Z(n1833) );
  XOR U4922 ( .A(n1833), .B(x[90]), .Z(n1832) );
  XNOR U4923 ( .A(n1834), .B(n1832), .Z(n1869) );
  XNOR U4924 ( .A(x[93]), .B(n1833), .Z(n1944) );
  XOR U4925 ( .A(n1944), .B(x[92]), .Z(n1912) );
  IV U4926 ( .A(n1912), .Z(n1843) );
  XNOR U4927 ( .A(x[95]), .B(x[92]), .Z(n1837) );
  XNOR U4928 ( .A(n1834), .B(n1837), .Z(n1897) );
  NOR U4929 ( .A(n1843), .B(n1897), .Z(n1836) );
  XNOR U4930 ( .A(n1944), .B(x[95]), .Z(n1930) );
  XNOR U4931 ( .A(x[90]), .B(n1930), .Z(n1852) );
  XNOR U4932 ( .A(x[89]), .B(n1852), .Z(n1847) );
  AND U4933 ( .A(x[88]), .B(n1847), .Z(n1835) );
  XNOR U4934 ( .A(n1836), .B(n1835), .Z(n1840) );
  XNOR U4935 ( .A(n1869), .B(n1930), .Z(n1859) );
  IV U4936 ( .A(n1869), .Z(n1854) );
  XNOR U4937 ( .A(x[88]), .B(n1854), .Z(n1874) );
  IV U4938 ( .A(n1837), .Z(n1902) );
  AND U4939 ( .A(n1874), .B(n1902), .Z(n1842) );
  IV U4940 ( .A(n1944), .Z(n1861) );
  XNOR U4941 ( .A(n1869), .B(n1861), .Z(n1891) );
  XOR U4942 ( .A(n1891), .B(n1897), .Z(n1894) );
  XOR U4943 ( .A(x[90]), .B(x[92]), .Z(n1904) );
  NAND U4944 ( .A(n1894), .B(n1904), .Z(n1838) );
  XNOR U4945 ( .A(n1842), .B(n1838), .Z(n1863) );
  XNOR U4946 ( .A(n1859), .B(n1863), .Z(n1839) );
  XNOR U4947 ( .A(n1840), .B(n1839), .Z(n1886) );
  XOR U4948 ( .A(x[90]), .B(x[95]), .Z(n1918) );
  XNOR U4949 ( .A(x[88]), .B(n1897), .Z(n1898) );
  XNOR U4950 ( .A(n1944), .B(n1898), .Z(n1889) );
  NAND U4951 ( .A(n1918), .B(n1889), .Z(n1841) );
  XNOR U4952 ( .A(n1842), .B(n1841), .Z(n1855) );
  IV U4953 ( .A(n1847), .Z(n1901) );
  XNOR U4954 ( .A(n1901), .B(n1843), .Z(n1908) );
  AND U4955 ( .A(n1897), .B(n1908), .Z(n1845) );
  AND U4956 ( .A(x[88]), .B(n1912), .Z(n1844) );
  XNOR U4957 ( .A(n1845), .B(n1844), .Z(n1846) );
  NANDN U4958 ( .A(n1898), .B(n1846), .Z(n1850) );
  NAND U4959 ( .A(x[88]), .B(n1897), .Z(n1848) );
  OR U4960 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U4961 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U4962 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U4963 ( .A(n1855), .B(n1853), .Z(n1875) );
  IV U4964 ( .A(n1875), .Z(n1882) );
  AND U4965 ( .A(n1930), .B(n1854), .Z(n1857) );
  XOR U4966 ( .A(x[89]), .B(x[95]), .Z(n1932) );
  AND U4967 ( .A(n1891), .B(n1932), .Z(n1860) );
  XNOR U4968 ( .A(n1860), .B(n1855), .Z(n1856) );
  XNOR U4969 ( .A(n1857), .B(n1856), .Z(n1881) );
  NANDN U4970 ( .A(n1882), .B(n1881), .Z(n1858) );
  NAND U4971 ( .A(n1886), .B(n1858), .Z(n1868) );
  XNOR U4972 ( .A(n1860), .B(n1859), .Z(n1865) );
  ANDN U4973 ( .B(n1861), .A(x[89]), .Z(n1862) );
  XNOR U4974 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U4975 ( .A(n1865), .B(n1864), .Z(n1878) );
  XOR U4976 ( .A(n1881), .B(n1878), .Z(n1866) );
  NAND U4977 ( .A(n1882), .B(n1866), .Z(n1867) );
  NAND U4978 ( .A(n1868), .B(n1867), .Z(n1929) );
  ANDN U4979 ( .B(n1869), .A(n1929), .Z(n1893) );
  IV U4980 ( .A(n1878), .Z(n1884) );
  XOR U4981 ( .A(n1886), .B(n1882), .Z(n1870) );
  NANDN U4982 ( .A(n1884), .B(n1870), .Z(n1873) );
  NANDN U4983 ( .A(n1882), .B(n1884), .Z(n1871) );
  NANDN U4984 ( .A(n1881), .B(n1871), .Z(n1872) );
  NAND U4985 ( .A(n1873), .B(n1872), .Z(n1939) );
  XNOR U4986 ( .A(n1929), .B(n1939), .Z(n1903) );
  AND U4987 ( .A(n1874), .B(n1903), .Z(n1896) );
  OR U4988 ( .A(n1881), .B(n1878), .Z(n1880) );
  ANDN U4989 ( .B(n1881), .A(n1875), .Z(n1876) );
  XNOR U4990 ( .A(n1876), .B(n1886), .Z(n1877) );
  NAND U4991 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U4992 ( .A(n1880), .B(n1879), .Z(n1900) );
  NAND U4993 ( .A(n1882), .B(n1886), .Z(n1888) );
  NAND U4994 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U4995 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U4996 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4997 ( .A(n1888), .B(n1887), .Z(n1946) );
  NAND U4998 ( .A(n1919), .B(n1889), .Z(n1890) );
  XNOR U4999 ( .A(n1896), .B(n1890), .Z(n1941) );
  XOR U5000 ( .A(n1929), .B(n1946), .Z(n1931) );
  AND U5001 ( .A(n1891), .B(n1931), .Z(n1914) );
  XNOR U5002 ( .A(n1941), .B(n1914), .Z(n1892) );
  XNOR U5003 ( .A(n1893), .B(n1892), .Z(n1949) );
  NAND U5004 ( .A(n1905), .B(n1894), .Z(n1895) );
  XNOR U5005 ( .A(n1896), .B(n1895), .Z(n1922) );
  AND U5006 ( .A(n1897), .B(n1907), .Z(n1940) );
  NANDN U5007 ( .A(n1898), .B(n1900), .Z(n1899) );
  XNOR U5008 ( .A(n1940), .B(n1899), .Z(n1928) );
  XNOR U5009 ( .A(n1922), .B(n1928), .Z(n1911) );
  XOR U5010 ( .A(n1949), .B(n1911), .Z(z[88]) );
  AND U5011 ( .A(n1901), .B(n1900), .Z(n1910) );
  AND U5012 ( .A(n1903), .B(n1902), .Z(n1921) );
  NAND U5013 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U5014 ( .A(n1921), .B(n1906), .Z(n1950) );
  AND U5015 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U5016 ( .A(n1950), .B(n1915), .Z(n1909) );
  XNOR U5017 ( .A(n1910), .B(n1909), .Z(n1937) );
  XNOR U5018 ( .A(n1937), .B(n1911), .Z(n1955) );
  AND U5019 ( .A(n1912), .B(n1939), .Z(n1917) );
  NANDN U5020 ( .A(n1946), .B(n1944), .Z(n1913) );
  XNOR U5021 ( .A(n1914), .B(n1913), .Z(n1927) );
  XNOR U5022 ( .A(n1915), .B(n1927), .Z(n1916) );
  XNOR U5023 ( .A(n1917), .B(n1916), .Z(n1924) );
  NAND U5024 ( .A(n1919), .B(n1918), .Z(n1920) );
  XNOR U5025 ( .A(n1921), .B(n1920), .Z(n1933) );
  XNOR U5026 ( .A(n1922), .B(n1933), .Z(n1923) );
  XNOR U5027 ( .A(n1924), .B(n1923), .Z(n1936) );
  XNOR U5028 ( .A(n1955), .B(n1936), .Z(z[89]) );
  XOR U5029 ( .A(n1926), .B(n1925), .Z(z[8]) );
  XNOR U5030 ( .A(n1928), .B(n1927), .Z(z[90]) );
  NOR U5031 ( .A(n1930), .B(n1929), .Z(n1935) );
  AND U5032 ( .A(n1932), .B(n1931), .Z(n1948) );
  XNOR U5033 ( .A(n1933), .B(n1948), .Z(n1934) );
  XNOR U5034 ( .A(n1935), .B(n1934), .Z(n1954) );
  XOR U5035 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U5036 ( .A(n1954), .B(n1938), .Z(z[91]) );
  XOR U5037 ( .A(n1949), .B(z[90]), .Z(z[92]) );
  AND U5038 ( .A(x[88]), .B(n1939), .Z(n1943) );
  XNOR U5039 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5040 ( .A(n1943), .B(n1942), .Z(n1956) );
  XOR U5041 ( .A(n1944), .B(x[89]), .Z(n1945) );
  NANDN U5042 ( .A(n1946), .B(n1945), .Z(n1947) );
  XNOR U5043 ( .A(n1948), .B(n1947), .Z(n1952) );
  XNOR U5044 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U5045 ( .A(n1952), .B(n1951), .Z(n1953) );
  XNOR U5046 ( .A(n1956), .B(n1953), .Z(z[93]) );
  XNOR U5047 ( .A(n1955), .B(n1954), .Z(z[94]) );
  XOR U5048 ( .A(n1956), .B(z[89]), .Z(z[95]) );
  XOR U5049 ( .A(n1958), .B(n1957), .Z(z[96]) );
  XOR U5050 ( .A(n1960), .B(n1959), .Z(n1961) );
  XNOR U5051 ( .A(n1962), .B(n1961), .Z(z[99]) );
endmodule


module SubBytes_2 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;

  XOR U2962 ( .A(n622), .B(n585), .Z(n592) );
  XOR U2963 ( .A(n1814), .B(n1777), .Z(n1784) );
  XOR U2964 ( .A(n1181), .B(n1144), .Z(n1151) );
  XOR U2965 ( .A(n1427), .B(n775), .Z(n782) );
  XOR U2966 ( .A(n467), .B(n430), .Z(n437) );
  XOR U2967 ( .A(n923), .B(n886), .Z(n893) );
  XOR U2968 ( .A(n1690), .B(n1653), .Z(n1660) );
  XOR U2969 ( .A(n1048), .B(n1011), .Z(n1018) );
  XOR U2970 ( .A(n290), .B(n253), .Z(n260) );
  XOR U2971 ( .A(n1565), .B(n1528), .Z(n1535) );
  XOR U2972 ( .A(n1442), .B(n1390), .Z(n1397) );
  XOR U2973 ( .A(n800), .B(n738), .Z(n745) );
  XOR U2974 ( .A(n1939), .B(n1900), .Z(n1907) );
  XOR U2975 ( .A(n1304), .B(n1267), .Z(n1274) );
  XNOR U2976 ( .A(n1777), .B(n1821), .Z(n1796) );
  XNOR U2977 ( .A(n585), .B(n629), .Z(n604) );
  XNOR U2978 ( .A(n1144), .B(n1188), .Z(n1163) );
  XNOR U2979 ( .A(n775), .B(n1434), .Z(n794) );
  XNOR U2980 ( .A(n886), .B(n930), .Z(n905) );
  XNOR U2981 ( .A(n430), .B(n474), .Z(n449) );
  XNOR U2982 ( .A(n1011), .B(n1055), .Z(n1030) );
  XNOR U2983 ( .A(n1528), .B(n1572), .Z(n1547) );
  XNOR U2984 ( .A(n1390), .B(n1449), .Z(n1409) );
  XNOR U2985 ( .A(n738), .B(n807), .Z(n757) );
  XNOR U2986 ( .A(n253), .B(n297), .Z(n272) );
  NOR U2987 ( .A(n654), .B(x[9]), .Z(n1) );
  XNOR U2988 ( .A(n329), .B(n328), .Z(n2) );
  XNOR U2989 ( .A(n1), .B(n2), .Z(n3) );
  XNOR U2990 ( .A(n312), .B(n3), .Z(n345) );
  XNOR U2991 ( .A(n1900), .B(n1946), .Z(n1919) );
  XNOR U2992 ( .A(n1267), .B(n1311), .Z(n1286) );
  XNOR U2993 ( .A(n1653), .B(n1697), .Z(n1672) );
  XOR U2994 ( .A(n163), .B(n134), .Z(n157) );
  XOR U2995 ( .A(n77), .B(n78), .Z(n129) );
  XNOR U2996 ( .A(x[9]), .B(n323), .Z(n318) );
  XOR U2997 ( .A(n794), .B(n778), .Z(n780) );
  XOR U2998 ( .A(n604), .B(n588), .Z(n590) );
  XOR U2999 ( .A(n1796), .B(n1780), .Z(n1782) );
  XOR U3000 ( .A(n1163), .B(n1147), .Z(n1149) );
  XOR U3001 ( .A(n1030), .B(n1014), .Z(n1016) );
  XOR U3002 ( .A(n1672), .B(n1656), .Z(n1658) );
  XOR U3003 ( .A(n905), .B(n889), .Z(n891) );
  XOR U3004 ( .A(n449), .B(n433), .Z(n435) );
  XOR U3005 ( .A(n757), .B(n741), .Z(n743) );
  XOR U3006 ( .A(n272), .B(n256), .Z(n258) );
  XOR U3007 ( .A(n1409), .B(n1393), .Z(n1395) );
  XOR U3008 ( .A(n1547), .B(n1531), .Z(n1533) );
  XOR U3009 ( .A(n1286), .B(n1270), .Z(n1272) );
  XOR U3010 ( .A(n1919), .B(n1903), .Z(n1905) );
  XOR U3011 ( .A(n643), .B(n508), .Z(n511) );
  NANDN U3012 ( .A(n116), .B(n121), .Z(n4) );
  XOR U3013 ( .A(n116), .B(n119), .Z(n5) );
  OR U3014 ( .A(n121), .B(n5), .Z(n6) );
  NANDN U3015 ( .A(n117), .B(n6), .Z(n7) );
  NAND U3016 ( .A(n4), .B(n7), .Z(n169) );
  XOR U3017 ( .A(x[3]), .B(x[1]), .Z(n10) );
  XNOR U3018 ( .A(x[0]), .B(x[6]), .Z(n9) );
  XOR U3019 ( .A(n9), .B(x[2]), .Z(n8) );
  XNOR U3020 ( .A(n10), .B(n8), .Z(n45) );
  XNOR U3021 ( .A(x[5]), .B(n9), .Z(n1432) );
  XOR U3022 ( .A(n1432), .B(x[4]), .Z(n787) );
  IV U3023 ( .A(n787), .Z(n19) );
  XNOR U3024 ( .A(x[7]), .B(x[4]), .Z(n13) );
  XNOR U3025 ( .A(n10), .B(n13), .Z(n73) );
  NOR U3026 ( .A(n19), .B(n73), .Z(n12) );
  XNOR U3027 ( .A(n1432), .B(x[7]), .Z(n1067) );
  XNOR U3028 ( .A(x[2]), .B(n1067), .Z(n28) );
  XNOR U3029 ( .A(x[1]), .B(n28), .Z(n23) );
  AND U3030 ( .A(x[0]), .B(n23), .Z(n11) );
  XNOR U3031 ( .A(n12), .B(n11), .Z(n16) );
  XNOR U3032 ( .A(n45), .B(n1067), .Z(n35) );
  IV U3033 ( .A(n45), .Z(n30) );
  XNOR U3034 ( .A(x[0]), .B(n30), .Z(n50) );
  IV U3035 ( .A(n13), .Z(n777) );
  AND U3036 ( .A(n50), .B(n777), .Z(n18) );
  IV U3037 ( .A(n1432), .Z(n37) );
  XNOR U3038 ( .A(n45), .B(n37), .Z(n67) );
  XOR U3039 ( .A(n67), .B(n73), .Z(n70) );
  XOR U3040 ( .A(x[2]), .B(x[4]), .Z(n779) );
  NAND U3041 ( .A(n70), .B(n779), .Z(n14) );
  XNOR U3042 ( .A(n18), .B(n14), .Z(n39) );
  XNOR U3043 ( .A(n35), .B(n39), .Z(n15) );
  XNOR U3044 ( .A(n16), .B(n15), .Z(n62) );
  XOR U3045 ( .A(x[2]), .B(x[7]), .Z(n793) );
  XNOR U3046 ( .A(x[0]), .B(n73), .Z(n74) );
  XNOR U3047 ( .A(n1432), .B(n74), .Z(n65) );
  NAND U3048 ( .A(n793), .B(n65), .Z(n17) );
  XNOR U3049 ( .A(n18), .B(n17), .Z(n31) );
  IV U3050 ( .A(n23), .Z(n776) );
  XNOR U3051 ( .A(n776), .B(n19), .Z(n783) );
  AND U3052 ( .A(n73), .B(n783), .Z(n21) );
  AND U3053 ( .A(x[0]), .B(n787), .Z(n20) );
  XNOR U3054 ( .A(n21), .B(n20), .Z(n22) );
  NANDN U3055 ( .A(n74), .B(n22), .Z(n26) );
  NAND U3056 ( .A(x[0]), .B(n73), .Z(n24) );
  OR U3057 ( .A(n24), .B(n23), .Z(n25) );
  NAND U3058 ( .A(n26), .B(n25), .Z(n27) );
  XNOR U3059 ( .A(n28), .B(n27), .Z(n29) );
  XNOR U3060 ( .A(n31), .B(n29), .Z(n51) );
  IV U3061 ( .A(n51), .Z(n58) );
  AND U3062 ( .A(n1067), .B(n30), .Z(n33) );
  XOR U3063 ( .A(x[1]), .B(x[7]), .Z(n1069) );
  AND U3064 ( .A(n67), .B(n1069), .Z(n36) );
  XNOR U3065 ( .A(n36), .B(n31), .Z(n32) );
  XNOR U3066 ( .A(n33), .B(n32), .Z(n57) );
  NANDN U3067 ( .A(n58), .B(n57), .Z(n34) );
  NAND U3068 ( .A(n62), .B(n34), .Z(n44) );
  XNOR U3069 ( .A(n36), .B(n35), .Z(n41) );
  ANDN U3070 ( .B(n37), .A(x[1]), .Z(n38) );
  XNOR U3071 ( .A(n39), .B(n38), .Z(n40) );
  XNOR U3072 ( .A(n41), .B(n40), .Z(n54) );
  XOR U3073 ( .A(n57), .B(n54), .Z(n42) );
  NAND U3074 ( .A(n58), .B(n42), .Z(n43) );
  NAND U3075 ( .A(n44), .B(n43), .Z(n1066) );
  ANDN U3076 ( .B(n45), .A(n1066), .Z(n69) );
  IV U3077 ( .A(n54), .Z(n60) );
  XOR U3078 ( .A(n62), .B(n58), .Z(n46) );
  NANDN U3079 ( .A(n60), .B(n46), .Z(n49) );
  NANDN U3080 ( .A(n58), .B(n60), .Z(n47) );
  NANDN U3081 ( .A(n57), .B(n47), .Z(n48) );
  NAND U3082 ( .A(n49), .B(n48), .Z(n1427) );
  XNOR U3083 ( .A(n1066), .B(n1427), .Z(n778) );
  AND U3084 ( .A(n50), .B(n778), .Z(n72) );
  OR U3085 ( .A(n57), .B(n54), .Z(n56) );
  ANDN U3086 ( .B(n57), .A(n51), .Z(n52) );
  XNOR U3087 ( .A(n52), .B(n62), .Z(n53) );
  NAND U3088 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3089 ( .A(n56), .B(n55), .Z(n775) );
  NAND U3090 ( .A(n58), .B(n62), .Z(n64) );
  NAND U3091 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U3092 ( .A(n60), .B(n59), .Z(n61) );
  NANDN U3093 ( .A(n62), .B(n61), .Z(n63) );
  NAND U3094 ( .A(n64), .B(n63), .Z(n1434) );
  NAND U3095 ( .A(n794), .B(n65), .Z(n66) );
  XNOR U3096 ( .A(n72), .B(n66), .Z(n1429) );
  XOR U3097 ( .A(n1066), .B(n1434), .Z(n1068) );
  AND U3098 ( .A(n67), .B(n1068), .Z(n789) );
  XNOR U3099 ( .A(n1429), .B(n789), .Z(n68) );
  XNOR U3100 ( .A(n69), .B(n68), .Z(n1437) );
  NAND U3101 ( .A(n780), .B(n70), .Z(n71) );
  XNOR U3102 ( .A(n72), .B(n71), .Z(n797) );
  AND U3103 ( .A(n73), .B(n782), .Z(n1428) );
  NANDN U3104 ( .A(n74), .B(n775), .Z(n75) );
  XNOR U3105 ( .A(n1428), .B(n75), .Z(n939) );
  XNOR U3106 ( .A(n797), .B(n939), .Z(n786) );
  XOR U3107 ( .A(n1437), .B(n786), .Z(z[0]) );
  XOR U3108 ( .A(x[99]), .B(x[97]), .Z(n76) );
  XNOR U3109 ( .A(n76), .B(x[98]), .Z(n77) );
  XNOR U3110 ( .A(x[101]), .B(n77), .Z(n114) );
  XOR U3111 ( .A(x[98]), .B(x[100]), .Z(n135) );
  XNOR U3112 ( .A(x[102]), .B(n77), .Z(n128) );
  XOR U3113 ( .A(x[103]), .B(x[100]), .Z(n133) );
  XOR U3114 ( .A(n76), .B(n133), .Z(n124) );
  XNOR U3115 ( .A(x[96]), .B(n124), .Z(n93) );
  IV U3116 ( .A(n93), .Z(n125) );
  XNOR U3117 ( .A(x[102]), .B(x[96]), .Z(n78) );
  XNOR U3118 ( .A(x[101]), .B(n78), .Z(n139) );
  XOR U3119 ( .A(n125), .B(n139), .Z(n127) );
  XOR U3120 ( .A(n128), .B(n127), .Z(n156) );
  AND U3121 ( .A(n135), .B(n156), .Z(n80) );
  AND U3122 ( .A(n128), .B(n133), .Z(n86) );
  IV U3123 ( .A(n139), .Z(n102) );
  XNOR U3124 ( .A(x[103]), .B(n102), .Z(n161) );
  XOR U3125 ( .A(n129), .B(n161), .Z(n84) );
  XNOR U3126 ( .A(n86), .B(n84), .Z(n79) );
  XNOR U3127 ( .A(n80), .B(n79), .Z(n103) );
  XOR U3128 ( .A(x[98]), .B(n161), .Z(n98) );
  XOR U3129 ( .A(x[97]), .B(n98), .Z(n150) );
  ANDN U3130 ( .B(x[96]), .A(n150), .Z(n82) );
  XNOR U3131 ( .A(x[100]), .B(n102), .Z(n170) );
  NANDN U3132 ( .A(n124), .B(n170), .Z(n81) );
  XNOR U3133 ( .A(n82), .B(n81), .Z(n83) );
  XOR U3134 ( .A(n103), .B(n83), .Z(n119) );
  XOR U3135 ( .A(x[97]), .B(x[103]), .Z(n138) );
  AND U3136 ( .A(n138), .B(n114), .Z(n104) );
  XOR U3137 ( .A(n84), .B(n104), .Z(n89) );
  XOR U3138 ( .A(x[98]), .B(x[103]), .Z(n162) );
  NAND U3139 ( .A(n162), .B(n127), .Z(n85) );
  XOR U3140 ( .A(n86), .B(n85), .Z(n99) );
  AND U3141 ( .A(n129), .B(n161), .Z(n87) );
  XOR U3142 ( .A(n99), .B(n87), .Z(n88) );
  XNOR U3143 ( .A(n89), .B(n88), .Z(n117) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n152) );
  AND U3145 ( .A(n124), .B(n152), .Z(n91) );
  AND U3146 ( .A(x[96]), .B(n170), .Z(n90) );
  XNOR U3147 ( .A(n91), .B(n90), .Z(n92) );
  NANDN U3148 ( .A(n93), .B(n92), .Z(n96) );
  NAND U3149 ( .A(n124), .B(x[96]), .Z(n94) );
  NANDN U3150 ( .A(n94), .B(n150), .Z(n95) );
  NAND U3151 ( .A(n96), .B(n95), .Z(n97) );
  XNOR U3152 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U3153 ( .A(n100), .B(n99), .Z(n116) );
  OR U3154 ( .A(n117), .B(n116), .Z(n101) );
  NANDN U3155 ( .A(n119), .B(n101), .Z(n109) );
  ANDN U3156 ( .B(n102), .A(x[97]), .Z(n106) );
  XNOR U3157 ( .A(n104), .B(n103), .Z(n105) );
  XNOR U3158 ( .A(n106), .B(n105), .Z(n121) );
  XOR U3159 ( .A(n117), .B(n121), .Z(n107) );
  NAND U3160 ( .A(n116), .B(n107), .Z(n108) );
  NAND U3161 ( .A(n109), .B(n108), .Z(n160) );
  OR U3162 ( .A(n119), .B(n116), .Z(n113) );
  ANDN U3163 ( .B(n116), .A(n117), .Z(n110) );
  XNOR U3164 ( .A(n110), .B(n121), .Z(n111) );
  NAND U3165 ( .A(n119), .B(n111), .Z(n112) );
  NAND U3166 ( .A(n113), .B(n112), .Z(n141) );
  XNOR U3167 ( .A(n160), .B(n141), .Z(n137) );
  AND U3168 ( .A(n114), .B(n137), .Z(n131) );
  NAND U3169 ( .A(n139), .B(n141), .Z(n115) );
  XNOR U3170 ( .A(n131), .B(n115), .Z(n172) );
  NANDN U3171 ( .A(n117), .B(n121), .Z(n123) );
  NANDN U3172 ( .A(n117), .B(n116), .Z(n118) );
  XOR U3173 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U3174 ( .A(n121), .B(n120), .Z(n122) );
  NAND U3175 ( .A(n123), .B(n122), .Z(n149) );
  XOR U3176 ( .A(n169), .B(n149), .Z(n151) );
  AND U3177 ( .A(n124), .B(n151), .Z(n144) );
  NANDN U3178 ( .A(n149), .B(n125), .Z(n126) );
  XNOR U3179 ( .A(n144), .B(n126), .Z(n159) );
  XNOR U3180 ( .A(n172), .B(n159), .Z(z[98]) );
  XNOR U3181 ( .A(n149), .B(n141), .Z(n163) );
  AND U3182 ( .A(n127), .B(n163), .Z(n183) );
  XOR U3183 ( .A(n169), .B(n160), .Z(n134) );
  AND U3184 ( .A(n128), .B(n134), .Z(n181) );
  NANDN U3185 ( .A(n160), .B(n129), .Z(n130) );
  XNOR U3186 ( .A(n131), .B(n130), .Z(n145) );
  XNOR U3187 ( .A(n181), .B(n145), .Z(n132) );
  XNOR U3188 ( .A(n183), .B(n132), .Z(n1958) );
  XOR U3189 ( .A(n1958), .B(z[98]), .Z(z[100]) );
  AND U3190 ( .A(n133), .B(n134), .Z(n165) );
  NAND U3191 ( .A(n157), .B(n135), .Z(n136) );
  XNOR U3192 ( .A(n165), .B(n136), .Z(n153) );
  AND U3193 ( .A(n138), .B(n137), .Z(n166) );
  XOR U3194 ( .A(x[97]), .B(n139), .Z(n140) );
  NAND U3195 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U3196 ( .A(n166), .B(n142), .Z(n147) );
  NANDN U3197 ( .A(n169), .B(x[96]), .Z(n143) );
  XNOR U3198 ( .A(n144), .B(n143), .Z(n180) );
  XNOR U3199 ( .A(n180), .B(n145), .Z(n146) );
  XNOR U3200 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U3201 ( .A(n153), .B(n148), .Z(z[101]) );
  ANDN U3202 ( .B(n150), .A(n149), .Z(n155) );
  AND U3203 ( .A(n152), .B(n151), .Z(n171) );
  XNOR U3204 ( .A(n171), .B(n153), .Z(n154) );
  XNOR U3205 ( .A(n155), .B(n154), .Z(n1959) );
  NAND U3206 ( .A(n157), .B(n156), .Z(n158) );
  XNOR U3207 ( .A(n181), .B(n158), .Z(n175) );
  XNOR U3208 ( .A(n175), .B(n159), .Z(n1957) );
  XNOR U3209 ( .A(n1959), .B(n1957), .Z(n179) );
  ANDN U3210 ( .B(n161), .A(n160), .Z(n168) );
  NAND U3211 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U3212 ( .A(n165), .B(n164), .Z(n176) );
  XNOR U3213 ( .A(n176), .B(n166), .Z(n167) );
  XNOR U3214 ( .A(n168), .B(n167), .Z(n1962) );
  XNOR U3215 ( .A(n179), .B(n1962), .Z(z[102]) );
  ANDN U3216 ( .B(n170), .A(n169), .Z(n174) );
  XNOR U3217 ( .A(n172), .B(n171), .Z(n173) );
  XNOR U3218 ( .A(n174), .B(n173), .Z(n178) );
  XNOR U3219 ( .A(n176), .B(n175), .Z(n177) );
  XNOR U3220 ( .A(n178), .B(n177), .Z(n1960) );
  XNOR U3221 ( .A(n1960), .B(n179), .Z(z[97]) );
  XNOR U3222 ( .A(n181), .B(n180), .Z(n182) );
  XNOR U3223 ( .A(n183), .B(n182), .Z(n184) );
  XOR U3224 ( .A(n184), .B(z[97]), .Z(z[103]) );
  XOR U3225 ( .A(x[107]), .B(x[105]), .Z(n187) );
  XNOR U3226 ( .A(x[104]), .B(x[110]), .Z(n186) );
  XOR U3227 ( .A(n186), .B(x[106]), .Z(n185) );
  XNOR U3228 ( .A(n187), .B(n185), .Z(n222) );
  XNOR U3229 ( .A(x[109]), .B(n186), .Z(n295) );
  XOR U3230 ( .A(n295), .B(x[108]), .Z(n265) );
  IV U3231 ( .A(n265), .Z(n196) );
  XNOR U3232 ( .A(x[111]), .B(x[108]), .Z(n190) );
  XNOR U3233 ( .A(n187), .B(n190), .Z(n250) );
  NOR U3234 ( .A(n196), .B(n250), .Z(n189) );
  XNOR U3235 ( .A(n295), .B(x[111]), .Z(n281) );
  XNOR U3236 ( .A(x[106]), .B(n281), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n205), .Z(n200) );
  AND U3238 ( .A(x[104]), .B(n200), .Z(n188) );
  XNOR U3239 ( .A(n189), .B(n188), .Z(n193) );
  XNOR U3240 ( .A(n222), .B(n281), .Z(n212) );
  IV U3241 ( .A(n222), .Z(n207) );
  XNOR U3242 ( .A(x[104]), .B(n207), .Z(n227) );
  IV U3243 ( .A(n190), .Z(n255) );
  AND U3244 ( .A(n227), .B(n255), .Z(n195) );
  IV U3245 ( .A(n295), .Z(n214) );
  XNOR U3246 ( .A(n222), .B(n214), .Z(n244) );
  XOR U3247 ( .A(n244), .B(n250), .Z(n247) );
  XOR U3248 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NAND U3249 ( .A(n247), .B(n257), .Z(n191) );
  XNOR U3250 ( .A(n195), .B(n191), .Z(n216) );
  XNOR U3251 ( .A(n212), .B(n216), .Z(n192) );
  XNOR U3252 ( .A(n193), .B(n192), .Z(n239) );
  XOR U3253 ( .A(x[106]), .B(x[111]), .Z(n271) );
  XNOR U3254 ( .A(x[104]), .B(n250), .Z(n251) );
  XNOR U3255 ( .A(n295), .B(n251), .Z(n242) );
  NAND U3256 ( .A(n271), .B(n242), .Z(n194) );
  XNOR U3257 ( .A(n195), .B(n194), .Z(n208) );
  IV U3258 ( .A(n200), .Z(n254) );
  XNOR U3259 ( .A(n254), .B(n196), .Z(n261) );
  AND U3260 ( .A(n250), .B(n261), .Z(n198) );
  AND U3261 ( .A(x[104]), .B(n265), .Z(n197) );
  XNOR U3262 ( .A(n198), .B(n197), .Z(n199) );
  NANDN U3263 ( .A(n251), .B(n199), .Z(n203) );
  NAND U3264 ( .A(x[104]), .B(n250), .Z(n201) );
  OR U3265 ( .A(n201), .B(n200), .Z(n202) );
  NAND U3266 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U3267 ( .A(n205), .B(n204), .Z(n206) );
  XNOR U3268 ( .A(n208), .B(n206), .Z(n228) );
  IV U3269 ( .A(n228), .Z(n235) );
  AND U3270 ( .A(n281), .B(n207), .Z(n210) );
  XOR U3271 ( .A(x[105]), .B(x[111]), .Z(n283) );
  AND U3272 ( .A(n244), .B(n283), .Z(n213) );
  XNOR U3273 ( .A(n213), .B(n208), .Z(n209) );
  XNOR U3274 ( .A(n210), .B(n209), .Z(n234) );
  NANDN U3275 ( .A(n235), .B(n234), .Z(n211) );
  NAND U3276 ( .A(n239), .B(n211), .Z(n221) );
  XNOR U3277 ( .A(n213), .B(n212), .Z(n218) );
  ANDN U3278 ( .B(n214), .A(x[105]), .Z(n215) );
  XNOR U3279 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3280 ( .A(n218), .B(n217), .Z(n231) );
  XOR U3281 ( .A(n234), .B(n231), .Z(n219) );
  NAND U3282 ( .A(n235), .B(n219), .Z(n220) );
  NAND U3283 ( .A(n221), .B(n220), .Z(n280) );
  ANDN U3284 ( .B(n222), .A(n280), .Z(n246) );
  IV U3285 ( .A(n231), .Z(n237) );
  XOR U3286 ( .A(n239), .B(n235), .Z(n223) );
  NANDN U3287 ( .A(n237), .B(n223), .Z(n226) );
  NANDN U3288 ( .A(n235), .B(n237), .Z(n224) );
  NANDN U3289 ( .A(n234), .B(n224), .Z(n225) );
  NAND U3290 ( .A(n226), .B(n225), .Z(n290) );
  XNOR U3291 ( .A(n280), .B(n290), .Z(n256) );
  AND U3292 ( .A(n227), .B(n256), .Z(n249) );
  OR U3293 ( .A(n234), .B(n231), .Z(n233) );
  ANDN U3294 ( .B(n234), .A(n228), .Z(n229) );
  XNOR U3295 ( .A(n229), .B(n239), .Z(n230) );
  NAND U3296 ( .A(n231), .B(n230), .Z(n232) );
  NAND U3297 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3298 ( .A(n235), .B(n239), .Z(n241) );
  NAND U3299 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U3300 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U3301 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3302 ( .A(n241), .B(n240), .Z(n297) );
  NAND U3303 ( .A(n272), .B(n242), .Z(n243) );
  XNOR U3304 ( .A(n249), .B(n243), .Z(n292) );
  XOR U3305 ( .A(n280), .B(n297), .Z(n282) );
  AND U3306 ( .A(n244), .B(n282), .Z(n267) );
  XNOR U3307 ( .A(n292), .B(n267), .Z(n245) );
  XNOR U3308 ( .A(n246), .B(n245), .Z(n300) );
  NAND U3309 ( .A(n258), .B(n247), .Z(n248) );
  XNOR U3310 ( .A(n249), .B(n248), .Z(n275) );
  AND U3311 ( .A(n250), .B(n260), .Z(n291) );
  NANDN U3312 ( .A(n251), .B(n253), .Z(n252) );
  XNOR U3313 ( .A(n291), .B(n252), .Z(n279) );
  XNOR U3314 ( .A(n275), .B(n279), .Z(n264) );
  XOR U3315 ( .A(n300), .B(n264), .Z(z[104]) );
  AND U3316 ( .A(n254), .B(n253), .Z(n263) );
  AND U3317 ( .A(n256), .B(n255), .Z(n274) );
  NAND U3318 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3319 ( .A(n274), .B(n259), .Z(n301) );
  AND U3320 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3321 ( .A(n301), .B(n268), .Z(n262) );
  XNOR U3322 ( .A(n263), .B(n262), .Z(n288) );
  XNOR U3323 ( .A(n288), .B(n264), .Z(n360) );
  AND U3324 ( .A(n265), .B(n290), .Z(n270) );
  NANDN U3325 ( .A(n297), .B(n295), .Z(n266) );
  XNOR U3326 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3327 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3328 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3329 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3330 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3331 ( .A(n275), .B(n284), .Z(n276) );
  XNOR U3332 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3333 ( .A(n360), .B(n287), .Z(z[105]) );
  XNOR U3334 ( .A(n279), .B(n278), .Z(z[106]) );
  NOR U3335 ( .A(n281), .B(n280), .Z(n286) );
  AND U3336 ( .A(n283), .B(n282), .Z(n299) );
  XNOR U3337 ( .A(n284), .B(n299), .Z(n285) );
  XNOR U3338 ( .A(n286), .B(n285), .Z(n359) );
  XOR U3339 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U3340 ( .A(n359), .B(n289), .Z(z[107]) );
  XOR U3341 ( .A(n300), .B(z[106]), .Z(z[108]) );
  AND U3342 ( .A(x[104]), .B(n290), .Z(n294) );
  XNOR U3343 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U3344 ( .A(n294), .B(n293), .Z(n361) );
  XOR U3345 ( .A(n295), .B(x[105]), .Z(n296) );
  NANDN U3346 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U3347 ( .A(n299), .B(n298), .Z(n303) );
  XNOR U3348 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U3349 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U3350 ( .A(n361), .B(n304), .Z(z[109]) );
  XOR U3351 ( .A(x[9]), .B(x[11]), .Z(n305) );
  XOR U3352 ( .A(x[15]), .B(x[12]), .Z(n486) );
  XOR U3353 ( .A(n305), .B(n486), .Z(n341) );
  XNOR U3354 ( .A(x[8]), .B(x[14]), .Z(n307) );
  XNOR U3355 ( .A(x[13]), .B(n307), .Z(n654) );
  XNOR U3356 ( .A(x[15]), .B(n654), .Z(n485) );
  XNOR U3357 ( .A(n305), .B(x[10]), .Z(n306) );
  XNOR U3358 ( .A(n307), .B(n306), .Z(n308) );
  AND U3359 ( .A(n485), .B(n308), .Z(n311) );
  IV U3360 ( .A(n308), .Z(n641) );
  XOR U3361 ( .A(n641), .B(n654), .Z(n357) );
  XOR U3362 ( .A(x[9]), .B(x[15]), .Z(n491) );
  AND U3363 ( .A(n357), .B(n491), .Z(n312) );
  XNOR U3364 ( .A(x[8]), .B(n308), .Z(n509) );
  AND U3365 ( .A(n486), .B(n509), .Z(n314) );
  XOR U3366 ( .A(x[15]), .B(x[10]), .Z(n488) );
  XNOR U3367 ( .A(n341), .B(x[8]), .Z(n342) );
  XNOR U3368 ( .A(n654), .B(n342), .Z(n642) );
  NAND U3369 ( .A(n488), .B(n642), .Z(n309) );
  XNOR U3370 ( .A(n314), .B(n309), .Z(n325) );
  XNOR U3371 ( .A(n312), .B(n325), .Z(n310) );
  XNOR U3372 ( .A(n311), .B(n310), .Z(n349) );
  XNOR U3373 ( .A(n641), .B(n485), .Z(n329) );
  XOR U3374 ( .A(x[12]), .B(x[10]), .Z(n496) );
  XOR U3375 ( .A(n341), .B(n357), .Z(n510) );
  NAND U3376 ( .A(n496), .B(n510), .Z(n313) );
  XNOR U3377 ( .A(n314), .B(n313), .Z(n328) );
  OR U3378 ( .A(n349), .B(n345), .Z(n335) );
  XNOR U3379 ( .A(x[10]), .B(n485), .Z(n323) );
  IV U3380 ( .A(n318), .Z(n495) );
  XNOR U3381 ( .A(x[12]), .B(n654), .Z(n503) );
  XNOR U3382 ( .A(n495), .B(n503), .Z(n500) );
  AND U3383 ( .A(n341), .B(n500), .Z(n316) );
  ANDN U3384 ( .B(x[8]), .A(n503), .Z(n315) );
  XNOR U3385 ( .A(n316), .B(n315), .Z(n317) );
  NANDN U3386 ( .A(n342), .B(n317), .Z(n321) );
  NAND U3387 ( .A(n341), .B(x[8]), .Z(n319) );
  OR U3388 ( .A(n319), .B(n318), .Z(n320) );
  NAND U3389 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U3390 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U3391 ( .A(n325), .B(n324), .Z(n336) );
  ANDN U3392 ( .B(n349), .A(n336), .Z(n332) );
  NOR U3393 ( .A(n503), .B(n341), .Z(n327) );
  ANDN U3394 ( .B(x[8]), .A(n495), .Z(n326) );
  XNOR U3395 ( .A(n327), .B(n326), .Z(n331) );
  XNOR U3396 ( .A(n329), .B(n328), .Z(n330) );
  XNOR U3397 ( .A(n331), .B(n330), .Z(n354) );
  XNOR U3398 ( .A(n332), .B(n354), .Z(n333) );
  NAND U3399 ( .A(n345), .B(n333), .Z(n334) );
  NAND U3400 ( .A(n335), .B(n334), .Z(n494) );
  IV U3401 ( .A(n494), .Z(n487) );
  IV U3402 ( .A(n345), .Z(n352) );
  IV U3403 ( .A(n336), .Z(n350) );
  XOR U3404 ( .A(n354), .B(n350), .Z(n337) );
  NANDN U3405 ( .A(n352), .B(n337), .Z(n340) );
  NANDN U3406 ( .A(n350), .B(n352), .Z(n338) );
  NANDN U3407 ( .A(n349), .B(n338), .Z(n339) );
  NAND U3408 ( .A(n340), .B(n339), .Z(n649) );
  XNOR U3409 ( .A(n487), .B(n649), .Z(n499) );
  AND U3410 ( .A(n341), .B(n499), .Z(n651) );
  NANDN U3411 ( .A(n342), .B(n494), .Z(n343) );
  XNOR U3412 ( .A(n651), .B(n343), .Z(n663) );
  NANDN U3413 ( .A(n350), .B(n349), .Z(n344) );
  NAND U3414 ( .A(n354), .B(n344), .Z(n348) );
  XOR U3415 ( .A(n349), .B(n345), .Z(n346) );
  NAND U3416 ( .A(n350), .B(n346), .Z(n347) );
  NAND U3417 ( .A(n348), .B(n347), .Z(n640) );
  NAND U3418 ( .A(n350), .B(n354), .Z(n356) );
  NAND U3419 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U3420 ( .A(n352), .B(n351), .Z(n353) );
  NANDN U3421 ( .A(n354), .B(n353), .Z(n355) );
  NAND U3422 ( .A(n356), .B(n355), .Z(n656) );
  XOR U3423 ( .A(n640), .B(n656), .Z(n490) );
  AND U3424 ( .A(n357), .B(n490), .Z(n646) );
  NANDN U3425 ( .A(n656), .B(n654), .Z(n358) );
  XNOR U3426 ( .A(n646), .B(n358), .Z(n513) );
  XNOR U3427 ( .A(n663), .B(n513), .Z(z[10]) );
  XNOR U3428 ( .A(n360), .B(n359), .Z(z[110]) );
  XOR U3429 ( .A(n361), .B(z[105]), .Z(z[111]) );
  XOR U3430 ( .A(x[115]), .B(x[113]), .Z(n364) );
  XNOR U3431 ( .A(x[112]), .B(x[118]), .Z(n363) );
  XOR U3432 ( .A(n363), .B(x[114]), .Z(n362) );
  XNOR U3433 ( .A(n364), .B(n362), .Z(n399) );
  XNOR U3434 ( .A(x[117]), .B(n363), .Z(n472) );
  XOR U3435 ( .A(n472), .B(x[116]), .Z(n442) );
  IV U3436 ( .A(n442), .Z(n373) );
  XNOR U3437 ( .A(x[119]), .B(x[116]), .Z(n367) );
  XNOR U3438 ( .A(n364), .B(n367), .Z(n427) );
  NOR U3439 ( .A(n373), .B(n427), .Z(n366) );
  XNOR U3440 ( .A(n472), .B(x[119]), .Z(n458) );
  XNOR U3441 ( .A(x[114]), .B(n458), .Z(n382) );
  XNOR U3442 ( .A(x[113]), .B(n382), .Z(n377) );
  AND U3443 ( .A(x[112]), .B(n377), .Z(n365) );
  XNOR U3444 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U3445 ( .A(n399), .B(n458), .Z(n389) );
  IV U3446 ( .A(n399), .Z(n384) );
  XNOR U3447 ( .A(x[112]), .B(n384), .Z(n404) );
  IV U3448 ( .A(n367), .Z(n432) );
  AND U3449 ( .A(n404), .B(n432), .Z(n372) );
  IV U3450 ( .A(n472), .Z(n391) );
  XNOR U3451 ( .A(n399), .B(n391), .Z(n421) );
  XOR U3452 ( .A(n421), .B(n427), .Z(n424) );
  XOR U3453 ( .A(x[114]), .B(x[116]), .Z(n434) );
  NAND U3454 ( .A(n424), .B(n434), .Z(n368) );
  XNOR U3455 ( .A(n372), .B(n368), .Z(n393) );
  XNOR U3456 ( .A(n389), .B(n393), .Z(n369) );
  XNOR U3457 ( .A(n370), .B(n369), .Z(n416) );
  XOR U3458 ( .A(x[114]), .B(x[119]), .Z(n448) );
  XNOR U3459 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3460 ( .A(n472), .B(n428), .Z(n419) );
  NAND U3461 ( .A(n448), .B(n419), .Z(n371) );
  XNOR U3462 ( .A(n372), .B(n371), .Z(n385) );
  IV U3463 ( .A(n377), .Z(n431) );
  XNOR U3464 ( .A(n431), .B(n373), .Z(n438) );
  AND U3465 ( .A(n427), .B(n438), .Z(n375) );
  AND U3466 ( .A(x[112]), .B(n442), .Z(n374) );
  XNOR U3467 ( .A(n375), .B(n374), .Z(n376) );
  NANDN U3468 ( .A(n428), .B(n376), .Z(n380) );
  NAND U3469 ( .A(x[112]), .B(n427), .Z(n378) );
  OR U3470 ( .A(n378), .B(n377), .Z(n379) );
  NAND U3471 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U3472 ( .A(n382), .B(n381), .Z(n383) );
  XNOR U3473 ( .A(n385), .B(n383), .Z(n405) );
  IV U3474 ( .A(n405), .Z(n412) );
  AND U3475 ( .A(n458), .B(n384), .Z(n387) );
  XOR U3476 ( .A(x[113]), .B(x[119]), .Z(n460) );
  AND U3477 ( .A(n421), .B(n460), .Z(n390) );
  XNOR U3478 ( .A(n390), .B(n385), .Z(n386) );
  XNOR U3479 ( .A(n387), .B(n386), .Z(n411) );
  NANDN U3480 ( .A(n412), .B(n411), .Z(n388) );
  NAND U3481 ( .A(n416), .B(n388), .Z(n398) );
  XNOR U3482 ( .A(n390), .B(n389), .Z(n395) );
  ANDN U3483 ( .B(n391), .A(x[113]), .Z(n392) );
  XNOR U3484 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U3485 ( .A(n395), .B(n394), .Z(n408) );
  XOR U3486 ( .A(n411), .B(n408), .Z(n396) );
  NAND U3487 ( .A(n412), .B(n396), .Z(n397) );
  NAND U3488 ( .A(n398), .B(n397), .Z(n457) );
  ANDN U3489 ( .B(n399), .A(n457), .Z(n423) );
  IV U3490 ( .A(n408), .Z(n414) );
  XOR U3491 ( .A(n416), .B(n412), .Z(n400) );
  NANDN U3492 ( .A(n414), .B(n400), .Z(n403) );
  NANDN U3493 ( .A(n412), .B(n414), .Z(n401) );
  NANDN U3494 ( .A(n411), .B(n401), .Z(n402) );
  NAND U3495 ( .A(n403), .B(n402), .Z(n467) );
  XNOR U3496 ( .A(n457), .B(n467), .Z(n433) );
  AND U3497 ( .A(n404), .B(n433), .Z(n426) );
  OR U3498 ( .A(n411), .B(n408), .Z(n410) );
  ANDN U3499 ( .B(n411), .A(n405), .Z(n406) );
  XNOR U3500 ( .A(n406), .B(n416), .Z(n407) );
  NAND U3501 ( .A(n408), .B(n407), .Z(n409) );
  NAND U3502 ( .A(n410), .B(n409), .Z(n430) );
  NAND U3503 ( .A(n412), .B(n416), .Z(n418) );
  NAND U3504 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U3505 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U3506 ( .A(n416), .B(n415), .Z(n417) );
  NAND U3507 ( .A(n418), .B(n417), .Z(n474) );
  NAND U3508 ( .A(n449), .B(n419), .Z(n420) );
  XNOR U3509 ( .A(n426), .B(n420), .Z(n469) );
  XOR U3510 ( .A(n457), .B(n474), .Z(n459) );
  AND U3511 ( .A(n421), .B(n459), .Z(n444) );
  XNOR U3512 ( .A(n469), .B(n444), .Z(n422) );
  XNOR U3513 ( .A(n423), .B(n422), .Z(n477) );
  NAND U3514 ( .A(n435), .B(n424), .Z(n425) );
  XNOR U3515 ( .A(n426), .B(n425), .Z(n452) );
  AND U3516 ( .A(n427), .B(n437), .Z(n468) );
  NANDN U3517 ( .A(n428), .B(n430), .Z(n429) );
  XNOR U3518 ( .A(n468), .B(n429), .Z(n456) );
  XNOR U3519 ( .A(n452), .B(n456), .Z(n441) );
  XOR U3520 ( .A(n477), .B(n441), .Z(z[112]) );
  AND U3521 ( .A(n431), .B(n430), .Z(n440) );
  AND U3522 ( .A(n433), .B(n432), .Z(n451) );
  NAND U3523 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U3524 ( .A(n451), .B(n436), .Z(n478) );
  AND U3525 ( .A(n438), .B(n437), .Z(n445) );
  XNOR U3526 ( .A(n478), .B(n445), .Z(n439) );
  XNOR U3527 ( .A(n440), .B(n439), .Z(n465) );
  XNOR U3528 ( .A(n465), .B(n441), .Z(n483) );
  AND U3529 ( .A(n442), .B(n467), .Z(n447) );
  NANDN U3530 ( .A(n474), .B(n472), .Z(n443) );
  XNOR U3531 ( .A(n444), .B(n443), .Z(n455) );
  XNOR U3532 ( .A(n445), .B(n455), .Z(n446) );
  XNOR U3533 ( .A(n447), .B(n446), .Z(n454) );
  NAND U3534 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U3535 ( .A(n451), .B(n450), .Z(n461) );
  XNOR U3536 ( .A(n452), .B(n461), .Z(n453) );
  XNOR U3537 ( .A(n454), .B(n453), .Z(n464) );
  XNOR U3538 ( .A(n483), .B(n464), .Z(z[113]) );
  XNOR U3539 ( .A(n456), .B(n455), .Z(z[114]) );
  NOR U3540 ( .A(n458), .B(n457), .Z(n463) );
  AND U3541 ( .A(n460), .B(n459), .Z(n476) );
  XNOR U3542 ( .A(n461), .B(n476), .Z(n462) );
  XNOR U3543 ( .A(n463), .B(n462), .Z(n482) );
  XOR U3544 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U3545 ( .A(n482), .B(n466), .Z(z[115]) );
  XOR U3546 ( .A(n477), .B(z[114]), .Z(z[116]) );
  AND U3547 ( .A(x[112]), .B(n467), .Z(n471) );
  XNOR U3548 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U3549 ( .A(n471), .B(n470), .Z(n484) );
  XOR U3550 ( .A(n472), .B(x[113]), .Z(n473) );
  NANDN U3551 ( .A(n474), .B(n473), .Z(n475) );
  XNOR U3552 ( .A(n476), .B(n475), .Z(n480) );
  XNOR U3553 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U3554 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U3555 ( .A(n484), .B(n481), .Z(z[117]) );
  XNOR U3556 ( .A(n483), .B(n482), .Z(z[118]) );
  XOR U3557 ( .A(n484), .B(z[113]), .Z(z[119]) );
  NOR U3558 ( .A(n485), .B(n640), .Z(n493) );
  XNOR U3559 ( .A(n640), .B(n649), .Z(n508) );
  AND U3560 ( .A(n486), .B(n508), .Z(n498) );
  XOR U3561 ( .A(n487), .B(n656), .Z(n643) );
  NAND U3562 ( .A(n643), .B(n488), .Z(n489) );
  XNOR U3563 ( .A(n498), .B(n489), .Z(n504) );
  AND U3564 ( .A(n491), .B(n490), .Z(n658) );
  XNOR U3565 ( .A(n504), .B(n658), .Z(n492) );
  XNOR U3566 ( .A(n493), .B(n492), .Z(n666) );
  AND U3567 ( .A(n495), .B(n494), .Z(n502) );
  NAND U3568 ( .A(n511), .B(n496), .Z(n497) );
  XNOR U3569 ( .A(n498), .B(n497), .Z(n659) );
  AND U3570 ( .A(n500), .B(n499), .Z(n505) );
  XNOR U3571 ( .A(n659), .B(n505), .Z(n501) );
  XNOR U3572 ( .A(n502), .B(n501), .Z(n665) );
  ANDN U3573 ( .B(n649), .A(n503), .Z(n507) );
  XNOR U3574 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U3575 ( .A(n507), .B(n506), .Z(n515) );
  AND U3576 ( .A(n509), .B(n508), .Z(n645) );
  NAND U3577 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U3578 ( .A(n645), .B(n512), .Z(n664) );
  XNOR U3579 ( .A(n664), .B(n513), .Z(n514) );
  XNOR U3580 ( .A(n515), .B(n514), .Z(n667) );
  XOR U3581 ( .A(n665), .B(n667), .Z(n516) );
  XNOR U3582 ( .A(n666), .B(n516), .Z(z[11]) );
  XOR U3583 ( .A(x[123]), .B(x[121]), .Z(n519) );
  XNOR U3584 ( .A(x[120]), .B(x[126]), .Z(n518) );
  XOR U3585 ( .A(n518), .B(x[122]), .Z(n517) );
  XNOR U3586 ( .A(n519), .B(n517), .Z(n554) );
  XNOR U3587 ( .A(x[125]), .B(n518), .Z(n627) );
  XOR U3588 ( .A(n627), .B(x[124]), .Z(n597) );
  IV U3589 ( .A(n597), .Z(n528) );
  XNOR U3590 ( .A(x[127]), .B(x[124]), .Z(n522) );
  XNOR U3591 ( .A(n519), .B(n522), .Z(n582) );
  NOR U3592 ( .A(n528), .B(n582), .Z(n521) );
  XNOR U3593 ( .A(n627), .B(x[127]), .Z(n613) );
  XNOR U3594 ( .A(x[122]), .B(n613), .Z(n537) );
  XNOR U3595 ( .A(x[121]), .B(n537), .Z(n532) );
  AND U3596 ( .A(x[120]), .B(n532), .Z(n520) );
  XNOR U3597 ( .A(n521), .B(n520), .Z(n525) );
  XNOR U3598 ( .A(n554), .B(n613), .Z(n544) );
  IV U3599 ( .A(n554), .Z(n539) );
  XNOR U3600 ( .A(x[120]), .B(n539), .Z(n559) );
  IV U3601 ( .A(n522), .Z(n587) );
  AND U3602 ( .A(n559), .B(n587), .Z(n527) );
  IV U3603 ( .A(n627), .Z(n546) );
  XNOR U3604 ( .A(n554), .B(n546), .Z(n576) );
  XOR U3605 ( .A(n576), .B(n582), .Z(n579) );
  XOR U3606 ( .A(x[122]), .B(x[124]), .Z(n589) );
  NAND U3607 ( .A(n579), .B(n589), .Z(n523) );
  XNOR U3608 ( .A(n527), .B(n523), .Z(n548) );
  XNOR U3609 ( .A(n544), .B(n548), .Z(n524) );
  XNOR U3610 ( .A(n525), .B(n524), .Z(n571) );
  XOR U3611 ( .A(x[122]), .B(x[127]), .Z(n603) );
  XNOR U3612 ( .A(x[120]), .B(n582), .Z(n583) );
  XNOR U3613 ( .A(n627), .B(n583), .Z(n574) );
  NAND U3614 ( .A(n603), .B(n574), .Z(n526) );
  XNOR U3615 ( .A(n527), .B(n526), .Z(n540) );
  IV U3616 ( .A(n532), .Z(n586) );
  XNOR U3617 ( .A(n586), .B(n528), .Z(n593) );
  AND U3618 ( .A(n582), .B(n593), .Z(n530) );
  AND U3619 ( .A(x[120]), .B(n597), .Z(n529) );
  XNOR U3620 ( .A(n530), .B(n529), .Z(n531) );
  NANDN U3621 ( .A(n583), .B(n531), .Z(n535) );
  NAND U3622 ( .A(x[120]), .B(n582), .Z(n533) );
  OR U3623 ( .A(n533), .B(n532), .Z(n534) );
  NAND U3624 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U3625 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U3626 ( .A(n540), .B(n538), .Z(n560) );
  IV U3627 ( .A(n560), .Z(n567) );
  AND U3628 ( .A(n613), .B(n539), .Z(n542) );
  XOR U3629 ( .A(x[121]), .B(x[127]), .Z(n615) );
  AND U3630 ( .A(n576), .B(n615), .Z(n545) );
  XNOR U3631 ( .A(n545), .B(n540), .Z(n541) );
  XNOR U3632 ( .A(n542), .B(n541), .Z(n566) );
  NANDN U3633 ( .A(n567), .B(n566), .Z(n543) );
  NAND U3634 ( .A(n571), .B(n543), .Z(n553) );
  XNOR U3635 ( .A(n545), .B(n544), .Z(n550) );
  ANDN U3636 ( .B(n546), .A(x[121]), .Z(n547) );
  XNOR U3637 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U3638 ( .A(n550), .B(n549), .Z(n563) );
  XOR U3639 ( .A(n566), .B(n563), .Z(n551) );
  NAND U3640 ( .A(n567), .B(n551), .Z(n552) );
  NAND U3641 ( .A(n553), .B(n552), .Z(n612) );
  ANDN U3642 ( .B(n554), .A(n612), .Z(n578) );
  IV U3643 ( .A(n563), .Z(n569) );
  XOR U3644 ( .A(n571), .B(n567), .Z(n555) );
  NANDN U3645 ( .A(n569), .B(n555), .Z(n558) );
  NANDN U3646 ( .A(n567), .B(n569), .Z(n556) );
  NANDN U3647 ( .A(n566), .B(n556), .Z(n557) );
  NAND U3648 ( .A(n558), .B(n557), .Z(n622) );
  XNOR U3649 ( .A(n612), .B(n622), .Z(n588) );
  AND U3650 ( .A(n559), .B(n588), .Z(n581) );
  OR U3651 ( .A(n566), .B(n563), .Z(n565) );
  ANDN U3652 ( .B(n566), .A(n560), .Z(n561) );
  XNOR U3653 ( .A(n561), .B(n571), .Z(n562) );
  NAND U3654 ( .A(n563), .B(n562), .Z(n564) );
  NAND U3655 ( .A(n565), .B(n564), .Z(n585) );
  NAND U3656 ( .A(n567), .B(n571), .Z(n573) );
  NAND U3657 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U3658 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U3659 ( .A(n571), .B(n570), .Z(n572) );
  NAND U3660 ( .A(n573), .B(n572), .Z(n629) );
  NAND U3661 ( .A(n604), .B(n574), .Z(n575) );
  XNOR U3662 ( .A(n581), .B(n575), .Z(n624) );
  XOR U3663 ( .A(n612), .B(n629), .Z(n614) );
  AND U3664 ( .A(n576), .B(n614), .Z(n599) );
  XNOR U3665 ( .A(n624), .B(n599), .Z(n577) );
  XNOR U3666 ( .A(n578), .B(n577), .Z(n632) );
  NAND U3667 ( .A(n590), .B(n579), .Z(n580) );
  XNOR U3668 ( .A(n581), .B(n580), .Z(n607) );
  AND U3669 ( .A(n582), .B(n592), .Z(n623) );
  NANDN U3670 ( .A(n583), .B(n585), .Z(n584) );
  XNOR U3671 ( .A(n623), .B(n584), .Z(n611) );
  XNOR U3672 ( .A(n607), .B(n611), .Z(n596) );
  XOR U3673 ( .A(n632), .B(n596), .Z(z[120]) );
  AND U3674 ( .A(n586), .B(n585), .Z(n595) );
  AND U3675 ( .A(n588), .B(n587), .Z(n606) );
  NAND U3676 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U3677 ( .A(n606), .B(n591), .Z(n633) );
  AND U3678 ( .A(n593), .B(n592), .Z(n600) );
  XNOR U3679 ( .A(n633), .B(n600), .Z(n594) );
  XNOR U3680 ( .A(n595), .B(n594), .Z(n620) );
  XNOR U3681 ( .A(n620), .B(n596), .Z(n638) );
  AND U3682 ( .A(n597), .B(n622), .Z(n602) );
  NANDN U3683 ( .A(n629), .B(n627), .Z(n598) );
  XNOR U3684 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U3685 ( .A(n600), .B(n610), .Z(n601) );
  XNOR U3686 ( .A(n602), .B(n601), .Z(n609) );
  NAND U3687 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U3688 ( .A(n606), .B(n605), .Z(n616) );
  XNOR U3689 ( .A(n607), .B(n616), .Z(n608) );
  XNOR U3690 ( .A(n609), .B(n608), .Z(n619) );
  XNOR U3691 ( .A(n638), .B(n619), .Z(z[121]) );
  XNOR U3692 ( .A(n611), .B(n610), .Z(z[122]) );
  NOR U3693 ( .A(n613), .B(n612), .Z(n618) );
  AND U3694 ( .A(n615), .B(n614), .Z(n631) );
  XNOR U3695 ( .A(n616), .B(n631), .Z(n617) );
  XNOR U3696 ( .A(n618), .B(n617), .Z(n637) );
  XOR U3697 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U3698 ( .A(n637), .B(n621), .Z(z[123]) );
  XOR U3699 ( .A(n632), .B(z[122]), .Z(z[124]) );
  AND U3700 ( .A(x[120]), .B(n622), .Z(n626) );
  XNOR U3701 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U3702 ( .A(n626), .B(n625), .Z(n639) );
  XOR U3703 ( .A(n627), .B(x[121]), .Z(n628) );
  NANDN U3704 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U3705 ( .A(n631), .B(n630), .Z(n635) );
  XNOR U3706 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U3707 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U3708 ( .A(n639), .B(n636), .Z(z[125]) );
  XNOR U3709 ( .A(n638), .B(n637), .Z(z[126]) );
  XOR U3710 ( .A(n639), .B(z[121]), .Z(z[127]) );
  ANDN U3711 ( .B(n641), .A(n640), .Z(n648) );
  NAND U3712 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U3713 ( .A(n645), .B(n644), .Z(n650) );
  XNOR U3714 ( .A(n650), .B(n646), .Z(n647) );
  XNOR U3715 ( .A(n648), .B(n647), .Z(n1926) );
  XOR U3716 ( .A(n1926), .B(z[10]), .Z(z[12]) );
  AND U3717 ( .A(x[8]), .B(n649), .Z(n653) );
  XNOR U3718 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U3719 ( .A(n653), .B(n652), .Z(n669) );
  XOR U3720 ( .A(n654), .B(x[9]), .Z(n655) );
  NANDN U3721 ( .A(n656), .B(n655), .Z(n657) );
  XNOR U3722 ( .A(n658), .B(n657), .Z(n661) );
  XNOR U3723 ( .A(n659), .B(n1926), .Z(n660) );
  XNOR U3724 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U3725 ( .A(n669), .B(n662), .Z(z[13]) );
  XNOR U3726 ( .A(n664), .B(n663), .Z(n1925) );
  XNOR U3727 ( .A(n665), .B(n1925), .Z(n668) );
  XNOR U3728 ( .A(n668), .B(n666), .Z(z[14]) );
  XNOR U3729 ( .A(n668), .B(n667), .Z(z[9]) );
  XOR U3730 ( .A(n669), .B(z[9]), .Z(z[15]) );
  XOR U3731 ( .A(x[19]), .B(x[17]), .Z(n672) );
  XNOR U3732 ( .A(x[16]), .B(x[22]), .Z(n671) );
  XOR U3733 ( .A(n671), .B(x[18]), .Z(n670) );
  XNOR U3734 ( .A(n672), .B(n670), .Z(n707) );
  XNOR U3735 ( .A(x[21]), .B(n671), .Z(n805) );
  XOR U3736 ( .A(n805), .B(x[20]), .Z(n750) );
  IV U3737 ( .A(n750), .Z(n681) );
  XNOR U3738 ( .A(x[23]), .B(x[20]), .Z(n675) );
  XNOR U3739 ( .A(n672), .B(n675), .Z(n735) );
  NOR U3740 ( .A(n681), .B(n735), .Z(n674) );
  XNOR U3741 ( .A(n805), .B(x[23]), .Z(n766) );
  XNOR U3742 ( .A(x[18]), .B(n766), .Z(n690) );
  XNOR U3743 ( .A(x[17]), .B(n690), .Z(n685) );
  AND U3744 ( .A(x[16]), .B(n685), .Z(n673) );
  XNOR U3745 ( .A(n674), .B(n673), .Z(n678) );
  XNOR U3746 ( .A(n707), .B(n766), .Z(n697) );
  IV U3747 ( .A(n707), .Z(n692) );
  XNOR U3748 ( .A(x[16]), .B(n692), .Z(n712) );
  IV U3749 ( .A(n675), .Z(n740) );
  AND U3750 ( .A(n712), .B(n740), .Z(n680) );
  IV U3751 ( .A(n805), .Z(n699) );
  XNOR U3752 ( .A(n707), .B(n699), .Z(n729) );
  XOR U3753 ( .A(n729), .B(n735), .Z(n732) );
  XOR U3754 ( .A(x[18]), .B(x[20]), .Z(n742) );
  NAND U3755 ( .A(n732), .B(n742), .Z(n676) );
  XNOR U3756 ( .A(n680), .B(n676), .Z(n701) );
  XNOR U3757 ( .A(n697), .B(n701), .Z(n677) );
  XNOR U3758 ( .A(n678), .B(n677), .Z(n724) );
  XOR U3759 ( .A(x[18]), .B(x[23]), .Z(n756) );
  XNOR U3760 ( .A(x[16]), .B(n735), .Z(n736) );
  XNOR U3761 ( .A(n805), .B(n736), .Z(n727) );
  NAND U3762 ( .A(n756), .B(n727), .Z(n679) );
  XNOR U3763 ( .A(n680), .B(n679), .Z(n693) );
  IV U3764 ( .A(n685), .Z(n739) );
  XNOR U3765 ( .A(n739), .B(n681), .Z(n746) );
  AND U3766 ( .A(n735), .B(n746), .Z(n683) );
  AND U3767 ( .A(x[16]), .B(n750), .Z(n682) );
  XNOR U3768 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U3769 ( .A(n736), .B(n684), .Z(n688) );
  NAND U3770 ( .A(x[16]), .B(n735), .Z(n686) );
  OR U3771 ( .A(n686), .B(n685), .Z(n687) );
  NAND U3772 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U3773 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U3774 ( .A(n693), .B(n691), .Z(n713) );
  IV U3775 ( .A(n713), .Z(n720) );
  AND U3776 ( .A(n766), .B(n692), .Z(n695) );
  XOR U3777 ( .A(x[17]), .B(x[23]), .Z(n768) );
  AND U3778 ( .A(n729), .B(n768), .Z(n698) );
  XNOR U3779 ( .A(n698), .B(n693), .Z(n694) );
  XNOR U3780 ( .A(n695), .B(n694), .Z(n719) );
  NANDN U3781 ( .A(n720), .B(n719), .Z(n696) );
  NAND U3782 ( .A(n724), .B(n696), .Z(n706) );
  XNOR U3783 ( .A(n698), .B(n697), .Z(n703) );
  ANDN U3784 ( .B(n699), .A(x[17]), .Z(n700) );
  XNOR U3785 ( .A(n701), .B(n700), .Z(n702) );
  XNOR U3786 ( .A(n703), .B(n702), .Z(n716) );
  XOR U3787 ( .A(n719), .B(n716), .Z(n704) );
  NAND U3788 ( .A(n720), .B(n704), .Z(n705) );
  NAND U3789 ( .A(n706), .B(n705), .Z(n765) );
  ANDN U3790 ( .B(n707), .A(n765), .Z(n731) );
  IV U3791 ( .A(n716), .Z(n722) );
  XOR U3792 ( .A(n724), .B(n720), .Z(n708) );
  NANDN U3793 ( .A(n722), .B(n708), .Z(n711) );
  NANDN U3794 ( .A(n720), .B(n722), .Z(n709) );
  NANDN U3795 ( .A(n719), .B(n709), .Z(n710) );
  NAND U3796 ( .A(n711), .B(n710), .Z(n800) );
  XNOR U3797 ( .A(n765), .B(n800), .Z(n741) );
  AND U3798 ( .A(n712), .B(n741), .Z(n734) );
  OR U3799 ( .A(n719), .B(n716), .Z(n718) );
  ANDN U3800 ( .B(n719), .A(n713), .Z(n714) );
  XNOR U3801 ( .A(n714), .B(n724), .Z(n715) );
  NAND U3802 ( .A(n716), .B(n715), .Z(n717) );
  NAND U3803 ( .A(n718), .B(n717), .Z(n738) );
  NAND U3804 ( .A(n720), .B(n724), .Z(n726) );
  NAND U3805 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U3806 ( .A(n722), .B(n721), .Z(n723) );
  NANDN U3807 ( .A(n724), .B(n723), .Z(n725) );
  NAND U3808 ( .A(n726), .B(n725), .Z(n807) );
  NAND U3809 ( .A(n757), .B(n727), .Z(n728) );
  XNOR U3810 ( .A(n734), .B(n728), .Z(n802) );
  XOR U3811 ( .A(n765), .B(n807), .Z(n767) );
  AND U3812 ( .A(n729), .B(n767), .Z(n752) );
  XNOR U3813 ( .A(n802), .B(n752), .Z(n730) );
  XNOR U3814 ( .A(n731), .B(n730), .Z(n810) );
  NAND U3815 ( .A(n743), .B(n732), .Z(n733) );
  XNOR U3816 ( .A(n734), .B(n733), .Z(n760) );
  AND U3817 ( .A(n735), .B(n745), .Z(n801) );
  NANDN U3818 ( .A(n736), .B(n738), .Z(n737) );
  XNOR U3819 ( .A(n801), .B(n737), .Z(n764) );
  XNOR U3820 ( .A(n760), .B(n764), .Z(n749) );
  XOR U3821 ( .A(n810), .B(n749), .Z(z[16]) );
  AND U3822 ( .A(n739), .B(n738), .Z(n748) );
  AND U3823 ( .A(n741), .B(n740), .Z(n759) );
  NAND U3824 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U3825 ( .A(n759), .B(n744), .Z(n811) );
  AND U3826 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U3827 ( .A(n811), .B(n753), .Z(n747) );
  XNOR U3828 ( .A(n748), .B(n747), .Z(n773) );
  XNOR U3829 ( .A(n773), .B(n749), .Z(n816) );
  AND U3830 ( .A(n750), .B(n800), .Z(n755) );
  NANDN U3831 ( .A(n807), .B(n805), .Z(n751) );
  XNOR U3832 ( .A(n752), .B(n751), .Z(n763) );
  XNOR U3833 ( .A(n753), .B(n763), .Z(n754) );
  XNOR U3834 ( .A(n755), .B(n754), .Z(n762) );
  NAND U3835 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U3836 ( .A(n759), .B(n758), .Z(n769) );
  XNOR U3837 ( .A(n760), .B(n769), .Z(n761) );
  XNOR U3838 ( .A(n762), .B(n761), .Z(n772) );
  XNOR U3839 ( .A(n816), .B(n772), .Z(z[17]) );
  XNOR U3840 ( .A(n764), .B(n763), .Z(z[18]) );
  NOR U3841 ( .A(n766), .B(n765), .Z(n771) );
  AND U3842 ( .A(n768), .B(n767), .Z(n809) );
  XNOR U3843 ( .A(n769), .B(n809), .Z(n770) );
  XNOR U3844 ( .A(n771), .B(n770), .Z(n815) );
  XOR U3845 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U3846 ( .A(n815), .B(n774), .Z(z[19]) );
  AND U3847 ( .A(n776), .B(n775), .Z(n785) );
  AND U3848 ( .A(n778), .B(n777), .Z(n796) );
  NAND U3849 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U3850 ( .A(n796), .B(n781), .Z(n1438) );
  AND U3851 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U3852 ( .A(n1438), .B(n790), .Z(n784) );
  XNOR U3853 ( .A(n785), .B(n784), .Z(n1074) );
  XNOR U3854 ( .A(n1074), .B(n786), .Z(n1581) );
  AND U3855 ( .A(n787), .B(n1427), .Z(n792) );
  NANDN U3856 ( .A(n1434), .B(n1432), .Z(n788) );
  XNOR U3857 ( .A(n789), .B(n788), .Z(n938) );
  XNOR U3858 ( .A(n790), .B(n938), .Z(n791) );
  XNOR U3859 ( .A(n792), .B(n791), .Z(n799) );
  NAND U3860 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U3861 ( .A(n796), .B(n795), .Z(n1070) );
  XNOR U3862 ( .A(n797), .B(n1070), .Z(n798) );
  XNOR U3863 ( .A(n799), .B(n798), .Z(n1073) );
  XNOR U3864 ( .A(n1581), .B(n1073), .Z(z[1]) );
  XOR U3865 ( .A(n810), .B(z[18]), .Z(z[20]) );
  AND U3866 ( .A(x[16]), .B(n800), .Z(n804) );
  XNOR U3867 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U3868 ( .A(n804), .B(n803), .Z(n817) );
  XOR U3869 ( .A(n805), .B(x[17]), .Z(n806) );
  NANDN U3870 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3871 ( .A(n809), .B(n808), .Z(n813) );
  XNOR U3872 ( .A(n811), .B(n810), .Z(n812) );
  XNOR U3873 ( .A(n813), .B(n812), .Z(n814) );
  XNOR U3874 ( .A(n817), .B(n814), .Z(z[21]) );
  XNOR U3875 ( .A(n816), .B(n815), .Z(z[22]) );
  XOR U3876 ( .A(n817), .B(z[17]), .Z(z[23]) );
  XOR U3877 ( .A(x[27]), .B(x[25]), .Z(n820) );
  XNOR U3878 ( .A(x[24]), .B(x[30]), .Z(n819) );
  XOR U3879 ( .A(n819), .B(x[26]), .Z(n818) );
  XNOR U3880 ( .A(n820), .B(n818), .Z(n855) );
  XNOR U3881 ( .A(x[29]), .B(n819), .Z(n928) );
  XOR U3882 ( .A(n928), .B(x[28]), .Z(n898) );
  IV U3883 ( .A(n898), .Z(n829) );
  XNOR U3884 ( .A(x[31]), .B(x[28]), .Z(n823) );
  XNOR U3885 ( .A(n820), .B(n823), .Z(n883) );
  NOR U3886 ( .A(n829), .B(n883), .Z(n822) );
  XNOR U3887 ( .A(n928), .B(x[31]), .Z(n914) );
  XNOR U3888 ( .A(x[26]), .B(n914), .Z(n838) );
  XNOR U3889 ( .A(x[25]), .B(n838), .Z(n833) );
  AND U3890 ( .A(x[24]), .B(n833), .Z(n821) );
  XNOR U3891 ( .A(n822), .B(n821), .Z(n826) );
  XNOR U3892 ( .A(n855), .B(n914), .Z(n845) );
  IV U3893 ( .A(n855), .Z(n840) );
  XNOR U3894 ( .A(x[24]), .B(n840), .Z(n860) );
  IV U3895 ( .A(n823), .Z(n888) );
  AND U3896 ( .A(n860), .B(n888), .Z(n828) );
  IV U3897 ( .A(n928), .Z(n847) );
  XNOR U3898 ( .A(n855), .B(n847), .Z(n877) );
  XOR U3899 ( .A(n877), .B(n883), .Z(n880) );
  XOR U3900 ( .A(x[26]), .B(x[28]), .Z(n890) );
  NAND U3901 ( .A(n880), .B(n890), .Z(n824) );
  XNOR U3902 ( .A(n828), .B(n824), .Z(n849) );
  XNOR U3903 ( .A(n845), .B(n849), .Z(n825) );
  XNOR U3904 ( .A(n826), .B(n825), .Z(n872) );
  XOR U3905 ( .A(x[26]), .B(x[31]), .Z(n904) );
  XNOR U3906 ( .A(x[24]), .B(n883), .Z(n884) );
  XNOR U3907 ( .A(n928), .B(n884), .Z(n875) );
  NAND U3908 ( .A(n904), .B(n875), .Z(n827) );
  XNOR U3909 ( .A(n828), .B(n827), .Z(n841) );
  IV U3910 ( .A(n833), .Z(n887) );
  XNOR U3911 ( .A(n887), .B(n829), .Z(n894) );
  AND U3912 ( .A(n883), .B(n894), .Z(n831) );
  AND U3913 ( .A(x[24]), .B(n898), .Z(n830) );
  XNOR U3914 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U3915 ( .A(n884), .B(n832), .Z(n836) );
  NAND U3916 ( .A(x[24]), .B(n883), .Z(n834) );
  OR U3917 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3918 ( .A(n836), .B(n835), .Z(n837) );
  XNOR U3919 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U3920 ( .A(n841), .B(n839), .Z(n861) );
  IV U3921 ( .A(n861), .Z(n868) );
  AND U3922 ( .A(n914), .B(n840), .Z(n843) );
  XOR U3923 ( .A(x[25]), .B(x[31]), .Z(n916) );
  AND U3924 ( .A(n877), .B(n916), .Z(n846) );
  XNOR U3925 ( .A(n846), .B(n841), .Z(n842) );
  XNOR U3926 ( .A(n843), .B(n842), .Z(n867) );
  NANDN U3927 ( .A(n868), .B(n867), .Z(n844) );
  NAND U3928 ( .A(n872), .B(n844), .Z(n854) );
  XNOR U3929 ( .A(n846), .B(n845), .Z(n851) );
  ANDN U3930 ( .B(n847), .A(x[25]), .Z(n848) );
  XNOR U3931 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U3932 ( .A(n851), .B(n850), .Z(n864) );
  XOR U3933 ( .A(n867), .B(n864), .Z(n852) );
  NAND U3934 ( .A(n868), .B(n852), .Z(n853) );
  NAND U3935 ( .A(n854), .B(n853), .Z(n913) );
  ANDN U3936 ( .B(n855), .A(n913), .Z(n879) );
  IV U3937 ( .A(n864), .Z(n870) );
  XOR U3938 ( .A(n872), .B(n868), .Z(n856) );
  NANDN U3939 ( .A(n870), .B(n856), .Z(n859) );
  NANDN U3940 ( .A(n868), .B(n870), .Z(n857) );
  NANDN U3941 ( .A(n867), .B(n857), .Z(n858) );
  NAND U3942 ( .A(n859), .B(n858), .Z(n923) );
  XNOR U3943 ( .A(n913), .B(n923), .Z(n889) );
  AND U3944 ( .A(n860), .B(n889), .Z(n882) );
  OR U3945 ( .A(n867), .B(n864), .Z(n866) );
  ANDN U3946 ( .B(n867), .A(n861), .Z(n862) );
  XNOR U3947 ( .A(n862), .B(n872), .Z(n863) );
  NAND U3948 ( .A(n864), .B(n863), .Z(n865) );
  NAND U3949 ( .A(n866), .B(n865), .Z(n886) );
  NAND U3950 ( .A(n868), .B(n872), .Z(n874) );
  NAND U3951 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U3952 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U3953 ( .A(n872), .B(n871), .Z(n873) );
  NAND U3954 ( .A(n874), .B(n873), .Z(n930) );
  NAND U3955 ( .A(n905), .B(n875), .Z(n876) );
  XNOR U3956 ( .A(n882), .B(n876), .Z(n925) );
  XOR U3957 ( .A(n913), .B(n930), .Z(n915) );
  AND U3958 ( .A(n877), .B(n915), .Z(n900) );
  XNOR U3959 ( .A(n925), .B(n900), .Z(n878) );
  XNOR U3960 ( .A(n879), .B(n878), .Z(n933) );
  NAND U3961 ( .A(n891), .B(n880), .Z(n881) );
  XNOR U3962 ( .A(n882), .B(n881), .Z(n908) );
  AND U3963 ( .A(n883), .B(n893), .Z(n924) );
  NANDN U3964 ( .A(n884), .B(n886), .Z(n885) );
  XNOR U3965 ( .A(n924), .B(n885), .Z(n912) );
  XNOR U3966 ( .A(n908), .B(n912), .Z(n897) );
  XOR U3967 ( .A(n933), .B(n897), .Z(z[24]) );
  AND U3968 ( .A(n887), .B(n886), .Z(n896) );
  AND U3969 ( .A(n889), .B(n888), .Z(n907) );
  NAND U3970 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U3971 ( .A(n907), .B(n892), .Z(n934) );
  AND U3972 ( .A(n894), .B(n893), .Z(n901) );
  XNOR U3973 ( .A(n934), .B(n901), .Z(n895) );
  XNOR U3974 ( .A(n896), .B(n895), .Z(n921) );
  XNOR U3975 ( .A(n921), .B(n897), .Z(n941) );
  AND U3976 ( .A(n898), .B(n923), .Z(n903) );
  NANDN U3977 ( .A(n930), .B(n928), .Z(n899) );
  XNOR U3978 ( .A(n900), .B(n899), .Z(n911) );
  XNOR U3979 ( .A(n901), .B(n911), .Z(n902) );
  XNOR U3980 ( .A(n903), .B(n902), .Z(n910) );
  NAND U3981 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3982 ( .A(n907), .B(n906), .Z(n917) );
  XNOR U3983 ( .A(n908), .B(n917), .Z(n909) );
  XNOR U3984 ( .A(n910), .B(n909), .Z(n920) );
  XNOR U3985 ( .A(n941), .B(n920), .Z(z[25]) );
  XNOR U3986 ( .A(n912), .B(n911), .Z(z[26]) );
  NOR U3987 ( .A(n914), .B(n913), .Z(n919) );
  AND U3988 ( .A(n916), .B(n915), .Z(n932) );
  XNOR U3989 ( .A(n917), .B(n932), .Z(n918) );
  XNOR U3990 ( .A(n919), .B(n918), .Z(n940) );
  XOR U3991 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U3992 ( .A(n940), .B(n922), .Z(z[27]) );
  XOR U3993 ( .A(n933), .B(z[26]), .Z(z[28]) );
  AND U3994 ( .A(x[24]), .B(n923), .Z(n927) );
  XNOR U3995 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U3996 ( .A(n927), .B(n926), .Z(n942) );
  XOR U3997 ( .A(n928), .B(x[25]), .Z(n929) );
  NANDN U3998 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U3999 ( .A(n932), .B(n931), .Z(n936) );
  XNOR U4000 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U4001 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U4002 ( .A(n942), .B(n937), .Z(z[29]) );
  XNOR U4003 ( .A(n939), .B(n938), .Z(z[2]) );
  XNOR U4004 ( .A(n941), .B(n940), .Z(z[30]) );
  XOR U4005 ( .A(n942), .B(z[25]), .Z(z[31]) );
  XOR U4006 ( .A(x[35]), .B(x[33]), .Z(n945) );
  XNOR U4007 ( .A(x[32]), .B(x[38]), .Z(n944) );
  XOR U4008 ( .A(n944), .B(x[34]), .Z(n943) );
  XNOR U4009 ( .A(n945), .B(n943), .Z(n980) );
  XNOR U4010 ( .A(x[37]), .B(n944), .Z(n1053) );
  XOR U4011 ( .A(n1053), .B(x[36]), .Z(n1023) );
  IV U4012 ( .A(n1023), .Z(n954) );
  XNOR U4013 ( .A(x[39]), .B(x[36]), .Z(n948) );
  XNOR U4014 ( .A(n945), .B(n948), .Z(n1008) );
  NOR U4015 ( .A(n954), .B(n1008), .Z(n947) );
  XNOR U4016 ( .A(n1053), .B(x[39]), .Z(n1039) );
  XNOR U4017 ( .A(x[34]), .B(n1039), .Z(n963) );
  XNOR U4018 ( .A(x[33]), .B(n963), .Z(n958) );
  AND U4019 ( .A(x[32]), .B(n958), .Z(n946) );
  XNOR U4020 ( .A(n947), .B(n946), .Z(n951) );
  XNOR U4021 ( .A(n980), .B(n1039), .Z(n970) );
  IV U4022 ( .A(n980), .Z(n965) );
  XNOR U4023 ( .A(x[32]), .B(n965), .Z(n985) );
  IV U4024 ( .A(n948), .Z(n1013) );
  AND U4025 ( .A(n985), .B(n1013), .Z(n953) );
  IV U4026 ( .A(n1053), .Z(n972) );
  XNOR U4027 ( .A(n980), .B(n972), .Z(n1002) );
  XOR U4028 ( .A(n1002), .B(n1008), .Z(n1005) );
  XOR U4029 ( .A(x[34]), .B(x[36]), .Z(n1015) );
  NAND U4030 ( .A(n1005), .B(n1015), .Z(n949) );
  XNOR U4031 ( .A(n953), .B(n949), .Z(n974) );
  XNOR U4032 ( .A(n970), .B(n974), .Z(n950) );
  XNOR U4033 ( .A(n951), .B(n950), .Z(n997) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1029) );
  XNOR U4035 ( .A(x[32]), .B(n1008), .Z(n1009) );
  XNOR U4036 ( .A(n1053), .B(n1009), .Z(n1000) );
  NAND U4037 ( .A(n1029), .B(n1000), .Z(n952) );
  XNOR U4038 ( .A(n953), .B(n952), .Z(n966) );
  IV U4039 ( .A(n958), .Z(n1012) );
  XNOR U4040 ( .A(n1012), .B(n954), .Z(n1019) );
  AND U4041 ( .A(n1008), .B(n1019), .Z(n956) );
  AND U4042 ( .A(x[32]), .B(n1023), .Z(n955) );
  XNOR U4043 ( .A(n956), .B(n955), .Z(n957) );
  NANDN U4044 ( .A(n1009), .B(n957), .Z(n961) );
  NAND U4045 ( .A(x[32]), .B(n1008), .Z(n959) );
  OR U4046 ( .A(n959), .B(n958), .Z(n960) );
  NAND U4047 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U4048 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U4049 ( .A(n966), .B(n964), .Z(n986) );
  IV U4050 ( .A(n986), .Z(n993) );
  AND U4051 ( .A(n1039), .B(n965), .Z(n968) );
  XOR U4052 ( .A(x[33]), .B(x[39]), .Z(n1041) );
  AND U4053 ( .A(n1002), .B(n1041), .Z(n971) );
  XNOR U4054 ( .A(n971), .B(n966), .Z(n967) );
  XNOR U4055 ( .A(n968), .B(n967), .Z(n992) );
  NANDN U4056 ( .A(n993), .B(n992), .Z(n969) );
  NAND U4057 ( .A(n997), .B(n969), .Z(n979) );
  XNOR U4058 ( .A(n971), .B(n970), .Z(n976) );
  ANDN U4059 ( .B(n972), .A(x[33]), .Z(n973) );
  XNOR U4060 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U4061 ( .A(n976), .B(n975), .Z(n989) );
  XOR U4062 ( .A(n992), .B(n989), .Z(n977) );
  NAND U4063 ( .A(n993), .B(n977), .Z(n978) );
  NAND U4064 ( .A(n979), .B(n978), .Z(n1038) );
  ANDN U4065 ( .B(n980), .A(n1038), .Z(n1004) );
  IV U4066 ( .A(n989), .Z(n995) );
  XOR U4067 ( .A(n997), .B(n993), .Z(n981) );
  NANDN U4068 ( .A(n995), .B(n981), .Z(n984) );
  NANDN U4069 ( .A(n993), .B(n995), .Z(n982) );
  NANDN U4070 ( .A(n992), .B(n982), .Z(n983) );
  NAND U4071 ( .A(n984), .B(n983), .Z(n1048) );
  XNOR U4072 ( .A(n1038), .B(n1048), .Z(n1014) );
  AND U4073 ( .A(n985), .B(n1014), .Z(n1007) );
  OR U4074 ( .A(n992), .B(n989), .Z(n991) );
  ANDN U4075 ( .B(n992), .A(n986), .Z(n987) );
  XNOR U4076 ( .A(n987), .B(n997), .Z(n988) );
  NAND U4077 ( .A(n989), .B(n988), .Z(n990) );
  NAND U4078 ( .A(n991), .B(n990), .Z(n1011) );
  NAND U4079 ( .A(n993), .B(n997), .Z(n999) );
  NAND U4080 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U4081 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U4082 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4083 ( .A(n999), .B(n998), .Z(n1055) );
  NAND U4084 ( .A(n1030), .B(n1000), .Z(n1001) );
  XNOR U4085 ( .A(n1007), .B(n1001), .Z(n1050) );
  XOR U4086 ( .A(n1038), .B(n1055), .Z(n1040) );
  AND U4087 ( .A(n1002), .B(n1040), .Z(n1025) );
  XNOR U4088 ( .A(n1050), .B(n1025), .Z(n1003) );
  XNOR U4089 ( .A(n1004), .B(n1003), .Z(n1058) );
  NAND U4090 ( .A(n1016), .B(n1005), .Z(n1006) );
  XNOR U4091 ( .A(n1007), .B(n1006), .Z(n1033) );
  AND U4092 ( .A(n1008), .B(n1018), .Z(n1049) );
  NANDN U4093 ( .A(n1009), .B(n1011), .Z(n1010) );
  XNOR U4094 ( .A(n1049), .B(n1010), .Z(n1037) );
  XNOR U4095 ( .A(n1033), .B(n1037), .Z(n1022) );
  XOR U4096 ( .A(n1058), .B(n1022), .Z(z[32]) );
  AND U4097 ( .A(n1012), .B(n1011), .Z(n1021) );
  AND U4098 ( .A(n1014), .B(n1013), .Z(n1032) );
  NAND U4099 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U4100 ( .A(n1032), .B(n1017), .Z(n1059) );
  AND U4101 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U4102 ( .A(n1059), .B(n1026), .Z(n1020) );
  XNOR U4103 ( .A(n1021), .B(n1020), .Z(n1046) );
  XNOR U4104 ( .A(n1046), .B(n1022), .Z(n1064) );
  AND U4105 ( .A(n1023), .B(n1048), .Z(n1028) );
  NANDN U4106 ( .A(n1055), .B(n1053), .Z(n1024) );
  XNOR U4107 ( .A(n1025), .B(n1024), .Z(n1036) );
  XNOR U4108 ( .A(n1026), .B(n1036), .Z(n1027) );
  XNOR U4109 ( .A(n1028), .B(n1027), .Z(n1035) );
  NAND U4110 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U4111 ( .A(n1032), .B(n1031), .Z(n1042) );
  XNOR U4112 ( .A(n1033), .B(n1042), .Z(n1034) );
  XNOR U4113 ( .A(n1035), .B(n1034), .Z(n1045) );
  XNOR U4114 ( .A(n1064), .B(n1045), .Z(z[33]) );
  XNOR U4115 ( .A(n1037), .B(n1036), .Z(z[34]) );
  NOR U4116 ( .A(n1039), .B(n1038), .Z(n1044) );
  AND U4117 ( .A(n1041), .B(n1040), .Z(n1057) );
  XNOR U4118 ( .A(n1042), .B(n1057), .Z(n1043) );
  XNOR U4119 ( .A(n1044), .B(n1043), .Z(n1063) );
  XOR U4120 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U4121 ( .A(n1063), .B(n1047), .Z(z[35]) );
  XOR U4122 ( .A(n1058), .B(z[34]), .Z(z[36]) );
  AND U4123 ( .A(x[32]), .B(n1048), .Z(n1052) );
  XNOR U4124 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U4125 ( .A(n1052), .B(n1051), .Z(n1065) );
  XOR U4126 ( .A(n1053), .B(x[33]), .Z(n1054) );
  NANDN U4127 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U4128 ( .A(n1057), .B(n1056), .Z(n1061) );
  XNOR U4129 ( .A(n1059), .B(n1058), .Z(n1060) );
  XNOR U4130 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U4131 ( .A(n1065), .B(n1062), .Z(z[37]) );
  XNOR U4132 ( .A(n1064), .B(n1063), .Z(z[38]) );
  XOR U4133 ( .A(n1065), .B(z[33]), .Z(z[39]) );
  NOR U4134 ( .A(n1067), .B(n1066), .Z(n1072) );
  AND U4135 ( .A(n1069), .B(n1068), .Z(n1436) );
  XNOR U4136 ( .A(n1070), .B(n1436), .Z(n1071) );
  XNOR U4137 ( .A(n1072), .B(n1071), .Z(n1580) );
  XOR U4138 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U4139 ( .A(n1580), .B(n1075), .Z(z[3]) );
  XOR U4140 ( .A(x[43]), .B(x[41]), .Z(n1078) );
  XNOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1077) );
  XOR U4142 ( .A(n1077), .B(x[42]), .Z(n1076) );
  XNOR U4143 ( .A(n1078), .B(n1076), .Z(n1113) );
  XNOR U4144 ( .A(x[45]), .B(n1077), .Z(n1186) );
  XOR U4145 ( .A(n1186), .B(x[44]), .Z(n1156) );
  IV U4146 ( .A(n1156), .Z(n1087) );
  XNOR U4147 ( .A(x[47]), .B(x[44]), .Z(n1081) );
  XNOR U4148 ( .A(n1078), .B(n1081), .Z(n1141) );
  NOR U4149 ( .A(n1087), .B(n1141), .Z(n1080) );
  XNOR U4150 ( .A(n1186), .B(x[47]), .Z(n1172) );
  XNOR U4151 ( .A(x[42]), .B(n1172), .Z(n1096) );
  XNOR U4152 ( .A(x[41]), .B(n1096), .Z(n1091) );
  AND U4153 ( .A(x[40]), .B(n1091), .Z(n1079) );
  XNOR U4154 ( .A(n1080), .B(n1079), .Z(n1084) );
  XNOR U4155 ( .A(n1113), .B(n1172), .Z(n1103) );
  IV U4156 ( .A(n1113), .Z(n1098) );
  XNOR U4157 ( .A(x[40]), .B(n1098), .Z(n1118) );
  IV U4158 ( .A(n1081), .Z(n1146) );
  AND U4159 ( .A(n1118), .B(n1146), .Z(n1086) );
  IV U4160 ( .A(n1186), .Z(n1105) );
  XNOR U4161 ( .A(n1113), .B(n1105), .Z(n1135) );
  XOR U4162 ( .A(n1135), .B(n1141), .Z(n1138) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1148) );
  NAND U4164 ( .A(n1138), .B(n1148), .Z(n1082) );
  XNOR U4165 ( .A(n1086), .B(n1082), .Z(n1107) );
  XNOR U4166 ( .A(n1103), .B(n1107), .Z(n1083) );
  XNOR U4167 ( .A(n1084), .B(n1083), .Z(n1130) );
  XOR U4168 ( .A(x[42]), .B(x[47]), .Z(n1162) );
  XNOR U4169 ( .A(x[40]), .B(n1141), .Z(n1142) );
  XNOR U4170 ( .A(n1186), .B(n1142), .Z(n1133) );
  NAND U4171 ( .A(n1162), .B(n1133), .Z(n1085) );
  XNOR U4172 ( .A(n1086), .B(n1085), .Z(n1099) );
  IV U4173 ( .A(n1091), .Z(n1145) );
  XNOR U4174 ( .A(n1145), .B(n1087), .Z(n1152) );
  AND U4175 ( .A(n1141), .B(n1152), .Z(n1089) );
  AND U4176 ( .A(x[40]), .B(n1156), .Z(n1088) );
  XNOR U4177 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U4178 ( .A(n1142), .B(n1090), .Z(n1094) );
  NAND U4179 ( .A(x[40]), .B(n1141), .Z(n1092) );
  OR U4180 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U4181 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U4182 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U4183 ( .A(n1099), .B(n1097), .Z(n1119) );
  IV U4184 ( .A(n1119), .Z(n1126) );
  AND U4185 ( .A(n1172), .B(n1098), .Z(n1101) );
  XOR U4186 ( .A(x[41]), .B(x[47]), .Z(n1174) );
  AND U4187 ( .A(n1135), .B(n1174), .Z(n1104) );
  XNOR U4188 ( .A(n1104), .B(n1099), .Z(n1100) );
  XNOR U4189 ( .A(n1101), .B(n1100), .Z(n1125) );
  NANDN U4190 ( .A(n1126), .B(n1125), .Z(n1102) );
  NAND U4191 ( .A(n1130), .B(n1102), .Z(n1112) );
  XNOR U4192 ( .A(n1104), .B(n1103), .Z(n1109) );
  ANDN U4193 ( .B(n1105), .A(x[41]), .Z(n1106) );
  XNOR U4194 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U4195 ( .A(n1109), .B(n1108), .Z(n1122) );
  XOR U4196 ( .A(n1125), .B(n1122), .Z(n1110) );
  NAND U4197 ( .A(n1126), .B(n1110), .Z(n1111) );
  NAND U4198 ( .A(n1112), .B(n1111), .Z(n1171) );
  ANDN U4199 ( .B(n1113), .A(n1171), .Z(n1137) );
  IV U4200 ( .A(n1122), .Z(n1128) );
  XOR U4201 ( .A(n1130), .B(n1126), .Z(n1114) );
  NANDN U4202 ( .A(n1128), .B(n1114), .Z(n1117) );
  NANDN U4203 ( .A(n1126), .B(n1128), .Z(n1115) );
  NANDN U4204 ( .A(n1125), .B(n1115), .Z(n1116) );
  NAND U4205 ( .A(n1117), .B(n1116), .Z(n1181) );
  XNOR U4206 ( .A(n1171), .B(n1181), .Z(n1147) );
  AND U4207 ( .A(n1118), .B(n1147), .Z(n1140) );
  OR U4208 ( .A(n1125), .B(n1122), .Z(n1124) );
  ANDN U4209 ( .B(n1125), .A(n1119), .Z(n1120) );
  XNOR U4210 ( .A(n1120), .B(n1130), .Z(n1121) );
  NAND U4211 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U4212 ( .A(n1124), .B(n1123), .Z(n1144) );
  NAND U4213 ( .A(n1126), .B(n1130), .Z(n1132) );
  NAND U4214 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U4215 ( .A(n1128), .B(n1127), .Z(n1129) );
  NANDN U4216 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U4217 ( .A(n1132), .B(n1131), .Z(n1188) );
  NAND U4218 ( .A(n1163), .B(n1133), .Z(n1134) );
  XNOR U4219 ( .A(n1140), .B(n1134), .Z(n1183) );
  XOR U4220 ( .A(n1171), .B(n1188), .Z(n1173) );
  AND U4221 ( .A(n1135), .B(n1173), .Z(n1158) );
  XNOR U4222 ( .A(n1183), .B(n1158), .Z(n1136) );
  XNOR U4223 ( .A(n1137), .B(n1136), .Z(n1191) );
  NAND U4224 ( .A(n1149), .B(n1138), .Z(n1139) );
  XNOR U4225 ( .A(n1140), .B(n1139), .Z(n1166) );
  AND U4226 ( .A(n1141), .B(n1151), .Z(n1182) );
  NANDN U4227 ( .A(n1142), .B(n1144), .Z(n1143) );
  XNOR U4228 ( .A(n1182), .B(n1143), .Z(n1170) );
  XNOR U4229 ( .A(n1166), .B(n1170), .Z(n1155) );
  XOR U4230 ( .A(n1191), .B(n1155), .Z(z[40]) );
  AND U4231 ( .A(n1145), .B(n1144), .Z(n1154) );
  AND U4232 ( .A(n1147), .B(n1146), .Z(n1165) );
  NAND U4233 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U4234 ( .A(n1165), .B(n1150), .Z(n1192) );
  AND U4235 ( .A(n1152), .B(n1151), .Z(n1159) );
  XNOR U4236 ( .A(n1192), .B(n1159), .Z(n1153) );
  XNOR U4237 ( .A(n1154), .B(n1153), .Z(n1179) );
  XNOR U4238 ( .A(n1179), .B(n1155), .Z(n1197) );
  AND U4239 ( .A(n1156), .B(n1181), .Z(n1161) );
  NANDN U4240 ( .A(n1188), .B(n1186), .Z(n1157) );
  XNOR U4241 ( .A(n1158), .B(n1157), .Z(n1169) );
  XNOR U4242 ( .A(n1159), .B(n1169), .Z(n1160) );
  XNOR U4243 ( .A(n1161), .B(n1160), .Z(n1168) );
  NAND U4244 ( .A(n1163), .B(n1162), .Z(n1164) );
  XNOR U4245 ( .A(n1165), .B(n1164), .Z(n1175) );
  XNOR U4246 ( .A(n1166), .B(n1175), .Z(n1167) );
  XNOR U4247 ( .A(n1168), .B(n1167), .Z(n1178) );
  XNOR U4248 ( .A(n1197), .B(n1178), .Z(z[41]) );
  XNOR U4249 ( .A(n1170), .B(n1169), .Z(z[42]) );
  NOR U4250 ( .A(n1172), .B(n1171), .Z(n1177) );
  AND U4251 ( .A(n1174), .B(n1173), .Z(n1190) );
  XNOR U4252 ( .A(n1175), .B(n1190), .Z(n1176) );
  XNOR U4253 ( .A(n1177), .B(n1176), .Z(n1196) );
  XOR U4254 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4255 ( .A(n1196), .B(n1180), .Z(z[43]) );
  XOR U4256 ( .A(n1191), .B(z[42]), .Z(z[44]) );
  AND U4257 ( .A(x[40]), .B(n1181), .Z(n1185) );
  XNOR U4258 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U4259 ( .A(n1185), .B(n1184), .Z(n1198) );
  XOR U4260 ( .A(n1186), .B(x[41]), .Z(n1187) );
  NANDN U4261 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U4262 ( .A(n1190), .B(n1189), .Z(n1194) );
  XNOR U4263 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U4264 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U4265 ( .A(n1198), .B(n1195), .Z(z[45]) );
  XNOR U4266 ( .A(n1197), .B(n1196), .Z(z[46]) );
  XOR U4267 ( .A(n1198), .B(z[41]), .Z(z[47]) );
  XOR U4268 ( .A(x[51]), .B(x[49]), .Z(n1201) );
  XNOR U4269 ( .A(x[48]), .B(x[54]), .Z(n1200) );
  XOR U4270 ( .A(n1200), .B(x[50]), .Z(n1199) );
  XNOR U4271 ( .A(n1201), .B(n1199), .Z(n1236) );
  XNOR U4272 ( .A(x[53]), .B(n1200), .Z(n1309) );
  XOR U4273 ( .A(n1309), .B(x[52]), .Z(n1279) );
  IV U4274 ( .A(n1279), .Z(n1210) );
  XNOR U4275 ( .A(x[55]), .B(x[52]), .Z(n1204) );
  XNOR U4276 ( .A(n1201), .B(n1204), .Z(n1264) );
  NOR U4277 ( .A(n1210), .B(n1264), .Z(n1203) );
  XNOR U4278 ( .A(n1309), .B(x[55]), .Z(n1295) );
  XNOR U4279 ( .A(x[50]), .B(n1295), .Z(n1219) );
  XNOR U4280 ( .A(x[49]), .B(n1219), .Z(n1214) );
  AND U4281 ( .A(x[48]), .B(n1214), .Z(n1202) );
  XNOR U4282 ( .A(n1203), .B(n1202), .Z(n1207) );
  XNOR U4283 ( .A(n1236), .B(n1295), .Z(n1226) );
  IV U4284 ( .A(n1236), .Z(n1221) );
  XNOR U4285 ( .A(x[48]), .B(n1221), .Z(n1241) );
  IV U4286 ( .A(n1204), .Z(n1269) );
  AND U4287 ( .A(n1241), .B(n1269), .Z(n1209) );
  IV U4288 ( .A(n1309), .Z(n1228) );
  XNOR U4289 ( .A(n1236), .B(n1228), .Z(n1258) );
  XOR U4290 ( .A(n1258), .B(n1264), .Z(n1261) );
  XOR U4291 ( .A(x[50]), .B(x[52]), .Z(n1271) );
  NAND U4292 ( .A(n1261), .B(n1271), .Z(n1205) );
  XNOR U4293 ( .A(n1209), .B(n1205), .Z(n1230) );
  XNOR U4294 ( .A(n1226), .B(n1230), .Z(n1206) );
  XNOR U4295 ( .A(n1207), .B(n1206), .Z(n1253) );
  XOR U4296 ( .A(x[50]), .B(x[55]), .Z(n1285) );
  XNOR U4297 ( .A(x[48]), .B(n1264), .Z(n1265) );
  XNOR U4298 ( .A(n1309), .B(n1265), .Z(n1256) );
  NAND U4299 ( .A(n1285), .B(n1256), .Z(n1208) );
  XNOR U4300 ( .A(n1209), .B(n1208), .Z(n1222) );
  IV U4301 ( .A(n1214), .Z(n1268) );
  XNOR U4302 ( .A(n1268), .B(n1210), .Z(n1275) );
  AND U4303 ( .A(n1264), .B(n1275), .Z(n1212) );
  AND U4304 ( .A(x[48]), .B(n1279), .Z(n1211) );
  XNOR U4305 ( .A(n1212), .B(n1211), .Z(n1213) );
  NANDN U4306 ( .A(n1265), .B(n1213), .Z(n1217) );
  NAND U4307 ( .A(x[48]), .B(n1264), .Z(n1215) );
  OR U4308 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4309 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U4310 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U4311 ( .A(n1222), .B(n1220), .Z(n1242) );
  IV U4312 ( .A(n1242), .Z(n1249) );
  AND U4313 ( .A(n1295), .B(n1221), .Z(n1224) );
  XOR U4314 ( .A(x[49]), .B(x[55]), .Z(n1297) );
  AND U4315 ( .A(n1258), .B(n1297), .Z(n1227) );
  XNOR U4316 ( .A(n1227), .B(n1222), .Z(n1223) );
  XNOR U4317 ( .A(n1224), .B(n1223), .Z(n1248) );
  NANDN U4318 ( .A(n1249), .B(n1248), .Z(n1225) );
  NAND U4319 ( .A(n1253), .B(n1225), .Z(n1235) );
  XNOR U4320 ( .A(n1227), .B(n1226), .Z(n1232) );
  ANDN U4321 ( .B(n1228), .A(x[49]), .Z(n1229) );
  XNOR U4322 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U4323 ( .A(n1232), .B(n1231), .Z(n1245) );
  XOR U4324 ( .A(n1248), .B(n1245), .Z(n1233) );
  NAND U4325 ( .A(n1249), .B(n1233), .Z(n1234) );
  NAND U4326 ( .A(n1235), .B(n1234), .Z(n1294) );
  ANDN U4327 ( .B(n1236), .A(n1294), .Z(n1260) );
  IV U4328 ( .A(n1245), .Z(n1251) );
  XOR U4329 ( .A(n1253), .B(n1249), .Z(n1237) );
  NANDN U4330 ( .A(n1251), .B(n1237), .Z(n1240) );
  NANDN U4331 ( .A(n1249), .B(n1251), .Z(n1238) );
  NANDN U4332 ( .A(n1248), .B(n1238), .Z(n1239) );
  NAND U4333 ( .A(n1240), .B(n1239), .Z(n1304) );
  XNOR U4334 ( .A(n1294), .B(n1304), .Z(n1270) );
  AND U4335 ( .A(n1241), .B(n1270), .Z(n1263) );
  OR U4336 ( .A(n1248), .B(n1245), .Z(n1247) );
  ANDN U4337 ( .B(n1248), .A(n1242), .Z(n1243) );
  XNOR U4338 ( .A(n1243), .B(n1253), .Z(n1244) );
  NAND U4339 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U4340 ( .A(n1247), .B(n1246), .Z(n1267) );
  NAND U4341 ( .A(n1249), .B(n1253), .Z(n1255) );
  NAND U4342 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U4343 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U4344 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U4345 ( .A(n1255), .B(n1254), .Z(n1311) );
  NAND U4346 ( .A(n1286), .B(n1256), .Z(n1257) );
  XNOR U4347 ( .A(n1263), .B(n1257), .Z(n1306) );
  XOR U4348 ( .A(n1294), .B(n1311), .Z(n1296) );
  AND U4349 ( .A(n1258), .B(n1296), .Z(n1281) );
  XNOR U4350 ( .A(n1306), .B(n1281), .Z(n1259) );
  XNOR U4351 ( .A(n1260), .B(n1259), .Z(n1314) );
  NAND U4352 ( .A(n1272), .B(n1261), .Z(n1262) );
  XNOR U4353 ( .A(n1263), .B(n1262), .Z(n1289) );
  AND U4354 ( .A(n1264), .B(n1274), .Z(n1305) );
  NANDN U4355 ( .A(n1265), .B(n1267), .Z(n1266) );
  XNOR U4356 ( .A(n1305), .B(n1266), .Z(n1293) );
  XNOR U4357 ( .A(n1289), .B(n1293), .Z(n1278) );
  XOR U4358 ( .A(n1314), .B(n1278), .Z(z[48]) );
  AND U4359 ( .A(n1268), .B(n1267), .Z(n1277) );
  AND U4360 ( .A(n1270), .B(n1269), .Z(n1288) );
  NAND U4361 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U4362 ( .A(n1288), .B(n1273), .Z(n1315) );
  AND U4363 ( .A(n1275), .B(n1274), .Z(n1282) );
  XNOR U4364 ( .A(n1315), .B(n1282), .Z(n1276) );
  XNOR U4365 ( .A(n1277), .B(n1276), .Z(n1302) );
  XNOR U4366 ( .A(n1302), .B(n1278), .Z(n1320) );
  AND U4367 ( .A(n1279), .B(n1304), .Z(n1284) );
  NANDN U4368 ( .A(n1311), .B(n1309), .Z(n1280) );
  XNOR U4369 ( .A(n1281), .B(n1280), .Z(n1292) );
  XNOR U4370 ( .A(n1282), .B(n1292), .Z(n1283) );
  XNOR U4371 ( .A(n1284), .B(n1283), .Z(n1291) );
  NAND U4372 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U4373 ( .A(n1288), .B(n1287), .Z(n1298) );
  XNOR U4374 ( .A(n1289), .B(n1298), .Z(n1290) );
  XNOR U4375 ( .A(n1291), .B(n1290), .Z(n1301) );
  XNOR U4376 ( .A(n1320), .B(n1301), .Z(z[49]) );
  XOR U4377 ( .A(n1437), .B(z[2]), .Z(z[4]) );
  XNOR U4378 ( .A(n1293), .B(n1292), .Z(z[50]) );
  NOR U4379 ( .A(n1295), .B(n1294), .Z(n1300) );
  AND U4380 ( .A(n1297), .B(n1296), .Z(n1313) );
  XNOR U4381 ( .A(n1298), .B(n1313), .Z(n1299) );
  XNOR U4382 ( .A(n1300), .B(n1299), .Z(n1319) );
  XOR U4383 ( .A(n1302), .B(n1301), .Z(n1303) );
  XNOR U4384 ( .A(n1319), .B(n1303), .Z(z[51]) );
  XOR U4385 ( .A(n1314), .B(z[50]), .Z(z[52]) );
  AND U4386 ( .A(x[48]), .B(n1304), .Z(n1308) );
  XNOR U4387 ( .A(n1306), .B(n1305), .Z(n1307) );
  XNOR U4388 ( .A(n1308), .B(n1307), .Z(n1321) );
  XOR U4389 ( .A(n1309), .B(x[49]), .Z(n1310) );
  NANDN U4390 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U4391 ( .A(n1313), .B(n1312), .Z(n1317) );
  XNOR U4392 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U4393 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U4394 ( .A(n1321), .B(n1318), .Z(z[53]) );
  XNOR U4395 ( .A(n1320), .B(n1319), .Z(z[54]) );
  XOR U4396 ( .A(n1321), .B(z[49]), .Z(z[55]) );
  XOR U4397 ( .A(x[59]), .B(x[57]), .Z(n1324) );
  XNOR U4398 ( .A(x[56]), .B(x[62]), .Z(n1323) );
  XOR U4399 ( .A(n1323), .B(x[58]), .Z(n1322) );
  XNOR U4400 ( .A(n1324), .B(n1322), .Z(n1359) );
  XNOR U4401 ( .A(x[61]), .B(n1323), .Z(n1447) );
  XOR U4402 ( .A(n1447), .B(x[60]), .Z(n1402) );
  IV U4403 ( .A(n1402), .Z(n1333) );
  XNOR U4404 ( .A(x[63]), .B(x[60]), .Z(n1327) );
  XNOR U4405 ( .A(n1324), .B(n1327), .Z(n1387) );
  NOR U4406 ( .A(n1333), .B(n1387), .Z(n1326) );
  XNOR U4407 ( .A(n1447), .B(x[63]), .Z(n1418) );
  XNOR U4408 ( .A(x[58]), .B(n1418), .Z(n1342) );
  XNOR U4409 ( .A(x[57]), .B(n1342), .Z(n1337) );
  AND U4410 ( .A(x[56]), .B(n1337), .Z(n1325) );
  XNOR U4411 ( .A(n1326), .B(n1325), .Z(n1330) );
  XNOR U4412 ( .A(n1359), .B(n1418), .Z(n1349) );
  IV U4413 ( .A(n1359), .Z(n1344) );
  XNOR U4414 ( .A(x[56]), .B(n1344), .Z(n1364) );
  IV U4415 ( .A(n1327), .Z(n1392) );
  AND U4416 ( .A(n1364), .B(n1392), .Z(n1332) );
  IV U4417 ( .A(n1447), .Z(n1351) );
  XNOR U4418 ( .A(n1359), .B(n1351), .Z(n1381) );
  XOR U4419 ( .A(n1381), .B(n1387), .Z(n1384) );
  XOR U4420 ( .A(x[58]), .B(x[60]), .Z(n1394) );
  NAND U4421 ( .A(n1384), .B(n1394), .Z(n1328) );
  XNOR U4422 ( .A(n1332), .B(n1328), .Z(n1353) );
  XNOR U4423 ( .A(n1349), .B(n1353), .Z(n1329) );
  XNOR U4424 ( .A(n1330), .B(n1329), .Z(n1376) );
  XOR U4425 ( .A(x[58]), .B(x[63]), .Z(n1408) );
  XNOR U4426 ( .A(x[56]), .B(n1387), .Z(n1388) );
  XNOR U4427 ( .A(n1447), .B(n1388), .Z(n1379) );
  NAND U4428 ( .A(n1408), .B(n1379), .Z(n1331) );
  XNOR U4429 ( .A(n1332), .B(n1331), .Z(n1345) );
  IV U4430 ( .A(n1337), .Z(n1391) );
  XNOR U4431 ( .A(n1391), .B(n1333), .Z(n1398) );
  AND U4432 ( .A(n1387), .B(n1398), .Z(n1335) );
  AND U4433 ( .A(x[56]), .B(n1402), .Z(n1334) );
  XNOR U4434 ( .A(n1335), .B(n1334), .Z(n1336) );
  NANDN U4435 ( .A(n1388), .B(n1336), .Z(n1340) );
  NAND U4436 ( .A(x[56]), .B(n1387), .Z(n1338) );
  OR U4437 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U4438 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4439 ( .A(n1342), .B(n1341), .Z(n1343) );
  XNOR U4440 ( .A(n1345), .B(n1343), .Z(n1365) );
  IV U4441 ( .A(n1365), .Z(n1372) );
  AND U4442 ( .A(n1418), .B(n1344), .Z(n1347) );
  XOR U4443 ( .A(x[57]), .B(x[63]), .Z(n1420) );
  AND U4444 ( .A(n1381), .B(n1420), .Z(n1350) );
  XNOR U4445 ( .A(n1350), .B(n1345), .Z(n1346) );
  XNOR U4446 ( .A(n1347), .B(n1346), .Z(n1371) );
  NANDN U4447 ( .A(n1372), .B(n1371), .Z(n1348) );
  NAND U4448 ( .A(n1376), .B(n1348), .Z(n1358) );
  XNOR U4449 ( .A(n1350), .B(n1349), .Z(n1355) );
  ANDN U4450 ( .B(n1351), .A(x[57]), .Z(n1352) );
  XNOR U4451 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U4452 ( .A(n1355), .B(n1354), .Z(n1368) );
  XOR U4453 ( .A(n1371), .B(n1368), .Z(n1356) );
  NAND U4454 ( .A(n1372), .B(n1356), .Z(n1357) );
  NAND U4455 ( .A(n1358), .B(n1357), .Z(n1417) );
  ANDN U4456 ( .B(n1359), .A(n1417), .Z(n1383) );
  IV U4457 ( .A(n1368), .Z(n1374) );
  XOR U4458 ( .A(n1376), .B(n1372), .Z(n1360) );
  NANDN U4459 ( .A(n1374), .B(n1360), .Z(n1363) );
  NANDN U4460 ( .A(n1372), .B(n1374), .Z(n1361) );
  NANDN U4461 ( .A(n1371), .B(n1361), .Z(n1362) );
  NAND U4462 ( .A(n1363), .B(n1362), .Z(n1442) );
  XNOR U4463 ( .A(n1417), .B(n1442), .Z(n1393) );
  AND U4464 ( .A(n1364), .B(n1393), .Z(n1386) );
  OR U4465 ( .A(n1371), .B(n1368), .Z(n1370) );
  ANDN U4466 ( .B(n1371), .A(n1365), .Z(n1366) );
  XNOR U4467 ( .A(n1366), .B(n1376), .Z(n1367) );
  NAND U4468 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U4469 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U4470 ( .A(n1372), .B(n1376), .Z(n1378) );
  NAND U4471 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4472 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U4473 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U4474 ( .A(n1378), .B(n1377), .Z(n1449) );
  NAND U4475 ( .A(n1409), .B(n1379), .Z(n1380) );
  XNOR U4476 ( .A(n1386), .B(n1380), .Z(n1444) );
  XOR U4477 ( .A(n1417), .B(n1449), .Z(n1419) );
  AND U4478 ( .A(n1381), .B(n1419), .Z(n1404) );
  XNOR U4479 ( .A(n1444), .B(n1404), .Z(n1382) );
  XNOR U4480 ( .A(n1383), .B(n1382), .Z(n1452) );
  NAND U4481 ( .A(n1395), .B(n1384), .Z(n1385) );
  XNOR U4482 ( .A(n1386), .B(n1385), .Z(n1412) );
  AND U4483 ( .A(n1387), .B(n1397), .Z(n1443) );
  NANDN U4484 ( .A(n1388), .B(n1390), .Z(n1389) );
  XNOR U4485 ( .A(n1443), .B(n1389), .Z(n1416) );
  XNOR U4486 ( .A(n1412), .B(n1416), .Z(n1401) );
  XOR U4487 ( .A(n1452), .B(n1401), .Z(z[56]) );
  AND U4488 ( .A(n1391), .B(n1390), .Z(n1400) );
  AND U4489 ( .A(n1393), .B(n1392), .Z(n1411) );
  NAND U4490 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U4491 ( .A(n1411), .B(n1396), .Z(n1453) );
  AND U4492 ( .A(n1398), .B(n1397), .Z(n1405) );
  XNOR U4493 ( .A(n1453), .B(n1405), .Z(n1399) );
  XNOR U4494 ( .A(n1400), .B(n1399), .Z(n1425) );
  XNOR U4495 ( .A(n1425), .B(n1401), .Z(n1458) );
  AND U4496 ( .A(n1402), .B(n1442), .Z(n1407) );
  NANDN U4497 ( .A(n1449), .B(n1447), .Z(n1403) );
  XNOR U4498 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U4499 ( .A(n1405), .B(n1415), .Z(n1406) );
  XNOR U4500 ( .A(n1407), .B(n1406), .Z(n1414) );
  NAND U4501 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U4502 ( .A(n1411), .B(n1410), .Z(n1421) );
  XNOR U4503 ( .A(n1412), .B(n1421), .Z(n1413) );
  XNOR U4504 ( .A(n1414), .B(n1413), .Z(n1424) );
  XNOR U4505 ( .A(n1458), .B(n1424), .Z(z[57]) );
  XNOR U4506 ( .A(n1416), .B(n1415), .Z(z[58]) );
  NOR U4507 ( .A(n1418), .B(n1417), .Z(n1423) );
  AND U4508 ( .A(n1420), .B(n1419), .Z(n1451) );
  XNOR U4509 ( .A(n1421), .B(n1451), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1457) );
  XOR U4511 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U4512 ( .A(n1457), .B(n1426), .Z(z[59]) );
  AND U4513 ( .A(x[0]), .B(n1427), .Z(n1431) );
  XNOR U4514 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U4515 ( .A(n1431), .B(n1430), .Z(n1708) );
  XOR U4516 ( .A(n1432), .B(x[1]), .Z(n1433) );
  NANDN U4517 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U4518 ( .A(n1436), .B(n1435), .Z(n1440) );
  XNOR U4519 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U4520 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U4521 ( .A(n1708), .B(n1441), .Z(z[5]) );
  XOR U4522 ( .A(n1452), .B(z[58]), .Z(z[60]) );
  AND U4523 ( .A(x[56]), .B(n1442), .Z(n1446) );
  XNOR U4524 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U4525 ( .A(n1446), .B(n1445), .Z(n1459) );
  XOR U4526 ( .A(n1447), .B(x[57]), .Z(n1448) );
  NANDN U4527 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U4528 ( .A(n1451), .B(n1450), .Z(n1455) );
  XNOR U4529 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U4530 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U4531 ( .A(n1459), .B(n1456), .Z(z[61]) );
  XNOR U4532 ( .A(n1458), .B(n1457), .Z(z[62]) );
  XOR U4533 ( .A(n1459), .B(z[57]), .Z(z[63]) );
  XOR U4534 ( .A(x[67]), .B(x[65]), .Z(n1462) );
  XNOR U4535 ( .A(x[64]), .B(x[70]), .Z(n1461) );
  XOR U4536 ( .A(n1461), .B(x[66]), .Z(n1460) );
  XNOR U4537 ( .A(n1462), .B(n1460), .Z(n1497) );
  XNOR U4538 ( .A(x[69]), .B(n1461), .Z(n1570) );
  XOR U4539 ( .A(n1570), .B(x[68]), .Z(n1540) );
  IV U4540 ( .A(n1540), .Z(n1471) );
  XNOR U4541 ( .A(x[71]), .B(x[68]), .Z(n1465) );
  XNOR U4542 ( .A(n1462), .B(n1465), .Z(n1525) );
  NOR U4543 ( .A(n1471), .B(n1525), .Z(n1464) );
  XNOR U4544 ( .A(n1570), .B(x[71]), .Z(n1556) );
  XNOR U4545 ( .A(x[66]), .B(n1556), .Z(n1480) );
  XNOR U4546 ( .A(x[65]), .B(n1480), .Z(n1475) );
  AND U4547 ( .A(x[64]), .B(n1475), .Z(n1463) );
  XNOR U4548 ( .A(n1464), .B(n1463), .Z(n1468) );
  XNOR U4549 ( .A(n1497), .B(n1556), .Z(n1487) );
  IV U4550 ( .A(n1497), .Z(n1482) );
  XNOR U4551 ( .A(x[64]), .B(n1482), .Z(n1502) );
  IV U4552 ( .A(n1465), .Z(n1530) );
  AND U4553 ( .A(n1502), .B(n1530), .Z(n1470) );
  IV U4554 ( .A(n1570), .Z(n1489) );
  XNOR U4555 ( .A(n1497), .B(n1489), .Z(n1519) );
  XOR U4556 ( .A(n1519), .B(n1525), .Z(n1522) );
  XOR U4557 ( .A(x[66]), .B(x[68]), .Z(n1532) );
  NAND U4558 ( .A(n1522), .B(n1532), .Z(n1466) );
  XNOR U4559 ( .A(n1470), .B(n1466), .Z(n1491) );
  XNOR U4560 ( .A(n1487), .B(n1491), .Z(n1467) );
  XNOR U4561 ( .A(n1468), .B(n1467), .Z(n1514) );
  XOR U4562 ( .A(x[66]), .B(x[71]), .Z(n1546) );
  XNOR U4563 ( .A(x[64]), .B(n1525), .Z(n1526) );
  XNOR U4564 ( .A(n1570), .B(n1526), .Z(n1517) );
  NAND U4565 ( .A(n1546), .B(n1517), .Z(n1469) );
  XNOR U4566 ( .A(n1470), .B(n1469), .Z(n1483) );
  IV U4567 ( .A(n1475), .Z(n1529) );
  XNOR U4568 ( .A(n1529), .B(n1471), .Z(n1536) );
  AND U4569 ( .A(n1525), .B(n1536), .Z(n1473) );
  AND U4570 ( .A(x[64]), .B(n1540), .Z(n1472) );
  XNOR U4571 ( .A(n1473), .B(n1472), .Z(n1474) );
  NANDN U4572 ( .A(n1526), .B(n1474), .Z(n1478) );
  NAND U4573 ( .A(x[64]), .B(n1525), .Z(n1476) );
  OR U4574 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U4575 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4576 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR U4577 ( .A(n1483), .B(n1481), .Z(n1503) );
  IV U4578 ( .A(n1503), .Z(n1510) );
  AND U4579 ( .A(n1556), .B(n1482), .Z(n1485) );
  XOR U4580 ( .A(x[65]), .B(x[71]), .Z(n1558) );
  AND U4581 ( .A(n1519), .B(n1558), .Z(n1488) );
  XNOR U4582 ( .A(n1488), .B(n1483), .Z(n1484) );
  XNOR U4583 ( .A(n1485), .B(n1484), .Z(n1509) );
  NANDN U4584 ( .A(n1510), .B(n1509), .Z(n1486) );
  NAND U4585 ( .A(n1514), .B(n1486), .Z(n1496) );
  XNOR U4586 ( .A(n1488), .B(n1487), .Z(n1493) );
  ANDN U4587 ( .B(n1489), .A(x[65]), .Z(n1490) );
  XNOR U4588 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U4589 ( .A(n1493), .B(n1492), .Z(n1506) );
  XOR U4590 ( .A(n1509), .B(n1506), .Z(n1494) );
  NAND U4591 ( .A(n1510), .B(n1494), .Z(n1495) );
  NAND U4592 ( .A(n1496), .B(n1495), .Z(n1555) );
  ANDN U4593 ( .B(n1497), .A(n1555), .Z(n1521) );
  IV U4594 ( .A(n1506), .Z(n1512) );
  XOR U4595 ( .A(n1514), .B(n1510), .Z(n1498) );
  NANDN U4596 ( .A(n1512), .B(n1498), .Z(n1501) );
  NANDN U4597 ( .A(n1510), .B(n1512), .Z(n1499) );
  NANDN U4598 ( .A(n1509), .B(n1499), .Z(n1500) );
  NAND U4599 ( .A(n1501), .B(n1500), .Z(n1565) );
  XNOR U4600 ( .A(n1555), .B(n1565), .Z(n1531) );
  AND U4601 ( .A(n1502), .B(n1531), .Z(n1524) );
  OR U4602 ( .A(n1509), .B(n1506), .Z(n1508) );
  ANDN U4603 ( .B(n1509), .A(n1503), .Z(n1504) );
  XNOR U4604 ( .A(n1504), .B(n1514), .Z(n1505) );
  NAND U4605 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U4606 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U4607 ( .A(n1510), .B(n1514), .Z(n1516) );
  NAND U4608 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4609 ( .A(n1512), .B(n1511), .Z(n1513) );
  NANDN U4610 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U4611 ( .A(n1516), .B(n1515), .Z(n1572) );
  NAND U4612 ( .A(n1547), .B(n1517), .Z(n1518) );
  XNOR U4613 ( .A(n1524), .B(n1518), .Z(n1567) );
  XOR U4614 ( .A(n1555), .B(n1572), .Z(n1557) );
  AND U4615 ( .A(n1519), .B(n1557), .Z(n1542) );
  XNOR U4616 ( .A(n1567), .B(n1542), .Z(n1520) );
  XNOR U4617 ( .A(n1521), .B(n1520), .Z(n1575) );
  NAND U4618 ( .A(n1533), .B(n1522), .Z(n1523) );
  XNOR U4619 ( .A(n1524), .B(n1523), .Z(n1550) );
  AND U4620 ( .A(n1525), .B(n1535), .Z(n1566) );
  NANDN U4621 ( .A(n1526), .B(n1528), .Z(n1527) );
  XNOR U4622 ( .A(n1566), .B(n1527), .Z(n1554) );
  XNOR U4623 ( .A(n1550), .B(n1554), .Z(n1539) );
  XOR U4624 ( .A(n1575), .B(n1539), .Z(z[64]) );
  AND U4625 ( .A(n1529), .B(n1528), .Z(n1538) );
  AND U4626 ( .A(n1531), .B(n1530), .Z(n1549) );
  NAND U4627 ( .A(n1533), .B(n1532), .Z(n1534) );
  XNOR U4628 ( .A(n1549), .B(n1534), .Z(n1576) );
  AND U4629 ( .A(n1536), .B(n1535), .Z(n1543) );
  XNOR U4630 ( .A(n1576), .B(n1543), .Z(n1537) );
  XNOR U4631 ( .A(n1538), .B(n1537), .Z(n1563) );
  XNOR U4632 ( .A(n1563), .B(n1539), .Z(n1583) );
  AND U4633 ( .A(n1540), .B(n1565), .Z(n1545) );
  NANDN U4634 ( .A(n1572), .B(n1570), .Z(n1541) );
  XNOR U4635 ( .A(n1542), .B(n1541), .Z(n1553) );
  XNOR U4636 ( .A(n1543), .B(n1553), .Z(n1544) );
  XNOR U4637 ( .A(n1545), .B(n1544), .Z(n1552) );
  NAND U4638 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U4639 ( .A(n1549), .B(n1548), .Z(n1559) );
  XNOR U4640 ( .A(n1550), .B(n1559), .Z(n1551) );
  XNOR U4641 ( .A(n1552), .B(n1551), .Z(n1562) );
  XNOR U4642 ( .A(n1583), .B(n1562), .Z(z[65]) );
  XNOR U4643 ( .A(n1554), .B(n1553), .Z(z[66]) );
  NOR U4644 ( .A(n1556), .B(n1555), .Z(n1561) );
  AND U4645 ( .A(n1558), .B(n1557), .Z(n1574) );
  XNOR U4646 ( .A(n1559), .B(n1574), .Z(n1560) );
  XNOR U4647 ( .A(n1561), .B(n1560), .Z(n1582) );
  XOR U4648 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U4649 ( .A(n1582), .B(n1564), .Z(z[67]) );
  XOR U4650 ( .A(n1575), .B(z[66]), .Z(z[68]) );
  AND U4651 ( .A(x[64]), .B(n1565), .Z(n1569) );
  XNOR U4652 ( .A(n1567), .B(n1566), .Z(n1568) );
  XNOR U4653 ( .A(n1569), .B(n1568), .Z(n1584) );
  XOR U4654 ( .A(n1570), .B(x[65]), .Z(n1571) );
  NANDN U4655 ( .A(n1572), .B(n1571), .Z(n1573) );
  XNOR U4656 ( .A(n1574), .B(n1573), .Z(n1578) );
  XNOR U4657 ( .A(n1576), .B(n1575), .Z(n1577) );
  XNOR U4658 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U4659 ( .A(n1584), .B(n1579), .Z(z[69]) );
  XNOR U4660 ( .A(n1581), .B(n1580), .Z(z[6]) );
  XNOR U4661 ( .A(n1583), .B(n1582), .Z(z[70]) );
  XOR U4662 ( .A(n1584), .B(z[65]), .Z(z[71]) );
  XOR U4663 ( .A(x[75]), .B(x[73]), .Z(n1587) );
  XNOR U4664 ( .A(x[72]), .B(x[78]), .Z(n1586) );
  XOR U4665 ( .A(n1586), .B(x[74]), .Z(n1585) );
  XNOR U4666 ( .A(n1587), .B(n1585), .Z(n1622) );
  XNOR U4667 ( .A(x[77]), .B(n1586), .Z(n1695) );
  XOR U4668 ( .A(n1695), .B(x[76]), .Z(n1665) );
  IV U4669 ( .A(n1665), .Z(n1596) );
  XNOR U4670 ( .A(x[79]), .B(x[76]), .Z(n1590) );
  XNOR U4671 ( .A(n1587), .B(n1590), .Z(n1650) );
  NOR U4672 ( .A(n1596), .B(n1650), .Z(n1589) );
  XNOR U4673 ( .A(n1695), .B(x[79]), .Z(n1681) );
  XNOR U4674 ( .A(x[74]), .B(n1681), .Z(n1605) );
  XNOR U4675 ( .A(x[73]), .B(n1605), .Z(n1600) );
  AND U4676 ( .A(x[72]), .B(n1600), .Z(n1588) );
  XNOR U4677 ( .A(n1589), .B(n1588), .Z(n1593) );
  XNOR U4678 ( .A(n1622), .B(n1681), .Z(n1612) );
  IV U4679 ( .A(n1622), .Z(n1607) );
  XNOR U4680 ( .A(x[72]), .B(n1607), .Z(n1627) );
  IV U4681 ( .A(n1590), .Z(n1655) );
  AND U4682 ( .A(n1627), .B(n1655), .Z(n1595) );
  IV U4683 ( .A(n1695), .Z(n1614) );
  XNOR U4684 ( .A(n1622), .B(n1614), .Z(n1644) );
  XOR U4685 ( .A(n1644), .B(n1650), .Z(n1647) );
  XOR U4686 ( .A(x[74]), .B(x[76]), .Z(n1657) );
  NAND U4687 ( .A(n1647), .B(n1657), .Z(n1591) );
  XNOR U4688 ( .A(n1595), .B(n1591), .Z(n1616) );
  XNOR U4689 ( .A(n1612), .B(n1616), .Z(n1592) );
  XNOR U4690 ( .A(n1593), .B(n1592), .Z(n1639) );
  XOR U4691 ( .A(x[74]), .B(x[79]), .Z(n1671) );
  XNOR U4692 ( .A(x[72]), .B(n1650), .Z(n1651) );
  XNOR U4693 ( .A(n1695), .B(n1651), .Z(n1642) );
  NAND U4694 ( .A(n1671), .B(n1642), .Z(n1594) );
  XNOR U4695 ( .A(n1595), .B(n1594), .Z(n1608) );
  IV U4696 ( .A(n1600), .Z(n1654) );
  XNOR U4697 ( .A(n1654), .B(n1596), .Z(n1661) );
  AND U4698 ( .A(n1650), .B(n1661), .Z(n1598) );
  AND U4699 ( .A(x[72]), .B(n1665), .Z(n1597) );
  XNOR U4700 ( .A(n1598), .B(n1597), .Z(n1599) );
  NANDN U4701 ( .A(n1651), .B(n1599), .Z(n1603) );
  NAND U4702 ( .A(x[72]), .B(n1650), .Z(n1601) );
  OR U4703 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U4704 ( .A(n1603), .B(n1602), .Z(n1604) );
  XNOR U4705 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U4706 ( .A(n1608), .B(n1606), .Z(n1628) );
  IV U4707 ( .A(n1628), .Z(n1635) );
  AND U4708 ( .A(n1681), .B(n1607), .Z(n1610) );
  XOR U4709 ( .A(x[73]), .B(x[79]), .Z(n1683) );
  AND U4710 ( .A(n1644), .B(n1683), .Z(n1613) );
  XNOR U4711 ( .A(n1613), .B(n1608), .Z(n1609) );
  XNOR U4712 ( .A(n1610), .B(n1609), .Z(n1634) );
  NANDN U4713 ( .A(n1635), .B(n1634), .Z(n1611) );
  NAND U4714 ( .A(n1639), .B(n1611), .Z(n1621) );
  XNOR U4715 ( .A(n1613), .B(n1612), .Z(n1618) );
  ANDN U4716 ( .B(n1614), .A(x[73]), .Z(n1615) );
  XNOR U4717 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4718 ( .A(n1618), .B(n1617), .Z(n1631) );
  XOR U4719 ( .A(n1634), .B(n1631), .Z(n1619) );
  NAND U4720 ( .A(n1635), .B(n1619), .Z(n1620) );
  NAND U4721 ( .A(n1621), .B(n1620), .Z(n1680) );
  ANDN U4722 ( .B(n1622), .A(n1680), .Z(n1646) );
  IV U4723 ( .A(n1631), .Z(n1637) );
  XOR U4724 ( .A(n1639), .B(n1635), .Z(n1623) );
  NANDN U4725 ( .A(n1637), .B(n1623), .Z(n1626) );
  NANDN U4726 ( .A(n1635), .B(n1637), .Z(n1624) );
  NANDN U4727 ( .A(n1634), .B(n1624), .Z(n1625) );
  NAND U4728 ( .A(n1626), .B(n1625), .Z(n1690) );
  XNOR U4729 ( .A(n1680), .B(n1690), .Z(n1656) );
  AND U4730 ( .A(n1627), .B(n1656), .Z(n1649) );
  OR U4731 ( .A(n1634), .B(n1631), .Z(n1633) );
  ANDN U4732 ( .B(n1634), .A(n1628), .Z(n1629) );
  XNOR U4733 ( .A(n1629), .B(n1639), .Z(n1630) );
  NAND U4734 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U4735 ( .A(n1633), .B(n1632), .Z(n1653) );
  NAND U4736 ( .A(n1635), .B(n1639), .Z(n1641) );
  NAND U4737 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U4738 ( .A(n1637), .B(n1636), .Z(n1638) );
  NANDN U4739 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U4740 ( .A(n1641), .B(n1640), .Z(n1697) );
  NAND U4741 ( .A(n1672), .B(n1642), .Z(n1643) );
  XNOR U4742 ( .A(n1649), .B(n1643), .Z(n1692) );
  XOR U4743 ( .A(n1680), .B(n1697), .Z(n1682) );
  AND U4744 ( .A(n1644), .B(n1682), .Z(n1667) );
  XNOR U4745 ( .A(n1692), .B(n1667), .Z(n1645) );
  XNOR U4746 ( .A(n1646), .B(n1645), .Z(n1700) );
  NAND U4747 ( .A(n1658), .B(n1647), .Z(n1648) );
  XNOR U4748 ( .A(n1649), .B(n1648), .Z(n1675) );
  AND U4749 ( .A(n1650), .B(n1660), .Z(n1691) );
  NANDN U4750 ( .A(n1651), .B(n1653), .Z(n1652) );
  XNOR U4751 ( .A(n1691), .B(n1652), .Z(n1679) );
  XNOR U4752 ( .A(n1675), .B(n1679), .Z(n1664) );
  XOR U4753 ( .A(n1700), .B(n1664), .Z(z[72]) );
  AND U4754 ( .A(n1654), .B(n1653), .Z(n1663) );
  AND U4755 ( .A(n1656), .B(n1655), .Z(n1674) );
  NAND U4756 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U4757 ( .A(n1674), .B(n1659), .Z(n1701) );
  AND U4758 ( .A(n1661), .B(n1660), .Z(n1668) );
  XNOR U4759 ( .A(n1701), .B(n1668), .Z(n1662) );
  XNOR U4760 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U4761 ( .A(n1688), .B(n1664), .Z(n1706) );
  AND U4762 ( .A(n1665), .B(n1690), .Z(n1670) );
  NANDN U4763 ( .A(n1697), .B(n1695), .Z(n1666) );
  XNOR U4764 ( .A(n1667), .B(n1666), .Z(n1678) );
  XNOR U4765 ( .A(n1668), .B(n1678), .Z(n1669) );
  XNOR U4766 ( .A(n1670), .B(n1669), .Z(n1677) );
  NAND U4767 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR U4768 ( .A(n1674), .B(n1673), .Z(n1684) );
  XNOR U4769 ( .A(n1675), .B(n1684), .Z(n1676) );
  XNOR U4770 ( .A(n1677), .B(n1676), .Z(n1687) );
  XNOR U4771 ( .A(n1706), .B(n1687), .Z(z[73]) );
  XNOR U4772 ( .A(n1679), .B(n1678), .Z(z[74]) );
  NOR U4773 ( .A(n1681), .B(n1680), .Z(n1686) );
  AND U4774 ( .A(n1683), .B(n1682), .Z(n1699) );
  XNOR U4775 ( .A(n1684), .B(n1699), .Z(n1685) );
  XNOR U4776 ( .A(n1686), .B(n1685), .Z(n1705) );
  XOR U4777 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4778 ( .A(n1705), .B(n1689), .Z(z[75]) );
  XOR U4779 ( .A(n1700), .B(z[74]), .Z(z[76]) );
  AND U4780 ( .A(x[72]), .B(n1690), .Z(n1694) );
  XNOR U4781 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4782 ( .A(n1694), .B(n1693), .Z(n1707) );
  XOR U4783 ( .A(n1695), .B(x[73]), .Z(n1696) );
  NANDN U4784 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U4785 ( .A(n1699), .B(n1698), .Z(n1703) );
  XNOR U4786 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U4787 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U4788 ( .A(n1707), .B(n1704), .Z(z[77]) );
  XNOR U4789 ( .A(n1706), .B(n1705), .Z(z[78]) );
  XOR U4790 ( .A(n1707), .B(z[73]), .Z(z[79]) );
  XOR U4791 ( .A(n1708), .B(z[1]), .Z(z[7]) );
  XOR U4792 ( .A(x[83]), .B(x[81]), .Z(n1711) );
  XNOR U4793 ( .A(x[80]), .B(x[86]), .Z(n1710) );
  XOR U4794 ( .A(n1710), .B(x[82]), .Z(n1709) );
  XNOR U4795 ( .A(n1711), .B(n1709), .Z(n1746) );
  XNOR U4796 ( .A(x[85]), .B(n1710), .Z(n1819) );
  XOR U4797 ( .A(n1819), .B(x[84]), .Z(n1789) );
  IV U4798 ( .A(n1789), .Z(n1720) );
  XNOR U4799 ( .A(x[87]), .B(x[84]), .Z(n1714) );
  XNOR U4800 ( .A(n1711), .B(n1714), .Z(n1774) );
  NOR U4801 ( .A(n1720), .B(n1774), .Z(n1713) );
  XNOR U4802 ( .A(n1819), .B(x[87]), .Z(n1805) );
  XNOR U4803 ( .A(x[82]), .B(n1805), .Z(n1729) );
  XNOR U4804 ( .A(x[81]), .B(n1729), .Z(n1724) );
  AND U4805 ( .A(x[80]), .B(n1724), .Z(n1712) );
  XNOR U4806 ( .A(n1713), .B(n1712), .Z(n1717) );
  XNOR U4807 ( .A(n1746), .B(n1805), .Z(n1736) );
  IV U4808 ( .A(n1746), .Z(n1731) );
  XNOR U4809 ( .A(x[80]), .B(n1731), .Z(n1751) );
  IV U4810 ( .A(n1714), .Z(n1779) );
  AND U4811 ( .A(n1751), .B(n1779), .Z(n1719) );
  IV U4812 ( .A(n1819), .Z(n1738) );
  XNOR U4813 ( .A(n1746), .B(n1738), .Z(n1768) );
  XOR U4814 ( .A(n1768), .B(n1774), .Z(n1771) );
  XOR U4815 ( .A(x[82]), .B(x[84]), .Z(n1781) );
  NAND U4816 ( .A(n1771), .B(n1781), .Z(n1715) );
  XNOR U4817 ( .A(n1719), .B(n1715), .Z(n1740) );
  XNOR U4818 ( .A(n1736), .B(n1740), .Z(n1716) );
  XNOR U4819 ( .A(n1717), .B(n1716), .Z(n1763) );
  XOR U4820 ( .A(x[82]), .B(x[87]), .Z(n1795) );
  XNOR U4821 ( .A(x[80]), .B(n1774), .Z(n1775) );
  XNOR U4822 ( .A(n1819), .B(n1775), .Z(n1766) );
  NAND U4823 ( .A(n1795), .B(n1766), .Z(n1718) );
  XNOR U4824 ( .A(n1719), .B(n1718), .Z(n1732) );
  IV U4825 ( .A(n1724), .Z(n1778) );
  XNOR U4826 ( .A(n1778), .B(n1720), .Z(n1785) );
  AND U4827 ( .A(n1774), .B(n1785), .Z(n1722) );
  AND U4828 ( .A(x[80]), .B(n1789), .Z(n1721) );
  XNOR U4829 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U4830 ( .A(n1775), .B(n1723), .Z(n1727) );
  NAND U4831 ( .A(x[80]), .B(n1774), .Z(n1725) );
  OR U4832 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U4833 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U4834 ( .A(n1729), .B(n1728), .Z(n1730) );
  XNOR U4835 ( .A(n1732), .B(n1730), .Z(n1752) );
  IV U4836 ( .A(n1752), .Z(n1759) );
  AND U4837 ( .A(n1805), .B(n1731), .Z(n1734) );
  XOR U4838 ( .A(x[81]), .B(x[87]), .Z(n1807) );
  AND U4839 ( .A(n1768), .B(n1807), .Z(n1737) );
  XNOR U4840 ( .A(n1737), .B(n1732), .Z(n1733) );
  XNOR U4841 ( .A(n1734), .B(n1733), .Z(n1758) );
  NANDN U4842 ( .A(n1759), .B(n1758), .Z(n1735) );
  NAND U4843 ( .A(n1763), .B(n1735), .Z(n1745) );
  XNOR U4844 ( .A(n1737), .B(n1736), .Z(n1742) );
  ANDN U4845 ( .B(n1738), .A(x[81]), .Z(n1739) );
  XNOR U4846 ( .A(n1740), .B(n1739), .Z(n1741) );
  XNOR U4847 ( .A(n1742), .B(n1741), .Z(n1755) );
  XOR U4848 ( .A(n1758), .B(n1755), .Z(n1743) );
  NAND U4849 ( .A(n1759), .B(n1743), .Z(n1744) );
  NAND U4850 ( .A(n1745), .B(n1744), .Z(n1804) );
  ANDN U4851 ( .B(n1746), .A(n1804), .Z(n1770) );
  IV U4852 ( .A(n1755), .Z(n1761) );
  XOR U4853 ( .A(n1763), .B(n1759), .Z(n1747) );
  NANDN U4854 ( .A(n1761), .B(n1747), .Z(n1750) );
  NANDN U4855 ( .A(n1759), .B(n1761), .Z(n1748) );
  NANDN U4856 ( .A(n1758), .B(n1748), .Z(n1749) );
  NAND U4857 ( .A(n1750), .B(n1749), .Z(n1814) );
  XNOR U4858 ( .A(n1804), .B(n1814), .Z(n1780) );
  AND U4859 ( .A(n1751), .B(n1780), .Z(n1773) );
  OR U4860 ( .A(n1758), .B(n1755), .Z(n1757) );
  ANDN U4861 ( .B(n1758), .A(n1752), .Z(n1753) );
  XNOR U4862 ( .A(n1753), .B(n1763), .Z(n1754) );
  NAND U4863 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U4864 ( .A(n1757), .B(n1756), .Z(n1777) );
  NAND U4865 ( .A(n1759), .B(n1763), .Z(n1765) );
  NAND U4866 ( .A(n1759), .B(n1758), .Z(n1760) );
  XNOR U4867 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U4868 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1821) );
  NAND U4870 ( .A(n1796), .B(n1766), .Z(n1767) );
  XNOR U4871 ( .A(n1773), .B(n1767), .Z(n1816) );
  XOR U4872 ( .A(n1804), .B(n1821), .Z(n1806) );
  AND U4873 ( .A(n1768), .B(n1806), .Z(n1791) );
  XNOR U4874 ( .A(n1816), .B(n1791), .Z(n1769) );
  XNOR U4875 ( .A(n1770), .B(n1769), .Z(n1824) );
  NAND U4876 ( .A(n1782), .B(n1771), .Z(n1772) );
  XNOR U4877 ( .A(n1773), .B(n1772), .Z(n1799) );
  AND U4878 ( .A(n1774), .B(n1784), .Z(n1815) );
  NANDN U4879 ( .A(n1775), .B(n1777), .Z(n1776) );
  XNOR U4880 ( .A(n1815), .B(n1776), .Z(n1803) );
  XNOR U4881 ( .A(n1799), .B(n1803), .Z(n1788) );
  XOR U4882 ( .A(n1824), .B(n1788), .Z(z[80]) );
  AND U4883 ( .A(n1778), .B(n1777), .Z(n1787) );
  AND U4884 ( .A(n1780), .B(n1779), .Z(n1798) );
  NAND U4885 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U4886 ( .A(n1798), .B(n1783), .Z(n1825) );
  AND U4887 ( .A(n1785), .B(n1784), .Z(n1792) );
  XNOR U4888 ( .A(n1825), .B(n1792), .Z(n1786) );
  XNOR U4889 ( .A(n1787), .B(n1786), .Z(n1812) );
  XNOR U4890 ( .A(n1812), .B(n1788), .Z(n1830) );
  AND U4891 ( .A(n1789), .B(n1814), .Z(n1794) );
  NANDN U4892 ( .A(n1821), .B(n1819), .Z(n1790) );
  XNOR U4893 ( .A(n1791), .B(n1790), .Z(n1802) );
  XNOR U4894 ( .A(n1792), .B(n1802), .Z(n1793) );
  XNOR U4895 ( .A(n1794), .B(n1793), .Z(n1801) );
  NAND U4896 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U4897 ( .A(n1798), .B(n1797), .Z(n1808) );
  XNOR U4898 ( .A(n1799), .B(n1808), .Z(n1800) );
  XNOR U4899 ( .A(n1801), .B(n1800), .Z(n1811) );
  XNOR U4900 ( .A(n1830), .B(n1811), .Z(z[81]) );
  XNOR U4901 ( .A(n1803), .B(n1802), .Z(z[82]) );
  NOR U4902 ( .A(n1805), .B(n1804), .Z(n1810) );
  AND U4903 ( .A(n1807), .B(n1806), .Z(n1823) );
  XNOR U4904 ( .A(n1808), .B(n1823), .Z(n1809) );
  XNOR U4905 ( .A(n1810), .B(n1809), .Z(n1829) );
  XOR U4906 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U4907 ( .A(n1829), .B(n1813), .Z(z[83]) );
  XOR U4908 ( .A(n1824), .B(z[82]), .Z(z[84]) );
  AND U4909 ( .A(x[80]), .B(n1814), .Z(n1818) );
  XNOR U4910 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U4911 ( .A(n1818), .B(n1817), .Z(n1831) );
  XOR U4912 ( .A(n1819), .B(x[81]), .Z(n1820) );
  NANDN U4913 ( .A(n1821), .B(n1820), .Z(n1822) );
  XNOR U4914 ( .A(n1823), .B(n1822), .Z(n1827) );
  XNOR U4915 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U4916 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U4917 ( .A(n1831), .B(n1828), .Z(z[85]) );
  XNOR U4918 ( .A(n1830), .B(n1829), .Z(z[86]) );
  XOR U4919 ( .A(n1831), .B(z[81]), .Z(z[87]) );
  XOR U4920 ( .A(x[91]), .B(x[89]), .Z(n1834) );
  XNOR U4921 ( .A(x[88]), .B(x[94]), .Z(n1833) );
  XOR U4922 ( .A(n1833), .B(x[90]), .Z(n1832) );
  XNOR U4923 ( .A(n1834), .B(n1832), .Z(n1869) );
  XNOR U4924 ( .A(x[93]), .B(n1833), .Z(n1944) );
  XOR U4925 ( .A(n1944), .B(x[92]), .Z(n1912) );
  IV U4926 ( .A(n1912), .Z(n1843) );
  XNOR U4927 ( .A(x[95]), .B(x[92]), .Z(n1837) );
  XNOR U4928 ( .A(n1834), .B(n1837), .Z(n1897) );
  NOR U4929 ( .A(n1843), .B(n1897), .Z(n1836) );
  XNOR U4930 ( .A(n1944), .B(x[95]), .Z(n1930) );
  XNOR U4931 ( .A(x[90]), .B(n1930), .Z(n1852) );
  XNOR U4932 ( .A(x[89]), .B(n1852), .Z(n1847) );
  AND U4933 ( .A(x[88]), .B(n1847), .Z(n1835) );
  XNOR U4934 ( .A(n1836), .B(n1835), .Z(n1840) );
  XNOR U4935 ( .A(n1869), .B(n1930), .Z(n1859) );
  IV U4936 ( .A(n1869), .Z(n1854) );
  XNOR U4937 ( .A(x[88]), .B(n1854), .Z(n1874) );
  IV U4938 ( .A(n1837), .Z(n1902) );
  AND U4939 ( .A(n1874), .B(n1902), .Z(n1842) );
  IV U4940 ( .A(n1944), .Z(n1861) );
  XNOR U4941 ( .A(n1869), .B(n1861), .Z(n1891) );
  XOR U4942 ( .A(n1891), .B(n1897), .Z(n1894) );
  XOR U4943 ( .A(x[90]), .B(x[92]), .Z(n1904) );
  NAND U4944 ( .A(n1894), .B(n1904), .Z(n1838) );
  XNOR U4945 ( .A(n1842), .B(n1838), .Z(n1863) );
  XNOR U4946 ( .A(n1859), .B(n1863), .Z(n1839) );
  XNOR U4947 ( .A(n1840), .B(n1839), .Z(n1886) );
  XOR U4948 ( .A(x[90]), .B(x[95]), .Z(n1918) );
  XNOR U4949 ( .A(x[88]), .B(n1897), .Z(n1898) );
  XNOR U4950 ( .A(n1944), .B(n1898), .Z(n1889) );
  NAND U4951 ( .A(n1918), .B(n1889), .Z(n1841) );
  XNOR U4952 ( .A(n1842), .B(n1841), .Z(n1855) );
  IV U4953 ( .A(n1847), .Z(n1901) );
  XNOR U4954 ( .A(n1901), .B(n1843), .Z(n1908) );
  AND U4955 ( .A(n1897), .B(n1908), .Z(n1845) );
  AND U4956 ( .A(x[88]), .B(n1912), .Z(n1844) );
  XNOR U4957 ( .A(n1845), .B(n1844), .Z(n1846) );
  NANDN U4958 ( .A(n1898), .B(n1846), .Z(n1850) );
  NAND U4959 ( .A(x[88]), .B(n1897), .Z(n1848) );
  OR U4960 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U4961 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U4962 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U4963 ( .A(n1855), .B(n1853), .Z(n1875) );
  IV U4964 ( .A(n1875), .Z(n1882) );
  AND U4965 ( .A(n1930), .B(n1854), .Z(n1857) );
  XOR U4966 ( .A(x[89]), .B(x[95]), .Z(n1932) );
  AND U4967 ( .A(n1891), .B(n1932), .Z(n1860) );
  XNOR U4968 ( .A(n1860), .B(n1855), .Z(n1856) );
  XNOR U4969 ( .A(n1857), .B(n1856), .Z(n1881) );
  NANDN U4970 ( .A(n1882), .B(n1881), .Z(n1858) );
  NAND U4971 ( .A(n1886), .B(n1858), .Z(n1868) );
  XNOR U4972 ( .A(n1860), .B(n1859), .Z(n1865) );
  ANDN U4973 ( .B(n1861), .A(x[89]), .Z(n1862) );
  XNOR U4974 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U4975 ( .A(n1865), .B(n1864), .Z(n1878) );
  XOR U4976 ( .A(n1881), .B(n1878), .Z(n1866) );
  NAND U4977 ( .A(n1882), .B(n1866), .Z(n1867) );
  NAND U4978 ( .A(n1868), .B(n1867), .Z(n1929) );
  ANDN U4979 ( .B(n1869), .A(n1929), .Z(n1893) );
  IV U4980 ( .A(n1878), .Z(n1884) );
  XOR U4981 ( .A(n1886), .B(n1882), .Z(n1870) );
  NANDN U4982 ( .A(n1884), .B(n1870), .Z(n1873) );
  NANDN U4983 ( .A(n1882), .B(n1884), .Z(n1871) );
  NANDN U4984 ( .A(n1881), .B(n1871), .Z(n1872) );
  NAND U4985 ( .A(n1873), .B(n1872), .Z(n1939) );
  XNOR U4986 ( .A(n1929), .B(n1939), .Z(n1903) );
  AND U4987 ( .A(n1874), .B(n1903), .Z(n1896) );
  OR U4988 ( .A(n1881), .B(n1878), .Z(n1880) );
  ANDN U4989 ( .B(n1881), .A(n1875), .Z(n1876) );
  XNOR U4990 ( .A(n1876), .B(n1886), .Z(n1877) );
  NAND U4991 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U4992 ( .A(n1880), .B(n1879), .Z(n1900) );
  NAND U4993 ( .A(n1882), .B(n1886), .Z(n1888) );
  NAND U4994 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U4995 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U4996 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4997 ( .A(n1888), .B(n1887), .Z(n1946) );
  NAND U4998 ( .A(n1919), .B(n1889), .Z(n1890) );
  XNOR U4999 ( .A(n1896), .B(n1890), .Z(n1941) );
  XOR U5000 ( .A(n1929), .B(n1946), .Z(n1931) );
  AND U5001 ( .A(n1891), .B(n1931), .Z(n1914) );
  XNOR U5002 ( .A(n1941), .B(n1914), .Z(n1892) );
  XNOR U5003 ( .A(n1893), .B(n1892), .Z(n1949) );
  NAND U5004 ( .A(n1905), .B(n1894), .Z(n1895) );
  XNOR U5005 ( .A(n1896), .B(n1895), .Z(n1922) );
  AND U5006 ( .A(n1897), .B(n1907), .Z(n1940) );
  NANDN U5007 ( .A(n1898), .B(n1900), .Z(n1899) );
  XNOR U5008 ( .A(n1940), .B(n1899), .Z(n1928) );
  XNOR U5009 ( .A(n1922), .B(n1928), .Z(n1911) );
  XOR U5010 ( .A(n1949), .B(n1911), .Z(z[88]) );
  AND U5011 ( .A(n1901), .B(n1900), .Z(n1910) );
  AND U5012 ( .A(n1903), .B(n1902), .Z(n1921) );
  NAND U5013 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U5014 ( .A(n1921), .B(n1906), .Z(n1950) );
  AND U5015 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U5016 ( .A(n1950), .B(n1915), .Z(n1909) );
  XNOR U5017 ( .A(n1910), .B(n1909), .Z(n1937) );
  XNOR U5018 ( .A(n1937), .B(n1911), .Z(n1955) );
  AND U5019 ( .A(n1912), .B(n1939), .Z(n1917) );
  NANDN U5020 ( .A(n1946), .B(n1944), .Z(n1913) );
  XNOR U5021 ( .A(n1914), .B(n1913), .Z(n1927) );
  XNOR U5022 ( .A(n1915), .B(n1927), .Z(n1916) );
  XNOR U5023 ( .A(n1917), .B(n1916), .Z(n1924) );
  NAND U5024 ( .A(n1919), .B(n1918), .Z(n1920) );
  XNOR U5025 ( .A(n1921), .B(n1920), .Z(n1933) );
  XNOR U5026 ( .A(n1922), .B(n1933), .Z(n1923) );
  XNOR U5027 ( .A(n1924), .B(n1923), .Z(n1936) );
  XNOR U5028 ( .A(n1955), .B(n1936), .Z(z[89]) );
  XOR U5029 ( .A(n1926), .B(n1925), .Z(z[8]) );
  XNOR U5030 ( .A(n1928), .B(n1927), .Z(z[90]) );
  NOR U5031 ( .A(n1930), .B(n1929), .Z(n1935) );
  AND U5032 ( .A(n1932), .B(n1931), .Z(n1948) );
  XNOR U5033 ( .A(n1933), .B(n1948), .Z(n1934) );
  XNOR U5034 ( .A(n1935), .B(n1934), .Z(n1954) );
  XOR U5035 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U5036 ( .A(n1954), .B(n1938), .Z(z[91]) );
  XOR U5037 ( .A(n1949), .B(z[90]), .Z(z[92]) );
  AND U5038 ( .A(x[88]), .B(n1939), .Z(n1943) );
  XNOR U5039 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5040 ( .A(n1943), .B(n1942), .Z(n1956) );
  XOR U5041 ( .A(n1944), .B(x[89]), .Z(n1945) );
  NANDN U5042 ( .A(n1946), .B(n1945), .Z(n1947) );
  XNOR U5043 ( .A(n1948), .B(n1947), .Z(n1952) );
  XNOR U5044 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U5045 ( .A(n1952), .B(n1951), .Z(n1953) );
  XNOR U5046 ( .A(n1956), .B(n1953), .Z(z[93]) );
  XNOR U5047 ( .A(n1955), .B(n1954), .Z(z[94]) );
  XOR U5048 ( .A(n1956), .B(z[89]), .Z(z[95]) );
  XOR U5049 ( .A(n1958), .B(n1957), .Z(z[96]) );
  XOR U5050 ( .A(n1960), .B(n1959), .Z(n1961) );
  XNOR U5051 ( .A(n1962), .B(n1961), .Z(z[99]) );
endmodule


module SubBytes_3 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;

  XNOR U2962 ( .A(n886), .B(n930), .Z(n905) );
  XNOR U2963 ( .A(n775), .B(n1434), .Z(n794) );
  XNOR U2964 ( .A(n1144), .B(n1188), .Z(n1163) );
  XOR U2965 ( .A(n1814), .B(n1777), .Z(n1784) );
  XNOR U2966 ( .A(n1390), .B(n1449), .Z(n1409) );
  XNOR U2967 ( .A(n738), .B(n807), .Z(n757) );
  XOR U2968 ( .A(n1565), .B(n1528), .Z(n1535) );
  XOR U2969 ( .A(n290), .B(n253), .Z(n260) );
  XNOR U2970 ( .A(n1900), .B(n1946), .Z(n1919) );
  XNOR U2971 ( .A(n1267), .B(n1311), .Z(n1286) );
  XOR U2972 ( .A(n622), .B(n585), .Z(n592) );
  XOR U2973 ( .A(n1048), .B(n1011), .Z(n1018) );
  XOR U2974 ( .A(n1690), .B(n1653), .Z(n1660) );
  XOR U2975 ( .A(n467), .B(n430), .Z(n437) );
  NOR U2976 ( .A(n654), .B(x[9]), .Z(n1) );
  XNOR U2977 ( .A(n329), .B(n328), .Z(n2) );
  XNOR U2978 ( .A(n1), .B(n2), .Z(n3) );
  XNOR U2979 ( .A(n312), .B(n3), .Z(n345) );
  XOR U2980 ( .A(n923), .B(n886), .Z(n893) );
  XOR U2981 ( .A(n1427), .B(n775), .Z(n782) );
  XNOR U2982 ( .A(n1777), .B(n1821), .Z(n1796) );
  XOR U2983 ( .A(n1181), .B(n1144), .Z(n1151) );
  XNOR U2984 ( .A(n1528), .B(n1572), .Z(n1547) );
  XOR U2985 ( .A(n800), .B(n738), .Z(n745) );
  XOR U2986 ( .A(n1442), .B(n1390), .Z(n1397) );
  XNOR U2987 ( .A(n253), .B(n297), .Z(n272) );
  XOR U2988 ( .A(n1304), .B(n1267), .Z(n1274) );
  XOR U2989 ( .A(n1939), .B(n1900), .Z(n1907) );
  XNOR U2990 ( .A(n585), .B(n629), .Z(n604) );
  XNOR U2991 ( .A(n1653), .B(n1697), .Z(n1672) );
  XNOR U2992 ( .A(n1011), .B(n1055), .Z(n1030) );
  XNOR U2993 ( .A(n430), .B(n474), .Z(n449) );
  XOR U2994 ( .A(n163), .B(n134), .Z(n157) );
  XOR U2995 ( .A(n77), .B(n78), .Z(n129) );
  XNOR U2996 ( .A(x[9]), .B(n323), .Z(n318) );
  XOR U2997 ( .A(n604), .B(n588), .Z(n590) );
  XOR U2998 ( .A(n905), .B(n889), .Z(n891) );
  XOR U2999 ( .A(n794), .B(n778), .Z(n780) );
  XOR U3000 ( .A(n643), .B(n508), .Z(n511) );
  XOR U3001 ( .A(n757), .B(n741), .Z(n743) );
  XOR U3002 ( .A(n1409), .B(n1393), .Z(n1395) );
  XOR U3003 ( .A(n1286), .B(n1270), .Z(n1272) );
  XOR U3004 ( .A(n1030), .B(n1014), .Z(n1016) );
  XOR U3005 ( .A(n1163), .B(n1147), .Z(n1149) );
  XOR U3006 ( .A(n1672), .B(n1656), .Z(n1658) );
  XOR U3007 ( .A(n1796), .B(n1780), .Z(n1782) );
  XOR U3008 ( .A(n1547), .B(n1531), .Z(n1533) );
  XOR U3009 ( .A(n1919), .B(n1903), .Z(n1905) );
  XOR U3010 ( .A(n272), .B(n256), .Z(n258) );
  NANDN U3011 ( .A(n116), .B(n121), .Z(n4) );
  XOR U3012 ( .A(n116), .B(n119), .Z(n5) );
  OR U3013 ( .A(n121), .B(n5), .Z(n6) );
  NANDN U3014 ( .A(n117), .B(n6), .Z(n7) );
  NAND U3015 ( .A(n4), .B(n7), .Z(n169) );
  XOR U3016 ( .A(n449), .B(n433), .Z(n435) );
  XOR U3017 ( .A(x[3]), .B(x[1]), .Z(n10) );
  XNOR U3018 ( .A(x[0]), .B(x[6]), .Z(n9) );
  XOR U3019 ( .A(n9), .B(x[2]), .Z(n8) );
  XNOR U3020 ( .A(n10), .B(n8), .Z(n45) );
  XNOR U3021 ( .A(x[5]), .B(n9), .Z(n1432) );
  XOR U3022 ( .A(n1432), .B(x[4]), .Z(n787) );
  IV U3023 ( .A(n787), .Z(n19) );
  XNOR U3024 ( .A(x[7]), .B(x[4]), .Z(n13) );
  XNOR U3025 ( .A(n10), .B(n13), .Z(n73) );
  NOR U3026 ( .A(n19), .B(n73), .Z(n12) );
  XNOR U3027 ( .A(n1432), .B(x[7]), .Z(n1067) );
  XNOR U3028 ( .A(x[2]), .B(n1067), .Z(n28) );
  XNOR U3029 ( .A(x[1]), .B(n28), .Z(n23) );
  AND U3030 ( .A(x[0]), .B(n23), .Z(n11) );
  XNOR U3031 ( .A(n12), .B(n11), .Z(n16) );
  XNOR U3032 ( .A(n45), .B(n1067), .Z(n35) );
  IV U3033 ( .A(n45), .Z(n30) );
  XNOR U3034 ( .A(x[0]), .B(n30), .Z(n50) );
  IV U3035 ( .A(n13), .Z(n777) );
  AND U3036 ( .A(n50), .B(n777), .Z(n18) );
  IV U3037 ( .A(n1432), .Z(n37) );
  XNOR U3038 ( .A(n45), .B(n37), .Z(n67) );
  XOR U3039 ( .A(n67), .B(n73), .Z(n70) );
  XOR U3040 ( .A(x[2]), .B(x[4]), .Z(n779) );
  NAND U3041 ( .A(n70), .B(n779), .Z(n14) );
  XNOR U3042 ( .A(n18), .B(n14), .Z(n39) );
  XNOR U3043 ( .A(n35), .B(n39), .Z(n15) );
  XNOR U3044 ( .A(n16), .B(n15), .Z(n62) );
  XOR U3045 ( .A(x[2]), .B(x[7]), .Z(n793) );
  XNOR U3046 ( .A(x[0]), .B(n73), .Z(n74) );
  XNOR U3047 ( .A(n1432), .B(n74), .Z(n65) );
  NAND U3048 ( .A(n793), .B(n65), .Z(n17) );
  XNOR U3049 ( .A(n18), .B(n17), .Z(n31) );
  IV U3050 ( .A(n23), .Z(n776) );
  XNOR U3051 ( .A(n776), .B(n19), .Z(n783) );
  AND U3052 ( .A(n73), .B(n783), .Z(n21) );
  AND U3053 ( .A(x[0]), .B(n787), .Z(n20) );
  XNOR U3054 ( .A(n21), .B(n20), .Z(n22) );
  NANDN U3055 ( .A(n74), .B(n22), .Z(n26) );
  NAND U3056 ( .A(x[0]), .B(n73), .Z(n24) );
  OR U3057 ( .A(n24), .B(n23), .Z(n25) );
  NAND U3058 ( .A(n26), .B(n25), .Z(n27) );
  XNOR U3059 ( .A(n28), .B(n27), .Z(n29) );
  XNOR U3060 ( .A(n31), .B(n29), .Z(n51) );
  IV U3061 ( .A(n51), .Z(n58) );
  AND U3062 ( .A(n1067), .B(n30), .Z(n33) );
  XOR U3063 ( .A(x[1]), .B(x[7]), .Z(n1069) );
  AND U3064 ( .A(n67), .B(n1069), .Z(n36) );
  XNOR U3065 ( .A(n36), .B(n31), .Z(n32) );
  XNOR U3066 ( .A(n33), .B(n32), .Z(n57) );
  NANDN U3067 ( .A(n58), .B(n57), .Z(n34) );
  NAND U3068 ( .A(n62), .B(n34), .Z(n44) );
  XNOR U3069 ( .A(n36), .B(n35), .Z(n41) );
  ANDN U3070 ( .B(n37), .A(x[1]), .Z(n38) );
  XNOR U3071 ( .A(n39), .B(n38), .Z(n40) );
  XNOR U3072 ( .A(n41), .B(n40), .Z(n54) );
  XOR U3073 ( .A(n57), .B(n54), .Z(n42) );
  NAND U3074 ( .A(n58), .B(n42), .Z(n43) );
  NAND U3075 ( .A(n44), .B(n43), .Z(n1066) );
  ANDN U3076 ( .B(n45), .A(n1066), .Z(n69) );
  IV U3077 ( .A(n54), .Z(n60) );
  XOR U3078 ( .A(n62), .B(n58), .Z(n46) );
  NANDN U3079 ( .A(n60), .B(n46), .Z(n49) );
  NANDN U3080 ( .A(n58), .B(n60), .Z(n47) );
  NANDN U3081 ( .A(n57), .B(n47), .Z(n48) );
  NAND U3082 ( .A(n49), .B(n48), .Z(n1427) );
  XNOR U3083 ( .A(n1066), .B(n1427), .Z(n778) );
  AND U3084 ( .A(n50), .B(n778), .Z(n72) );
  OR U3085 ( .A(n57), .B(n54), .Z(n56) );
  ANDN U3086 ( .B(n57), .A(n51), .Z(n52) );
  XNOR U3087 ( .A(n52), .B(n62), .Z(n53) );
  NAND U3088 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3089 ( .A(n56), .B(n55), .Z(n775) );
  NAND U3090 ( .A(n58), .B(n62), .Z(n64) );
  NAND U3091 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U3092 ( .A(n60), .B(n59), .Z(n61) );
  NANDN U3093 ( .A(n62), .B(n61), .Z(n63) );
  NAND U3094 ( .A(n64), .B(n63), .Z(n1434) );
  NAND U3095 ( .A(n794), .B(n65), .Z(n66) );
  XNOR U3096 ( .A(n72), .B(n66), .Z(n1429) );
  XOR U3097 ( .A(n1066), .B(n1434), .Z(n1068) );
  AND U3098 ( .A(n67), .B(n1068), .Z(n789) );
  XNOR U3099 ( .A(n1429), .B(n789), .Z(n68) );
  XNOR U3100 ( .A(n69), .B(n68), .Z(n1437) );
  NAND U3101 ( .A(n780), .B(n70), .Z(n71) );
  XNOR U3102 ( .A(n72), .B(n71), .Z(n797) );
  AND U3103 ( .A(n73), .B(n782), .Z(n1428) );
  NANDN U3104 ( .A(n74), .B(n775), .Z(n75) );
  XNOR U3105 ( .A(n1428), .B(n75), .Z(n939) );
  XNOR U3106 ( .A(n797), .B(n939), .Z(n786) );
  XOR U3107 ( .A(n1437), .B(n786), .Z(z[0]) );
  XOR U3108 ( .A(x[99]), .B(x[97]), .Z(n76) );
  XNOR U3109 ( .A(n76), .B(x[98]), .Z(n77) );
  XNOR U3110 ( .A(x[101]), .B(n77), .Z(n114) );
  XOR U3111 ( .A(x[98]), .B(x[100]), .Z(n135) );
  XNOR U3112 ( .A(x[102]), .B(n77), .Z(n128) );
  XOR U3113 ( .A(x[103]), .B(x[100]), .Z(n133) );
  XOR U3114 ( .A(n76), .B(n133), .Z(n124) );
  XNOR U3115 ( .A(x[96]), .B(n124), .Z(n93) );
  IV U3116 ( .A(n93), .Z(n125) );
  XNOR U3117 ( .A(x[102]), .B(x[96]), .Z(n78) );
  XNOR U3118 ( .A(x[101]), .B(n78), .Z(n139) );
  XOR U3119 ( .A(n125), .B(n139), .Z(n127) );
  XOR U3120 ( .A(n128), .B(n127), .Z(n156) );
  AND U3121 ( .A(n135), .B(n156), .Z(n80) );
  AND U3122 ( .A(n128), .B(n133), .Z(n86) );
  IV U3123 ( .A(n139), .Z(n102) );
  XNOR U3124 ( .A(x[103]), .B(n102), .Z(n161) );
  XOR U3125 ( .A(n129), .B(n161), .Z(n84) );
  XNOR U3126 ( .A(n86), .B(n84), .Z(n79) );
  XNOR U3127 ( .A(n80), .B(n79), .Z(n103) );
  XOR U3128 ( .A(x[98]), .B(n161), .Z(n98) );
  XOR U3129 ( .A(x[97]), .B(n98), .Z(n150) );
  ANDN U3130 ( .B(x[96]), .A(n150), .Z(n82) );
  XNOR U3131 ( .A(x[100]), .B(n102), .Z(n170) );
  NANDN U3132 ( .A(n124), .B(n170), .Z(n81) );
  XNOR U3133 ( .A(n82), .B(n81), .Z(n83) );
  XOR U3134 ( .A(n103), .B(n83), .Z(n119) );
  XOR U3135 ( .A(x[97]), .B(x[103]), .Z(n138) );
  AND U3136 ( .A(n138), .B(n114), .Z(n104) );
  XOR U3137 ( .A(n84), .B(n104), .Z(n89) );
  XOR U3138 ( .A(x[98]), .B(x[103]), .Z(n162) );
  NAND U3139 ( .A(n162), .B(n127), .Z(n85) );
  XOR U3140 ( .A(n86), .B(n85), .Z(n99) );
  AND U3141 ( .A(n129), .B(n161), .Z(n87) );
  XOR U3142 ( .A(n99), .B(n87), .Z(n88) );
  XNOR U3143 ( .A(n89), .B(n88), .Z(n117) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n152) );
  AND U3145 ( .A(n124), .B(n152), .Z(n91) );
  AND U3146 ( .A(x[96]), .B(n170), .Z(n90) );
  XNOR U3147 ( .A(n91), .B(n90), .Z(n92) );
  NANDN U3148 ( .A(n93), .B(n92), .Z(n96) );
  NAND U3149 ( .A(n124), .B(x[96]), .Z(n94) );
  NANDN U3150 ( .A(n94), .B(n150), .Z(n95) );
  NAND U3151 ( .A(n96), .B(n95), .Z(n97) );
  XNOR U3152 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U3153 ( .A(n100), .B(n99), .Z(n116) );
  OR U3154 ( .A(n117), .B(n116), .Z(n101) );
  NANDN U3155 ( .A(n119), .B(n101), .Z(n109) );
  ANDN U3156 ( .B(n102), .A(x[97]), .Z(n106) );
  XNOR U3157 ( .A(n104), .B(n103), .Z(n105) );
  XNOR U3158 ( .A(n106), .B(n105), .Z(n121) );
  XOR U3159 ( .A(n117), .B(n121), .Z(n107) );
  NAND U3160 ( .A(n116), .B(n107), .Z(n108) );
  NAND U3161 ( .A(n109), .B(n108), .Z(n160) );
  OR U3162 ( .A(n119), .B(n116), .Z(n113) );
  ANDN U3163 ( .B(n116), .A(n117), .Z(n110) );
  XNOR U3164 ( .A(n110), .B(n121), .Z(n111) );
  NAND U3165 ( .A(n119), .B(n111), .Z(n112) );
  NAND U3166 ( .A(n113), .B(n112), .Z(n141) );
  XNOR U3167 ( .A(n160), .B(n141), .Z(n137) );
  AND U3168 ( .A(n114), .B(n137), .Z(n131) );
  NAND U3169 ( .A(n139), .B(n141), .Z(n115) );
  XNOR U3170 ( .A(n131), .B(n115), .Z(n172) );
  NANDN U3171 ( .A(n117), .B(n121), .Z(n123) );
  NANDN U3172 ( .A(n117), .B(n116), .Z(n118) );
  XOR U3173 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U3174 ( .A(n121), .B(n120), .Z(n122) );
  NAND U3175 ( .A(n123), .B(n122), .Z(n149) );
  XOR U3176 ( .A(n169), .B(n149), .Z(n151) );
  AND U3177 ( .A(n124), .B(n151), .Z(n144) );
  NANDN U3178 ( .A(n149), .B(n125), .Z(n126) );
  XNOR U3179 ( .A(n144), .B(n126), .Z(n159) );
  XNOR U3180 ( .A(n172), .B(n159), .Z(z[98]) );
  XNOR U3181 ( .A(n149), .B(n141), .Z(n163) );
  AND U3182 ( .A(n127), .B(n163), .Z(n183) );
  XOR U3183 ( .A(n169), .B(n160), .Z(n134) );
  AND U3184 ( .A(n128), .B(n134), .Z(n181) );
  NANDN U3185 ( .A(n160), .B(n129), .Z(n130) );
  XNOR U3186 ( .A(n131), .B(n130), .Z(n145) );
  XNOR U3187 ( .A(n181), .B(n145), .Z(n132) );
  XNOR U3188 ( .A(n183), .B(n132), .Z(n1958) );
  XOR U3189 ( .A(n1958), .B(z[98]), .Z(z[100]) );
  AND U3190 ( .A(n133), .B(n134), .Z(n165) );
  NAND U3191 ( .A(n157), .B(n135), .Z(n136) );
  XNOR U3192 ( .A(n165), .B(n136), .Z(n153) );
  AND U3193 ( .A(n138), .B(n137), .Z(n166) );
  XOR U3194 ( .A(x[97]), .B(n139), .Z(n140) );
  NAND U3195 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U3196 ( .A(n166), .B(n142), .Z(n147) );
  NANDN U3197 ( .A(n169), .B(x[96]), .Z(n143) );
  XNOR U3198 ( .A(n144), .B(n143), .Z(n180) );
  XNOR U3199 ( .A(n180), .B(n145), .Z(n146) );
  XNOR U3200 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U3201 ( .A(n153), .B(n148), .Z(z[101]) );
  ANDN U3202 ( .B(n150), .A(n149), .Z(n155) );
  AND U3203 ( .A(n152), .B(n151), .Z(n171) );
  XNOR U3204 ( .A(n171), .B(n153), .Z(n154) );
  XNOR U3205 ( .A(n155), .B(n154), .Z(n1959) );
  NAND U3206 ( .A(n157), .B(n156), .Z(n158) );
  XNOR U3207 ( .A(n181), .B(n158), .Z(n175) );
  XNOR U3208 ( .A(n175), .B(n159), .Z(n1957) );
  XNOR U3209 ( .A(n1959), .B(n1957), .Z(n179) );
  ANDN U3210 ( .B(n161), .A(n160), .Z(n168) );
  NAND U3211 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U3212 ( .A(n165), .B(n164), .Z(n176) );
  XNOR U3213 ( .A(n176), .B(n166), .Z(n167) );
  XNOR U3214 ( .A(n168), .B(n167), .Z(n1962) );
  XNOR U3215 ( .A(n179), .B(n1962), .Z(z[102]) );
  ANDN U3216 ( .B(n170), .A(n169), .Z(n174) );
  XNOR U3217 ( .A(n172), .B(n171), .Z(n173) );
  XNOR U3218 ( .A(n174), .B(n173), .Z(n178) );
  XNOR U3219 ( .A(n176), .B(n175), .Z(n177) );
  XNOR U3220 ( .A(n178), .B(n177), .Z(n1960) );
  XNOR U3221 ( .A(n1960), .B(n179), .Z(z[97]) );
  XNOR U3222 ( .A(n181), .B(n180), .Z(n182) );
  XNOR U3223 ( .A(n183), .B(n182), .Z(n184) );
  XOR U3224 ( .A(n184), .B(z[97]), .Z(z[103]) );
  XOR U3225 ( .A(x[107]), .B(x[105]), .Z(n187) );
  XNOR U3226 ( .A(x[104]), .B(x[110]), .Z(n186) );
  XOR U3227 ( .A(n186), .B(x[106]), .Z(n185) );
  XNOR U3228 ( .A(n187), .B(n185), .Z(n222) );
  XNOR U3229 ( .A(x[109]), .B(n186), .Z(n295) );
  XOR U3230 ( .A(n295), .B(x[108]), .Z(n265) );
  IV U3231 ( .A(n265), .Z(n196) );
  XNOR U3232 ( .A(x[111]), .B(x[108]), .Z(n190) );
  XNOR U3233 ( .A(n187), .B(n190), .Z(n250) );
  NOR U3234 ( .A(n196), .B(n250), .Z(n189) );
  XNOR U3235 ( .A(n295), .B(x[111]), .Z(n281) );
  XNOR U3236 ( .A(x[106]), .B(n281), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n205), .Z(n200) );
  AND U3238 ( .A(x[104]), .B(n200), .Z(n188) );
  XNOR U3239 ( .A(n189), .B(n188), .Z(n193) );
  XNOR U3240 ( .A(n222), .B(n281), .Z(n212) );
  IV U3241 ( .A(n222), .Z(n207) );
  XNOR U3242 ( .A(x[104]), .B(n207), .Z(n227) );
  IV U3243 ( .A(n190), .Z(n255) );
  AND U3244 ( .A(n227), .B(n255), .Z(n195) );
  IV U3245 ( .A(n295), .Z(n214) );
  XNOR U3246 ( .A(n222), .B(n214), .Z(n244) );
  XOR U3247 ( .A(n244), .B(n250), .Z(n247) );
  XOR U3248 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NAND U3249 ( .A(n247), .B(n257), .Z(n191) );
  XNOR U3250 ( .A(n195), .B(n191), .Z(n216) );
  XNOR U3251 ( .A(n212), .B(n216), .Z(n192) );
  XNOR U3252 ( .A(n193), .B(n192), .Z(n239) );
  XOR U3253 ( .A(x[106]), .B(x[111]), .Z(n271) );
  XNOR U3254 ( .A(x[104]), .B(n250), .Z(n251) );
  XNOR U3255 ( .A(n295), .B(n251), .Z(n242) );
  NAND U3256 ( .A(n271), .B(n242), .Z(n194) );
  XNOR U3257 ( .A(n195), .B(n194), .Z(n208) );
  IV U3258 ( .A(n200), .Z(n254) );
  XNOR U3259 ( .A(n254), .B(n196), .Z(n261) );
  AND U3260 ( .A(n250), .B(n261), .Z(n198) );
  AND U3261 ( .A(x[104]), .B(n265), .Z(n197) );
  XNOR U3262 ( .A(n198), .B(n197), .Z(n199) );
  NANDN U3263 ( .A(n251), .B(n199), .Z(n203) );
  NAND U3264 ( .A(x[104]), .B(n250), .Z(n201) );
  OR U3265 ( .A(n201), .B(n200), .Z(n202) );
  NAND U3266 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U3267 ( .A(n205), .B(n204), .Z(n206) );
  XNOR U3268 ( .A(n208), .B(n206), .Z(n228) );
  IV U3269 ( .A(n228), .Z(n235) );
  AND U3270 ( .A(n281), .B(n207), .Z(n210) );
  XOR U3271 ( .A(x[105]), .B(x[111]), .Z(n283) );
  AND U3272 ( .A(n244), .B(n283), .Z(n213) );
  XNOR U3273 ( .A(n213), .B(n208), .Z(n209) );
  XNOR U3274 ( .A(n210), .B(n209), .Z(n234) );
  NANDN U3275 ( .A(n235), .B(n234), .Z(n211) );
  NAND U3276 ( .A(n239), .B(n211), .Z(n221) );
  XNOR U3277 ( .A(n213), .B(n212), .Z(n218) );
  ANDN U3278 ( .B(n214), .A(x[105]), .Z(n215) );
  XNOR U3279 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3280 ( .A(n218), .B(n217), .Z(n231) );
  XOR U3281 ( .A(n234), .B(n231), .Z(n219) );
  NAND U3282 ( .A(n235), .B(n219), .Z(n220) );
  NAND U3283 ( .A(n221), .B(n220), .Z(n280) );
  ANDN U3284 ( .B(n222), .A(n280), .Z(n246) );
  IV U3285 ( .A(n231), .Z(n237) );
  XOR U3286 ( .A(n239), .B(n235), .Z(n223) );
  NANDN U3287 ( .A(n237), .B(n223), .Z(n226) );
  NANDN U3288 ( .A(n235), .B(n237), .Z(n224) );
  NANDN U3289 ( .A(n234), .B(n224), .Z(n225) );
  NAND U3290 ( .A(n226), .B(n225), .Z(n290) );
  XNOR U3291 ( .A(n280), .B(n290), .Z(n256) );
  AND U3292 ( .A(n227), .B(n256), .Z(n249) );
  OR U3293 ( .A(n234), .B(n231), .Z(n233) );
  ANDN U3294 ( .B(n234), .A(n228), .Z(n229) );
  XNOR U3295 ( .A(n229), .B(n239), .Z(n230) );
  NAND U3296 ( .A(n231), .B(n230), .Z(n232) );
  NAND U3297 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3298 ( .A(n235), .B(n239), .Z(n241) );
  NAND U3299 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U3300 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U3301 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3302 ( .A(n241), .B(n240), .Z(n297) );
  NAND U3303 ( .A(n272), .B(n242), .Z(n243) );
  XNOR U3304 ( .A(n249), .B(n243), .Z(n292) );
  XOR U3305 ( .A(n280), .B(n297), .Z(n282) );
  AND U3306 ( .A(n244), .B(n282), .Z(n267) );
  XNOR U3307 ( .A(n292), .B(n267), .Z(n245) );
  XNOR U3308 ( .A(n246), .B(n245), .Z(n300) );
  NAND U3309 ( .A(n258), .B(n247), .Z(n248) );
  XNOR U3310 ( .A(n249), .B(n248), .Z(n275) );
  AND U3311 ( .A(n250), .B(n260), .Z(n291) );
  NANDN U3312 ( .A(n251), .B(n253), .Z(n252) );
  XNOR U3313 ( .A(n291), .B(n252), .Z(n279) );
  XNOR U3314 ( .A(n275), .B(n279), .Z(n264) );
  XOR U3315 ( .A(n300), .B(n264), .Z(z[104]) );
  AND U3316 ( .A(n254), .B(n253), .Z(n263) );
  AND U3317 ( .A(n256), .B(n255), .Z(n274) );
  NAND U3318 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3319 ( .A(n274), .B(n259), .Z(n301) );
  AND U3320 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3321 ( .A(n301), .B(n268), .Z(n262) );
  XNOR U3322 ( .A(n263), .B(n262), .Z(n288) );
  XNOR U3323 ( .A(n288), .B(n264), .Z(n360) );
  AND U3324 ( .A(n265), .B(n290), .Z(n270) );
  NANDN U3325 ( .A(n297), .B(n295), .Z(n266) );
  XNOR U3326 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3327 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3328 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3329 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3330 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3331 ( .A(n275), .B(n284), .Z(n276) );
  XNOR U3332 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3333 ( .A(n360), .B(n287), .Z(z[105]) );
  XNOR U3334 ( .A(n279), .B(n278), .Z(z[106]) );
  NOR U3335 ( .A(n281), .B(n280), .Z(n286) );
  AND U3336 ( .A(n283), .B(n282), .Z(n299) );
  XNOR U3337 ( .A(n284), .B(n299), .Z(n285) );
  XNOR U3338 ( .A(n286), .B(n285), .Z(n359) );
  XOR U3339 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U3340 ( .A(n359), .B(n289), .Z(z[107]) );
  XOR U3341 ( .A(n300), .B(z[106]), .Z(z[108]) );
  AND U3342 ( .A(x[104]), .B(n290), .Z(n294) );
  XNOR U3343 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U3344 ( .A(n294), .B(n293), .Z(n361) );
  XOR U3345 ( .A(n295), .B(x[105]), .Z(n296) );
  NANDN U3346 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U3347 ( .A(n299), .B(n298), .Z(n303) );
  XNOR U3348 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U3349 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U3350 ( .A(n361), .B(n304), .Z(z[109]) );
  XOR U3351 ( .A(x[9]), .B(x[11]), .Z(n305) );
  XOR U3352 ( .A(x[15]), .B(x[12]), .Z(n486) );
  XOR U3353 ( .A(n305), .B(n486), .Z(n341) );
  XNOR U3354 ( .A(x[8]), .B(x[14]), .Z(n307) );
  XNOR U3355 ( .A(x[13]), .B(n307), .Z(n654) );
  XNOR U3356 ( .A(x[15]), .B(n654), .Z(n485) );
  XNOR U3357 ( .A(n305), .B(x[10]), .Z(n306) );
  XNOR U3358 ( .A(n307), .B(n306), .Z(n308) );
  AND U3359 ( .A(n485), .B(n308), .Z(n311) );
  IV U3360 ( .A(n308), .Z(n641) );
  XOR U3361 ( .A(n641), .B(n654), .Z(n357) );
  XOR U3362 ( .A(x[9]), .B(x[15]), .Z(n491) );
  AND U3363 ( .A(n357), .B(n491), .Z(n312) );
  XNOR U3364 ( .A(x[8]), .B(n308), .Z(n509) );
  AND U3365 ( .A(n486), .B(n509), .Z(n314) );
  XOR U3366 ( .A(x[15]), .B(x[10]), .Z(n488) );
  XNOR U3367 ( .A(n341), .B(x[8]), .Z(n342) );
  XNOR U3368 ( .A(n654), .B(n342), .Z(n642) );
  NAND U3369 ( .A(n488), .B(n642), .Z(n309) );
  XNOR U3370 ( .A(n314), .B(n309), .Z(n325) );
  XNOR U3371 ( .A(n312), .B(n325), .Z(n310) );
  XNOR U3372 ( .A(n311), .B(n310), .Z(n349) );
  XNOR U3373 ( .A(n641), .B(n485), .Z(n329) );
  XOR U3374 ( .A(x[12]), .B(x[10]), .Z(n496) );
  XOR U3375 ( .A(n341), .B(n357), .Z(n510) );
  NAND U3376 ( .A(n496), .B(n510), .Z(n313) );
  XNOR U3377 ( .A(n314), .B(n313), .Z(n328) );
  OR U3378 ( .A(n349), .B(n345), .Z(n335) );
  XNOR U3379 ( .A(x[10]), .B(n485), .Z(n323) );
  IV U3380 ( .A(n318), .Z(n495) );
  XNOR U3381 ( .A(x[12]), .B(n654), .Z(n503) );
  XNOR U3382 ( .A(n495), .B(n503), .Z(n500) );
  AND U3383 ( .A(n341), .B(n500), .Z(n316) );
  ANDN U3384 ( .B(x[8]), .A(n503), .Z(n315) );
  XNOR U3385 ( .A(n316), .B(n315), .Z(n317) );
  NANDN U3386 ( .A(n342), .B(n317), .Z(n321) );
  NAND U3387 ( .A(n341), .B(x[8]), .Z(n319) );
  OR U3388 ( .A(n319), .B(n318), .Z(n320) );
  NAND U3389 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U3390 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U3391 ( .A(n325), .B(n324), .Z(n336) );
  ANDN U3392 ( .B(n349), .A(n336), .Z(n332) );
  NOR U3393 ( .A(n503), .B(n341), .Z(n327) );
  ANDN U3394 ( .B(x[8]), .A(n495), .Z(n326) );
  XNOR U3395 ( .A(n327), .B(n326), .Z(n331) );
  XNOR U3396 ( .A(n329), .B(n328), .Z(n330) );
  XNOR U3397 ( .A(n331), .B(n330), .Z(n354) );
  XNOR U3398 ( .A(n332), .B(n354), .Z(n333) );
  NAND U3399 ( .A(n345), .B(n333), .Z(n334) );
  NAND U3400 ( .A(n335), .B(n334), .Z(n494) );
  IV U3401 ( .A(n494), .Z(n487) );
  IV U3402 ( .A(n345), .Z(n352) );
  IV U3403 ( .A(n336), .Z(n350) );
  XOR U3404 ( .A(n354), .B(n350), .Z(n337) );
  NANDN U3405 ( .A(n352), .B(n337), .Z(n340) );
  NANDN U3406 ( .A(n350), .B(n352), .Z(n338) );
  NANDN U3407 ( .A(n349), .B(n338), .Z(n339) );
  NAND U3408 ( .A(n340), .B(n339), .Z(n649) );
  XNOR U3409 ( .A(n487), .B(n649), .Z(n499) );
  AND U3410 ( .A(n341), .B(n499), .Z(n651) );
  NANDN U3411 ( .A(n342), .B(n494), .Z(n343) );
  XNOR U3412 ( .A(n651), .B(n343), .Z(n663) );
  NANDN U3413 ( .A(n350), .B(n349), .Z(n344) );
  NAND U3414 ( .A(n354), .B(n344), .Z(n348) );
  XOR U3415 ( .A(n349), .B(n345), .Z(n346) );
  NAND U3416 ( .A(n350), .B(n346), .Z(n347) );
  NAND U3417 ( .A(n348), .B(n347), .Z(n640) );
  NAND U3418 ( .A(n350), .B(n354), .Z(n356) );
  NAND U3419 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U3420 ( .A(n352), .B(n351), .Z(n353) );
  NANDN U3421 ( .A(n354), .B(n353), .Z(n355) );
  NAND U3422 ( .A(n356), .B(n355), .Z(n656) );
  XOR U3423 ( .A(n640), .B(n656), .Z(n490) );
  AND U3424 ( .A(n357), .B(n490), .Z(n646) );
  NANDN U3425 ( .A(n656), .B(n654), .Z(n358) );
  XNOR U3426 ( .A(n646), .B(n358), .Z(n513) );
  XNOR U3427 ( .A(n663), .B(n513), .Z(z[10]) );
  XNOR U3428 ( .A(n360), .B(n359), .Z(z[110]) );
  XOR U3429 ( .A(n361), .B(z[105]), .Z(z[111]) );
  XOR U3430 ( .A(x[115]), .B(x[113]), .Z(n364) );
  XNOR U3431 ( .A(x[112]), .B(x[118]), .Z(n363) );
  XOR U3432 ( .A(n363), .B(x[114]), .Z(n362) );
  XNOR U3433 ( .A(n364), .B(n362), .Z(n399) );
  XNOR U3434 ( .A(x[117]), .B(n363), .Z(n472) );
  XOR U3435 ( .A(n472), .B(x[116]), .Z(n442) );
  IV U3436 ( .A(n442), .Z(n373) );
  XNOR U3437 ( .A(x[119]), .B(x[116]), .Z(n367) );
  XNOR U3438 ( .A(n364), .B(n367), .Z(n427) );
  NOR U3439 ( .A(n373), .B(n427), .Z(n366) );
  XNOR U3440 ( .A(n472), .B(x[119]), .Z(n458) );
  XNOR U3441 ( .A(x[114]), .B(n458), .Z(n382) );
  XNOR U3442 ( .A(x[113]), .B(n382), .Z(n377) );
  AND U3443 ( .A(x[112]), .B(n377), .Z(n365) );
  XNOR U3444 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U3445 ( .A(n399), .B(n458), .Z(n389) );
  IV U3446 ( .A(n399), .Z(n384) );
  XNOR U3447 ( .A(x[112]), .B(n384), .Z(n404) );
  IV U3448 ( .A(n367), .Z(n432) );
  AND U3449 ( .A(n404), .B(n432), .Z(n372) );
  IV U3450 ( .A(n472), .Z(n391) );
  XNOR U3451 ( .A(n399), .B(n391), .Z(n421) );
  XOR U3452 ( .A(n421), .B(n427), .Z(n424) );
  XOR U3453 ( .A(x[114]), .B(x[116]), .Z(n434) );
  NAND U3454 ( .A(n424), .B(n434), .Z(n368) );
  XNOR U3455 ( .A(n372), .B(n368), .Z(n393) );
  XNOR U3456 ( .A(n389), .B(n393), .Z(n369) );
  XNOR U3457 ( .A(n370), .B(n369), .Z(n416) );
  XOR U3458 ( .A(x[114]), .B(x[119]), .Z(n448) );
  XNOR U3459 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3460 ( .A(n472), .B(n428), .Z(n419) );
  NAND U3461 ( .A(n448), .B(n419), .Z(n371) );
  XNOR U3462 ( .A(n372), .B(n371), .Z(n385) );
  IV U3463 ( .A(n377), .Z(n431) );
  XNOR U3464 ( .A(n431), .B(n373), .Z(n438) );
  AND U3465 ( .A(n427), .B(n438), .Z(n375) );
  AND U3466 ( .A(x[112]), .B(n442), .Z(n374) );
  XNOR U3467 ( .A(n375), .B(n374), .Z(n376) );
  NANDN U3468 ( .A(n428), .B(n376), .Z(n380) );
  NAND U3469 ( .A(x[112]), .B(n427), .Z(n378) );
  OR U3470 ( .A(n378), .B(n377), .Z(n379) );
  NAND U3471 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U3472 ( .A(n382), .B(n381), .Z(n383) );
  XNOR U3473 ( .A(n385), .B(n383), .Z(n405) );
  IV U3474 ( .A(n405), .Z(n412) );
  AND U3475 ( .A(n458), .B(n384), .Z(n387) );
  XOR U3476 ( .A(x[113]), .B(x[119]), .Z(n460) );
  AND U3477 ( .A(n421), .B(n460), .Z(n390) );
  XNOR U3478 ( .A(n390), .B(n385), .Z(n386) );
  XNOR U3479 ( .A(n387), .B(n386), .Z(n411) );
  NANDN U3480 ( .A(n412), .B(n411), .Z(n388) );
  NAND U3481 ( .A(n416), .B(n388), .Z(n398) );
  XNOR U3482 ( .A(n390), .B(n389), .Z(n395) );
  ANDN U3483 ( .B(n391), .A(x[113]), .Z(n392) );
  XNOR U3484 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U3485 ( .A(n395), .B(n394), .Z(n408) );
  XOR U3486 ( .A(n411), .B(n408), .Z(n396) );
  NAND U3487 ( .A(n412), .B(n396), .Z(n397) );
  NAND U3488 ( .A(n398), .B(n397), .Z(n457) );
  ANDN U3489 ( .B(n399), .A(n457), .Z(n423) );
  IV U3490 ( .A(n408), .Z(n414) );
  XOR U3491 ( .A(n416), .B(n412), .Z(n400) );
  NANDN U3492 ( .A(n414), .B(n400), .Z(n403) );
  NANDN U3493 ( .A(n412), .B(n414), .Z(n401) );
  NANDN U3494 ( .A(n411), .B(n401), .Z(n402) );
  NAND U3495 ( .A(n403), .B(n402), .Z(n467) );
  XNOR U3496 ( .A(n457), .B(n467), .Z(n433) );
  AND U3497 ( .A(n404), .B(n433), .Z(n426) );
  OR U3498 ( .A(n411), .B(n408), .Z(n410) );
  ANDN U3499 ( .B(n411), .A(n405), .Z(n406) );
  XNOR U3500 ( .A(n406), .B(n416), .Z(n407) );
  NAND U3501 ( .A(n408), .B(n407), .Z(n409) );
  NAND U3502 ( .A(n410), .B(n409), .Z(n430) );
  NAND U3503 ( .A(n412), .B(n416), .Z(n418) );
  NAND U3504 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U3505 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U3506 ( .A(n416), .B(n415), .Z(n417) );
  NAND U3507 ( .A(n418), .B(n417), .Z(n474) );
  NAND U3508 ( .A(n449), .B(n419), .Z(n420) );
  XNOR U3509 ( .A(n426), .B(n420), .Z(n469) );
  XOR U3510 ( .A(n457), .B(n474), .Z(n459) );
  AND U3511 ( .A(n421), .B(n459), .Z(n444) );
  XNOR U3512 ( .A(n469), .B(n444), .Z(n422) );
  XNOR U3513 ( .A(n423), .B(n422), .Z(n477) );
  NAND U3514 ( .A(n435), .B(n424), .Z(n425) );
  XNOR U3515 ( .A(n426), .B(n425), .Z(n452) );
  AND U3516 ( .A(n427), .B(n437), .Z(n468) );
  NANDN U3517 ( .A(n428), .B(n430), .Z(n429) );
  XNOR U3518 ( .A(n468), .B(n429), .Z(n456) );
  XNOR U3519 ( .A(n452), .B(n456), .Z(n441) );
  XOR U3520 ( .A(n477), .B(n441), .Z(z[112]) );
  AND U3521 ( .A(n431), .B(n430), .Z(n440) );
  AND U3522 ( .A(n433), .B(n432), .Z(n451) );
  NAND U3523 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U3524 ( .A(n451), .B(n436), .Z(n478) );
  AND U3525 ( .A(n438), .B(n437), .Z(n445) );
  XNOR U3526 ( .A(n478), .B(n445), .Z(n439) );
  XNOR U3527 ( .A(n440), .B(n439), .Z(n465) );
  XNOR U3528 ( .A(n465), .B(n441), .Z(n483) );
  AND U3529 ( .A(n442), .B(n467), .Z(n447) );
  NANDN U3530 ( .A(n474), .B(n472), .Z(n443) );
  XNOR U3531 ( .A(n444), .B(n443), .Z(n455) );
  XNOR U3532 ( .A(n445), .B(n455), .Z(n446) );
  XNOR U3533 ( .A(n447), .B(n446), .Z(n454) );
  NAND U3534 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U3535 ( .A(n451), .B(n450), .Z(n461) );
  XNOR U3536 ( .A(n452), .B(n461), .Z(n453) );
  XNOR U3537 ( .A(n454), .B(n453), .Z(n464) );
  XNOR U3538 ( .A(n483), .B(n464), .Z(z[113]) );
  XNOR U3539 ( .A(n456), .B(n455), .Z(z[114]) );
  NOR U3540 ( .A(n458), .B(n457), .Z(n463) );
  AND U3541 ( .A(n460), .B(n459), .Z(n476) );
  XNOR U3542 ( .A(n461), .B(n476), .Z(n462) );
  XNOR U3543 ( .A(n463), .B(n462), .Z(n482) );
  XOR U3544 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U3545 ( .A(n482), .B(n466), .Z(z[115]) );
  XOR U3546 ( .A(n477), .B(z[114]), .Z(z[116]) );
  AND U3547 ( .A(x[112]), .B(n467), .Z(n471) );
  XNOR U3548 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U3549 ( .A(n471), .B(n470), .Z(n484) );
  XOR U3550 ( .A(n472), .B(x[113]), .Z(n473) );
  NANDN U3551 ( .A(n474), .B(n473), .Z(n475) );
  XNOR U3552 ( .A(n476), .B(n475), .Z(n480) );
  XNOR U3553 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U3554 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U3555 ( .A(n484), .B(n481), .Z(z[117]) );
  XNOR U3556 ( .A(n483), .B(n482), .Z(z[118]) );
  XOR U3557 ( .A(n484), .B(z[113]), .Z(z[119]) );
  NOR U3558 ( .A(n485), .B(n640), .Z(n493) );
  XNOR U3559 ( .A(n640), .B(n649), .Z(n508) );
  AND U3560 ( .A(n486), .B(n508), .Z(n498) );
  XOR U3561 ( .A(n487), .B(n656), .Z(n643) );
  NAND U3562 ( .A(n643), .B(n488), .Z(n489) );
  XNOR U3563 ( .A(n498), .B(n489), .Z(n504) );
  AND U3564 ( .A(n491), .B(n490), .Z(n658) );
  XNOR U3565 ( .A(n504), .B(n658), .Z(n492) );
  XNOR U3566 ( .A(n493), .B(n492), .Z(n666) );
  AND U3567 ( .A(n495), .B(n494), .Z(n502) );
  NAND U3568 ( .A(n511), .B(n496), .Z(n497) );
  XNOR U3569 ( .A(n498), .B(n497), .Z(n659) );
  AND U3570 ( .A(n500), .B(n499), .Z(n505) );
  XNOR U3571 ( .A(n659), .B(n505), .Z(n501) );
  XNOR U3572 ( .A(n502), .B(n501), .Z(n665) );
  ANDN U3573 ( .B(n649), .A(n503), .Z(n507) );
  XNOR U3574 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U3575 ( .A(n507), .B(n506), .Z(n515) );
  AND U3576 ( .A(n509), .B(n508), .Z(n645) );
  NAND U3577 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U3578 ( .A(n645), .B(n512), .Z(n664) );
  XNOR U3579 ( .A(n664), .B(n513), .Z(n514) );
  XNOR U3580 ( .A(n515), .B(n514), .Z(n667) );
  XOR U3581 ( .A(n665), .B(n667), .Z(n516) );
  XNOR U3582 ( .A(n666), .B(n516), .Z(z[11]) );
  XOR U3583 ( .A(x[123]), .B(x[121]), .Z(n519) );
  XNOR U3584 ( .A(x[120]), .B(x[126]), .Z(n518) );
  XOR U3585 ( .A(n518), .B(x[122]), .Z(n517) );
  XNOR U3586 ( .A(n519), .B(n517), .Z(n554) );
  XNOR U3587 ( .A(x[125]), .B(n518), .Z(n627) );
  XOR U3588 ( .A(n627), .B(x[124]), .Z(n597) );
  IV U3589 ( .A(n597), .Z(n528) );
  XNOR U3590 ( .A(x[127]), .B(x[124]), .Z(n522) );
  XNOR U3591 ( .A(n519), .B(n522), .Z(n582) );
  NOR U3592 ( .A(n528), .B(n582), .Z(n521) );
  XNOR U3593 ( .A(n627), .B(x[127]), .Z(n613) );
  XNOR U3594 ( .A(x[122]), .B(n613), .Z(n537) );
  XNOR U3595 ( .A(x[121]), .B(n537), .Z(n532) );
  AND U3596 ( .A(x[120]), .B(n532), .Z(n520) );
  XNOR U3597 ( .A(n521), .B(n520), .Z(n525) );
  XNOR U3598 ( .A(n554), .B(n613), .Z(n544) );
  IV U3599 ( .A(n554), .Z(n539) );
  XNOR U3600 ( .A(x[120]), .B(n539), .Z(n559) );
  IV U3601 ( .A(n522), .Z(n587) );
  AND U3602 ( .A(n559), .B(n587), .Z(n527) );
  IV U3603 ( .A(n627), .Z(n546) );
  XNOR U3604 ( .A(n554), .B(n546), .Z(n576) );
  XOR U3605 ( .A(n576), .B(n582), .Z(n579) );
  XOR U3606 ( .A(x[122]), .B(x[124]), .Z(n589) );
  NAND U3607 ( .A(n579), .B(n589), .Z(n523) );
  XNOR U3608 ( .A(n527), .B(n523), .Z(n548) );
  XNOR U3609 ( .A(n544), .B(n548), .Z(n524) );
  XNOR U3610 ( .A(n525), .B(n524), .Z(n571) );
  XOR U3611 ( .A(x[122]), .B(x[127]), .Z(n603) );
  XNOR U3612 ( .A(x[120]), .B(n582), .Z(n583) );
  XNOR U3613 ( .A(n627), .B(n583), .Z(n574) );
  NAND U3614 ( .A(n603), .B(n574), .Z(n526) );
  XNOR U3615 ( .A(n527), .B(n526), .Z(n540) );
  IV U3616 ( .A(n532), .Z(n586) );
  XNOR U3617 ( .A(n586), .B(n528), .Z(n593) );
  AND U3618 ( .A(n582), .B(n593), .Z(n530) );
  AND U3619 ( .A(x[120]), .B(n597), .Z(n529) );
  XNOR U3620 ( .A(n530), .B(n529), .Z(n531) );
  NANDN U3621 ( .A(n583), .B(n531), .Z(n535) );
  NAND U3622 ( .A(x[120]), .B(n582), .Z(n533) );
  OR U3623 ( .A(n533), .B(n532), .Z(n534) );
  NAND U3624 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U3625 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U3626 ( .A(n540), .B(n538), .Z(n560) );
  IV U3627 ( .A(n560), .Z(n567) );
  AND U3628 ( .A(n613), .B(n539), .Z(n542) );
  XOR U3629 ( .A(x[121]), .B(x[127]), .Z(n615) );
  AND U3630 ( .A(n576), .B(n615), .Z(n545) );
  XNOR U3631 ( .A(n545), .B(n540), .Z(n541) );
  XNOR U3632 ( .A(n542), .B(n541), .Z(n566) );
  NANDN U3633 ( .A(n567), .B(n566), .Z(n543) );
  NAND U3634 ( .A(n571), .B(n543), .Z(n553) );
  XNOR U3635 ( .A(n545), .B(n544), .Z(n550) );
  ANDN U3636 ( .B(n546), .A(x[121]), .Z(n547) );
  XNOR U3637 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U3638 ( .A(n550), .B(n549), .Z(n563) );
  XOR U3639 ( .A(n566), .B(n563), .Z(n551) );
  NAND U3640 ( .A(n567), .B(n551), .Z(n552) );
  NAND U3641 ( .A(n553), .B(n552), .Z(n612) );
  ANDN U3642 ( .B(n554), .A(n612), .Z(n578) );
  IV U3643 ( .A(n563), .Z(n569) );
  XOR U3644 ( .A(n571), .B(n567), .Z(n555) );
  NANDN U3645 ( .A(n569), .B(n555), .Z(n558) );
  NANDN U3646 ( .A(n567), .B(n569), .Z(n556) );
  NANDN U3647 ( .A(n566), .B(n556), .Z(n557) );
  NAND U3648 ( .A(n558), .B(n557), .Z(n622) );
  XNOR U3649 ( .A(n612), .B(n622), .Z(n588) );
  AND U3650 ( .A(n559), .B(n588), .Z(n581) );
  OR U3651 ( .A(n566), .B(n563), .Z(n565) );
  ANDN U3652 ( .B(n566), .A(n560), .Z(n561) );
  XNOR U3653 ( .A(n561), .B(n571), .Z(n562) );
  NAND U3654 ( .A(n563), .B(n562), .Z(n564) );
  NAND U3655 ( .A(n565), .B(n564), .Z(n585) );
  NAND U3656 ( .A(n567), .B(n571), .Z(n573) );
  NAND U3657 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U3658 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U3659 ( .A(n571), .B(n570), .Z(n572) );
  NAND U3660 ( .A(n573), .B(n572), .Z(n629) );
  NAND U3661 ( .A(n604), .B(n574), .Z(n575) );
  XNOR U3662 ( .A(n581), .B(n575), .Z(n624) );
  XOR U3663 ( .A(n612), .B(n629), .Z(n614) );
  AND U3664 ( .A(n576), .B(n614), .Z(n599) );
  XNOR U3665 ( .A(n624), .B(n599), .Z(n577) );
  XNOR U3666 ( .A(n578), .B(n577), .Z(n632) );
  NAND U3667 ( .A(n590), .B(n579), .Z(n580) );
  XNOR U3668 ( .A(n581), .B(n580), .Z(n607) );
  AND U3669 ( .A(n582), .B(n592), .Z(n623) );
  NANDN U3670 ( .A(n583), .B(n585), .Z(n584) );
  XNOR U3671 ( .A(n623), .B(n584), .Z(n611) );
  XNOR U3672 ( .A(n607), .B(n611), .Z(n596) );
  XOR U3673 ( .A(n632), .B(n596), .Z(z[120]) );
  AND U3674 ( .A(n586), .B(n585), .Z(n595) );
  AND U3675 ( .A(n588), .B(n587), .Z(n606) );
  NAND U3676 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U3677 ( .A(n606), .B(n591), .Z(n633) );
  AND U3678 ( .A(n593), .B(n592), .Z(n600) );
  XNOR U3679 ( .A(n633), .B(n600), .Z(n594) );
  XNOR U3680 ( .A(n595), .B(n594), .Z(n620) );
  XNOR U3681 ( .A(n620), .B(n596), .Z(n638) );
  AND U3682 ( .A(n597), .B(n622), .Z(n602) );
  NANDN U3683 ( .A(n629), .B(n627), .Z(n598) );
  XNOR U3684 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U3685 ( .A(n600), .B(n610), .Z(n601) );
  XNOR U3686 ( .A(n602), .B(n601), .Z(n609) );
  NAND U3687 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U3688 ( .A(n606), .B(n605), .Z(n616) );
  XNOR U3689 ( .A(n607), .B(n616), .Z(n608) );
  XNOR U3690 ( .A(n609), .B(n608), .Z(n619) );
  XNOR U3691 ( .A(n638), .B(n619), .Z(z[121]) );
  XNOR U3692 ( .A(n611), .B(n610), .Z(z[122]) );
  NOR U3693 ( .A(n613), .B(n612), .Z(n618) );
  AND U3694 ( .A(n615), .B(n614), .Z(n631) );
  XNOR U3695 ( .A(n616), .B(n631), .Z(n617) );
  XNOR U3696 ( .A(n618), .B(n617), .Z(n637) );
  XOR U3697 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U3698 ( .A(n637), .B(n621), .Z(z[123]) );
  XOR U3699 ( .A(n632), .B(z[122]), .Z(z[124]) );
  AND U3700 ( .A(x[120]), .B(n622), .Z(n626) );
  XNOR U3701 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U3702 ( .A(n626), .B(n625), .Z(n639) );
  XOR U3703 ( .A(n627), .B(x[121]), .Z(n628) );
  NANDN U3704 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U3705 ( .A(n631), .B(n630), .Z(n635) );
  XNOR U3706 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U3707 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U3708 ( .A(n639), .B(n636), .Z(z[125]) );
  XNOR U3709 ( .A(n638), .B(n637), .Z(z[126]) );
  XOR U3710 ( .A(n639), .B(z[121]), .Z(z[127]) );
  ANDN U3711 ( .B(n641), .A(n640), .Z(n648) );
  NAND U3712 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U3713 ( .A(n645), .B(n644), .Z(n650) );
  XNOR U3714 ( .A(n650), .B(n646), .Z(n647) );
  XNOR U3715 ( .A(n648), .B(n647), .Z(n1926) );
  XOR U3716 ( .A(n1926), .B(z[10]), .Z(z[12]) );
  AND U3717 ( .A(x[8]), .B(n649), .Z(n653) );
  XNOR U3718 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U3719 ( .A(n653), .B(n652), .Z(n669) );
  XOR U3720 ( .A(n654), .B(x[9]), .Z(n655) );
  NANDN U3721 ( .A(n656), .B(n655), .Z(n657) );
  XNOR U3722 ( .A(n658), .B(n657), .Z(n661) );
  XNOR U3723 ( .A(n659), .B(n1926), .Z(n660) );
  XNOR U3724 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U3725 ( .A(n669), .B(n662), .Z(z[13]) );
  XNOR U3726 ( .A(n664), .B(n663), .Z(n1925) );
  XNOR U3727 ( .A(n665), .B(n1925), .Z(n668) );
  XNOR U3728 ( .A(n668), .B(n666), .Z(z[14]) );
  XNOR U3729 ( .A(n668), .B(n667), .Z(z[9]) );
  XOR U3730 ( .A(n669), .B(z[9]), .Z(z[15]) );
  XOR U3731 ( .A(x[19]), .B(x[17]), .Z(n672) );
  XNOR U3732 ( .A(x[16]), .B(x[22]), .Z(n671) );
  XOR U3733 ( .A(n671), .B(x[18]), .Z(n670) );
  XNOR U3734 ( .A(n672), .B(n670), .Z(n707) );
  XNOR U3735 ( .A(x[21]), .B(n671), .Z(n805) );
  XOR U3736 ( .A(n805), .B(x[20]), .Z(n750) );
  IV U3737 ( .A(n750), .Z(n681) );
  XNOR U3738 ( .A(x[23]), .B(x[20]), .Z(n675) );
  XNOR U3739 ( .A(n672), .B(n675), .Z(n735) );
  NOR U3740 ( .A(n681), .B(n735), .Z(n674) );
  XNOR U3741 ( .A(n805), .B(x[23]), .Z(n766) );
  XNOR U3742 ( .A(x[18]), .B(n766), .Z(n690) );
  XNOR U3743 ( .A(x[17]), .B(n690), .Z(n685) );
  AND U3744 ( .A(x[16]), .B(n685), .Z(n673) );
  XNOR U3745 ( .A(n674), .B(n673), .Z(n678) );
  XNOR U3746 ( .A(n707), .B(n766), .Z(n697) );
  IV U3747 ( .A(n707), .Z(n692) );
  XNOR U3748 ( .A(x[16]), .B(n692), .Z(n712) );
  IV U3749 ( .A(n675), .Z(n740) );
  AND U3750 ( .A(n712), .B(n740), .Z(n680) );
  IV U3751 ( .A(n805), .Z(n699) );
  XNOR U3752 ( .A(n707), .B(n699), .Z(n729) );
  XOR U3753 ( .A(n729), .B(n735), .Z(n732) );
  XOR U3754 ( .A(x[18]), .B(x[20]), .Z(n742) );
  NAND U3755 ( .A(n732), .B(n742), .Z(n676) );
  XNOR U3756 ( .A(n680), .B(n676), .Z(n701) );
  XNOR U3757 ( .A(n697), .B(n701), .Z(n677) );
  XNOR U3758 ( .A(n678), .B(n677), .Z(n724) );
  XOR U3759 ( .A(x[18]), .B(x[23]), .Z(n756) );
  XNOR U3760 ( .A(x[16]), .B(n735), .Z(n736) );
  XNOR U3761 ( .A(n805), .B(n736), .Z(n727) );
  NAND U3762 ( .A(n756), .B(n727), .Z(n679) );
  XNOR U3763 ( .A(n680), .B(n679), .Z(n693) );
  IV U3764 ( .A(n685), .Z(n739) );
  XNOR U3765 ( .A(n739), .B(n681), .Z(n746) );
  AND U3766 ( .A(n735), .B(n746), .Z(n683) );
  AND U3767 ( .A(x[16]), .B(n750), .Z(n682) );
  XNOR U3768 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U3769 ( .A(n736), .B(n684), .Z(n688) );
  NAND U3770 ( .A(x[16]), .B(n735), .Z(n686) );
  OR U3771 ( .A(n686), .B(n685), .Z(n687) );
  NAND U3772 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U3773 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U3774 ( .A(n693), .B(n691), .Z(n713) );
  IV U3775 ( .A(n713), .Z(n720) );
  AND U3776 ( .A(n766), .B(n692), .Z(n695) );
  XOR U3777 ( .A(x[17]), .B(x[23]), .Z(n768) );
  AND U3778 ( .A(n729), .B(n768), .Z(n698) );
  XNOR U3779 ( .A(n698), .B(n693), .Z(n694) );
  XNOR U3780 ( .A(n695), .B(n694), .Z(n719) );
  NANDN U3781 ( .A(n720), .B(n719), .Z(n696) );
  NAND U3782 ( .A(n724), .B(n696), .Z(n706) );
  XNOR U3783 ( .A(n698), .B(n697), .Z(n703) );
  ANDN U3784 ( .B(n699), .A(x[17]), .Z(n700) );
  XNOR U3785 ( .A(n701), .B(n700), .Z(n702) );
  XNOR U3786 ( .A(n703), .B(n702), .Z(n716) );
  XOR U3787 ( .A(n719), .B(n716), .Z(n704) );
  NAND U3788 ( .A(n720), .B(n704), .Z(n705) );
  NAND U3789 ( .A(n706), .B(n705), .Z(n765) );
  ANDN U3790 ( .B(n707), .A(n765), .Z(n731) );
  IV U3791 ( .A(n716), .Z(n722) );
  XOR U3792 ( .A(n724), .B(n720), .Z(n708) );
  NANDN U3793 ( .A(n722), .B(n708), .Z(n711) );
  NANDN U3794 ( .A(n720), .B(n722), .Z(n709) );
  NANDN U3795 ( .A(n719), .B(n709), .Z(n710) );
  NAND U3796 ( .A(n711), .B(n710), .Z(n800) );
  XNOR U3797 ( .A(n765), .B(n800), .Z(n741) );
  AND U3798 ( .A(n712), .B(n741), .Z(n734) );
  OR U3799 ( .A(n719), .B(n716), .Z(n718) );
  ANDN U3800 ( .B(n719), .A(n713), .Z(n714) );
  XNOR U3801 ( .A(n714), .B(n724), .Z(n715) );
  NAND U3802 ( .A(n716), .B(n715), .Z(n717) );
  NAND U3803 ( .A(n718), .B(n717), .Z(n738) );
  NAND U3804 ( .A(n720), .B(n724), .Z(n726) );
  NAND U3805 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U3806 ( .A(n722), .B(n721), .Z(n723) );
  NANDN U3807 ( .A(n724), .B(n723), .Z(n725) );
  NAND U3808 ( .A(n726), .B(n725), .Z(n807) );
  NAND U3809 ( .A(n757), .B(n727), .Z(n728) );
  XNOR U3810 ( .A(n734), .B(n728), .Z(n802) );
  XOR U3811 ( .A(n765), .B(n807), .Z(n767) );
  AND U3812 ( .A(n729), .B(n767), .Z(n752) );
  XNOR U3813 ( .A(n802), .B(n752), .Z(n730) );
  XNOR U3814 ( .A(n731), .B(n730), .Z(n810) );
  NAND U3815 ( .A(n743), .B(n732), .Z(n733) );
  XNOR U3816 ( .A(n734), .B(n733), .Z(n760) );
  AND U3817 ( .A(n735), .B(n745), .Z(n801) );
  NANDN U3818 ( .A(n736), .B(n738), .Z(n737) );
  XNOR U3819 ( .A(n801), .B(n737), .Z(n764) );
  XNOR U3820 ( .A(n760), .B(n764), .Z(n749) );
  XOR U3821 ( .A(n810), .B(n749), .Z(z[16]) );
  AND U3822 ( .A(n739), .B(n738), .Z(n748) );
  AND U3823 ( .A(n741), .B(n740), .Z(n759) );
  NAND U3824 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U3825 ( .A(n759), .B(n744), .Z(n811) );
  AND U3826 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U3827 ( .A(n811), .B(n753), .Z(n747) );
  XNOR U3828 ( .A(n748), .B(n747), .Z(n773) );
  XNOR U3829 ( .A(n773), .B(n749), .Z(n816) );
  AND U3830 ( .A(n750), .B(n800), .Z(n755) );
  NANDN U3831 ( .A(n807), .B(n805), .Z(n751) );
  XNOR U3832 ( .A(n752), .B(n751), .Z(n763) );
  XNOR U3833 ( .A(n753), .B(n763), .Z(n754) );
  XNOR U3834 ( .A(n755), .B(n754), .Z(n762) );
  NAND U3835 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U3836 ( .A(n759), .B(n758), .Z(n769) );
  XNOR U3837 ( .A(n760), .B(n769), .Z(n761) );
  XNOR U3838 ( .A(n762), .B(n761), .Z(n772) );
  XNOR U3839 ( .A(n816), .B(n772), .Z(z[17]) );
  XNOR U3840 ( .A(n764), .B(n763), .Z(z[18]) );
  NOR U3841 ( .A(n766), .B(n765), .Z(n771) );
  AND U3842 ( .A(n768), .B(n767), .Z(n809) );
  XNOR U3843 ( .A(n769), .B(n809), .Z(n770) );
  XNOR U3844 ( .A(n771), .B(n770), .Z(n815) );
  XOR U3845 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U3846 ( .A(n815), .B(n774), .Z(z[19]) );
  AND U3847 ( .A(n776), .B(n775), .Z(n785) );
  AND U3848 ( .A(n778), .B(n777), .Z(n796) );
  NAND U3849 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U3850 ( .A(n796), .B(n781), .Z(n1438) );
  AND U3851 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U3852 ( .A(n1438), .B(n790), .Z(n784) );
  XNOR U3853 ( .A(n785), .B(n784), .Z(n1074) );
  XNOR U3854 ( .A(n1074), .B(n786), .Z(n1581) );
  AND U3855 ( .A(n787), .B(n1427), .Z(n792) );
  NANDN U3856 ( .A(n1434), .B(n1432), .Z(n788) );
  XNOR U3857 ( .A(n789), .B(n788), .Z(n938) );
  XNOR U3858 ( .A(n790), .B(n938), .Z(n791) );
  XNOR U3859 ( .A(n792), .B(n791), .Z(n799) );
  NAND U3860 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U3861 ( .A(n796), .B(n795), .Z(n1070) );
  XNOR U3862 ( .A(n797), .B(n1070), .Z(n798) );
  XNOR U3863 ( .A(n799), .B(n798), .Z(n1073) );
  XNOR U3864 ( .A(n1581), .B(n1073), .Z(z[1]) );
  XOR U3865 ( .A(n810), .B(z[18]), .Z(z[20]) );
  AND U3866 ( .A(x[16]), .B(n800), .Z(n804) );
  XNOR U3867 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U3868 ( .A(n804), .B(n803), .Z(n817) );
  XOR U3869 ( .A(n805), .B(x[17]), .Z(n806) );
  NANDN U3870 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3871 ( .A(n809), .B(n808), .Z(n813) );
  XNOR U3872 ( .A(n811), .B(n810), .Z(n812) );
  XNOR U3873 ( .A(n813), .B(n812), .Z(n814) );
  XNOR U3874 ( .A(n817), .B(n814), .Z(z[21]) );
  XNOR U3875 ( .A(n816), .B(n815), .Z(z[22]) );
  XOR U3876 ( .A(n817), .B(z[17]), .Z(z[23]) );
  XOR U3877 ( .A(x[27]), .B(x[25]), .Z(n820) );
  XNOR U3878 ( .A(x[24]), .B(x[30]), .Z(n819) );
  XOR U3879 ( .A(n819), .B(x[26]), .Z(n818) );
  XNOR U3880 ( .A(n820), .B(n818), .Z(n855) );
  XNOR U3881 ( .A(x[29]), .B(n819), .Z(n928) );
  XOR U3882 ( .A(n928), .B(x[28]), .Z(n898) );
  IV U3883 ( .A(n898), .Z(n829) );
  XNOR U3884 ( .A(x[31]), .B(x[28]), .Z(n823) );
  XNOR U3885 ( .A(n820), .B(n823), .Z(n883) );
  NOR U3886 ( .A(n829), .B(n883), .Z(n822) );
  XNOR U3887 ( .A(n928), .B(x[31]), .Z(n914) );
  XNOR U3888 ( .A(x[26]), .B(n914), .Z(n838) );
  XNOR U3889 ( .A(x[25]), .B(n838), .Z(n833) );
  AND U3890 ( .A(x[24]), .B(n833), .Z(n821) );
  XNOR U3891 ( .A(n822), .B(n821), .Z(n826) );
  XNOR U3892 ( .A(n855), .B(n914), .Z(n845) );
  IV U3893 ( .A(n855), .Z(n840) );
  XNOR U3894 ( .A(x[24]), .B(n840), .Z(n860) );
  IV U3895 ( .A(n823), .Z(n888) );
  AND U3896 ( .A(n860), .B(n888), .Z(n828) );
  IV U3897 ( .A(n928), .Z(n847) );
  XNOR U3898 ( .A(n855), .B(n847), .Z(n877) );
  XOR U3899 ( .A(n877), .B(n883), .Z(n880) );
  XOR U3900 ( .A(x[26]), .B(x[28]), .Z(n890) );
  NAND U3901 ( .A(n880), .B(n890), .Z(n824) );
  XNOR U3902 ( .A(n828), .B(n824), .Z(n849) );
  XNOR U3903 ( .A(n845), .B(n849), .Z(n825) );
  XNOR U3904 ( .A(n826), .B(n825), .Z(n872) );
  XOR U3905 ( .A(x[26]), .B(x[31]), .Z(n904) );
  XNOR U3906 ( .A(x[24]), .B(n883), .Z(n884) );
  XNOR U3907 ( .A(n928), .B(n884), .Z(n875) );
  NAND U3908 ( .A(n904), .B(n875), .Z(n827) );
  XNOR U3909 ( .A(n828), .B(n827), .Z(n841) );
  IV U3910 ( .A(n833), .Z(n887) );
  XNOR U3911 ( .A(n887), .B(n829), .Z(n894) );
  AND U3912 ( .A(n883), .B(n894), .Z(n831) );
  AND U3913 ( .A(x[24]), .B(n898), .Z(n830) );
  XNOR U3914 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U3915 ( .A(n884), .B(n832), .Z(n836) );
  NAND U3916 ( .A(x[24]), .B(n883), .Z(n834) );
  OR U3917 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3918 ( .A(n836), .B(n835), .Z(n837) );
  XNOR U3919 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U3920 ( .A(n841), .B(n839), .Z(n861) );
  IV U3921 ( .A(n861), .Z(n868) );
  AND U3922 ( .A(n914), .B(n840), .Z(n843) );
  XOR U3923 ( .A(x[25]), .B(x[31]), .Z(n916) );
  AND U3924 ( .A(n877), .B(n916), .Z(n846) );
  XNOR U3925 ( .A(n846), .B(n841), .Z(n842) );
  XNOR U3926 ( .A(n843), .B(n842), .Z(n867) );
  NANDN U3927 ( .A(n868), .B(n867), .Z(n844) );
  NAND U3928 ( .A(n872), .B(n844), .Z(n854) );
  XNOR U3929 ( .A(n846), .B(n845), .Z(n851) );
  ANDN U3930 ( .B(n847), .A(x[25]), .Z(n848) );
  XNOR U3931 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U3932 ( .A(n851), .B(n850), .Z(n864) );
  XOR U3933 ( .A(n867), .B(n864), .Z(n852) );
  NAND U3934 ( .A(n868), .B(n852), .Z(n853) );
  NAND U3935 ( .A(n854), .B(n853), .Z(n913) );
  ANDN U3936 ( .B(n855), .A(n913), .Z(n879) );
  IV U3937 ( .A(n864), .Z(n870) );
  XOR U3938 ( .A(n872), .B(n868), .Z(n856) );
  NANDN U3939 ( .A(n870), .B(n856), .Z(n859) );
  NANDN U3940 ( .A(n868), .B(n870), .Z(n857) );
  NANDN U3941 ( .A(n867), .B(n857), .Z(n858) );
  NAND U3942 ( .A(n859), .B(n858), .Z(n923) );
  XNOR U3943 ( .A(n913), .B(n923), .Z(n889) );
  AND U3944 ( .A(n860), .B(n889), .Z(n882) );
  OR U3945 ( .A(n867), .B(n864), .Z(n866) );
  ANDN U3946 ( .B(n867), .A(n861), .Z(n862) );
  XNOR U3947 ( .A(n862), .B(n872), .Z(n863) );
  NAND U3948 ( .A(n864), .B(n863), .Z(n865) );
  NAND U3949 ( .A(n866), .B(n865), .Z(n886) );
  NAND U3950 ( .A(n868), .B(n872), .Z(n874) );
  NAND U3951 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U3952 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U3953 ( .A(n872), .B(n871), .Z(n873) );
  NAND U3954 ( .A(n874), .B(n873), .Z(n930) );
  NAND U3955 ( .A(n905), .B(n875), .Z(n876) );
  XNOR U3956 ( .A(n882), .B(n876), .Z(n925) );
  XOR U3957 ( .A(n913), .B(n930), .Z(n915) );
  AND U3958 ( .A(n877), .B(n915), .Z(n900) );
  XNOR U3959 ( .A(n925), .B(n900), .Z(n878) );
  XNOR U3960 ( .A(n879), .B(n878), .Z(n933) );
  NAND U3961 ( .A(n891), .B(n880), .Z(n881) );
  XNOR U3962 ( .A(n882), .B(n881), .Z(n908) );
  AND U3963 ( .A(n883), .B(n893), .Z(n924) );
  NANDN U3964 ( .A(n884), .B(n886), .Z(n885) );
  XNOR U3965 ( .A(n924), .B(n885), .Z(n912) );
  XNOR U3966 ( .A(n908), .B(n912), .Z(n897) );
  XOR U3967 ( .A(n933), .B(n897), .Z(z[24]) );
  AND U3968 ( .A(n887), .B(n886), .Z(n896) );
  AND U3969 ( .A(n889), .B(n888), .Z(n907) );
  NAND U3970 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U3971 ( .A(n907), .B(n892), .Z(n934) );
  AND U3972 ( .A(n894), .B(n893), .Z(n901) );
  XNOR U3973 ( .A(n934), .B(n901), .Z(n895) );
  XNOR U3974 ( .A(n896), .B(n895), .Z(n921) );
  XNOR U3975 ( .A(n921), .B(n897), .Z(n941) );
  AND U3976 ( .A(n898), .B(n923), .Z(n903) );
  NANDN U3977 ( .A(n930), .B(n928), .Z(n899) );
  XNOR U3978 ( .A(n900), .B(n899), .Z(n911) );
  XNOR U3979 ( .A(n901), .B(n911), .Z(n902) );
  XNOR U3980 ( .A(n903), .B(n902), .Z(n910) );
  NAND U3981 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3982 ( .A(n907), .B(n906), .Z(n917) );
  XNOR U3983 ( .A(n908), .B(n917), .Z(n909) );
  XNOR U3984 ( .A(n910), .B(n909), .Z(n920) );
  XNOR U3985 ( .A(n941), .B(n920), .Z(z[25]) );
  XNOR U3986 ( .A(n912), .B(n911), .Z(z[26]) );
  NOR U3987 ( .A(n914), .B(n913), .Z(n919) );
  AND U3988 ( .A(n916), .B(n915), .Z(n932) );
  XNOR U3989 ( .A(n917), .B(n932), .Z(n918) );
  XNOR U3990 ( .A(n919), .B(n918), .Z(n940) );
  XOR U3991 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U3992 ( .A(n940), .B(n922), .Z(z[27]) );
  XOR U3993 ( .A(n933), .B(z[26]), .Z(z[28]) );
  AND U3994 ( .A(x[24]), .B(n923), .Z(n927) );
  XNOR U3995 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U3996 ( .A(n927), .B(n926), .Z(n942) );
  XOR U3997 ( .A(n928), .B(x[25]), .Z(n929) );
  NANDN U3998 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U3999 ( .A(n932), .B(n931), .Z(n936) );
  XNOR U4000 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U4001 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U4002 ( .A(n942), .B(n937), .Z(z[29]) );
  XNOR U4003 ( .A(n939), .B(n938), .Z(z[2]) );
  XNOR U4004 ( .A(n941), .B(n940), .Z(z[30]) );
  XOR U4005 ( .A(n942), .B(z[25]), .Z(z[31]) );
  XOR U4006 ( .A(x[35]), .B(x[33]), .Z(n945) );
  XNOR U4007 ( .A(x[32]), .B(x[38]), .Z(n944) );
  XOR U4008 ( .A(n944), .B(x[34]), .Z(n943) );
  XNOR U4009 ( .A(n945), .B(n943), .Z(n980) );
  XNOR U4010 ( .A(x[37]), .B(n944), .Z(n1053) );
  XOR U4011 ( .A(n1053), .B(x[36]), .Z(n1023) );
  IV U4012 ( .A(n1023), .Z(n954) );
  XNOR U4013 ( .A(x[39]), .B(x[36]), .Z(n948) );
  XNOR U4014 ( .A(n945), .B(n948), .Z(n1008) );
  NOR U4015 ( .A(n954), .B(n1008), .Z(n947) );
  XNOR U4016 ( .A(n1053), .B(x[39]), .Z(n1039) );
  XNOR U4017 ( .A(x[34]), .B(n1039), .Z(n963) );
  XNOR U4018 ( .A(x[33]), .B(n963), .Z(n958) );
  AND U4019 ( .A(x[32]), .B(n958), .Z(n946) );
  XNOR U4020 ( .A(n947), .B(n946), .Z(n951) );
  XNOR U4021 ( .A(n980), .B(n1039), .Z(n970) );
  IV U4022 ( .A(n980), .Z(n965) );
  XNOR U4023 ( .A(x[32]), .B(n965), .Z(n985) );
  IV U4024 ( .A(n948), .Z(n1013) );
  AND U4025 ( .A(n985), .B(n1013), .Z(n953) );
  IV U4026 ( .A(n1053), .Z(n972) );
  XNOR U4027 ( .A(n980), .B(n972), .Z(n1002) );
  XOR U4028 ( .A(n1002), .B(n1008), .Z(n1005) );
  XOR U4029 ( .A(x[34]), .B(x[36]), .Z(n1015) );
  NAND U4030 ( .A(n1005), .B(n1015), .Z(n949) );
  XNOR U4031 ( .A(n953), .B(n949), .Z(n974) );
  XNOR U4032 ( .A(n970), .B(n974), .Z(n950) );
  XNOR U4033 ( .A(n951), .B(n950), .Z(n997) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1029) );
  XNOR U4035 ( .A(x[32]), .B(n1008), .Z(n1009) );
  XNOR U4036 ( .A(n1053), .B(n1009), .Z(n1000) );
  NAND U4037 ( .A(n1029), .B(n1000), .Z(n952) );
  XNOR U4038 ( .A(n953), .B(n952), .Z(n966) );
  IV U4039 ( .A(n958), .Z(n1012) );
  XNOR U4040 ( .A(n1012), .B(n954), .Z(n1019) );
  AND U4041 ( .A(n1008), .B(n1019), .Z(n956) );
  AND U4042 ( .A(x[32]), .B(n1023), .Z(n955) );
  XNOR U4043 ( .A(n956), .B(n955), .Z(n957) );
  NANDN U4044 ( .A(n1009), .B(n957), .Z(n961) );
  NAND U4045 ( .A(x[32]), .B(n1008), .Z(n959) );
  OR U4046 ( .A(n959), .B(n958), .Z(n960) );
  NAND U4047 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U4048 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U4049 ( .A(n966), .B(n964), .Z(n986) );
  IV U4050 ( .A(n986), .Z(n993) );
  AND U4051 ( .A(n1039), .B(n965), .Z(n968) );
  XOR U4052 ( .A(x[33]), .B(x[39]), .Z(n1041) );
  AND U4053 ( .A(n1002), .B(n1041), .Z(n971) );
  XNOR U4054 ( .A(n971), .B(n966), .Z(n967) );
  XNOR U4055 ( .A(n968), .B(n967), .Z(n992) );
  NANDN U4056 ( .A(n993), .B(n992), .Z(n969) );
  NAND U4057 ( .A(n997), .B(n969), .Z(n979) );
  XNOR U4058 ( .A(n971), .B(n970), .Z(n976) );
  ANDN U4059 ( .B(n972), .A(x[33]), .Z(n973) );
  XNOR U4060 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U4061 ( .A(n976), .B(n975), .Z(n989) );
  XOR U4062 ( .A(n992), .B(n989), .Z(n977) );
  NAND U4063 ( .A(n993), .B(n977), .Z(n978) );
  NAND U4064 ( .A(n979), .B(n978), .Z(n1038) );
  ANDN U4065 ( .B(n980), .A(n1038), .Z(n1004) );
  IV U4066 ( .A(n989), .Z(n995) );
  XOR U4067 ( .A(n997), .B(n993), .Z(n981) );
  NANDN U4068 ( .A(n995), .B(n981), .Z(n984) );
  NANDN U4069 ( .A(n993), .B(n995), .Z(n982) );
  NANDN U4070 ( .A(n992), .B(n982), .Z(n983) );
  NAND U4071 ( .A(n984), .B(n983), .Z(n1048) );
  XNOR U4072 ( .A(n1038), .B(n1048), .Z(n1014) );
  AND U4073 ( .A(n985), .B(n1014), .Z(n1007) );
  OR U4074 ( .A(n992), .B(n989), .Z(n991) );
  ANDN U4075 ( .B(n992), .A(n986), .Z(n987) );
  XNOR U4076 ( .A(n987), .B(n997), .Z(n988) );
  NAND U4077 ( .A(n989), .B(n988), .Z(n990) );
  NAND U4078 ( .A(n991), .B(n990), .Z(n1011) );
  NAND U4079 ( .A(n993), .B(n997), .Z(n999) );
  NAND U4080 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U4081 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U4082 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4083 ( .A(n999), .B(n998), .Z(n1055) );
  NAND U4084 ( .A(n1030), .B(n1000), .Z(n1001) );
  XNOR U4085 ( .A(n1007), .B(n1001), .Z(n1050) );
  XOR U4086 ( .A(n1038), .B(n1055), .Z(n1040) );
  AND U4087 ( .A(n1002), .B(n1040), .Z(n1025) );
  XNOR U4088 ( .A(n1050), .B(n1025), .Z(n1003) );
  XNOR U4089 ( .A(n1004), .B(n1003), .Z(n1058) );
  NAND U4090 ( .A(n1016), .B(n1005), .Z(n1006) );
  XNOR U4091 ( .A(n1007), .B(n1006), .Z(n1033) );
  AND U4092 ( .A(n1008), .B(n1018), .Z(n1049) );
  NANDN U4093 ( .A(n1009), .B(n1011), .Z(n1010) );
  XNOR U4094 ( .A(n1049), .B(n1010), .Z(n1037) );
  XNOR U4095 ( .A(n1033), .B(n1037), .Z(n1022) );
  XOR U4096 ( .A(n1058), .B(n1022), .Z(z[32]) );
  AND U4097 ( .A(n1012), .B(n1011), .Z(n1021) );
  AND U4098 ( .A(n1014), .B(n1013), .Z(n1032) );
  NAND U4099 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U4100 ( .A(n1032), .B(n1017), .Z(n1059) );
  AND U4101 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U4102 ( .A(n1059), .B(n1026), .Z(n1020) );
  XNOR U4103 ( .A(n1021), .B(n1020), .Z(n1046) );
  XNOR U4104 ( .A(n1046), .B(n1022), .Z(n1064) );
  AND U4105 ( .A(n1023), .B(n1048), .Z(n1028) );
  NANDN U4106 ( .A(n1055), .B(n1053), .Z(n1024) );
  XNOR U4107 ( .A(n1025), .B(n1024), .Z(n1036) );
  XNOR U4108 ( .A(n1026), .B(n1036), .Z(n1027) );
  XNOR U4109 ( .A(n1028), .B(n1027), .Z(n1035) );
  NAND U4110 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U4111 ( .A(n1032), .B(n1031), .Z(n1042) );
  XNOR U4112 ( .A(n1033), .B(n1042), .Z(n1034) );
  XNOR U4113 ( .A(n1035), .B(n1034), .Z(n1045) );
  XNOR U4114 ( .A(n1064), .B(n1045), .Z(z[33]) );
  XNOR U4115 ( .A(n1037), .B(n1036), .Z(z[34]) );
  NOR U4116 ( .A(n1039), .B(n1038), .Z(n1044) );
  AND U4117 ( .A(n1041), .B(n1040), .Z(n1057) );
  XNOR U4118 ( .A(n1042), .B(n1057), .Z(n1043) );
  XNOR U4119 ( .A(n1044), .B(n1043), .Z(n1063) );
  XOR U4120 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U4121 ( .A(n1063), .B(n1047), .Z(z[35]) );
  XOR U4122 ( .A(n1058), .B(z[34]), .Z(z[36]) );
  AND U4123 ( .A(x[32]), .B(n1048), .Z(n1052) );
  XNOR U4124 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U4125 ( .A(n1052), .B(n1051), .Z(n1065) );
  XOR U4126 ( .A(n1053), .B(x[33]), .Z(n1054) );
  NANDN U4127 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U4128 ( .A(n1057), .B(n1056), .Z(n1061) );
  XNOR U4129 ( .A(n1059), .B(n1058), .Z(n1060) );
  XNOR U4130 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U4131 ( .A(n1065), .B(n1062), .Z(z[37]) );
  XNOR U4132 ( .A(n1064), .B(n1063), .Z(z[38]) );
  XOR U4133 ( .A(n1065), .B(z[33]), .Z(z[39]) );
  NOR U4134 ( .A(n1067), .B(n1066), .Z(n1072) );
  AND U4135 ( .A(n1069), .B(n1068), .Z(n1436) );
  XNOR U4136 ( .A(n1070), .B(n1436), .Z(n1071) );
  XNOR U4137 ( .A(n1072), .B(n1071), .Z(n1580) );
  XOR U4138 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U4139 ( .A(n1580), .B(n1075), .Z(z[3]) );
  XOR U4140 ( .A(x[43]), .B(x[41]), .Z(n1078) );
  XNOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1077) );
  XOR U4142 ( .A(n1077), .B(x[42]), .Z(n1076) );
  XNOR U4143 ( .A(n1078), .B(n1076), .Z(n1113) );
  XNOR U4144 ( .A(x[45]), .B(n1077), .Z(n1186) );
  XOR U4145 ( .A(n1186), .B(x[44]), .Z(n1156) );
  IV U4146 ( .A(n1156), .Z(n1087) );
  XNOR U4147 ( .A(x[47]), .B(x[44]), .Z(n1081) );
  XNOR U4148 ( .A(n1078), .B(n1081), .Z(n1141) );
  NOR U4149 ( .A(n1087), .B(n1141), .Z(n1080) );
  XNOR U4150 ( .A(n1186), .B(x[47]), .Z(n1172) );
  XNOR U4151 ( .A(x[42]), .B(n1172), .Z(n1096) );
  XNOR U4152 ( .A(x[41]), .B(n1096), .Z(n1091) );
  AND U4153 ( .A(x[40]), .B(n1091), .Z(n1079) );
  XNOR U4154 ( .A(n1080), .B(n1079), .Z(n1084) );
  XNOR U4155 ( .A(n1113), .B(n1172), .Z(n1103) );
  IV U4156 ( .A(n1113), .Z(n1098) );
  XNOR U4157 ( .A(x[40]), .B(n1098), .Z(n1118) );
  IV U4158 ( .A(n1081), .Z(n1146) );
  AND U4159 ( .A(n1118), .B(n1146), .Z(n1086) );
  IV U4160 ( .A(n1186), .Z(n1105) );
  XNOR U4161 ( .A(n1113), .B(n1105), .Z(n1135) );
  XOR U4162 ( .A(n1135), .B(n1141), .Z(n1138) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1148) );
  NAND U4164 ( .A(n1138), .B(n1148), .Z(n1082) );
  XNOR U4165 ( .A(n1086), .B(n1082), .Z(n1107) );
  XNOR U4166 ( .A(n1103), .B(n1107), .Z(n1083) );
  XNOR U4167 ( .A(n1084), .B(n1083), .Z(n1130) );
  XOR U4168 ( .A(x[42]), .B(x[47]), .Z(n1162) );
  XNOR U4169 ( .A(x[40]), .B(n1141), .Z(n1142) );
  XNOR U4170 ( .A(n1186), .B(n1142), .Z(n1133) );
  NAND U4171 ( .A(n1162), .B(n1133), .Z(n1085) );
  XNOR U4172 ( .A(n1086), .B(n1085), .Z(n1099) );
  IV U4173 ( .A(n1091), .Z(n1145) );
  XNOR U4174 ( .A(n1145), .B(n1087), .Z(n1152) );
  AND U4175 ( .A(n1141), .B(n1152), .Z(n1089) );
  AND U4176 ( .A(x[40]), .B(n1156), .Z(n1088) );
  XNOR U4177 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U4178 ( .A(n1142), .B(n1090), .Z(n1094) );
  NAND U4179 ( .A(x[40]), .B(n1141), .Z(n1092) );
  OR U4180 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U4181 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U4182 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U4183 ( .A(n1099), .B(n1097), .Z(n1119) );
  IV U4184 ( .A(n1119), .Z(n1126) );
  AND U4185 ( .A(n1172), .B(n1098), .Z(n1101) );
  XOR U4186 ( .A(x[41]), .B(x[47]), .Z(n1174) );
  AND U4187 ( .A(n1135), .B(n1174), .Z(n1104) );
  XNOR U4188 ( .A(n1104), .B(n1099), .Z(n1100) );
  XNOR U4189 ( .A(n1101), .B(n1100), .Z(n1125) );
  NANDN U4190 ( .A(n1126), .B(n1125), .Z(n1102) );
  NAND U4191 ( .A(n1130), .B(n1102), .Z(n1112) );
  XNOR U4192 ( .A(n1104), .B(n1103), .Z(n1109) );
  ANDN U4193 ( .B(n1105), .A(x[41]), .Z(n1106) );
  XNOR U4194 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U4195 ( .A(n1109), .B(n1108), .Z(n1122) );
  XOR U4196 ( .A(n1125), .B(n1122), .Z(n1110) );
  NAND U4197 ( .A(n1126), .B(n1110), .Z(n1111) );
  NAND U4198 ( .A(n1112), .B(n1111), .Z(n1171) );
  ANDN U4199 ( .B(n1113), .A(n1171), .Z(n1137) );
  IV U4200 ( .A(n1122), .Z(n1128) );
  XOR U4201 ( .A(n1130), .B(n1126), .Z(n1114) );
  NANDN U4202 ( .A(n1128), .B(n1114), .Z(n1117) );
  NANDN U4203 ( .A(n1126), .B(n1128), .Z(n1115) );
  NANDN U4204 ( .A(n1125), .B(n1115), .Z(n1116) );
  NAND U4205 ( .A(n1117), .B(n1116), .Z(n1181) );
  XNOR U4206 ( .A(n1171), .B(n1181), .Z(n1147) );
  AND U4207 ( .A(n1118), .B(n1147), .Z(n1140) );
  OR U4208 ( .A(n1125), .B(n1122), .Z(n1124) );
  ANDN U4209 ( .B(n1125), .A(n1119), .Z(n1120) );
  XNOR U4210 ( .A(n1120), .B(n1130), .Z(n1121) );
  NAND U4211 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U4212 ( .A(n1124), .B(n1123), .Z(n1144) );
  NAND U4213 ( .A(n1126), .B(n1130), .Z(n1132) );
  NAND U4214 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U4215 ( .A(n1128), .B(n1127), .Z(n1129) );
  NANDN U4216 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U4217 ( .A(n1132), .B(n1131), .Z(n1188) );
  NAND U4218 ( .A(n1163), .B(n1133), .Z(n1134) );
  XNOR U4219 ( .A(n1140), .B(n1134), .Z(n1183) );
  XOR U4220 ( .A(n1171), .B(n1188), .Z(n1173) );
  AND U4221 ( .A(n1135), .B(n1173), .Z(n1158) );
  XNOR U4222 ( .A(n1183), .B(n1158), .Z(n1136) );
  XNOR U4223 ( .A(n1137), .B(n1136), .Z(n1191) );
  NAND U4224 ( .A(n1149), .B(n1138), .Z(n1139) );
  XNOR U4225 ( .A(n1140), .B(n1139), .Z(n1166) );
  AND U4226 ( .A(n1141), .B(n1151), .Z(n1182) );
  NANDN U4227 ( .A(n1142), .B(n1144), .Z(n1143) );
  XNOR U4228 ( .A(n1182), .B(n1143), .Z(n1170) );
  XNOR U4229 ( .A(n1166), .B(n1170), .Z(n1155) );
  XOR U4230 ( .A(n1191), .B(n1155), .Z(z[40]) );
  AND U4231 ( .A(n1145), .B(n1144), .Z(n1154) );
  AND U4232 ( .A(n1147), .B(n1146), .Z(n1165) );
  NAND U4233 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U4234 ( .A(n1165), .B(n1150), .Z(n1192) );
  AND U4235 ( .A(n1152), .B(n1151), .Z(n1159) );
  XNOR U4236 ( .A(n1192), .B(n1159), .Z(n1153) );
  XNOR U4237 ( .A(n1154), .B(n1153), .Z(n1179) );
  XNOR U4238 ( .A(n1179), .B(n1155), .Z(n1197) );
  AND U4239 ( .A(n1156), .B(n1181), .Z(n1161) );
  NANDN U4240 ( .A(n1188), .B(n1186), .Z(n1157) );
  XNOR U4241 ( .A(n1158), .B(n1157), .Z(n1169) );
  XNOR U4242 ( .A(n1159), .B(n1169), .Z(n1160) );
  XNOR U4243 ( .A(n1161), .B(n1160), .Z(n1168) );
  NAND U4244 ( .A(n1163), .B(n1162), .Z(n1164) );
  XNOR U4245 ( .A(n1165), .B(n1164), .Z(n1175) );
  XNOR U4246 ( .A(n1166), .B(n1175), .Z(n1167) );
  XNOR U4247 ( .A(n1168), .B(n1167), .Z(n1178) );
  XNOR U4248 ( .A(n1197), .B(n1178), .Z(z[41]) );
  XNOR U4249 ( .A(n1170), .B(n1169), .Z(z[42]) );
  NOR U4250 ( .A(n1172), .B(n1171), .Z(n1177) );
  AND U4251 ( .A(n1174), .B(n1173), .Z(n1190) );
  XNOR U4252 ( .A(n1175), .B(n1190), .Z(n1176) );
  XNOR U4253 ( .A(n1177), .B(n1176), .Z(n1196) );
  XOR U4254 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4255 ( .A(n1196), .B(n1180), .Z(z[43]) );
  XOR U4256 ( .A(n1191), .B(z[42]), .Z(z[44]) );
  AND U4257 ( .A(x[40]), .B(n1181), .Z(n1185) );
  XNOR U4258 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U4259 ( .A(n1185), .B(n1184), .Z(n1198) );
  XOR U4260 ( .A(n1186), .B(x[41]), .Z(n1187) );
  NANDN U4261 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U4262 ( .A(n1190), .B(n1189), .Z(n1194) );
  XNOR U4263 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U4264 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U4265 ( .A(n1198), .B(n1195), .Z(z[45]) );
  XNOR U4266 ( .A(n1197), .B(n1196), .Z(z[46]) );
  XOR U4267 ( .A(n1198), .B(z[41]), .Z(z[47]) );
  XOR U4268 ( .A(x[51]), .B(x[49]), .Z(n1201) );
  XNOR U4269 ( .A(x[48]), .B(x[54]), .Z(n1200) );
  XOR U4270 ( .A(n1200), .B(x[50]), .Z(n1199) );
  XNOR U4271 ( .A(n1201), .B(n1199), .Z(n1236) );
  XNOR U4272 ( .A(x[53]), .B(n1200), .Z(n1309) );
  XOR U4273 ( .A(n1309), .B(x[52]), .Z(n1279) );
  IV U4274 ( .A(n1279), .Z(n1210) );
  XNOR U4275 ( .A(x[55]), .B(x[52]), .Z(n1204) );
  XNOR U4276 ( .A(n1201), .B(n1204), .Z(n1264) );
  NOR U4277 ( .A(n1210), .B(n1264), .Z(n1203) );
  XNOR U4278 ( .A(n1309), .B(x[55]), .Z(n1295) );
  XNOR U4279 ( .A(x[50]), .B(n1295), .Z(n1219) );
  XNOR U4280 ( .A(x[49]), .B(n1219), .Z(n1214) );
  AND U4281 ( .A(x[48]), .B(n1214), .Z(n1202) );
  XNOR U4282 ( .A(n1203), .B(n1202), .Z(n1207) );
  XNOR U4283 ( .A(n1236), .B(n1295), .Z(n1226) );
  IV U4284 ( .A(n1236), .Z(n1221) );
  XNOR U4285 ( .A(x[48]), .B(n1221), .Z(n1241) );
  IV U4286 ( .A(n1204), .Z(n1269) );
  AND U4287 ( .A(n1241), .B(n1269), .Z(n1209) );
  IV U4288 ( .A(n1309), .Z(n1228) );
  XNOR U4289 ( .A(n1236), .B(n1228), .Z(n1258) );
  XOR U4290 ( .A(n1258), .B(n1264), .Z(n1261) );
  XOR U4291 ( .A(x[50]), .B(x[52]), .Z(n1271) );
  NAND U4292 ( .A(n1261), .B(n1271), .Z(n1205) );
  XNOR U4293 ( .A(n1209), .B(n1205), .Z(n1230) );
  XNOR U4294 ( .A(n1226), .B(n1230), .Z(n1206) );
  XNOR U4295 ( .A(n1207), .B(n1206), .Z(n1253) );
  XOR U4296 ( .A(x[50]), .B(x[55]), .Z(n1285) );
  XNOR U4297 ( .A(x[48]), .B(n1264), .Z(n1265) );
  XNOR U4298 ( .A(n1309), .B(n1265), .Z(n1256) );
  NAND U4299 ( .A(n1285), .B(n1256), .Z(n1208) );
  XNOR U4300 ( .A(n1209), .B(n1208), .Z(n1222) );
  IV U4301 ( .A(n1214), .Z(n1268) );
  XNOR U4302 ( .A(n1268), .B(n1210), .Z(n1275) );
  AND U4303 ( .A(n1264), .B(n1275), .Z(n1212) );
  AND U4304 ( .A(x[48]), .B(n1279), .Z(n1211) );
  XNOR U4305 ( .A(n1212), .B(n1211), .Z(n1213) );
  NANDN U4306 ( .A(n1265), .B(n1213), .Z(n1217) );
  NAND U4307 ( .A(x[48]), .B(n1264), .Z(n1215) );
  OR U4308 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4309 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U4310 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U4311 ( .A(n1222), .B(n1220), .Z(n1242) );
  IV U4312 ( .A(n1242), .Z(n1249) );
  AND U4313 ( .A(n1295), .B(n1221), .Z(n1224) );
  XOR U4314 ( .A(x[49]), .B(x[55]), .Z(n1297) );
  AND U4315 ( .A(n1258), .B(n1297), .Z(n1227) );
  XNOR U4316 ( .A(n1227), .B(n1222), .Z(n1223) );
  XNOR U4317 ( .A(n1224), .B(n1223), .Z(n1248) );
  NANDN U4318 ( .A(n1249), .B(n1248), .Z(n1225) );
  NAND U4319 ( .A(n1253), .B(n1225), .Z(n1235) );
  XNOR U4320 ( .A(n1227), .B(n1226), .Z(n1232) );
  ANDN U4321 ( .B(n1228), .A(x[49]), .Z(n1229) );
  XNOR U4322 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U4323 ( .A(n1232), .B(n1231), .Z(n1245) );
  XOR U4324 ( .A(n1248), .B(n1245), .Z(n1233) );
  NAND U4325 ( .A(n1249), .B(n1233), .Z(n1234) );
  NAND U4326 ( .A(n1235), .B(n1234), .Z(n1294) );
  ANDN U4327 ( .B(n1236), .A(n1294), .Z(n1260) );
  IV U4328 ( .A(n1245), .Z(n1251) );
  XOR U4329 ( .A(n1253), .B(n1249), .Z(n1237) );
  NANDN U4330 ( .A(n1251), .B(n1237), .Z(n1240) );
  NANDN U4331 ( .A(n1249), .B(n1251), .Z(n1238) );
  NANDN U4332 ( .A(n1248), .B(n1238), .Z(n1239) );
  NAND U4333 ( .A(n1240), .B(n1239), .Z(n1304) );
  XNOR U4334 ( .A(n1294), .B(n1304), .Z(n1270) );
  AND U4335 ( .A(n1241), .B(n1270), .Z(n1263) );
  OR U4336 ( .A(n1248), .B(n1245), .Z(n1247) );
  ANDN U4337 ( .B(n1248), .A(n1242), .Z(n1243) );
  XNOR U4338 ( .A(n1243), .B(n1253), .Z(n1244) );
  NAND U4339 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U4340 ( .A(n1247), .B(n1246), .Z(n1267) );
  NAND U4341 ( .A(n1249), .B(n1253), .Z(n1255) );
  NAND U4342 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U4343 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U4344 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U4345 ( .A(n1255), .B(n1254), .Z(n1311) );
  NAND U4346 ( .A(n1286), .B(n1256), .Z(n1257) );
  XNOR U4347 ( .A(n1263), .B(n1257), .Z(n1306) );
  XOR U4348 ( .A(n1294), .B(n1311), .Z(n1296) );
  AND U4349 ( .A(n1258), .B(n1296), .Z(n1281) );
  XNOR U4350 ( .A(n1306), .B(n1281), .Z(n1259) );
  XNOR U4351 ( .A(n1260), .B(n1259), .Z(n1314) );
  NAND U4352 ( .A(n1272), .B(n1261), .Z(n1262) );
  XNOR U4353 ( .A(n1263), .B(n1262), .Z(n1289) );
  AND U4354 ( .A(n1264), .B(n1274), .Z(n1305) );
  NANDN U4355 ( .A(n1265), .B(n1267), .Z(n1266) );
  XNOR U4356 ( .A(n1305), .B(n1266), .Z(n1293) );
  XNOR U4357 ( .A(n1289), .B(n1293), .Z(n1278) );
  XOR U4358 ( .A(n1314), .B(n1278), .Z(z[48]) );
  AND U4359 ( .A(n1268), .B(n1267), .Z(n1277) );
  AND U4360 ( .A(n1270), .B(n1269), .Z(n1288) );
  NAND U4361 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U4362 ( .A(n1288), .B(n1273), .Z(n1315) );
  AND U4363 ( .A(n1275), .B(n1274), .Z(n1282) );
  XNOR U4364 ( .A(n1315), .B(n1282), .Z(n1276) );
  XNOR U4365 ( .A(n1277), .B(n1276), .Z(n1302) );
  XNOR U4366 ( .A(n1302), .B(n1278), .Z(n1320) );
  AND U4367 ( .A(n1279), .B(n1304), .Z(n1284) );
  NANDN U4368 ( .A(n1311), .B(n1309), .Z(n1280) );
  XNOR U4369 ( .A(n1281), .B(n1280), .Z(n1292) );
  XNOR U4370 ( .A(n1282), .B(n1292), .Z(n1283) );
  XNOR U4371 ( .A(n1284), .B(n1283), .Z(n1291) );
  NAND U4372 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U4373 ( .A(n1288), .B(n1287), .Z(n1298) );
  XNOR U4374 ( .A(n1289), .B(n1298), .Z(n1290) );
  XNOR U4375 ( .A(n1291), .B(n1290), .Z(n1301) );
  XNOR U4376 ( .A(n1320), .B(n1301), .Z(z[49]) );
  XOR U4377 ( .A(n1437), .B(z[2]), .Z(z[4]) );
  XNOR U4378 ( .A(n1293), .B(n1292), .Z(z[50]) );
  NOR U4379 ( .A(n1295), .B(n1294), .Z(n1300) );
  AND U4380 ( .A(n1297), .B(n1296), .Z(n1313) );
  XNOR U4381 ( .A(n1298), .B(n1313), .Z(n1299) );
  XNOR U4382 ( .A(n1300), .B(n1299), .Z(n1319) );
  XOR U4383 ( .A(n1302), .B(n1301), .Z(n1303) );
  XNOR U4384 ( .A(n1319), .B(n1303), .Z(z[51]) );
  XOR U4385 ( .A(n1314), .B(z[50]), .Z(z[52]) );
  AND U4386 ( .A(x[48]), .B(n1304), .Z(n1308) );
  XNOR U4387 ( .A(n1306), .B(n1305), .Z(n1307) );
  XNOR U4388 ( .A(n1308), .B(n1307), .Z(n1321) );
  XOR U4389 ( .A(n1309), .B(x[49]), .Z(n1310) );
  NANDN U4390 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U4391 ( .A(n1313), .B(n1312), .Z(n1317) );
  XNOR U4392 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U4393 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U4394 ( .A(n1321), .B(n1318), .Z(z[53]) );
  XNOR U4395 ( .A(n1320), .B(n1319), .Z(z[54]) );
  XOR U4396 ( .A(n1321), .B(z[49]), .Z(z[55]) );
  XOR U4397 ( .A(x[59]), .B(x[57]), .Z(n1324) );
  XNOR U4398 ( .A(x[56]), .B(x[62]), .Z(n1323) );
  XOR U4399 ( .A(n1323), .B(x[58]), .Z(n1322) );
  XNOR U4400 ( .A(n1324), .B(n1322), .Z(n1359) );
  XNOR U4401 ( .A(x[61]), .B(n1323), .Z(n1447) );
  XOR U4402 ( .A(n1447), .B(x[60]), .Z(n1402) );
  IV U4403 ( .A(n1402), .Z(n1333) );
  XNOR U4404 ( .A(x[63]), .B(x[60]), .Z(n1327) );
  XNOR U4405 ( .A(n1324), .B(n1327), .Z(n1387) );
  NOR U4406 ( .A(n1333), .B(n1387), .Z(n1326) );
  XNOR U4407 ( .A(n1447), .B(x[63]), .Z(n1418) );
  XNOR U4408 ( .A(x[58]), .B(n1418), .Z(n1342) );
  XNOR U4409 ( .A(x[57]), .B(n1342), .Z(n1337) );
  AND U4410 ( .A(x[56]), .B(n1337), .Z(n1325) );
  XNOR U4411 ( .A(n1326), .B(n1325), .Z(n1330) );
  XNOR U4412 ( .A(n1359), .B(n1418), .Z(n1349) );
  IV U4413 ( .A(n1359), .Z(n1344) );
  XNOR U4414 ( .A(x[56]), .B(n1344), .Z(n1364) );
  IV U4415 ( .A(n1327), .Z(n1392) );
  AND U4416 ( .A(n1364), .B(n1392), .Z(n1332) );
  IV U4417 ( .A(n1447), .Z(n1351) );
  XNOR U4418 ( .A(n1359), .B(n1351), .Z(n1381) );
  XOR U4419 ( .A(n1381), .B(n1387), .Z(n1384) );
  XOR U4420 ( .A(x[58]), .B(x[60]), .Z(n1394) );
  NAND U4421 ( .A(n1384), .B(n1394), .Z(n1328) );
  XNOR U4422 ( .A(n1332), .B(n1328), .Z(n1353) );
  XNOR U4423 ( .A(n1349), .B(n1353), .Z(n1329) );
  XNOR U4424 ( .A(n1330), .B(n1329), .Z(n1376) );
  XOR U4425 ( .A(x[58]), .B(x[63]), .Z(n1408) );
  XNOR U4426 ( .A(x[56]), .B(n1387), .Z(n1388) );
  XNOR U4427 ( .A(n1447), .B(n1388), .Z(n1379) );
  NAND U4428 ( .A(n1408), .B(n1379), .Z(n1331) );
  XNOR U4429 ( .A(n1332), .B(n1331), .Z(n1345) );
  IV U4430 ( .A(n1337), .Z(n1391) );
  XNOR U4431 ( .A(n1391), .B(n1333), .Z(n1398) );
  AND U4432 ( .A(n1387), .B(n1398), .Z(n1335) );
  AND U4433 ( .A(x[56]), .B(n1402), .Z(n1334) );
  XNOR U4434 ( .A(n1335), .B(n1334), .Z(n1336) );
  NANDN U4435 ( .A(n1388), .B(n1336), .Z(n1340) );
  NAND U4436 ( .A(x[56]), .B(n1387), .Z(n1338) );
  OR U4437 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U4438 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4439 ( .A(n1342), .B(n1341), .Z(n1343) );
  XNOR U4440 ( .A(n1345), .B(n1343), .Z(n1365) );
  IV U4441 ( .A(n1365), .Z(n1372) );
  AND U4442 ( .A(n1418), .B(n1344), .Z(n1347) );
  XOR U4443 ( .A(x[57]), .B(x[63]), .Z(n1420) );
  AND U4444 ( .A(n1381), .B(n1420), .Z(n1350) );
  XNOR U4445 ( .A(n1350), .B(n1345), .Z(n1346) );
  XNOR U4446 ( .A(n1347), .B(n1346), .Z(n1371) );
  NANDN U4447 ( .A(n1372), .B(n1371), .Z(n1348) );
  NAND U4448 ( .A(n1376), .B(n1348), .Z(n1358) );
  XNOR U4449 ( .A(n1350), .B(n1349), .Z(n1355) );
  ANDN U4450 ( .B(n1351), .A(x[57]), .Z(n1352) );
  XNOR U4451 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U4452 ( .A(n1355), .B(n1354), .Z(n1368) );
  XOR U4453 ( .A(n1371), .B(n1368), .Z(n1356) );
  NAND U4454 ( .A(n1372), .B(n1356), .Z(n1357) );
  NAND U4455 ( .A(n1358), .B(n1357), .Z(n1417) );
  ANDN U4456 ( .B(n1359), .A(n1417), .Z(n1383) );
  IV U4457 ( .A(n1368), .Z(n1374) );
  XOR U4458 ( .A(n1376), .B(n1372), .Z(n1360) );
  NANDN U4459 ( .A(n1374), .B(n1360), .Z(n1363) );
  NANDN U4460 ( .A(n1372), .B(n1374), .Z(n1361) );
  NANDN U4461 ( .A(n1371), .B(n1361), .Z(n1362) );
  NAND U4462 ( .A(n1363), .B(n1362), .Z(n1442) );
  XNOR U4463 ( .A(n1417), .B(n1442), .Z(n1393) );
  AND U4464 ( .A(n1364), .B(n1393), .Z(n1386) );
  OR U4465 ( .A(n1371), .B(n1368), .Z(n1370) );
  ANDN U4466 ( .B(n1371), .A(n1365), .Z(n1366) );
  XNOR U4467 ( .A(n1366), .B(n1376), .Z(n1367) );
  NAND U4468 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U4469 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U4470 ( .A(n1372), .B(n1376), .Z(n1378) );
  NAND U4471 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4472 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U4473 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U4474 ( .A(n1378), .B(n1377), .Z(n1449) );
  NAND U4475 ( .A(n1409), .B(n1379), .Z(n1380) );
  XNOR U4476 ( .A(n1386), .B(n1380), .Z(n1444) );
  XOR U4477 ( .A(n1417), .B(n1449), .Z(n1419) );
  AND U4478 ( .A(n1381), .B(n1419), .Z(n1404) );
  XNOR U4479 ( .A(n1444), .B(n1404), .Z(n1382) );
  XNOR U4480 ( .A(n1383), .B(n1382), .Z(n1452) );
  NAND U4481 ( .A(n1395), .B(n1384), .Z(n1385) );
  XNOR U4482 ( .A(n1386), .B(n1385), .Z(n1412) );
  AND U4483 ( .A(n1387), .B(n1397), .Z(n1443) );
  NANDN U4484 ( .A(n1388), .B(n1390), .Z(n1389) );
  XNOR U4485 ( .A(n1443), .B(n1389), .Z(n1416) );
  XNOR U4486 ( .A(n1412), .B(n1416), .Z(n1401) );
  XOR U4487 ( .A(n1452), .B(n1401), .Z(z[56]) );
  AND U4488 ( .A(n1391), .B(n1390), .Z(n1400) );
  AND U4489 ( .A(n1393), .B(n1392), .Z(n1411) );
  NAND U4490 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U4491 ( .A(n1411), .B(n1396), .Z(n1453) );
  AND U4492 ( .A(n1398), .B(n1397), .Z(n1405) );
  XNOR U4493 ( .A(n1453), .B(n1405), .Z(n1399) );
  XNOR U4494 ( .A(n1400), .B(n1399), .Z(n1425) );
  XNOR U4495 ( .A(n1425), .B(n1401), .Z(n1458) );
  AND U4496 ( .A(n1402), .B(n1442), .Z(n1407) );
  NANDN U4497 ( .A(n1449), .B(n1447), .Z(n1403) );
  XNOR U4498 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U4499 ( .A(n1405), .B(n1415), .Z(n1406) );
  XNOR U4500 ( .A(n1407), .B(n1406), .Z(n1414) );
  NAND U4501 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U4502 ( .A(n1411), .B(n1410), .Z(n1421) );
  XNOR U4503 ( .A(n1412), .B(n1421), .Z(n1413) );
  XNOR U4504 ( .A(n1414), .B(n1413), .Z(n1424) );
  XNOR U4505 ( .A(n1458), .B(n1424), .Z(z[57]) );
  XNOR U4506 ( .A(n1416), .B(n1415), .Z(z[58]) );
  NOR U4507 ( .A(n1418), .B(n1417), .Z(n1423) );
  AND U4508 ( .A(n1420), .B(n1419), .Z(n1451) );
  XNOR U4509 ( .A(n1421), .B(n1451), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1457) );
  XOR U4511 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U4512 ( .A(n1457), .B(n1426), .Z(z[59]) );
  AND U4513 ( .A(x[0]), .B(n1427), .Z(n1431) );
  XNOR U4514 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U4515 ( .A(n1431), .B(n1430), .Z(n1708) );
  XOR U4516 ( .A(n1432), .B(x[1]), .Z(n1433) );
  NANDN U4517 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U4518 ( .A(n1436), .B(n1435), .Z(n1440) );
  XNOR U4519 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U4520 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U4521 ( .A(n1708), .B(n1441), .Z(z[5]) );
  XOR U4522 ( .A(n1452), .B(z[58]), .Z(z[60]) );
  AND U4523 ( .A(x[56]), .B(n1442), .Z(n1446) );
  XNOR U4524 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U4525 ( .A(n1446), .B(n1445), .Z(n1459) );
  XOR U4526 ( .A(n1447), .B(x[57]), .Z(n1448) );
  NANDN U4527 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U4528 ( .A(n1451), .B(n1450), .Z(n1455) );
  XNOR U4529 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U4530 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U4531 ( .A(n1459), .B(n1456), .Z(z[61]) );
  XNOR U4532 ( .A(n1458), .B(n1457), .Z(z[62]) );
  XOR U4533 ( .A(n1459), .B(z[57]), .Z(z[63]) );
  XOR U4534 ( .A(x[67]), .B(x[65]), .Z(n1462) );
  XNOR U4535 ( .A(x[64]), .B(x[70]), .Z(n1461) );
  XOR U4536 ( .A(n1461), .B(x[66]), .Z(n1460) );
  XNOR U4537 ( .A(n1462), .B(n1460), .Z(n1497) );
  XNOR U4538 ( .A(x[69]), .B(n1461), .Z(n1570) );
  XOR U4539 ( .A(n1570), .B(x[68]), .Z(n1540) );
  IV U4540 ( .A(n1540), .Z(n1471) );
  XNOR U4541 ( .A(x[71]), .B(x[68]), .Z(n1465) );
  XNOR U4542 ( .A(n1462), .B(n1465), .Z(n1525) );
  NOR U4543 ( .A(n1471), .B(n1525), .Z(n1464) );
  XNOR U4544 ( .A(n1570), .B(x[71]), .Z(n1556) );
  XNOR U4545 ( .A(x[66]), .B(n1556), .Z(n1480) );
  XNOR U4546 ( .A(x[65]), .B(n1480), .Z(n1475) );
  AND U4547 ( .A(x[64]), .B(n1475), .Z(n1463) );
  XNOR U4548 ( .A(n1464), .B(n1463), .Z(n1468) );
  XNOR U4549 ( .A(n1497), .B(n1556), .Z(n1487) );
  IV U4550 ( .A(n1497), .Z(n1482) );
  XNOR U4551 ( .A(x[64]), .B(n1482), .Z(n1502) );
  IV U4552 ( .A(n1465), .Z(n1530) );
  AND U4553 ( .A(n1502), .B(n1530), .Z(n1470) );
  IV U4554 ( .A(n1570), .Z(n1489) );
  XNOR U4555 ( .A(n1497), .B(n1489), .Z(n1519) );
  XOR U4556 ( .A(n1519), .B(n1525), .Z(n1522) );
  XOR U4557 ( .A(x[66]), .B(x[68]), .Z(n1532) );
  NAND U4558 ( .A(n1522), .B(n1532), .Z(n1466) );
  XNOR U4559 ( .A(n1470), .B(n1466), .Z(n1491) );
  XNOR U4560 ( .A(n1487), .B(n1491), .Z(n1467) );
  XNOR U4561 ( .A(n1468), .B(n1467), .Z(n1514) );
  XOR U4562 ( .A(x[66]), .B(x[71]), .Z(n1546) );
  XNOR U4563 ( .A(x[64]), .B(n1525), .Z(n1526) );
  XNOR U4564 ( .A(n1570), .B(n1526), .Z(n1517) );
  NAND U4565 ( .A(n1546), .B(n1517), .Z(n1469) );
  XNOR U4566 ( .A(n1470), .B(n1469), .Z(n1483) );
  IV U4567 ( .A(n1475), .Z(n1529) );
  XNOR U4568 ( .A(n1529), .B(n1471), .Z(n1536) );
  AND U4569 ( .A(n1525), .B(n1536), .Z(n1473) );
  AND U4570 ( .A(x[64]), .B(n1540), .Z(n1472) );
  XNOR U4571 ( .A(n1473), .B(n1472), .Z(n1474) );
  NANDN U4572 ( .A(n1526), .B(n1474), .Z(n1478) );
  NAND U4573 ( .A(x[64]), .B(n1525), .Z(n1476) );
  OR U4574 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U4575 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4576 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR U4577 ( .A(n1483), .B(n1481), .Z(n1503) );
  IV U4578 ( .A(n1503), .Z(n1510) );
  AND U4579 ( .A(n1556), .B(n1482), .Z(n1485) );
  XOR U4580 ( .A(x[65]), .B(x[71]), .Z(n1558) );
  AND U4581 ( .A(n1519), .B(n1558), .Z(n1488) );
  XNOR U4582 ( .A(n1488), .B(n1483), .Z(n1484) );
  XNOR U4583 ( .A(n1485), .B(n1484), .Z(n1509) );
  NANDN U4584 ( .A(n1510), .B(n1509), .Z(n1486) );
  NAND U4585 ( .A(n1514), .B(n1486), .Z(n1496) );
  XNOR U4586 ( .A(n1488), .B(n1487), .Z(n1493) );
  ANDN U4587 ( .B(n1489), .A(x[65]), .Z(n1490) );
  XNOR U4588 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U4589 ( .A(n1493), .B(n1492), .Z(n1506) );
  XOR U4590 ( .A(n1509), .B(n1506), .Z(n1494) );
  NAND U4591 ( .A(n1510), .B(n1494), .Z(n1495) );
  NAND U4592 ( .A(n1496), .B(n1495), .Z(n1555) );
  ANDN U4593 ( .B(n1497), .A(n1555), .Z(n1521) );
  IV U4594 ( .A(n1506), .Z(n1512) );
  XOR U4595 ( .A(n1514), .B(n1510), .Z(n1498) );
  NANDN U4596 ( .A(n1512), .B(n1498), .Z(n1501) );
  NANDN U4597 ( .A(n1510), .B(n1512), .Z(n1499) );
  NANDN U4598 ( .A(n1509), .B(n1499), .Z(n1500) );
  NAND U4599 ( .A(n1501), .B(n1500), .Z(n1565) );
  XNOR U4600 ( .A(n1555), .B(n1565), .Z(n1531) );
  AND U4601 ( .A(n1502), .B(n1531), .Z(n1524) );
  OR U4602 ( .A(n1509), .B(n1506), .Z(n1508) );
  ANDN U4603 ( .B(n1509), .A(n1503), .Z(n1504) );
  XNOR U4604 ( .A(n1504), .B(n1514), .Z(n1505) );
  NAND U4605 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U4606 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U4607 ( .A(n1510), .B(n1514), .Z(n1516) );
  NAND U4608 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4609 ( .A(n1512), .B(n1511), .Z(n1513) );
  NANDN U4610 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U4611 ( .A(n1516), .B(n1515), .Z(n1572) );
  NAND U4612 ( .A(n1547), .B(n1517), .Z(n1518) );
  XNOR U4613 ( .A(n1524), .B(n1518), .Z(n1567) );
  XOR U4614 ( .A(n1555), .B(n1572), .Z(n1557) );
  AND U4615 ( .A(n1519), .B(n1557), .Z(n1542) );
  XNOR U4616 ( .A(n1567), .B(n1542), .Z(n1520) );
  XNOR U4617 ( .A(n1521), .B(n1520), .Z(n1575) );
  NAND U4618 ( .A(n1533), .B(n1522), .Z(n1523) );
  XNOR U4619 ( .A(n1524), .B(n1523), .Z(n1550) );
  AND U4620 ( .A(n1525), .B(n1535), .Z(n1566) );
  NANDN U4621 ( .A(n1526), .B(n1528), .Z(n1527) );
  XNOR U4622 ( .A(n1566), .B(n1527), .Z(n1554) );
  XNOR U4623 ( .A(n1550), .B(n1554), .Z(n1539) );
  XOR U4624 ( .A(n1575), .B(n1539), .Z(z[64]) );
  AND U4625 ( .A(n1529), .B(n1528), .Z(n1538) );
  AND U4626 ( .A(n1531), .B(n1530), .Z(n1549) );
  NAND U4627 ( .A(n1533), .B(n1532), .Z(n1534) );
  XNOR U4628 ( .A(n1549), .B(n1534), .Z(n1576) );
  AND U4629 ( .A(n1536), .B(n1535), .Z(n1543) );
  XNOR U4630 ( .A(n1576), .B(n1543), .Z(n1537) );
  XNOR U4631 ( .A(n1538), .B(n1537), .Z(n1563) );
  XNOR U4632 ( .A(n1563), .B(n1539), .Z(n1583) );
  AND U4633 ( .A(n1540), .B(n1565), .Z(n1545) );
  NANDN U4634 ( .A(n1572), .B(n1570), .Z(n1541) );
  XNOR U4635 ( .A(n1542), .B(n1541), .Z(n1553) );
  XNOR U4636 ( .A(n1543), .B(n1553), .Z(n1544) );
  XNOR U4637 ( .A(n1545), .B(n1544), .Z(n1552) );
  NAND U4638 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U4639 ( .A(n1549), .B(n1548), .Z(n1559) );
  XNOR U4640 ( .A(n1550), .B(n1559), .Z(n1551) );
  XNOR U4641 ( .A(n1552), .B(n1551), .Z(n1562) );
  XNOR U4642 ( .A(n1583), .B(n1562), .Z(z[65]) );
  XNOR U4643 ( .A(n1554), .B(n1553), .Z(z[66]) );
  NOR U4644 ( .A(n1556), .B(n1555), .Z(n1561) );
  AND U4645 ( .A(n1558), .B(n1557), .Z(n1574) );
  XNOR U4646 ( .A(n1559), .B(n1574), .Z(n1560) );
  XNOR U4647 ( .A(n1561), .B(n1560), .Z(n1582) );
  XOR U4648 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U4649 ( .A(n1582), .B(n1564), .Z(z[67]) );
  XOR U4650 ( .A(n1575), .B(z[66]), .Z(z[68]) );
  AND U4651 ( .A(x[64]), .B(n1565), .Z(n1569) );
  XNOR U4652 ( .A(n1567), .B(n1566), .Z(n1568) );
  XNOR U4653 ( .A(n1569), .B(n1568), .Z(n1584) );
  XOR U4654 ( .A(n1570), .B(x[65]), .Z(n1571) );
  NANDN U4655 ( .A(n1572), .B(n1571), .Z(n1573) );
  XNOR U4656 ( .A(n1574), .B(n1573), .Z(n1578) );
  XNOR U4657 ( .A(n1576), .B(n1575), .Z(n1577) );
  XNOR U4658 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U4659 ( .A(n1584), .B(n1579), .Z(z[69]) );
  XNOR U4660 ( .A(n1581), .B(n1580), .Z(z[6]) );
  XNOR U4661 ( .A(n1583), .B(n1582), .Z(z[70]) );
  XOR U4662 ( .A(n1584), .B(z[65]), .Z(z[71]) );
  XOR U4663 ( .A(x[75]), .B(x[73]), .Z(n1587) );
  XNOR U4664 ( .A(x[72]), .B(x[78]), .Z(n1586) );
  XOR U4665 ( .A(n1586), .B(x[74]), .Z(n1585) );
  XNOR U4666 ( .A(n1587), .B(n1585), .Z(n1622) );
  XNOR U4667 ( .A(x[77]), .B(n1586), .Z(n1695) );
  XOR U4668 ( .A(n1695), .B(x[76]), .Z(n1665) );
  IV U4669 ( .A(n1665), .Z(n1596) );
  XNOR U4670 ( .A(x[79]), .B(x[76]), .Z(n1590) );
  XNOR U4671 ( .A(n1587), .B(n1590), .Z(n1650) );
  NOR U4672 ( .A(n1596), .B(n1650), .Z(n1589) );
  XNOR U4673 ( .A(n1695), .B(x[79]), .Z(n1681) );
  XNOR U4674 ( .A(x[74]), .B(n1681), .Z(n1605) );
  XNOR U4675 ( .A(x[73]), .B(n1605), .Z(n1600) );
  AND U4676 ( .A(x[72]), .B(n1600), .Z(n1588) );
  XNOR U4677 ( .A(n1589), .B(n1588), .Z(n1593) );
  XNOR U4678 ( .A(n1622), .B(n1681), .Z(n1612) );
  IV U4679 ( .A(n1622), .Z(n1607) );
  XNOR U4680 ( .A(x[72]), .B(n1607), .Z(n1627) );
  IV U4681 ( .A(n1590), .Z(n1655) );
  AND U4682 ( .A(n1627), .B(n1655), .Z(n1595) );
  IV U4683 ( .A(n1695), .Z(n1614) );
  XNOR U4684 ( .A(n1622), .B(n1614), .Z(n1644) );
  XOR U4685 ( .A(n1644), .B(n1650), .Z(n1647) );
  XOR U4686 ( .A(x[74]), .B(x[76]), .Z(n1657) );
  NAND U4687 ( .A(n1647), .B(n1657), .Z(n1591) );
  XNOR U4688 ( .A(n1595), .B(n1591), .Z(n1616) );
  XNOR U4689 ( .A(n1612), .B(n1616), .Z(n1592) );
  XNOR U4690 ( .A(n1593), .B(n1592), .Z(n1639) );
  XOR U4691 ( .A(x[74]), .B(x[79]), .Z(n1671) );
  XNOR U4692 ( .A(x[72]), .B(n1650), .Z(n1651) );
  XNOR U4693 ( .A(n1695), .B(n1651), .Z(n1642) );
  NAND U4694 ( .A(n1671), .B(n1642), .Z(n1594) );
  XNOR U4695 ( .A(n1595), .B(n1594), .Z(n1608) );
  IV U4696 ( .A(n1600), .Z(n1654) );
  XNOR U4697 ( .A(n1654), .B(n1596), .Z(n1661) );
  AND U4698 ( .A(n1650), .B(n1661), .Z(n1598) );
  AND U4699 ( .A(x[72]), .B(n1665), .Z(n1597) );
  XNOR U4700 ( .A(n1598), .B(n1597), .Z(n1599) );
  NANDN U4701 ( .A(n1651), .B(n1599), .Z(n1603) );
  NAND U4702 ( .A(x[72]), .B(n1650), .Z(n1601) );
  OR U4703 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U4704 ( .A(n1603), .B(n1602), .Z(n1604) );
  XNOR U4705 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U4706 ( .A(n1608), .B(n1606), .Z(n1628) );
  IV U4707 ( .A(n1628), .Z(n1635) );
  AND U4708 ( .A(n1681), .B(n1607), .Z(n1610) );
  XOR U4709 ( .A(x[73]), .B(x[79]), .Z(n1683) );
  AND U4710 ( .A(n1644), .B(n1683), .Z(n1613) );
  XNOR U4711 ( .A(n1613), .B(n1608), .Z(n1609) );
  XNOR U4712 ( .A(n1610), .B(n1609), .Z(n1634) );
  NANDN U4713 ( .A(n1635), .B(n1634), .Z(n1611) );
  NAND U4714 ( .A(n1639), .B(n1611), .Z(n1621) );
  XNOR U4715 ( .A(n1613), .B(n1612), .Z(n1618) );
  ANDN U4716 ( .B(n1614), .A(x[73]), .Z(n1615) );
  XNOR U4717 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4718 ( .A(n1618), .B(n1617), .Z(n1631) );
  XOR U4719 ( .A(n1634), .B(n1631), .Z(n1619) );
  NAND U4720 ( .A(n1635), .B(n1619), .Z(n1620) );
  NAND U4721 ( .A(n1621), .B(n1620), .Z(n1680) );
  ANDN U4722 ( .B(n1622), .A(n1680), .Z(n1646) );
  IV U4723 ( .A(n1631), .Z(n1637) );
  XOR U4724 ( .A(n1639), .B(n1635), .Z(n1623) );
  NANDN U4725 ( .A(n1637), .B(n1623), .Z(n1626) );
  NANDN U4726 ( .A(n1635), .B(n1637), .Z(n1624) );
  NANDN U4727 ( .A(n1634), .B(n1624), .Z(n1625) );
  NAND U4728 ( .A(n1626), .B(n1625), .Z(n1690) );
  XNOR U4729 ( .A(n1680), .B(n1690), .Z(n1656) );
  AND U4730 ( .A(n1627), .B(n1656), .Z(n1649) );
  OR U4731 ( .A(n1634), .B(n1631), .Z(n1633) );
  ANDN U4732 ( .B(n1634), .A(n1628), .Z(n1629) );
  XNOR U4733 ( .A(n1629), .B(n1639), .Z(n1630) );
  NAND U4734 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U4735 ( .A(n1633), .B(n1632), .Z(n1653) );
  NAND U4736 ( .A(n1635), .B(n1639), .Z(n1641) );
  NAND U4737 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U4738 ( .A(n1637), .B(n1636), .Z(n1638) );
  NANDN U4739 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U4740 ( .A(n1641), .B(n1640), .Z(n1697) );
  NAND U4741 ( .A(n1672), .B(n1642), .Z(n1643) );
  XNOR U4742 ( .A(n1649), .B(n1643), .Z(n1692) );
  XOR U4743 ( .A(n1680), .B(n1697), .Z(n1682) );
  AND U4744 ( .A(n1644), .B(n1682), .Z(n1667) );
  XNOR U4745 ( .A(n1692), .B(n1667), .Z(n1645) );
  XNOR U4746 ( .A(n1646), .B(n1645), .Z(n1700) );
  NAND U4747 ( .A(n1658), .B(n1647), .Z(n1648) );
  XNOR U4748 ( .A(n1649), .B(n1648), .Z(n1675) );
  AND U4749 ( .A(n1650), .B(n1660), .Z(n1691) );
  NANDN U4750 ( .A(n1651), .B(n1653), .Z(n1652) );
  XNOR U4751 ( .A(n1691), .B(n1652), .Z(n1679) );
  XNOR U4752 ( .A(n1675), .B(n1679), .Z(n1664) );
  XOR U4753 ( .A(n1700), .B(n1664), .Z(z[72]) );
  AND U4754 ( .A(n1654), .B(n1653), .Z(n1663) );
  AND U4755 ( .A(n1656), .B(n1655), .Z(n1674) );
  NAND U4756 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U4757 ( .A(n1674), .B(n1659), .Z(n1701) );
  AND U4758 ( .A(n1661), .B(n1660), .Z(n1668) );
  XNOR U4759 ( .A(n1701), .B(n1668), .Z(n1662) );
  XNOR U4760 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U4761 ( .A(n1688), .B(n1664), .Z(n1706) );
  AND U4762 ( .A(n1665), .B(n1690), .Z(n1670) );
  NANDN U4763 ( .A(n1697), .B(n1695), .Z(n1666) );
  XNOR U4764 ( .A(n1667), .B(n1666), .Z(n1678) );
  XNOR U4765 ( .A(n1668), .B(n1678), .Z(n1669) );
  XNOR U4766 ( .A(n1670), .B(n1669), .Z(n1677) );
  NAND U4767 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR U4768 ( .A(n1674), .B(n1673), .Z(n1684) );
  XNOR U4769 ( .A(n1675), .B(n1684), .Z(n1676) );
  XNOR U4770 ( .A(n1677), .B(n1676), .Z(n1687) );
  XNOR U4771 ( .A(n1706), .B(n1687), .Z(z[73]) );
  XNOR U4772 ( .A(n1679), .B(n1678), .Z(z[74]) );
  NOR U4773 ( .A(n1681), .B(n1680), .Z(n1686) );
  AND U4774 ( .A(n1683), .B(n1682), .Z(n1699) );
  XNOR U4775 ( .A(n1684), .B(n1699), .Z(n1685) );
  XNOR U4776 ( .A(n1686), .B(n1685), .Z(n1705) );
  XOR U4777 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4778 ( .A(n1705), .B(n1689), .Z(z[75]) );
  XOR U4779 ( .A(n1700), .B(z[74]), .Z(z[76]) );
  AND U4780 ( .A(x[72]), .B(n1690), .Z(n1694) );
  XNOR U4781 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4782 ( .A(n1694), .B(n1693), .Z(n1707) );
  XOR U4783 ( .A(n1695), .B(x[73]), .Z(n1696) );
  NANDN U4784 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U4785 ( .A(n1699), .B(n1698), .Z(n1703) );
  XNOR U4786 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U4787 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U4788 ( .A(n1707), .B(n1704), .Z(z[77]) );
  XNOR U4789 ( .A(n1706), .B(n1705), .Z(z[78]) );
  XOR U4790 ( .A(n1707), .B(z[73]), .Z(z[79]) );
  XOR U4791 ( .A(n1708), .B(z[1]), .Z(z[7]) );
  XOR U4792 ( .A(x[83]), .B(x[81]), .Z(n1711) );
  XNOR U4793 ( .A(x[80]), .B(x[86]), .Z(n1710) );
  XOR U4794 ( .A(n1710), .B(x[82]), .Z(n1709) );
  XNOR U4795 ( .A(n1711), .B(n1709), .Z(n1746) );
  XNOR U4796 ( .A(x[85]), .B(n1710), .Z(n1819) );
  XOR U4797 ( .A(n1819), .B(x[84]), .Z(n1789) );
  IV U4798 ( .A(n1789), .Z(n1720) );
  XNOR U4799 ( .A(x[87]), .B(x[84]), .Z(n1714) );
  XNOR U4800 ( .A(n1711), .B(n1714), .Z(n1774) );
  NOR U4801 ( .A(n1720), .B(n1774), .Z(n1713) );
  XNOR U4802 ( .A(n1819), .B(x[87]), .Z(n1805) );
  XNOR U4803 ( .A(x[82]), .B(n1805), .Z(n1729) );
  XNOR U4804 ( .A(x[81]), .B(n1729), .Z(n1724) );
  AND U4805 ( .A(x[80]), .B(n1724), .Z(n1712) );
  XNOR U4806 ( .A(n1713), .B(n1712), .Z(n1717) );
  XNOR U4807 ( .A(n1746), .B(n1805), .Z(n1736) );
  IV U4808 ( .A(n1746), .Z(n1731) );
  XNOR U4809 ( .A(x[80]), .B(n1731), .Z(n1751) );
  IV U4810 ( .A(n1714), .Z(n1779) );
  AND U4811 ( .A(n1751), .B(n1779), .Z(n1719) );
  IV U4812 ( .A(n1819), .Z(n1738) );
  XNOR U4813 ( .A(n1746), .B(n1738), .Z(n1768) );
  XOR U4814 ( .A(n1768), .B(n1774), .Z(n1771) );
  XOR U4815 ( .A(x[82]), .B(x[84]), .Z(n1781) );
  NAND U4816 ( .A(n1771), .B(n1781), .Z(n1715) );
  XNOR U4817 ( .A(n1719), .B(n1715), .Z(n1740) );
  XNOR U4818 ( .A(n1736), .B(n1740), .Z(n1716) );
  XNOR U4819 ( .A(n1717), .B(n1716), .Z(n1763) );
  XOR U4820 ( .A(x[82]), .B(x[87]), .Z(n1795) );
  XNOR U4821 ( .A(x[80]), .B(n1774), .Z(n1775) );
  XNOR U4822 ( .A(n1819), .B(n1775), .Z(n1766) );
  NAND U4823 ( .A(n1795), .B(n1766), .Z(n1718) );
  XNOR U4824 ( .A(n1719), .B(n1718), .Z(n1732) );
  IV U4825 ( .A(n1724), .Z(n1778) );
  XNOR U4826 ( .A(n1778), .B(n1720), .Z(n1785) );
  AND U4827 ( .A(n1774), .B(n1785), .Z(n1722) );
  AND U4828 ( .A(x[80]), .B(n1789), .Z(n1721) );
  XNOR U4829 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U4830 ( .A(n1775), .B(n1723), .Z(n1727) );
  NAND U4831 ( .A(x[80]), .B(n1774), .Z(n1725) );
  OR U4832 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U4833 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U4834 ( .A(n1729), .B(n1728), .Z(n1730) );
  XNOR U4835 ( .A(n1732), .B(n1730), .Z(n1752) );
  IV U4836 ( .A(n1752), .Z(n1759) );
  AND U4837 ( .A(n1805), .B(n1731), .Z(n1734) );
  XOR U4838 ( .A(x[81]), .B(x[87]), .Z(n1807) );
  AND U4839 ( .A(n1768), .B(n1807), .Z(n1737) );
  XNOR U4840 ( .A(n1737), .B(n1732), .Z(n1733) );
  XNOR U4841 ( .A(n1734), .B(n1733), .Z(n1758) );
  NANDN U4842 ( .A(n1759), .B(n1758), .Z(n1735) );
  NAND U4843 ( .A(n1763), .B(n1735), .Z(n1745) );
  XNOR U4844 ( .A(n1737), .B(n1736), .Z(n1742) );
  ANDN U4845 ( .B(n1738), .A(x[81]), .Z(n1739) );
  XNOR U4846 ( .A(n1740), .B(n1739), .Z(n1741) );
  XNOR U4847 ( .A(n1742), .B(n1741), .Z(n1755) );
  XOR U4848 ( .A(n1758), .B(n1755), .Z(n1743) );
  NAND U4849 ( .A(n1759), .B(n1743), .Z(n1744) );
  NAND U4850 ( .A(n1745), .B(n1744), .Z(n1804) );
  ANDN U4851 ( .B(n1746), .A(n1804), .Z(n1770) );
  IV U4852 ( .A(n1755), .Z(n1761) );
  XOR U4853 ( .A(n1763), .B(n1759), .Z(n1747) );
  NANDN U4854 ( .A(n1761), .B(n1747), .Z(n1750) );
  NANDN U4855 ( .A(n1759), .B(n1761), .Z(n1748) );
  NANDN U4856 ( .A(n1758), .B(n1748), .Z(n1749) );
  NAND U4857 ( .A(n1750), .B(n1749), .Z(n1814) );
  XNOR U4858 ( .A(n1804), .B(n1814), .Z(n1780) );
  AND U4859 ( .A(n1751), .B(n1780), .Z(n1773) );
  OR U4860 ( .A(n1758), .B(n1755), .Z(n1757) );
  ANDN U4861 ( .B(n1758), .A(n1752), .Z(n1753) );
  XNOR U4862 ( .A(n1753), .B(n1763), .Z(n1754) );
  NAND U4863 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U4864 ( .A(n1757), .B(n1756), .Z(n1777) );
  NAND U4865 ( .A(n1759), .B(n1763), .Z(n1765) );
  NAND U4866 ( .A(n1759), .B(n1758), .Z(n1760) );
  XNOR U4867 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U4868 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1821) );
  NAND U4870 ( .A(n1796), .B(n1766), .Z(n1767) );
  XNOR U4871 ( .A(n1773), .B(n1767), .Z(n1816) );
  XOR U4872 ( .A(n1804), .B(n1821), .Z(n1806) );
  AND U4873 ( .A(n1768), .B(n1806), .Z(n1791) );
  XNOR U4874 ( .A(n1816), .B(n1791), .Z(n1769) );
  XNOR U4875 ( .A(n1770), .B(n1769), .Z(n1824) );
  NAND U4876 ( .A(n1782), .B(n1771), .Z(n1772) );
  XNOR U4877 ( .A(n1773), .B(n1772), .Z(n1799) );
  AND U4878 ( .A(n1774), .B(n1784), .Z(n1815) );
  NANDN U4879 ( .A(n1775), .B(n1777), .Z(n1776) );
  XNOR U4880 ( .A(n1815), .B(n1776), .Z(n1803) );
  XNOR U4881 ( .A(n1799), .B(n1803), .Z(n1788) );
  XOR U4882 ( .A(n1824), .B(n1788), .Z(z[80]) );
  AND U4883 ( .A(n1778), .B(n1777), .Z(n1787) );
  AND U4884 ( .A(n1780), .B(n1779), .Z(n1798) );
  NAND U4885 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U4886 ( .A(n1798), .B(n1783), .Z(n1825) );
  AND U4887 ( .A(n1785), .B(n1784), .Z(n1792) );
  XNOR U4888 ( .A(n1825), .B(n1792), .Z(n1786) );
  XNOR U4889 ( .A(n1787), .B(n1786), .Z(n1812) );
  XNOR U4890 ( .A(n1812), .B(n1788), .Z(n1830) );
  AND U4891 ( .A(n1789), .B(n1814), .Z(n1794) );
  NANDN U4892 ( .A(n1821), .B(n1819), .Z(n1790) );
  XNOR U4893 ( .A(n1791), .B(n1790), .Z(n1802) );
  XNOR U4894 ( .A(n1792), .B(n1802), .Z(n1793) );
  XNOR U4895 ( .A(n1794), .B(n1793), .Z(n1801) );
  NAND U4896 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U4897 ( .A(n1798), .B(n1797), .Z(n1808) );
  XNOR U4898 ( .A(n1799), .B(n1808), .Z(n1800) );
  XNOR U4899 ( .A(n1801), .B(n1800), .Z(n1811) );
  XNOR U4900 ( .A(n1830), .B(n1811), .Z(z[81]) );
  XNOR U4901 ( .A(n1803), .B(n1802), .Z(z[82]) );
  NOR U4902 ( .A(n1805), .B(n1804), .Z(n1810) );
  AND U4903 ( .A(n1807), .B(n1806), .Z(n1823) );
  XNOR U4904 ( .A(n1808), .B(n1823), .Z(n1809) );
  XNOR U4905 ( .A(n1810), .B(n1809), .Z(n1829) );
  XOR U4906 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U4907 ( .A(n1829), .B(n1813), .Z(z[83]) );
  XOR U4908 ( .A(n1824), .B(z[82]), .Z(z[84]) );
  AND U4909 ( .A(x[80]), .B(n1814), .Z(n1818) );
  XNOR U4910 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U4911 ( .A(n1818), .B(n1817), .Z(n1831) );
  XOR U4912 ( .A(n1819), .B(x[81]), .Z(n1820) );
  NANDN U4913 ( .A(n1821), .B(n1820), .Z(n1822) );
  XNOR U4914 ( .A(n1823), .B(n1822), .Z(n1827) );
  XNOR U4915 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U4916 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U4917 ( .A(n1831), .B(n1828), .Z(z[85]) );
  XNOR U4918 ( .A(n1830), .B(n1829), .Z(z[86]) );
  XOR U4919 ( .A(n1831), .B(z[81]), .Z(z[87]) );
  XOR U4920 ( .A(x[91]), .B(x[89]), .Z(n1834) );
  XNOR U4921 ( .A(x[88]), .B(x[94]), .Z(n1833) );
  XOR U4922 ( .A(n1833), .B(x[90]), .Z(n1832) );
  XNOR U4923 ( .A(n1834), .B(n1832), .Z(n1869) );
  XNOR U4924 ( .A(x[93]), .B(n1833), .Z(n1944) );
  XOR U4925 ( .A(n1944), .B(x[92]), .Z(n1912) );
  IV U4926 ( .A(n1912), .Z(n1843) );
  XNOR U4927 ( .A(x[95]), .B(x[92]), .Z(n1837) );
  XNOR U4928 ( .A(n1834), .B(n1837), .Z(n1897) );
  NOR U4929 ( .A(n1843), .B(n1897), .Z(n1836) );
  XNOR U4930 ( .A(n1944), .B(x[95]), .Z(n1930) );
  XNOR U4931 ( .A(x[90]), .B(n1930), .Z(n1852) );
  XNOR U4932 ( .A(x[89]), .B(n1852), .Z(n1847) );
  AND U4933 ( .A(x[88]), .B(n1847), .Z(n1835) );
  XNOR U4934 ( .A(n1836), .B(n1835), .Z(n1840) );
  XNOR U4935 ( .A(n1869), .B(n1930), .Z(n1859) );
  IV U4936 ( .A(n1869), .Z(n1854) );
  XNOR U4937 ( .A(x[88]), .B(n1854), .Z(n1874) );
  IV U4938 ( .A(n1837), .Z(n1902) );
  AND U4939 ( .A(n1874), .B(n1902), .Z(n1842) );
  IV U4940 ( .A(n1944), .Z(n1861) );
  XNOR U4941 ( .A(n1869), .B(n1861), .Z(n1891) );
  XOR U4942 ( .A(n1891), .B(n1897), .Z(n1894) );
  XOR U4943 ( .A(x[90]), .B(x[92]), .Z(n1904) );
  NAND U4944 ( .A(n1894), .B(n1904), .Z(n1838) );
  XNOR U4945 ( .A(n1842), .B(n1838), .Z(n1863) );
  XNOR U4946 ( .A(n1859), .B(n1863), .Z(n1839) );
  XNOR U4947 ( .A(n1840), .B(n1839), .Z(n1886) );
  XOR U4948 ( .A(x[90]), .B(x[95]), .Z(n1918) );
  XNOR U4949 ( .A(x[88]), .B(n1897), .Z(n1898) );
  XNOR U4950 ( .A(n1944), .B(n1898), .Z(n1889) );
  NAND U4951 ( .A(n1918), .B(n1889), .Z(n1841) );
  XNOR U4952 ( .A(n1842), .B(n1841), .Z(n1855) );
  IV U4953 ( .A(n1847), .Z(n1901) );
  XNOR U4954 ( .A(n1901), .B(n1843), .Z(n1908) );
  AND U4955 ( .A(n1897), .B(n1908), .Z(n1845) );
  AND U4956 ( .A(x[88]), .B(n1912), .Z(n1844) );
  XNOR U4957 ( .A(n1845), .B(n1844), .Z(n1846) );
  NANDN U4958 ( .A(n1898), .B(n1846), .Z(n1850) );
  NAND U4959 ( .A(x[88]), .B(n1897), .Z(n1848) );
  OR U4960 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U4961 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U4962 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U4963 ( .A(n1855), .B(n1853), .Z(n1875) );
  IV U4964 ( .A(n1875), .Z(n1882) );
  AND U4965 ( .A(n1930), .B(n1854), .Z(n1857) );
  XOR U4966 ( .A(x[89]), .B(x[95]), .Z(n1932) );
  AND U4967 ( .A(n1891), .B(n1932), .Z(n1860) );
  XNOR U4968 ( .A(n1860), .B(n1855), .Z(n1856) );
  XNOR U4969 ( .A(n1857), .B(n1856), .Z(n1881) );
  NANDN U4970 ( .A(n1882), .B(n1881), .Z(n1858) );
  NAND U4971 ( .A(n1886), .B(n1858), .Z(n1868) );
  XNOR U4972 ( .A(n1860), .B(n1859), .Z(n1865) );
  ANDN U4973 ( .B(n1861), .A(x[89]), .Z(n1862) );
  XNOR U4974 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U4975 ( .A(n1865), .B(n1864), .Z(n1878) );
  XOR U4976 ( .A(n1881), .B(n1878), .Z(n1866) );
  NAND U4977 ( .A(n1882), .B(n1866), .Z(n1867) );
  NAND U4978 ( .A(n1868), .B(n1867), .Z(n1929) );
  ANDN U4979 ( .B(n1869), .A(n1929), .Z(n1893) );
  IV U4980 ( .A(n1878), .Z(n1884) );
  XOR U4981 ( .A(n1886), .B(n1882), .Z(n1870) );
  NANDN U4982 ( .A(n1884), .B(n1870), .Z(n1873) );
  NANDN U4983 ( .A(n1882), .B(n1884), .Z(n1871) );
  NANDN U4984 ( .A(n1881), .B(n1871), .Z(n1872) );
  NAND U4985 ( .A(n1873), .B(n1872), .Z(n1939) );
  XNOR U4986 ( .A(n1929), .B(n1939), .Z(n1903) );
  AND U4987 ( .A(n1874), .B(n1903), .Z(n1896) );
  OR U4988 ( .A(n1881), .B(n1878), .Z(n1880) );
  ANDN U4989 ( .B(n1881), .A(n1875), .Z(n1876) );
  XNOR U4990 ( .A(n1876), .B(n1886), .Z(n1877) );
  NAND U4991 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U4992 ( .A(n1880), .B(n1879), .Z(n1900) );
  NAND U4993 ( .A(n1882), .B(n1886), .Z(n1888) );
  NAND U4994 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U4995 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U4996 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4997 ( .A(n1888), .B(n1887), .Z(n1946) );
  NAND U4998 ( .A(n1919), .B(n1889), .Z(n1890) );
  XNOR U4999 ( .A(n1896), .B(n1890), .Z(n1941) );
  XOR U5000 ( .A(n1929), .B(n1946), .Z(n1931) );
  AND U5001 ( .A(n1891), .B(n1931), .Z(n1914) );
  XNOR U5002 ( .A(n1941), .B(n1914), .Z(n1892) );
  XNOR U5003 ( .A(n1893), .B(n1892), .Z(n1949) );
  NAND U5004 ( .A(n1905), .B(n1894), .Z(n1895) );
  XNOR U5005 ( .A(n1896), .B(n1895), .Z(n1922) );
  AND U5006 ( .A(n1897), .B(n1907), .Z(n1940) );
  NANDN U5007 ( .A(n1898), .B(n1900), .Z(n1899) );
  XNOR U5008 ( .A(n1940), .B(n1899), .Z(n1928) );
  XNOR U5009 ( .A(n1922), .B(n1928), .Z(n1911) );
  XOR U5010 ( .A(n1949), .B(n1911), .Z(z[88]) );
  AND U5011 ( .A(n1901), .B(n1900), .Z(n1910) );
  AND U5012 ( .A(n1903), .B(n1902), .Z(n1921) );
  NAND U5013 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U5014 ( .A(n1921), .B(n1906), .Z(n1950) );
  AND U5015 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U5016 ( .A(n1950), .B(n1915), .Z(n1909) );
  XNOR U5017 ( .A(n1910), .B(n1909), .Z(n1937) );
  XNOR U5018 ( .A(n1937), .B(n1911), .Z(n1955) );
  AND U5019 ( .A(n1912), .B(n1939), .Z(n1917) );
  NANDN U5020 ( .A(n1946), .B(n1944), .Z(n1913) );
  XNOR U5021 ( .A(n1914), .B(n1913), .Z(n1927) );
  XNOR U5022 ( .A(n1915), .B(n1927), .Z(n1916) );
  XNOR U5023 ( .A(n1917), .B(n1916), .Z(n1924) );
  NAND U5024 ( .A(n1919), .B(n1918), .Z(n1920) );
  XNOR U5025 ( .A(n1921), .B(n1920), .Z(n1933) );
  XNOR U5026 ( .A(n1922), .B(n1933), .Z(n1923) );
  XNOR U5027 ( .A(n1924), .B(n1923), .Z(n1936) );
  XNOR U5028 ( .A(n1955), .B(n1936), .Z(z[89]) );
  XOR U5029 ( .A(n1926), .B(n1925), .Z(z[8]) );
  XNOR U5030 ( .A(n1928), .B(n1927), .Z(z[90]) );
  NOR U5031 ( .A(n1930), .B(n1929), .Z(n1935) );
  AND U5032 ( .A(n1932), .B(n1931), .Z(n1948) );
  XNOR U5033 ( .A(n1933), .B(n1948), .Z(n1934) );
  XNOR U5034 ( .A(n1935), .B(n1934), .Z(n1954) );
  XOR U5035 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U5036 ( .A(n1954), .B(n1938), .Z(z[91]) );
  XOR U5037 ( .A(n1949), .B(z[90]), .Z(z[92]) );
  AND U5038 ( .A(x[88]), .B(n1939), .Z(n1943) );
  XNOR U5039 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5040 ( .A(n1943), .B(n1942), .Z(n1956) );
  XOR U5041 ( .A(n1944), .B(x[89]), .Z(n1945) );
  NANDN U5042 ( .A(n1946), .B(n1945), .Z(n1947) );
  XNOR U5043 ( .A(n1948), .B(n1947), .Z(n1952) );
  XNOR U5044 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U5045 ( .A(n1952), .B(n1951), .Z(n1953) );
  XNOR U5046 ( .A(n1956), .B(n1953), .Z(z[93]) );
  XNOR U5047 ( .A(n1955), .B(n1954), .Z(z[94]) );
  XOR U5048 ( .A(n1956), .B(z[89]), .Z(z[95]) );
  XOR U5049 ( .A(n1958), .B(n1957), .Z(z[96]) );
  XOR U5050 ( .A(n1960), .B(n1959), .Z(n1961) );
  XNOR U5051 ( .A(n1962), .B(n1961), .Z(z[99]) );
endmodule


module SubBytes_4 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;

  XOR U2962 ( .A(n923), .B(n886), .Z(n893) );
  XOR U2963 ( .A(n1048), .B(n1011), .Z(n1018) );
  XNOR U2964 ( .A(n430), .B(n474), .Z(n449) );
  XOR U2965 ( .A(n1690), .B(n1653), .Z(n1660) );
  XOR U2966 ( .A(n1442), .B(n1390), .Z(n1397) );
  XNOR U2967 ( .A(n1528), .B(n1572), .Z(n1547) );
  XNOR U2968 ( .A(n253), .B(n297), .Z(n272) );
  XOR U2969 ( .A(n800), .B(n738), .Z(n745) );
  XNOR U2970 ( .A(n1900), .B(n1946), .Z(n1919) );
  XNOR U2971 ( .A(n1267), .B(n1311), .Z(n1286) );
  XNOR U2972 ( .A(n775), .B(n1434), .Z(n794) );
  XOR U2973 ( .A(n1814), .B(n1777), .Z(n1784) );
  XOR U2974 ( .A(n1181), .B(n1144), .Z(n1151) );
  XOR U2975 ( .A(n622), .B(n585), .Z(n592) );
  XNOR U2976 ( .A(n886), .B(n930), .Z(n905) );
  XNOR U2977 ( .A(n1011), .B(n1055), .Z(n1030) );
  XOR U2978 ( .A(n467), .B(n430), .Z(n437) );
  XNOR U2979 ( .A(n1653), .B(n1697), .Z(n1672) );
  XNOR U2980 ( .A(n1390), .B(n1449), .Z(n1409) );
  XOR U2981 ( .A(n290), .B(n253), .Z(n260) );
  XOR U2982 ( .A(n1565), .B(n1528), .Z(n1535) );
  XNOR U2983 ( .A(n738), .B(n807), .Z(n757) );
  NOR U2984 ( .A(n654), .B(x[9]), .Z(n1) );
  XNOR U2985 ( .A(n329), .B(n328), .Z(n2) );
  XNOR U2986 ( .A(n1), .B(n2), .Z(n3) );
  XNOR U2987 ( .A(n312), .B(n3), .Z(n345) );
  XOR U2988 ( .A(n1304), .B(n1267), .Z(n1274) );
  XOR U2989 ( .A(n1939), .B(n1900), .Z(n1907) );
  XOR U2990 ( .A(n1427), .B(n775), .Z(n782) );
  XNOR U2991 ( .A(n1777), .B(n1821), .Z(n1796) );
  XNOR U2992 ( .A(n1144), .B(n1188), .Z(n1163) );
  XNOR U2993 ( .A(n585), .B(n629), .Z(n604) );
  XOR U2994 ( .A(n163), .B(n134), .Z(n157) );
  XOR U2995 ( .A(n77), .B(n78), .Z(n129) );
  XNOR U2996 ( .A(x[9]), .B(n323), .Z(n318) );
  XOR U2997 ( .A(n794), .B(n778), .Z(n780) );
  XOR U2998 ( .A(n604), .B(n588), .Z(n590) );
  XOR U2999 ( .A(n1030), .B(n1014), .Z(n1016) );
  XOR U3000 ( .A(n905), .B(n889), .Z(n891) );
  XOR U3001 ( .A(n449), .B(n433), .Z(n435) );
  XOR U3002 ( .A(n1672), .B(n1656), .Z(n1658) );
  XOR U3003 ( .A(n1547), .B(n1531), .Z(n1533) );
  XOR U3004 ( .A(n272), .B(n256), .Z(n258) );
  XOR U3005 ( .A(n1409), .B(n1393), .Z(n1395) );
  XOR U3006 ( .A(n757), .B(n741), .Z(n743) );
  XOR U3007 ( .A(n1286), .B(n1270), .Z(n1272) );
  XOR U3008 ( .A(n643), .B(n508), .Z(n511) );
  XOR U3009 ( .A(n1919), .B(n1903), .Z(n1905) );
  NANDN U3010 ( .A(n116), .B(n121), .Z(n4) );
  XOR U3011 ( .A(n116), .B(n119), .Z(n5) );
  OR U3012 ( .A(n121), .B(n5), .Z(n6) );
  NANDN U3013 ( .A(n117), .B(n6), .Z(n7) );
  NAND U3014 ( .A(n4), .B(n7), .Z(n169) );
  XOR U3015 ( .A(n1796), .B(n1780), .Z(n1782) );
  XOR U3016 ( .A(n1163), .B(n1147), .Z(n1149) );
  XOR U3017 ( .A(x[3]), .B(x[1]), .Z(n10) );
  XNOR U3018 ( .A(x[0]), .B(x[6]), .Z(n9) );
  XOR U3019 ( .A(n9), .B(x[2]), .Z(n8) );
  XNOR U3020 ( .A(n10), .B(n8), .Z(n45) );
  XNOR U3021 ( .A(x[5]), .B(n9), .Z(n1432) );
  XOR U3022 ( .A(n1432), .B(x[4]), .Z(n787) );
  IV U3023 ( .A(n787), .Z(n19) );
  XNOR U3024 ( .A(x[7]), .B(x[4]), .Z(n13) );
  XNOR U3025 ( .A(n10), .B(n13), .Z(n73) );
  NOR U3026 ( .A(n19), .B(n73), .Z(n12) );
  XNOR U3027 ( .A(n1432), .B(x[7]), .Z(n1067) );
  XNOR U3028 ( .A(x[2]), .B(n1067), .Z(n28) );
  XNOR U3029 ( .A(x[1]), .B(n28), .Z(n23) );
  AND U3030 ( .A(x[0]), .B(n23), .Z(n11) );
  XNOR U3031 ( .A(n12), .B(n11), .Z(n16) );
  XNOR U3032 ( .A(n45), .B(n1067), .Z(n35) );
  IV U3033 ( .A(n45), .Z(n30) );
  XNOR U3034 ( .A(x[0]), .B(n30), .Z(n50) );
  IV U3035 ( .A(n13), .Z(n777) );
  AND U3036 ( .A(n50), .B(n777), .Z(n18) );
  IV U3037 ( .A(n1432), .Z(n37) );
  XNOR U3038 ( .A(n45), .B(n37), .Z(n67) );
  XOR U3039 ( .A(n67), .B(n73), .Z(n70) );
  XOR U3040 ( .A(x[2]), .B(x[4]), .Z(n779) );
  NAND U3041 ( .A(n70), .B(n779), .Z(n14) );
  XNOR U3042 ( .A(n18), .B(n14), .Z(n39) );
  XNOR U3043 ( .A(n35), .B(n39), .Z(n15) );
  XNOR U3044 ( .A(n16), .B(n15), .Z(n62) );
  XOR U3045 ( .A(x[2]), .B(x[7]), .Z(n793) );
  XNOR U3046 ( .A(x[0]), .B(n73), .Z(n74) );
  XNOR U3047 ( .A(n1432), .B(n74), .Z(n65) );
  NAND U3048 ( .A(n793), .B(n65), .Z(n17) );
  XNOR U3049 ( .A(n18), .B(n17), .Z(n31) );
  IV U3050 ( .A(n23), .Z(n776) );
  XNOR U3051 ( .A(n776), .B(n19), .Z(n783) );
  AND U3052 ( .A(n73), .B(n783), .Z(n21) );
  AND U3053 ( .A(x[0]), .B(n787), .Z(n20) );
  XNOR U3054 ( .A(n21), .B(n20), .Z(n22) );
  NANDN U3055 ( .A(n74), .B(n22), .Z(n26) );
  NAND U3056 ( .A(x[0]), .B(n73), .Z(n24) );
  OR U3057 ( .A(n24), .B(n23), .Z(n25) );
  NAND U3058 ( .A(n26), .B(n25), .Z(n27) );
  XNOR U3059 ( .A(n28), .B(n27), .Z(n29) );
  XNOR U3060 ( .A(n31), .B(n29), .Z(n51) );
  IV U3061 ( .A(n51), .Z(n58) );
  AND U3062 ( .A(n1067), .B(n30), .Z(n33) );
  XOR U3063 ( .A(x[1]), .B(x[7]), .Z(n1069) );
  AND U3064 ( .A(n67), .B(n1069), .Z(n36) );
  XNOR U3065 ( .A(n36), .B(n31), .Z(n32) );
  XNOR U3066 ( .A(n33), .B(n32), .Z(n57) );
  NANDN U3067 ( .A(n58), .B(n57), .Z(n34) );
  NAND U3068 ( .A(n62), .B(n34), .Z(n44) );
  XNOR U3069 ( .A(n36), .B(n35), .Z(n41) );
  ANDN U3070 ( .B(n37), .A(x[1]), .Z(n38) );
  XNOR U3071 ( .A(n39), .B(n38), .Z(n40) );
  XNOR U3072 ( .A(n41), .B(n40), .Z(n54) );
  XOR U3073 ( .A(n57), .B(n54), .Z(n42) );
  NAND U3074 ( .A(n58), .B(n42), .Z(n43) );
  NAND U3075 ( .A(n44), .B(n43), .Z(n1066) );
  ANDN U3076 ( .B(n45), .A(n1066), .Z(n69) );
  IV U3077 ( .A(n54), .Z(n60) );
  XOR U3078 ( .A(n62), .B(n58), .Z(n46) );
  NANDN U3079 ( .A(n60), .B(n46), .Z(n49) );
  NANDN U3080 ( .A(n58), .B(n60), .Z(n47) );
  NANDN U3081 ( .A(n57), .B(n47), .Z(n48) );
  NAND U3082 ( .A(n49), .B(n48), .Z(n1427) );
  XNOR U3083 ( .A(n1066), .B(n1427), .Z(n778) );
  AND U3084 ( .A(n50), .B(n778), .Z(n72) );
  OR U3085 ( .A(n57), .B(n54), .Z(n56) );
  ANDN U3086 ( .B(n57), .A(n51), .Z(n52) );
  XNOR U3087 ( .A(n52), .B(n62), .Z(n53) );
  NAND U3088 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3089 ( .A(n56), .B(n55), .Z(n775) );
  NAND U3090 ( .A(n58), .B(n62), .Z(n64) );
  NAND U3091 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U3092 ( .A(n60), .B(n59), .Z(n61) );
  NANDN U3093 ( .A(n62), .B(n61), .Z(n63) );
  NAND U3094 ( .A(n64), .B(n63), .Z(n1434) );
  NAND U3095 ( .A(n794), .B(n65), .Z(n66) );
  XNOR U3096 ( .A(n72), .B(n66), .Z(n1429) );
  XOR U3097 ( .A(n1066), .B(n1434), .Z(n1068) );
  AND U3098 ( .A(n67), .B(n1068), .Z(n789) );
  XNOR U3099 ( .A(n1429), .B(n789), .Z(n68) );
  XNOR U3100 ( .A(n69), .B(n68), .Z(n1437) );
  NAND U3101 ( .A(n780), .B(n70), .Z(n71) );
  XNOR U3102 ( .A(n72), .B(n71), .Z(n797) );
  AND U3103 ( .A(n73), .B(n782), .Z(n1428) );
  NANDN U3104 ( .A(n74), .B(n775), .Z(n75) );
  XNOR U3105 ( .A(n1428), .B(n75), .Z(n939) );
  XNOR U3106 ( .A(n797), .B(n939), .Z(n786) );
  XOR U3107 ( .A(n1437), .B(n786), .Z(z[0]) );
  XOR U3108 ( .A(x[99]), .B(x[97]), .Z(n76) );
  XNOR U3109 ( .A(n76), .B(x[98]), .Z(n77) );
  XNOR U3110 ( .A(x[101]), .B(n77), .Z(n114) );
  XOR U3111 ( .A(x[98]), .B(x[100]), .Z(n135) );
  XNOR U3112 ( .A(x[102]), .B(n77), .Z(n128) );
  XOR U3113 ( .A(x[103]), .B(x[100]), .Z(n133) );
  XOR U3114 ( .A(n76), .B(n133), .Z(n124) );
  XNOR U3115 ( .A(x[96]), .B(n124), .Z(n93) );
  IV U3116 ( .A(n93), .Z(n125) );
  XNOR U3117 ( .A(x[102]), .B(x[96]), .Z(n78) );
  XNOR U3118 ( .A(x[101]), .B(n78), .Z(n139) );
  XOR U3119 ( .A(n125), .B(n139), .Z(n127) );
  XOR U3120 ( .A(n128), .B(n127), .Z(n156) );
  AND U3121 ( .A(n135), .B(n156), .Z(n80) );
  AND U3122 ( .A(n128), .B(n133), .Z(n86) );
  IV U3123 ( .A(n139), .Z(n102) );
  XNOR U3124 ( .A(x[103]), .B(n102), .Z(n161) );
  XOR U3125 ( .A(n129), .B(n161), .Z(n84) );
  XNOR U3126 ( .A(n86), .B(n84), .Z(n79) );
  XNOR U3127 ( .A(n80), .B(n79), .Z(n103) );
  XOR U3128 ( .A(x[98]), .B(n161), .Z(n98) );
  XOR U3129 ( .A(x[97]), .B(n98), .Z(n150) );
  ANDN U3130 ( .B(x[96]), .A(n150), .Z(n82) );
  XNOR U3131 ( .A(x[100]), .B(n102), .Z(n170) );
  NANDN U3132 ( .A(n124), .B(n170), .Z(n81) );
  XNOR U3133 ( .A(n82), .B(n81), .Z(n83) );
  XOR U3134 ( .A(n103), .B(n83), .Z(n119) );
  XOR U3135 ( .A(x[97]), .B(x[103]), .Z(n138) );
  AND U3136 ( .A(n138), .B(n114), .Z(n104) );
  XOR U3137 ( .A(n84), .B(n104), .Z(n89) );
  XOR U3138 ( .A(x[98]), .B(x[103]), .Z(n162) );
  NAND U3139 ( .A(n162), .B(n127), .Z(n85) );
  XOR U3140 ( .A(n86), .B(n85), .Z(n99) );
  AND U3141 ( .A(n129), .B(n161), .Z(n87) );
  XOR U3142 ( .A(n99), .B(n87), .Z(n88) );
  XNOR U3143 ( .A(n89), .B(n88), .Z(n117) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n152) );
  AND U3145 ( .A(n124), .B(n152), .Z(n91) );
  AND U3146 ( .A(x[96]), .B(n170), .Z(n90) );
  XNOR U3147 ( .A(n91), .B(n90), .Z(n92) );
  NANDN U3148 ( .A(n93), .B(n92), .Z(n96) );
  NAND U3149 ( .A(n124), .B(x[96]), .Z(n94) );
  NANDN U3150 ( .A(n94), .B(n150), .Z(n95) );
  NAND U3151 ( .A(n96), .B(n95), .Z(n97) );
  XNOR U3152 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U3153 ( .A(n100), .B(n99), .Z(n116) );
  OR U3154 ( .A(n117), .B(n116), .Z(n101) );
  NANDN U3155 ( .A(n119), .B(n101), .Z(n109) );
  ANDN U3156 ( .B(n102), .A(x[97]), .Z(n106) );
  XNOR U3157 ( .A(n104), .B(n103), .Z(n105) );
  XNOR U3158 ( .A(n106), .B(n105), .Z(n121) );
  XOR U3159 ( .A(n117), .B(n121), .Z(n107) );
  NAND U3160 ( .A(n116), .B(n107), .Z(n108) );
  NAND U3161 ( .A(n109), .B(n108), .Z(n160) );
  OR U3162 ( .A(n119), .B(n116), .Z(n113) );
  ANDN U3163 ( .B(n116), .A(n117), .Z(n110) );
  XNOR U3164 ( .A(n110), .B(n121), .Z(n111) );
  NAND U3165 ( .A(n119), .B(n111), .Z(n112) );
  NAND U3166 ( .A(n113), .B(n112), .Z(n141) );
  XNOR U3167 ( .A(n160), .B(n141), .Z(n137) );
  AND U3168 ( .A(n114), .B(n137), .Z(n131) );
  NAND U3169 ( .A(n139), .B(n141), .Z(n115) );
  XNOR U3170 ( .A(n131), .B(n115), .Z(n172) );
  NANDN U3171 ( .A(n117), .B(n121), .Z(n123) );
  NANDN U3172 ( .A(n117), .B(n116), .Z(n118) );
  XOR U3173 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U3174 ( .A(n121), .B(n120), .Z(n122) );
  NAND U3175 ( .A(n123), .B(n122), .Z(n149) );
  XOR U3176 ( .A(n169), .B(n149), .Z(n151) );
  AND U3177 ( .A(n124), .B(n151), .Z(n144) );
  NANDN U3178 ( .A(n149), .B(n125), .Z(n126) );
  XNOR U3179 ( .A(n144), .B(n126), .Z(n159) );
  XNOR U3180 ( .A(n172), .B(n159), .Z(z[98]) );
  XNOR U3181 ( .A(n149), .B(n141), .Z(n163) );
  AND U3182 ( .A(n127), .B(n163), .Z(n183) );
  XOR U3183 ( .A(n169), .B(n160), .Z(n134) );
  AND U3184 ( .A(n128), .B(n134), .Z(n181) );
  NANDN U3185 ( .A(n160), .B(n129), .Z(n130) );
  XNOR U3186 ( .A(n131), .B(n130), .Z(n145) );
  XNOR U3187 ( .A(n181), .B(n145), .Z(n132) );
  XNOR U3188 ( .A(n183), .B(n132), .Z(n1958) );
  XOR U3189 ( .A(n1958), .B(z[98]), .Z(z[100]) );
  AND U3190 ( .A(n133), .B(n134), .Z(n165) );
  NAND U3191 ( .A(n157), .B(n135), .Z(n136) );
  XNOR U3192 ( .A(n165), .B(n136), .Z(n153) );
  AND U3193 ( .A(n138), .B(n137), .Z(n166) );
  XOR U3194 ( .A(x[97]), .B(n139), .Z(n140) );
  NAND U3195 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U3196 ( .A(n166), .B(n142), .Z(n147) );
  NANDN U3197 ( .A(n169), .B(x[96]), .Z(n143) );
  XNOR U3198 ( .A(n144), .B(n143), .Z(n180) );
  XNOR U3199 ( .A(n180), .B(n145), .Z(n146) );
  XNOR U3200 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U3201 ( .A(n153), .B(n148), .Z(z[101]) );
  ANDN U3202 ( .B(n150), .A(n149), .Z(n155) );
  AND U3203 ( .A(n152), .B(n151), .Z(n171) );
  XNOR U3204 ( .A(n171), .B(n153), .Z(n154) );
  XNOR U3205 ( .A(n155), .B(n154), .Z(n1959) );
  NAND U3206 ( .A(n157), .B(n156), .Z(n158) );
  XNOR U3207 ( .A(n181), .B(n158), .Z(n175) );
  XNOR U3208 ( .A(n175), .B(n159), .Z(n1957) );
  XNOR U3209 ( .A(n1959), .B(n1957), .Z(n179) );
  ANDN U3210 ( .B(n161), .A(n160), .Z(n168) );
  NAND U3211 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U3212 ( .A(n165), .B(n164), .Z(n176) );
  XNOR U3213 ( .A(n176), .B(n166), .Z(n167) );
  XNOR U3214 ( .A(n168), .B(n167), .Z(n1962) );
  XNOR U3215 ( .A(n179), .B(n1962), .Z(z[102]) );
  ANDN U3216 ( .B(n170), .A(n169), .Z(n174) );
  XNOR U3217 ( .A(n172), .B(n171), .Z(n173) );
  XNOR U3218 ( .A(n174), .B(n173), .Z(n178) );
  XNOR U3219 ( .A(n176), .B(n175), .Z(n177) );
  XNOR U3220 ( .A(n178), .B(n177), .Z(n1960) );
  XNOR U3221 ( .A(n1960), .B(n179), .Z(z[97]) );
  XNOR U3222 ( .A(n181), .B(n180), .Z(n182) );
  XNOR U3223 ( .A(n183), .B(n182), .Z(n184) );
  XOR U3224 ( .A(n184), .B(z[97]), .Z(z[103]) );
  XOR U3225 ( .A(x[107]), .B(x[105]), .Z(n187) );
  XNOR U3226 ( .A(x[104]), .B(x[110]), .Z(n186) );
  XOR U3227 ( .A(n186), .B(x[106]), .Z(n185) );
  XNOR U3228 ( .A(n187), .B(n185), .Z(n222) );
  XNOR U3229 ( .A(x[109]), .B(n186), .Z(n295) );
  XOR U3230 ( .A(n295), .B(x[108]), .Z(n265) );
  IV U3231 ( .A(n265), .Z(n196) );
  XNOR U3232 ( .A(x[111]), .B(x[108]), .Z(n190) );
  XNOR U3233 ( .A(n187), .B(n190), .Z(n250) );
  NOR U3234 ( .A(n196), .B(n250), .Z(n189) );
  XNOR U3235 ( .A(n295), .B(x[111]), .Z(n281) );
  XNOR U3236 ( .A(x[106]), .B(n281), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n205), .Z(n200) );
  AND U3238 ( .A(x[104]), .B(n200), .Z(n188) );
  XNOR U3239 ( .A(n189), .B(n188), .Z(n193) );
  XNOR U3240 ( .A(n222), .B(n281), .Z(n212) );
  IV U3241 ( .A(n222), .Z(n207) );
  XNOR U3242 ( .A(x[104]), .B(n207), .Z(n227) );
  IV U3243 ( .A(n190), .Z(n255) );
  AND U3244 ( .A(n227), .B(n255), .Z(n195) );
  IV U3245 ( .A(n295), .Z(n214) );
  XNOR U3246 ( .A(n222), .B(n214), .Z(n244) );
  XOR U3247 ( .A(n244), .B(n250), .Z(n247) );
  XOR U3248 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NAND U3249 ( .A(n247), .B(n257), .Z(n191) );
  XNOR U3250 ( .A(n195), .B(n191), .Z(n216) );
  XNOR U3251 ( .A(n212), .B(n216), .Z(n192) );
  XNOR U3252 ( .A(n193), .B(n192), .Z(n239) );
  XOR U3253 ( .A(x[106]), .B(x[111]), .Z(n271) );
  XNOR U3254 ( .A(x[104]), .B(n250), .Z(n251) );
  XNOR U3255 ( .A(n295), .B(n251), .Z(n242) );
  NAND U3256 ( .A(n271), .B(n242), .Z(n194) );
  XNOR U3257 ( .A(n195), .B(n194), .Z(n208) );
  IV U3258 ( .A(n200), .Z(n254) );
  XNOR U3259 ( .A(n254), .B(n196), .Z(n261) );
  AND U3260 ( .A(n250), .B(n261), .Z(n198) );
  AND U3261 ( .A(x[104]), .B(n265), .Z(n197) );
  XNOR U3262 ( .A(n198), .B(n197), .Z(n199) );
  NANDN U3263 ( .A(n251), .B(n199), .Z(n203) );
  NAND U3264 ( .A(x[104]), .B(n250), .Z(n201) );
  OR U3265 ( .A(n201), .B(n200), .Z(n202) );
  NAND U3266 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U3267 ( .A(n205), .B(n204), .Z(n206) );
  XNOR U3268 ( .A(n208), .B(n206), .Z(n228) );
  IV U3269 ( .A(n228), .Z(n235) );
  AND U3270 ( .A(n281), .B(n207), .Z(n210) );
  XOR U3271 ( .A(x[105]), .B(x[111]), .Z(n283) );
  AND U3272 ( .A(n244), .B(n283), .Z(n213) );
  XNOR U3273 ( .A(n213), .B(n208), .Z(n209) );
  XNOR U3274 ( .A(n210), .B(n209), .Z(n234) );
  NANDN U3275 ( .A(n235), .B(n234), .Z(n211) );
  NAND U3276 ( .A(n239), .B(n211), .Z(n221) );
  XNOR U3277 ( .A(n213), .B(n212), .Z(n218) );
  ANDN U3278 ( .B(n214), .A(x[105]), .Z(n215) );
  XNOR U3279 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3280 ( .A(n218), .B(n217), .Z(n231) );
  XOR U3281 ( .A(n234), .B(n231), .Z(n219) );
  NAND U3282 ( .A(n235), .B(n219), .Z(n220) );
  NAND U3283 ( .A(n221), .B(n220), .Z(n280) );
  ANDN U3284 ( .B(n222), .A(n280), .Z(n246) );
  IV U3285 ( .A(n231), .Z(n237) );
  XOR U3286 ( .A(n239), .B(n235), .Z(n223) );
  NANDN U3287 ( .A(n237), .B(n223), .Z(n226) );
  NANDN U3288 ( .A(n235), .B(n237), .Z(n224) );
  NANDN U3289 ( .A(n234), .B(n224), .Z(n225) );
  NAND U3290 ( .A(n226), .B(n225), .Z(n290) );
  XNOR U3291 ( .A(n280), .B(n290), .Z(n256) );
  AND U3292 ( .A(n227), .B(n256), .Z(n249) );
  OR U3293 ( .A(n234), .B(n231), .Z(n233) );
  ANDN U3294 ( .B(n234), .A(n228), .Z(n229) );
  XNOR U3295 ( .A(n229), .B(n239), .Z(n230) );
  NAND U3296 ( .A(n231), .B(n230), .Z(n232) );
  NAND U3297 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3298 ( .A(n235), .B(n239), .Z(n241) );
  NAND U3299 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U3300 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U3301 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3302 ( .A(n241), .B(n240), .Z(n297) );
  NAND U3303 ( .A(n272), .B(n242), .Z(n243) );
  XNOR U3304 ( .A(n249), .B(n243), .Z(n292) );
  XOR U3305 ( .A(n280), .B(n297), .Z(n282) );
  AND U3306 ( .A(n244), .B(n282), .Z(n267) );
  XNOR U3307 ( .A(n292), .B(n267), .Z(n245) );
  XNOR U3308 ( .A(n246), .B(n245), .Z(n300) );
  NAND U3309 ( .A(n258), .B(n247), .Z(n248) );
  XNOR U3310 ( .A(n249), .B(n248), .Z(n275) );
  AND U3311 ( .A(n250), .B(n260), .Z(n291) );
  NANDN U3312 ( .A(n251), .B(n253), .Z(n252) );
  XNOR U3313 ( .A(n291), .B(n252), .Z(n279) );
  XNOR U3314 ( .A(n275), .B(n279), .Z(n264) );
  XOR U3315 ( .A(n300), .B(n264), .Z(z[104]) );
  AND U3316 ( .A(n254), .B(n253), .Z(n263) );
  AND U3317 ( .A(n256), .B(n255), .Z(n274) );
  NAND U3318 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3319 ( .A(n274), .B(n259), .Z(n301) );
  AND U3320 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3321 ( .A(n301), .B(n268), .Z(n262) );
  XNOR U3322 ( .A(n263), .B(n262), .Z(n288) );
  XNOR U3323 ( .A(n288), .B(n264), .Z(n360) );
  AND U3324 ( .A(n265), .B(n290), .Z(n270) );
  NANDN U3325 ( .A(n297), .B(n295), .Z(n266) );
  XNOR U3326 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3327 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3328 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3329 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3330 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3331 ( .A(n275), .B(n284), .Z(n276) );
  XNOR U3332 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3333 ( .A(n360), .B(n287), .Z(z[105]) );
  XNOR U3334 ( .A(n279), .B(n278), .Z(z[106]) );
  NOR U3335 ( .A(n281), .B(n280), .Z(n286) );
  AND U3336 ( .A(n283), .B(n282), .Z(n299) );
  XNOR U3337 ( .A(n284), .B(n299), .Z(n285) );
  XNOR U3338 ( .A(n286), .B(n285), .Z(n359) );
  XOR U3339 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U3340 ( .A(n359), .B(n289), .Z(z[107]) );
  XOR U3341 ( .A(n300), .B(z[106]), .Z(z[108]) );
  AND U3342 ( .A(x[104]), .B(n290), .Z(n294) );
  XNOR U3343 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U3344 ( .A(n294), .B(n293), .Z(n361) );
  XOR U3345 ( .A(n295), .B(x[105]), .Z(n296) );
  NANDN U3346 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U3347 ( .A(n299), .B(n298), .Z(n303) );
  XNOR U3348 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U3349 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U3350 ( .A(n361), .B(n304), .Z(z[109]) );
  XOR U3351 ( .A(x[9]), .B(x[11]), .Z(n305) );
  XOR U3352 ( .A(x[15]), .B(x[12]), .Z(n486) );
  XOR U3353 ( .A(n305), .B(n486), .Z(n341) );
  XNOR U3354 ( .A(x[8]), .B(x[14]), .Z(n307) );
  XNOR U3355 ( .A(x[13]), .B(n307), .Z(n654) );
  XNOR U3356 ( .A(x[15]), .B(n654), .Z(n485) );
  XNOR U3357 ( .A(n305), .B(x[10]), .Z(n306) );
  XNOR U3358 ( .A(n307), .B(n306), .Z(n308) );
  AND U3359 ( .A(n485), .B(n308), .Z(n311) );
  IV U3360 ( .A(n308), .Z(n641) );
  XOR U3361 ( .A(n641), .B(n654), .Z(n357) );
  XOR U3362 ( .A(x[9]), .B(x[15]), .Z(n491) );
  AND U3363 ( .A(n357), .B(n491), .Z(n312) );
  XNOR U3364 ( .A(x[8]), .B(n308), .Z(n509) );
  AND U3365 ( .A(n486), .B(n509), .Z(n314) );
  XOR U3366 ( .A(x[15]), .B(x[10]), .Z(n488) );
  XNOR U3367 ( .A(n341), .B(x[8]), .Z(n342) );
  XNOR U3368 ( .A(n654), .B(n342), .Z(n642) );
  NAND U3369 ( .A(n488), .B(n642), .Z(n309) );
  XNOR U3370 ( .A(n314), .B(n309), .Z(n325) );
  XNOR U3371 ( .A(n312), .B(n325), .Z(n310) );
  XNOR U3372 ( .A(n311), .B(n310), .Z(n349) );
  XNOR U3373 ( .A(n641), .B(n485), .Z(n329) );
  XOR U3374 ( .A(x[12]), .B(x[10]), .Z(n496) );
  XOR U3375 ( .A(n341), .B(n357), .Z(n510) );
  NAND U3376 ( .A(n496), .B(n510), .Z(n313) );
  XNOR U3377 ( .A(n314), .B(n313), .Z(n328) );
  OR U3378 ( .A(n349), .B(n345), .Z(n335) );
  XNOR U3379 ( .A(x[10]), .B(n485), .Z(n323) );
  IV U3380 ( .A(n318), .Z(n495) );
  XNOR U3381 ( .A(x[12]), .B(n654), .Z(n503) );
  XNOR U3382 ( .A(n495), .B(n503), .Z(n500) );
  AND U3383 ( .A(n341), .B(n500), .Z(n316) );
  ANDN U3384 ( .B(x[8]), .A(n503), .Z(n315) );
  XNOR U3385 ( .A(n316), .B(n315), .Z(n317) );
  NANDN U3386 ( .A(n342), .B(n317), .Z(n321) );
  NAND U3387 ( .A(n341), .B(x[8]), .Z(n319) );
  OR U3388 ( .A(n319), .B(n318), .Z(n320) );
  NAND U3389 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U3390 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U3391 ( .A(n325), .B(n324), .Z(n336) );
  ANDN U3392 ( .B(n349), .A(n336), .Z(n332) );
  NOR U3393 ( .A(n503), .B(n341), .Z(n327) );
  ANDN U3394 ( .B(x[8]), .A(n495), .Z(n326) );
  XNOR U3395 ( .A(n327), .B(n326), .Z(n331) );
  XNOR U3396 ( .A(n329), .B(n328), .Z(n330) );
  XNOR U3397 ( .A(n331), .B(n330), .Z(n354) );
  XNOR U3398 ( .A(n332), .B(n354), .Z(n333) );
  NAND U3399 ( .A(n345), .B(n333), .Z(n334) );
  NAND U3400 ( .A(n335), .B(n334), .Z(n494) );
  IV U3401 ( .A(n494), .Z(n487) );
  IV U3402 ( .A(n345), .Z(n352) );
  IV U3403 ( .A(n336), .Z(n350) );
  XOR U3404 ( .A(n354), .B(n350), .Z(n337) );
  NANDN U3405 ( .A(n352), .B(n337), .Z(n340) );
  NANDN U3406 ( .A(n350), .B(n352), .Z(n338) );
  NANDN U3407 ( .A(n349), .B(n338), .Z(n339) );
  NAND U3408 ( .A(n340), .B(n339), .Z(n649) );
  XNOR U3409 ( .A(n487), .B(n649), .Z(n499) );
  AND U3410 ( .A(n341), .B(n499), .Z(n651) );
  NANDN U3411 ( .A(n342), .B(n494), .Z(n343) );
  XNOR U3412 ( .A(n651), .B(n343), .Z(n663) );
  NANDN U3413 ( .A(n350), .B(n349), .Z(n344) );
  NAND U3414 ( .A(n354), .B(n344), .Z(n348) );
  XOR U3415 ( .A(n349), .B(n345), .Z(n346) );
  NAND U3416 ( .A(n350), .B(n346), .Z(n347) );
  NAND U3417 ( .A(n348), .B(n347), .Z(n640) );
  NAND U3418 ( .A(n350), .B(n354), .Z(n356) );
  NAND U3419 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U3420 ( .A(n352), .B(n351), .Z(n353) );
  NANDN U3421 ( .A(n354), .B(n353), .Z(n355) );
  NAND U3422 ( .A(n356), .B(n355), .Z(n656) );
  XOR U3423 ( .A(n640), .B(n656), .Z(n490) );
  AND U3424 ( .A(n357), .B(n490), .Z(n646) );
  NANDN U3425 ( .A(n656), .B(n654), .Z(n358) );
  XNOR U3426 ( .A(n646), .B(n358), .Z(n513) );
  XNOR U3427 ( .A(n663), .B(n513), .Z(z[10]) );
  XNOR U3428 ( .A(n360), .B(n359), .Z(z[110]) );
  XOR U3429 ( .A(n361), .B(z[105]), .Z(z[111]) );
  XOR U3430 ( .A(x[115]), .B(x[113]), .Z(n364) );
  XNOR U3431 ( .A(x[112]), .B(x[118]), .Z(n363) );
  XOR U3432 ( .A(n363), .B(x[114]), .Z(n362) );
  XNOR U3433 ( .A(n364), .B(n362), .Z(n399) );
  XNOR U3434 ( .A(x[117]), .B(n363), .Z(n472) );
  XOR U3435 ( .A(n472), .B(x[116]), .Z(n442) );
  IV U3436 ( .A(n442), .Z(n373) );
  XNOR U3437 ( .A(x[119]), .B(x[116]), .Z(n367) );
  XNOR U3438 ( .A(n364), .B(n367), .Z(n427) );
  NOR U3439 ( .A(n373), .B(n427), .Z(n366) );
  XNOR U3440 ( .A(n472), .B(x[119]), .Z(n458) );
  XNOR U3441 ( .A(x[114]), .B(n458), .Z(n382) );
  XNOR U3442 ( .A(x[113]), .B(n382), .Z(n377) );
  AND U3443 ( .A(x[112]), .B(n377), .Z(n365) );
  XNOR U3444 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U3445 ( .A(n399), .B(n458), .Z(n389) );
  IV U3446 ( .A(n399), .Z(n384) );
  XNOR U3447 ( .A(x[112]), .B(n384), .Z(n404) );
  IV U3448 ( .A(n367), .Z(n432) );
  AND U3449 ( .A(n404), .B(n432), .Z(n372) );
  IV U3450 ( .A(n472), .Z(n391) );
  XNOR U3451 ( .A(n399), .B(n391), .Z(n421) );
  XOR U3452 ( .A(n421), .B(n427), .Z(n424) );
  XOR U3453 ( .A(x[114]), .B(x[116]), .Z(n434) );
  NAND U3454 ( .A(n424), .B(n434), .Z(n368) );
  XNOR U3455 ( .A(n372), .B(n368), .Z(n393) );
  XNOR U3456 ( .A(n389), .B(n393), .Z(n369) );
  XNOR U3457 ( .A(n370), .B(n369), .Z(n416) );
  XOR U3458 ( .A(x[114]), .B(x[119]), .Z(n448) );
  XNOR U3459 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3460 ( .A(n472), .B(n428), .Z(n419) );
  NAND U3461 ( .A(n448), .B(n419), .Z(n371) );
  XNOR U3462 ( .A(n372), .B(n371), .Z(n385) );
  IV U3463 ( .A(n377), .Z(n431) );
  XNOR U3464 ( .A(n431), .B(n373), .Z(n438) );
  AND U3465 ( .A(n427), .B(n438), .Z(n375) );
  AND U3466 ( .A(x[112]), .B(n442), .Z(n374) );
  XNOR U3467 ( .A(n375), .B(n374), .Z(n376) );
  NANDN U3468 ( .A(n428), .B(n376), .Z(n380) );
  NAND U3469 ( .A(x[112]), .B(n427), .Z(n378) );
  OR U3470 ( .A(n378), .B(n377), .Z(n379) );
  NAND U3471 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U3472 ( .A(n382), .B(n381), .Z(n383) );
  XNOR U3473 ( .A(n385), .B(n383), .Z(n405) );
  IV U3474 ( .A(n405), .Z(n412) );
  AND U3475 ( .A(n458), .B(n384), .Z(n387) );
  XOR U3476 ( .A(x[113]), .B(x[119]), .Z(n460) );
  AND U3477 ( .A(n421), .B(n460), .Z(n390) );
  XNOR U3478 ( .A(n390), .B(n385), .Z(n386) );
  XNOR U3479 ( .A(n387), .B(n386), .Z(n411) );
  NANDN U3480 ( .A(n412), .B(n411), .Z(n388) );
  NAND U3481 ( .A(n416), .B(n388), .Z(n398) );
  XNOR U3482 ( .A(n390), .B(n389), .Z(n395) );
  ANDN U3483 ( .B(n391), .A(x[113]), .Z(n392) );
  XNOR U3484 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U3485 ( .A(n395), .B(n394), .Z(n408) );
  XOR U3486 ( .A(n411), .B(n408), .Z(n396) );
  NAND U3487 ( .A(n412), .B(n396), .Z(n397) );
  NAND U3488 ( .A(n398), .B(n397), .Z(n457) );
  ANDN U3489 ( .B(n399), .A(n457), .Z(n423) );
  IV U3490 ( .A(n408), .Z(n414) );
  XOR U3491 ( .A(n416), .B(n412), .Z(n400) );
  NANDN U3492 ( .A(n414), .B(n400), .Z(n403) );
  NANDN U3493 ( .A(n412), .B(n414), .Z(n401) );
  NANDN U3494 ( .A(n411), .B(n401), .Z(n402) );
  NAND U3495 ( .A(n403), .B(n402), .Z(n467) );
  XNOR U3496 ( .A(n457), .B(n467), .Z(n433) );
  AND U3497 ( .A(n404), .B(n433), .Z(n426) );
  OR U3498 ( .A(n411), .B(n408), .Z(n410) );
  ANDN U3499 ( .B(n411), .A(n405), .Z(n406) );
  XNOR U3500 ( .A(n406), .B(n416), .Z(n407) );
  NAND U3501 ( .A(n408), .B(n407), .Z(n409) );
  NAND U3502 ( .A(n410), .B(n409), .Z(n430) );
  NAND U3503 ( .A(n412), .B(n416), .Z(n418) );
  NAND U3504 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U3505 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U3506 ( .A(n416), .B(n415), .Z(n417) );
  NAND U3507 ( .A(n418), .B(n417), .Z(n474) );
  NAND U3508 ( .A(n449), .B(n419), .Z(n420) );
  XNOR U3509 ( .A(n426), .B(n420), .Z(n469) );
  XOR U3510 ( .A(n457), .B(n474), .Z(n459) );
  AND U3511 ( .A(n421), .B(n459), .Z(n444) );
  XNOR U3512 ( .A(n469), .B(n444), .Z(n422) );
  XNOR U3513 ( .A(n423), .B(n422), .Z(n477) );
  NAND U3514 ( .A(n435), .B(n424), .Z(n425) );
  XNOR U3515 ( .A(n426), .B(n425), .Z(n452) );
  AND U3516 ( .A(n427), .B(n437), .Z(n468) );
  NANDN U3517 ( .A(n428), .B(n430), .Z(n429) );
  XNOR U3518 ( .A(n468), .B(n429), .Z(n456) );
  XNOR U3519 ( .A(n452), .B(n456), .Z(n441) );
  XOR U3520 ( .A(n477), .B(n441), .Z(z[112]) );
  AND U3521 ( .A(n431), .B(n430), .Z(n440) );
  AND U3522 ( .A(n433), .B(n432), .Z(n451) );
  NAND U3523 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U3524 ( .A(n451), .B(n436), .Z(n478) );
  AND U3525 ( .A(n438), .B(n437), .Z(n445) );
  XNOR U3526 ( .A(n478), .B(n445), .Z(n439) );
  XNOR U3527 ( .A(n440), .B(n439), .Z(n465) );
  XNOR U3528 ( .A(n465), .B(n441), .Z(n483) );
  AND U3529 ( .A(n442), .B(n467), .Z(n447) );
  NANDN U3530 ( .A(n474), .B(n472), .Z(n443) );
  XNOR U3531 ( .A(n444), .B(n443), .Z(n455) );
  XNOR U3532 ( .A(n445), .B(n455), .Z(n446) );
  XNOR U3533 ( .A(n447), .B(n446), .Z(n454) );
  NAND U3534 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U3535 ( .A(n451), .B(n450), .Z(n461) );
  XNOR U3536 ( .A(n452), .B(n461), .Z(n453) );
  XNOR U3537 ( .A(n454), .B(n453), .Z(n464) );
  XNOR U3538 ( .A(n483), .B(n464), .Z(z[113]) );
  XNOR U3539 ( .A(n456), .B(n455), .Z(z[114]) );
  NOR U3540 ( .A(n458), .B(n457), .Z(n463) );
  AND U3541 ( .A(n460), .B(n459), .Z(n476) );
  XNOR U3542 ( .A(n461), .B(n476), .Z(n462) );
  XNOR U3543 ( .A(n463), .B(n462), .Z(n482) );
  XOR U3544 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U3545 ( .A(n482), .B(n466), .Z(z[115]) );
  XOR U3546 ( .A(n477), .B(z[114]), .Z(z[116]) );
  AND U3547 ( .A(x[112]), .B(n467), .Z(n471) );
  XNOR U3548 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U3549 ( .A(n471), .B(n470), .Z(n484) );
  XOR U3550 ( .A(n472), .B(x[113]), .Z(n473) );
  NANDN U3551 ( .A(n474), .B(n473), .Z(n475) );
  XNOR U3552 ( .A(n476), .B(n475), .Z(n480) );
  XNOR U3553 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U3554 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U3555 ( .A(n484), .B(n481), .Z(z[117]) );
  XNOR U3556 ( .A(n483), .B(n482), .Z(z[118]) );
  XOR U3557 ( .A(n484), .B(z[113]), .Z(z[119]) );
  NOR U3558 ( .A(n485), .B(n640), .Z(n493) );
  XNOR U3559 ( .A(n640), .B(n649), .Z(n508) );
  AND U3560 ( .A(n486), .B(n508), .Z(n498) );
  XOR U3561 ( .A(n487), .B(n656), .Z(n643) );
  NAND U3562 ( .A(n643), .B(n488), .Z(n489) );
  XNOR U3563 ( .A(n498), .B(n489), .Z(n504) );
  AND U3564 ( .A(n491), .B(n490), .Z(n658) );
  XNOR U3565 ( .A(n504), .B(n658), .Z(n492) );
  XNOR U3566 ( .A(n493), .B(n492), .Z(n666) );
  AND U3567 ( .A(n495), .B(n494), .Z(n502) );
  NAND U3568 ( .A(n511), .B(n496), .Z(n497) );
  XNOR U3569 ( .A(n498), .B(n497), .Z(n659) );
  AND U3570 ( .A(n500), .B(n499), .Z(n505) );
  XNOR U3571 ( .A(n659), .B(n505), .Z(n501) );
  XNOR U3572 ( .A(n502), .B(n501), .Z(n665) );
  ANDN U3573 ( .B(n649), .A(n503), .Z(n507) );
  XNOR U3574 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U3575 ( .A(n507), .B(n506), .Z(n515) );
  AND U3576 ( .A(n509), .B(n508), .Z(n645) );
  NAND U3577 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U3578 ( .A(n645), .B(n512), .Z(n664) );
  XNOR U3579 ( .A(n664), .B(n513), .Z(n514) );
  XNOR U3580 ( .A(n515), .B(n514), .Z(n667) );
  XOR U3581 ( .A(n665), .B(n667), .Z(n516) );
  XNOR U3582 ( .A(n666), .B(n516), .Z(z[11]) );
  XOR U3583 ( .A(x[123]), .B(x[121]), .Z(n519) );
  XNOR U3584 ( .A(x[120]), .B(x[126]), .Z(n518) );
  XOR U3585 ( .A(n518), .B(x[122]), .Z(n517) );
  XNOR U3586 ( .A(n519), .B(n517), .Z(n554) );
  XNOR U3587 ( .A(x[125]), .B(n518), .Z(n627) );
  XOR U3588 ( .A(n627), .B(x[124]), .Z(n597) );
  IV U3589 ( .A(n597), .Z(n528) );
  XNOR U3590 ( .A(x[127]), .B(x[124]), .Z(n522) );
  XNOR U3591 ( .A(n519), .B(n522), .Z(n582) );
  NOR U3592 ( .A(n528), .B(n582), .Z(n521) );
  XNOR U3593 ( .A(n627), .B(x[127]), .Z(n613) );
  XNOR U3594 ( .A(x[122]), .B(n613), .Z(n537) );
  XNOR U3595 ( .A(x[121]), .B(n537), .Z(n532) );
  AND U3596 ( .A(x[120]), .B(n532), .Z(n520) );
  XNOR U3597 ( .A(n521), .B(n520), .Z(n525) );
  XNOR U3598 ( .A(n554), .B(n613), .Z(n544) );
  IV U3599 ( .A(n554), .Z(n539) );
  XNOR U3600 ( .A(x[120]), .B(n539), .Z(n559) );
  IV U3601 ( .A(n522), .Z(n587) );
  AND U3602 ( .A(n559), .B(n587), .Z(n527) );
  IV U3603 ( .A(n627), .Z(n546) );
  XNOR U3604 ( .A(n554), .B(n546), .Z(n576) );
  XOR U3605 ( .A(n576), .B(n582), .Z(n579) );
  XOR U3606 ( .A(x[122]), .B(x[124]), .Z(n589) );
  NAND U3607 ( .A(n579), .B(n589), .Z(n523) );
  XNOR U3608 ( .A(n527), .B(n523), .Z(n548) );
  XNOR U3609 ( .A(n544), .B(n548), .Z(n524) );
  XNOR U3610 ( .A(n525), .B(n524), .Z(n571) );
  XOR U3611 ( .A(x[122]), .B(x[127]), .Z(n603) );
  XNOR U3612 ( .A(x[120]), .B(n582), .Z(n583) );
  XNOR U3613 ( .A(n627), .B(n583), .Z(n574) );
  NAND U3614 ( .A(n603), .B(n574), .Z(n526) );
  XNOR U3615 ( .A(n527), .B(n526), .Z(n540) );
  IV U3616 ( .A(n532), .Z(n586) );
  XNOR U3617 ( .A(n586), .B(n528), .Z(n593) );
  AND U3618 ( .A(n582), .B(n593), .Z(n530) );
  AND U3619 ( .A(x[120]), .B(n597), .Z(n529) );
  XNOR U3620 ( .A(n530), .B(n529), .Z(n531) );
  NANDN U3621 ( .A(n583), .B(n531), .Z(n535) );
  NAND U3622 ( .A(x[120]), .B(n582), .Z(n533) );
  OR U3623 ( .A(n533), .B(n532), .Z(n534) );
  NAND U3624 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U3625 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U3626 ( .A(n540), .B(n538), .Z(n560) );
  IV U3627 ( .A(n560), .Z(n567) );
  AND U3628 ( .A(n613), .B(n539), .Z(n542) );
  XOR U3629 ( .A(x[121]), .B(x[127]), .Z(n615) );
  AND U3630 ( .A(n576), .B(n615), .Z(n545) );
  XNOR U3631 ( .A(n545), .B(n540), .Z(n541) );
  XNOR U3632 ( .A(n542), .B(n541), .Z(n566) );
  NANDN U3633 ( .A(n567), .B(n566), .Z(n543) );
  NAND U3634 ( .A(n571), .B(n543), .Z(n553) );
  XNOR U3635 ( .A(n545), .B(n544), .Z(n550) );
  ANDN U3636 ( .B(n546), .A(x[121]), .Z(n547) );
  XNOR U3637 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U3638 ( .A(n550), .B(n549), .Z(n563) );
  XOR U3639 ( .A(n566), .B(n563), .Z(n551) );
  NAND U3640 ( .A(n567), .B(n551), .Z(n552) );
  NAND U3641 ( .A(n553), .B(n552), .Z(n612) );
  ANDN U3642 ( .B(n554), .A(n612), .Z(n578) );
  IV U3643 ( .A(n563), .Z(n569) );
  XOR U3644 ( .A(n571), .B(n567), .Z(n555) );
  NANDN U3645 ( .A(n569), .B(n555), .Z(n558) );
  NANDN U3646 ( .A(n567), .B(n569), .Z(n556) );
  NANDN U3647 ( .A(n566), .B(n556), .Z(n557) );
  NAND U3648 ( .A(n558), .B(n557), .Z(n622) );
  XNOR U3649 ( .A(n612), .B(n622), .Z(n588) );
  AND U3650 ( .A(n559), .B(n588), .Z(n581) );
  OR U3651 ( .A(n566), .B(n563), .Z(n565) );
  ANDN U3652 ( .B(n566), .A(n560), .Z(n561) );
  XNOR U3653 ( .A(n561), .B(n571), .Z(n562) );
  NAND U3654 ( .A(n563), .B(n562), .Z(n564) );
  NAND U3655 ( .A(n565), .B(n564), .Z(n585) );
  NAND U3656 ( .A(n567), .B(n571), .Z(n573) );
  NAND U3657 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U3658 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U3659 ( .A(n571), .B(n570), .Z(n572) );
  NAND U3660 ( .A(n573), .B(n572), .Z(n629) );
  NAND U3661 ( .A(n604), .B(n574), .Z(n575) );
  XNOR U3662 ( .A(n581), .B(n575), .Z(n624) );
  XOR U3663 ( .A(n612), .B(n629), .Z(n614) );
  AND U3664 ( .A(n576), .B(n614), .Z(n599) );
  XNOR U3665 ( .A(n624), .B(n599), .Z(n577) );
  XNOR U3666 ( .A(n578), .B(n577), .Z(n632) );
  NAND U3667 ( .A(n590), .B(n579), .Z(n580) );
  XNOR U3668 ( .A(n581), .B(n580), .Z(n607) );
  AND U3669 ( .A(n582), .B(n592), .Z(n623) );
  NANDN U3670 ( .A(n583), .B(n585), .Z(n584) );
  XNOR U3671 ( .A(n623), .B(n584), .Z(n611) );
  XNOR U3672 ( .A(n607), .B(n611), .Z(n596) );
  XOR U3673 ( .A(n632), .B(n596), .Z(z[120]) );
  AND U3674 ( .A(n586), .B(n585), .Z(n595) );
  AND U3675 ( .A(n588), .B(n587), .Z(n606) );
  NAND U3676 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U3677 ( .A(n606), .B(n591), .Z(n633) );
  AND U3678 ( .A(n593), .B(n592), .Z(n600) );
  XNOR U3679 ( .A(n633), .B(n600), .Z(n594) );
  XNOR U3680 ( .A(n595), .B(n594), .Z(n620) );
  XNOR U3681 ( .A(n620), .B(n596), .Z(n638) );
  AND U3682 ( .A(n597), .B(n622), .Z(n602) );
  NANDN U3683 ( .A(n629), .B(n627), .Z(n598) );
  XNOR U3684 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U3685 ( .A(n600), .B(n610), .Z(n601) );
  XNOR U3686 ( .A(n602), .B(n601), .Z(n609) );
  NAND U3687 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U3688 ( .A(n606), .B(n605), .Z(n616) );
  XNOR U3689 ( .A(n607), .B(n616), .Z(n608) );
  XNOR U3690 ( .A(n609), .B(n608), .Z(n619) );
  XNOR U3691 ( .A(n638), .B(n619), .Z(z[121]) );
  XNOR U3692 ( .A(n611), .B(n610), .Z(z[122]) );
  NOR U3693 ( .A(n613), .B(n612), .Z(n618) );
  AND U3694 ( .A(n615), .B(n614), .Z(n631) );
  XNOR U3695 ( .A(n616), .B(n631), .Z(n617) );
  XNOR U3696 ( .A(n618), .B(n617), .Z(n637) );
  XOR U3697 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U3698 ( .A(n637), .B(n621), .Z(z[123]) );
  XOR U3699 ( .A(n632), .B(z[122]), .Z(z[124]) );
  AND U3700 ( .A(x[120]), .B(n622), .Z(n626) );
  XNOR U3701 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U3702 ( .A(n626), .B(n625), .Z(n639) );
  XOR U3703 ( .A(n627), .B(x[121]), .Z(n628) );
  NANDN U3704 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U3705 ( .A(n631), .B(n630), .Z(n635) );
  XNOR U3706 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U3707 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U3708 ( .A(n639), .B(n636), .Z(z[125]) );
  XNOR U3709 ( .A(n638), .B(n637), .Z(z[126]) );
  XOR U3710 ( .A(n639), .B(z[121]), .Z(z[127]) );
  ANDN U3711 ( .B(n641), .A(n640), .Z(n648) );
  NAND U3712 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U3713 ( .A(n645), .B(n644), .Z(n650) );
  XNOR U3714 ( .A(n650), .B(n646), .Z(n647) );
  XNOR U3715 ( .A(n648), .B(n647), .Z(n1926) );
  XOR U3716 ( .A(n1926), .B(z[10]), .Z(z[12]) );
  AND U3717 ( .A(x[8]), .B(n649), .Z(n653) );
  XNOR U3718 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U3719 ( .A(n653), .B(n652), .Z(n669) );
  XOR U3720 ( .A(n654), .B(x[9]), .Z(n655) );
  NANDN U3721 ( .A(n656), .B(n655), .Z(n657) );
  XNOR U3722 ( .A(n658), .B(n657), .Z(n661) );
  XNOR U3723 ( .A(n659), .B(n1926), .Z(n660) );
  XNOR U3724 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U3725 ( .A(n669), .B(n662), .Z(z[13]) );
  XNOR U3726 ( .A(n664), .B(n663), .Z(n1925) );
  XNOR U3727 ( .A(n665), .B(n1925), .Z(n668) );
  XNOR U3728 ( .A(n668), .B(n666), .Z(z[14]) );
  XNOR U3729 ( .A(n668), .B(n667), .Z(z[9]) );
  XOR U3730 ( .A(n669), .B(z[9]), .Z(z[15]) );
  XOR U3731 ( .A(x[19]), .B(x[17]), .Z(n672) );
  XNOR U3732 ( .A(x[16]), .B(x[22]), .Z(n671) );
  XOR U3733 ( .A(n671), .B(x[18]), .Z(n670) );
  XNOR U3734 ( .A(n672), .B(n670), .Z(n707) );
  XNOR U3735 ( .A(x[21]), .B(n671), .Z(n805) );
  XOR U3736 ( .A(n805), .B(x[20]), .Z(n750) );
  IV U3737 ( .A(n750), .Z(n681) );
  XNOR U3738 ( .A(x[23]), .B(x[20]), .Z(n675) );
  XNOR U3739 ( .A(n672), .B(n675), .Z(n735) );
  NOR U3740 ( .A(n681), .B(n735), .Z(n674) );
  XNOR U3741 ( .A(n805), .B(x[23]), .Z(n766) );
  XNOR U3742 ( .A(x[18]), .B(n766), .Z(n690) );
  XNOR U3743 ( .A(x[17]), .B(n690), .Z(n685) );
  AND U3744 ( .A(x[16]), .B(n685), .Z(n673) );
  XNOR U3745 ( .A(n674), .B(n673), .Z(n678) );
  XNOR U3746 ( .A(n707), .B(n766), .Z(n697) );
  IV U3747 ( .A(n707), .Z(n692) );
  XNOR U3748 ( .A(x[16]), .B(n692), .Z(n712) );
  IV U3749 ( .A(n675), .Z(n740) );
  AND U3750 ( .A(n712), .B(n740), .Z(n680) );
  IV U3751 ( .A(n805), .Z(n699) );
  XNOR U3752 ( .A(n707), .B(n699), .Z(n729) );
  XOR U3753 ( .A(n729), .B(n735), .Z(n732) );
  XOR U3754 ( .A(x[18]), .B(x[20]), .Z(n742) );
  NAND U3755 ( .A(n732), .B(n742), .Z(n676) );
  XNOR U3756 ( .A(n680), .B(n676), .Z(n701) );
  XNOR U3757 ( .A(n697), .B(n701), .Z(n677) );
  XNOR U3758 ( .A(n678), .B(n677), .Z(n724) );
  XOR U3759 ( .A(x[18]), .B(x[23]), .Z(n756) );
  XNOR U3760 ( .A(x[16]), .B(n735), .Z(n736) );
  XNOR U3761 ( .A(n805), .B(n736), .Z(n727) );
  NAND U3762 ( .A(n756), .B(n727), .Z(n679) );
  XNOR U3763 ( .A(n680), .B(n679), .Z(n693) );
  IV U3764 ( .A(n685), .Z(n739) );
  XNOR U3765 ( .A(n739), .B(n681), .Z(n746) );
  AND U3766 ( .A(n735), .B(n746), .Z(n683) );
  AND U3767 ( .A(x[16]), .B(n750), .Z(n682) );
  XNOR U3768 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U3769 ( .A(n736), .B(n684), .Z(n688) );
  NAND U3770 ( .A(x[16]), .B(n735), .Z(n686) );
  OR U3771 ( .A(n686), .B(n685), .Z(n687) );
  NAND U3772 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U3773 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U3774 ( .A(n693), .B(n691), .Z(n713) );
  IV U3775 ( .A(n713), .Z(n720) );
  AND U3776 ( .A(n766), .B(n692), .Z(n695) );
  XOR U3777 ( .A(x[17]), .B(x[23]), .Z(n768) );
  AND U3778 ( .A(n729), .B(n768), .Z(n698) );
  XNOR U3779 ( .A(n698), .B(n693), .Z(n694) );
  XNOR U3780 ( .A(n695), .B(n694), .Z(n719) );
  NANDN U3781 ( .A(n720), .B(n719), .Z(n696) );
  NAND U3782 ( .A(n724), .B(n696), .Z(n706) );
  XNOR U3783 ( .A(n698), .B(n697), .Z(n703) );
  ANDN U3784 ( .B(n699), .A(x[17]), .Z(n700) );
  XNOR U3785 ( .A(n701), .B(n700), .Z(n702) );
  XNOR U3786 ( .A(n703), .B(n702), .Z(n716) );
  XOR U3787 ( .A(n719), .B(n716), .Z(n704) );
  NAND U3788 ( .A(n720), .B(n704), .Z(n705) );
  NAND U3789 ( .A(n706), .B(n705), .Z(n765) );
  ANDN U3790 ( .B(n707), .A(n765), .Z(n731) );
  IV U3791 ( .A(n716), .Z(n722) );
  XOR U3792 ( .A(n724), .B(n720), .Z(n708) );
  NANDN U3793 ( .A(n722), .B(n708), .Z(n711) );
  NANDN U3794 ( .A(n720), .B(n722), .Z(n709) );
  NANDN U3795 ( .A(n719), .B(n709), .Z(n710) );
  NAND U3796 ( .A(n711), .B(n710), .Z(n800) );
  XNOR U3797 ( .A(n765), .B(n800), .Z(n741) );
  AND U3798 ( .A(n712), .B(n741), .Z(n734) );
  OR U3799 ( .A(n719), .B(n716), .Z(n718) );
  ANDN U3800 ( .B(n719), .A(n713), .Z(n714) );
  XNOR U3801 ( .A(n714), .B(n724), .Z(n715) );
  NAND U3802 ( .A(n716), .B(n715), .Z(n717) );
  NAND U3803 ( .A(n718), .B(n717), .Z(n738) );
  NAND U3804 ( .A(n720), .B(n724), .Z(n726) );
  NAND U3805 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U3806 ( .A(n722), .B(n721), .Z(n723) );
  NANDN U3807 ( .A(n724), .B(n723), .Z(n725) );
  NAND U3808 ( .A(n726), .B(n725), .Z(n807) );
  NAND U3809 ( .A(n757), .B(n727), .Z(n728) );
  XNOR U3810 ( .A(n734), .B(n728), .Z(n802) );
  XOR U3811 ( .A(n765), .B(n807), .Z(n767) );
  AND U3812 ( .A(n729), .B(n767), .Z(n752) );
  XNOR U3813 ( .A(n802), .B(n752), .Z(n730) );
  XNOR U3814 ( .A(n731), .B(n730), .Z(n810) );
  NAND U3815 ( .A(n743), .B(n732), .Z(n733) );
  XNOR U3816 ( .A(n734), .B(n733), .Z(n760) );
  AND U3817 ( .A(n735), .B(n745), .Z(n801) );
  NANDN U3818 ( .A(n736), .B(n738), .Z(n737) );
  XNOR U3819 ( .A(n801), .B(n737), .Z(n764) );
  XNOR U3820 ( .A(n760), .B(n764), .Z(n749) );
  XOR U3821 ( .A(n810), .B(n749), .Z(z[16]) );
  AND U3822 ( .A(n739), .B(n738), .Z(n748) );
  AND U3823 ( .A(n741), .B(n740), .Z(n759) );
  NAND U3824 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U3825 ( .A(n759), .B(n744), .Z(n811) );
  AND U3826 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U3827 ( .A(n811), .B(n753), .Z(n747) );
  XNOR U3828 ( .A(n748), .B(n747), .Z(n773) );
  XNOR U3829 ( .A(n773), .B(n749), .Z(n816) );
  AND U3830 ( .A(n750), .B(n800), .Z(n755) );
  NANDN U3831 ( .A(n807), .B(n805), .Z(n751) );
  XNOR U3832 ( .A(n752), .B(n751), .Z(n763) );
  XNOR U3833 ( .A(n753), .B(n763), .Z(n754) );
  XNOR U3834 ( .A(n755), .B(n754), .Z(n762) );
  NAND U3835 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U3836 ( .A(n759), .B(n758), .Z(n769) );
  XNOR U3837 ( .A(n760), .B(n769), .Z(n761) );
  XNOR U3838 ( .A(n762), .B(n761), .Z(n772) );
  XNOR U3839 ( .A(n816), .B(n772), .Z(z[17]) );
  XNOR U3840 ( .A(n764), .B(n763), .Z(z[18]) );
  NOR U3841 ( .A(n766), .B(n765), .Z(n771) );
  AND U3842 ( .A(n768), .B(n767), .Z(n809) );
  XNOR U3843 ( .A(n769), .B(n809), .Z(n770) );
  XNOR U3844 ( .A(n771), .B(n770), .Z(n815) );
  XOR U3845 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U3846 ( .A(n815), .B(n774), .Z(z[19]) );
  AND U3847 ( .A(n776), .B(n775), .Z(n785) );
  AND U3848 ( .A(n778), .B(n777), .Z(n796) );
  NAND U3849 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U3850 ( .A(n796), .B(n781), .Z(n1438) );
  AND U3851 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U3852 ( .A(n1438), .B(n790), .Z(n784) );
  XNOR U3853 ( .A(n785), .B(n784), .Z(n1074) );
  XNOR U3854 ( .A(n1074), .B(n786), .Z(n1581) );
  AND U3855 ( .A(n787), .B(n1427), .Z(n792) );
  NANDN U3856 ( .A(n1434), .B(n1432), .Z(n788) );
  XNOR U3857 ( .A(n789), .B(n788), .Z(n938) );
  XNOR U3858 ( .A(n790), .B(n938), .Z(n791) );
  XNOR U3859 ( .A(n792), .B(n791), .Z(n799) );
  NAND U3860 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U3861 ( .A(n796), .B(n795), .Z(n1070) );
  XNOR U3862 ( .A(n797), .B(n1070), .Z(n798) );
  XNOR U3863 ( .A(n799), .B(n798), .Z(n1073) );
  XNOR U3864 ( .A(n1581), .B(n1073), .Z(z[1]) );
  XOR U3865 ( .A(n810), .B(z[18]), .Z(z[20]) );
  AND U3866 ( .A(x[16]), .B(n800), .Z(n804) );
  XNOR U3867 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U3868 ( .A(n804), .B(n803), .Z(n817) );
  XOR U3869 ( .A(n805), .B(x[17]), .Z(n806) );
  NANDN U3870 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3871 ( .A(n809), .B(n808), .Z(n813) );
  XNOR U3872 ( .A(n811), .B(n810), .Z(n812) );
  XNOR U3873 ( .A(n813), .B(n812), .Z(n814) );
  XNOR U3874 ( .A(n817), .B(n814), .Z(z[21]) );
  XNOR U3875 ( .A(n816), .B(n815), .Z(z[22]) );
  XOR U3876 ( .A(n817), .B(z[17]), .Z(z[23]) );
  XOR U3877 ( .A(x[27]), .B(x[25]), .Z(n820) );
  XNOR U3878 ( .A(x[24]), .B(x[30]), .Z(n819) );
  XOR U3879 ( .A(n819), .B(x[26]), .Z(n818) );
  XNOR U3880 ( .A(n820), .B(n818), .Z(n855) );
  XNOR U3881 ( .A(x[29]), .B(n819), .Z(n928) );
  XOR U3882 ( .A(n928), .B(x[28]), .Z(n898) );
  IV U3883 ( .A(n898), .Z(n829) );
  XNOR U3884 ( .A(x[31]), .B(x[28]), .Z(n823) );
  XNOR U3885 ( .A(n820), .B(n823), .Z(n883) );
  NOR U3886 ( .A(n829), .B(n883), .Z(n822) );
  XNOR U3887 ( .A(n928), .B(x[31]), .Z(n914) );
  XNOR U3888 ( .A(x[26]), .B(n914), .Z(n838) );
  XNOR U3889 ( .A(x[25]), .B(n838), .Z(n833) );
  AND U3890 ( .A(x[24]), .B(n833), .Z(n821) );
  XNOR U3891 ( .A(n822), .B(n821), .Z(n826) );
  XNOR U3892 ( .A(n855), .B(n914), .Z(n845) );
  IV U3893 ( .A(n855), .Z(n840) );
  XNOR U3894 ( .A(x[24]), .B(n840), .Z(n860) );
  IV U3895 ( .A(n823), .Z(n888) );
  AND U3896 ( .A(n860), .B(n888), .Z(n828) );
  IV U3897 ( .A(n928), .Z(n847) );
  XNOR U3898 ( .A(n855), .B(n847), .Z(n877) );
  XOR U3899 ( .A(n877), .B(n883), .Z(n880) );
  XOR U3900 ( .A(x[26]), .B(x[28]), .Z(n890) );
  NAND U3901 ( .A(n880), .B(n890), .Z(n824) );
  XNOR U3902 ( .A(n828), .B(n824), .Z(n849) );
  XNOR U3903 ( .A(n845), .B(n849), .Z(n825) );
  XNOR U3904 ( .A(n826), .B(n825), .Z(n872) );
  XOR U3905 ( .A(x[26]), .B(x[31]), .Z(n904) );
  XNOR U3906 ( .A(x[24]), .B(n883), .Z(n884) );
  XNOR U3907 ( .A(n928), .B(n884), .Z(n875) );
  NAND U3908 ( .A(n904), .B(n875), .Z(n827) );
  XNOR U3909 ( .A(n828), .B(n827), .Z(n841) );
  IV U3910 ( .A(n833), .Z(n887) );
  XNOR U3911 ( .A(n887), .B(n829), .Z(n894) );
  AND U3912 ( .A(n883), .B(n894), .Z(n831) );
  AND U3913 ( .A(x[24]), .B(n898), .Z(n830) );
  XNOR U3914 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U3915 ( .A(n884), .B(n832), .Z(n836) );
  NAND U3916 ( .A(x[24]), .B(n883), .Z(n834) );
  OR U3917 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3918 ( .A(n836), .B(n835), .Z(n837) );
  XNOR U3919 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U3920 ( .A(n841), .B(n839), .Z(n861) );
  IV U3921 ( .A(n861), .Z(n868) );
  AND U3922 ( .A(n914), .B(n840), .Z(n843) );
  XOR U3923 ( .A(x[25]), .B(x[31]), .Z(n916) );
  AND U3924 ( .A(n877), .B(n916), .Z(n846) );
  XNOR U3925 ( .A(n846), .B(n841), .Z(n842) );
  XNOR U3926 ( .A(n843), .B(n842), .Z(n867) );
  NANDN U3927 ( .A(n868), .B(n867), .Z(n844) );
  NAND U3928 ( .A(n872), .B(n844), .Z(n854) );
  XNOR U3929 ( .A(n846), .B(n845), .Z(n851) );
  ANDN U3930 ( .B(n847), .A(x[25]), .Z(n848) );
  XNOR U3931 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U3932 ( .A(n851), .B(n850), .Z(n864) );
  XOR U3933 ( .A(n867), .B(n864), .Z(n852) );
  NAND U3934 ( .A(n868), .B(n852), .Z(n853) );
  NAND U3935 ( .A(n854), .B(n853), .Z(n913) );
  ANDN U3936 ( .B(n855), .A(n913), .Z(n879) );
  IV U3937 ( .A(n864), .Z(n870) );
  XOR U3938 ( .A(n872), .B(n868), .Z(n856) );
  NANDN U3939 ( .A(n870), .B(n856), .Z(n859) );
  NANDN U3940 ( .A(n868), .B(n870), .Z(n857) );
  NANDN U3941 ( .A(n867), .B(n857), .Z(n858) );
  NAND U3942 ( .A(n859), .B(n858), .Z(n923) );
  XNOR U3943 ( .A(n913), .B(n923), .Z(n889) );
  AND U3944 ( .A(n860), .B(n889), .Z(n882) );
  OR U3945 ( .A(n867), .B(n864), .Z(n866) );
  ANDN U3946 ( .B(n867), .A(n861), .Z(n862) );
  XNOR U3947 ( .A(n862), .B(n872), .Z(n863) );
  NAND U3948 ( .A(n864), .B(n863), .Z(n865) );
  NAND U3949 ( .A(n866), .B(n865), .Z(n886) );
  NAND U3950 ( .A(n868), .B(n872), .Z(n874) );
  NAND U3951 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U3952 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U3953 ( .A(n872), .B(n871), .Z(n873) );
  NAND U3954 ( .A(n874), .B(n873), .Z(n930) );
  NAND U3955 ( .A(n905), .B(n875), .Z(n876) );
  XNOR U3956 ( .A(n882), .B(n876), .Z(n925) );
  XOR U3957 ( .A(n913), .B(n930), .Z(n915) );
  AND U3958 ( .A(n877), .B(n915), .Z(n900) );
  XNOR U3959 ( .A(n925), .B(n900), .Z(n878) );
  XNOR U3960 ( .A(n879), .B(n878), .Z(n933) );
  NAND U3961 ( .A(n891), .B(n880), .Z(n881) );
  XNOR U3962 ( .A(n882), .B(n881), .Z(n908) );
  AND U3963 ( .A(n883), .B(n893), .Z(n924) );
  NANDN U3964 ( .A(n884), .B(n886), .Z(n885) );
  XNOR U3965 ( .A(n924), .B(n885), .Z(n912) );
  XNOR U3966 ( .A(n908), .B(n912), .Z(n897) );
  XOR U3967 ( .A(n933), .B(n897), .Z(z[24]) );
  AND U3968 ( .A(n887), .B(n886), .Z(n896) );
  AND U3969 ( .A(n889), .B(n888), .Z(n907) );
  NAND U3970 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U3971 ( .A(n907), .B(n892), .Z(n934) );
  AND U3972 ( .A(n894), .B(n893), .Z(n901) );
  XNOR U3973 ( .A(n934), .B(n901), .Z(n895) );
  XNOR U3974 ( .A(n896), .B(n895), .Z(n921) );
  XNOR U3975 ( .A(n921), .B(n897), .Z(n941) );
  AND U3976 ( .A(n898), .B(n923), .Z(n903) );
  NANDN U3977 ( .A(n930), .B(n928), .Z(n899) );
  XNOR U3978 ( .A(n900), .B(n899), .Z(n911) );
  XNOR U3979 ( .A(n901), .B(n911), .Z(n902) );
  XNOR U3980 ( .A(n903), .B(n902), .Z(n910) );
  NAND U3981 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3982 ( .A(n907), .B(n906), .Z(n917) );
  XNOR U3983 ( .A(n908), .B(n917), .Z(n909) );
  XNOR U3984 ( .A(n910), .B(n909), .Z(n920) );
  XNOR U3985 ( .A(n941), .B(n920), .Z(z[25]) );
  XNOR U3986 ( .A(n912), .B(n911), .Z(z[26]) );
  NOR U3987 ( .A(n914), .B(n913), .Z(n919) );
  AND U3988 ( .A(n916), .B(n915), .Z(n932) );
  XNOR U3989 ( .A(n917), .B(n932), .Z(n918) );
  XNOR U3990 ( .A(n919), .B(n918), .Z(n940) );
  XOR U3991 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U3992 ( .A(n940), .B(n922), .Z(z[27]) );
  XOR U3993 ( .A(n933), .B(z[26]), .Z(z[28]) );
  AND U3994 ( .A(x[24]), .B(n923), .Z(n927) );
  XNOR U3995 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U3996 ( .A(n927), .B(n926), .Z(n942) );
  XOR U3997 ( .A(n928), .B(x[25]), .Z(n929) );
  NANDN U3998 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U3999 ( .A(n932), .B(n931), .Z(n936) );
  XNOR U4000 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U4001 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U4002 ( .A(n942), .B(n937), .Z(z[29]) );
  XNOR U4003 ( .A(n939), .B(n938), .Z(z[2]) );
  XNOR U4004 ( .A(n941), .B(n940), .Z(z[30]) );
  XOR U4005 ( .A(n942), .B(z[25]), .Z(z[31]) );
  XOR U4006 ( .A(x[35]), .B(x[33]), .Z(n945) );
  XNOR U4007 ( .A(x[32]), .B(x[38]), .Z(n944) );
  XOR U4008 ( .A(n944), .B(x[34]), .Z(n943) );
  XNOR U4009 ( .A(n945), .B(n943), .Z(n980) );
  XNOR U4010 ( .A(x[37]), .B(n944), .Z(n1053) );
  XOR U4011 ( .A(n1053), .B(x[36]), .Z(n1023) );
  IV U4012 ( .A(n1023), .Z(n954) );
  XNOR U4013 ( .A(x[39]), .B(x[36]), .Z(n948) );
  XNOR U4014 ( .A(n945), .B(n948), .Z(n1008) );
  NOR U4015 ( .A(n954), .B(n1008), .Z(n947) );
  XNOR U4016 ( .A(n1053), .B(x[39]), .Z(n1039) );
  XNOR U4017 ( .A(x[34]), .B(n1039), .Z(n963) );
  XNOR U4018 ( .A(x[33]), .B(n963), .Z(n958) );
  AND U4019 ( .A(x[32]), .B(n958), .Z(n946) );
  XNOR U4020 ( .A(n947), .B(n946), .Z(n951) );
  XNOR U4021 ( .A(n980), .B(n1039), .Z(n970) );
  IV U4022 ( .A(n980), .Z(n965) );
  XNOR U4023 ( .A(x[32]), .B(n965), .Z(n985) );
  IV U4024 ( .A(n948), .Z(n1013) );
  AND U4025 ( .A(n985), .B(n1013), .Z(n953) );
  IV U4026 ( .A(n1053), .Z(n972) );
  XNOR U4027 ( .A(n980), .B(n972), .Z(n1002) );
  XOR U4028 ( .A(n1002), .B(n1008), .Z(n1005) );
  XOR U4029 ( .A(x[34]), .B(x[36]), .Z(n1015) );
  NAND U4030 ( .A(n1005), .B(n1015), .Z(n949) );
  XNOR U4031 ( .A(n953), .B(n949), .Z(n974) );
  XNOR U4032 ( .A(n970), .B(n974), .Z(n950) );
  XNOR U4033 ( .A(n951), .B(n950), .Z(n997) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1029) );
  XNOR U4035 ( .A(x[32]), .B(n1008), .Z(n1009) );
  XNOR U4036 ( .A(n1053), .B(n1009), .Z(n1000) );
  NAND U4037 ( .A(n1029), .B(n1000), .Z(n952) );
  XNOR U4038 ( .A(n953), .B(n952), .Z(n966) );
  IV U4039 ( .A(n958), .Z(n1012) );
  XNOR U4040 ( .A(n1012), .B(n954), .Z(n1019) );
  AND U4041 ( .A(n1008), .B(n1019), .Z(n956) );
  AND U4042 ( .A(x[32]), .B(n1023), .Z(n955) );
  XNOR U4043 ( .A(n956), .B(n955), .Z(n957) );
  NANDN U4044 ( .A(n1009), .B(n957), .Z(n961) );
  NAND U4045 ( .A(x[32]), .B(n1008), .Z(n959) );
  OR U4046 ( .A(n959), .B(n958), .Z(n960) );
  NAND U4047 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U4048 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U4049 ( .A(n966), .B(n964), .Z(n986) );
  IV U4050 ( .A(n986), .Z(n993) );
  AND U4051 ( .A(n1039), .B(n965), .Z(n968) );
  XOR U4052 ( .A(x[33]), .B(x[39]), .Z(n1041) );
  AND U4053 ( .A(n1002), .B(n1041), .Z(n971) );
  XNOR U4054 ( .A(n971), .B(n966), .Z(n967) );
  XNOR U4055 ( .A(n968), .B(n967), .Z(n992) );
  NANDN U4056 ( .A(n993), .B(n992), .Z(n969) );
  NAND U4057 ( .A(n997), .B(n969), .Z(n979) );
  XNOR U4058 ( .A(n971), .B(n970), .Z(n976) );
  ANDN U4059 ( .B(n972), .A(x[33]), .Z(n973) );
  XNOR U4060 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U4061 ( .A(n976), .B(n975), .Z(n989) );
  XOR U4062 ( .A(n992), .B(n989), .Z(n977) );
  NAND U4063 ( .A(n993), .B(n977), .Z(n978) );
  NAND U4064 ( .A(n979), .B(n978), .Z(n1038) );
  ANDN U4065 ( .B(n980), .A(n1038), .Z(n1004) );
  IV U4066 ( .A(n989), .Z(n995) );
  XOR U4067 ( .A(n997), .B(n993), .Z(n981) );
  NANDN U4068 ( .A(n995), .B(n981), .Z(n984) );
  NANDN U4069 ( .A(n993), .B(n995), .Z(n982) );
  NANDN U4070 ( .A(n992), .B(n982), .Z(n983) );
  NAND U4071 ( .A(n984), .B(n983), .Z(n1048) );
  XNOR U4072 ( .A(n1038), .B(n1048), .Z(n1014) );
  AND U4073 ( .A(n985), .B(n1014), .Z(n1007) );
  OR U4074 ( .A(n992), .B(n989), .Z(n991) );
  ANDN U4075 ( .B(n992), .A(n986), .Z(n987) );
  XNOR U4076 ( .A(n987), .B(n997), .Z(n988) );
  NAND U4077 ( .A(n989), .B(n988), .Z(n990) );
  NAND U4078 ( .A(n991), .B(n990), .Z(n1011) );
  NAND U4079 ( .A(n993), .B(n997), .Z(n999) );
  NAND U4080 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U4081 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U4082 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4083 ( .A(n999), .B(n998), .Z(n1055) );
  NAND U4084 ( .A(n1030), .B(n1000), .Z(n1001) );
  XNOR U4085 ( .A(n1007), .B(n1001), .Z(n1050) );
  XOR U4086 ( .A(n1038), .B(n1055), .Z(n1040) );
  AND U4087 ( .A(n1002), .B(n1040), .Z(n1025) );
  XNOR U4088 ( .A(n1050), .B(n1025), .Z(n1003) );
  XNOR U4089 ( .A(n1004), .B(n1003), .Z(n1058) );
  NAND U4090 ( .A(n1016), .B(n1005), .Z(n1006) );
  XNOR U4091 ( .A(n1007), .B(n1006), .Z(n1033) );
  AND U4092 ( .A(n1008), .B(n1018), .Z(n1049) );
  NANDN U4093 ( .A(n1009), .B(n1011), .Z(n1010) );
  XNOR U4094 ( .A(n1049), .B(n1010), .Z(n1037) );
  XNOR U4095 ( .A(n1033), .B(n1037), .Z(n1022) );
  XOR U4096 ( .A(n1058), .B(n1022), .Z(z[32]) );
  AND U4097 ( .A(n1012), .B(n1011), .Z(n1021) );
  AND U4098 ( .A(n1014), .B(n1013), .Z(n1032) );
  NAND U4099 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U4100 ( .A(n1032), .B(n1017), .Z(n1059) );
  AND U4101 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U4102 ( .A(n1059), .B(n1026), .Z(n1020) );
  XNOR U4103 ( .A(n1021), .B(n1020), .Z(n1046) );
  XNOR U4104 ( .A(n1046), .B(n1022), .Z(n1064) );
  AND U4105 ( .A(n1023), .B(n1048), .Z(n1028) );
  NANDN U4106 ( .A(n1055), .B(n1053), .Z(n1024) );
  XNOR U4107 ( .A(n1025), .B(n1024), .Z(n1036) );
  XNOR U4108 ( .A(n1026), .B(n1036), .Z(n1027) );
  XNOR U4109 ( .A(n1028), .B(n1027), .Z(n1035) );
  NAND U4110 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U4111 ( .A(n1032), .B(n1031), .Z(n1042) );
  XNOR U4112 ( .A(n1033), .B(n1042), .Z(n1034) );
  XNOR U4113 ( .A(n1035), .B(n1034), .Z(n1045) );
  XNOR U4114 ( .A(n1064), .B(n1045), .Z(z[33]) );
  XNOR U4115 ( .A(n1037), .B(n1036), .Z(z[34]) );
  NOR U4116 ( .A(n1039), .B(n1038), .Z(n1044) );
  AND U4117 ( .A(n1041), .B(n1040), .Z(n1057) );
  XNOR U4118 ( .A(n1042), .B(n1057), .Z(n1043) );
  XNOR U4119 ( .A(n1044), .B(n1043), .Z(n1063) );
  XOR U4120 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U4121 ( .A(n1063), .B(n1047), .Z(z[35]) );
  XOR U4122 ( .A(n1058), .B(z[34]), .Z(z[36]) );
  AND U4123 ( .A(x[32]), .B(n1048), .Z(n1052) );
  XNOR U4124 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U4125 ( .A(n1052), .B(n1051), .Z(n1065) );
  XOR U4126 ( .A(n1053), .B(x[33]), .Z(n1054) );
  NANDN U4127 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U4128 ( .A(n1057), .B(n1056), .Z(n1061) );
  XNOR U4129 ( .A(n1059), .B(n1058), .Z(n1060) );
  XNOR U4130 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U4131 ( .A(n1065), .B(n1062), .Z(z[37]) );
  XNOR U4132 ( .A(n1064), .B(n1063), .Z(z[38]) );
  XOR U4133 ( .A(n1065), .B(z[33]), .Z(z[39]) );
  NOR U4134 ( .A(n1067), .B(n1066), .Z(n1072) );
  AND U4135 ( .A(n1069), .B(n1068), .Z(n1436) );
  XNOR U4136 ( .A(n1070), .B(n1436), .Z(n1071) );
  XNOR U4137 ( .A(n1072), .B(n1071), .Z(n1580) );
  XOR U4138 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U4139 ( .A(n1580), .B(n1075), .Z(z[3]) );
  XOR U4140 ( .A(x[43]), .B(x[41]), .Z(n1078) );
  XNOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1077) );
  XOR U4142 ( .A(n1077), .B(x[42]), .Z(n1076) );
  XNOR U4143 ( .A(n1078), .B(n1076), .Z(n1113) );
  XNOR U4144 ( .A(x[45]), .B(n1077), .Z(n1186) );
  XOR U4145 ( .A(n1186), .B(x[44]), .Z(n1156) );
  IV U4146 ( .A(n1156), .Z(n1087) );
  XNOR U4147 ( .A(x[47]), .B(x[44]), .Z(n1081) );
  XNOR U4148 ( .A(n1078), .B(n1081), .Z(n1141) );
  NOR U4149 ( .A(n1087), .B(n1141), .Z(n1080) );
  XNOR U4150 ( .A(n1186), .B(x[47]), .Z(n1172) );
  XNOR U4151 ( .A(x[42]), .B(n1172), .Z(n1096) );
  XNOR U4152 ( .A(x[41]), .B(n1096), .Z(n1091) );
  AND U4153 ( .A(x[40]), .B(n1091), .Z(n1079) );
  XNOR U4154 ( .A(n1080), .B(n1079), .Z(n1084) );
  XNOR U4155 ( .A(n1113), .B(n1172), .Z(n1103) );
  IV U4156 ( .A(n1113), .Z(n1098) );
  XNOR U4157 ( .A(x[40]), .B(n1098), .Z(n1118) );
  IV U4158 ( .A(n1081), .Z(n1146) );
  AND U4159 ( .A(n1118), .B(n1146), .Z(n1086) );
  IV U4160 ( .A(n1186), .Z(n1105) );
  XNOR U4161 ( .A(n1113), .B(n1105), .Z(n1135) );
  XOR U4162 ( .A(n1135), .B(n1141), .Z(n1138) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1148) );
  NAND U4164 ( .A(n1138), .B(n1148), .Z(n1082) );
  XNOR U4165 ( .A(n1086), .B(n1082), .Z(n1107) );
  XNOR U4166 ( .A(n1103), .B(n1107), .Z(n1083) );
  XNOR U4167 ( .A(n1084), .B(n1083), .Z(n1130) );
  XOR U4168 ( .A(x[42]), .B(x[47]), .Z(n1162) );
  XNOR U4169 ( .A(x[40]), .B(n1141), .Z(n1142) );
  XNOR U4170 ( .A(n1186), .B(n1142), .Z(n1133) );
  NAND U4171 ( .A(n1162), .B(n1133), .Z(n1085) );
  XNOR U4172 ( .A(n1086), .B(n1085), .Z(n1099) );
  IV U4173 ( .A(n1091), .Z(n1145) );
  XNOR U4174 ( .A(n1145), .B(n1087), .Z(n1152) );
  AND U4175 ( .A(n1141), .B(n1152), .Z(n1089) );
  AND U4176 ( .A(x[40]), .B(n1156), .Z(n1088) );
  XNOR U4177 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U4178 ( .A(n1142), .B(n1090), .Z(n1094) );
  NAND U4179 ( .A(x[40]), .B(n1141), .Z(n1092) );
  OR U4180 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U4181 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U4182 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U4183 ( .A(n1099), .B(n1097), .Z(n1119) );
  IV U4184 ( .A(n1119), .Z(n1126) );
  AND U4185 ( .A(n1172), .B(n1098), .Z(n1101) );
  XOR U4186 ( .A(x[41]), .B(x[47]), .Z(n1174) );
  AND U4187 ( .A(n1135), .B(n1174), .Z(n1104) );
  XNOR U4188 ( .A(n1104), .B(n1099), .Z(n1100) );
  XNOR U4189 ( .A(n1101), .B(n1100), .Z(n1125) );
  NANDN U4190 ( .A(n1126), .B(n1125), .Z(n1102) );
  NAND U4191 ( .A(n1130), .B(n1102), .Z(n1112) );
  XNOR U4192 ( .A(n1104), .B(n1103), .Z(n1109) );
  ANDN U4193 ( .B(n1105), .A(x[41]), .Z(n1106) );
  XNOR U4194 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U4195 ( .A(n1109), .B(n1108), .Z(n1122) );
  XOR U4196 ( .A(n1125), .B(n1122), .Z(n1110) );
  NAND U4197 ( .A(n1126), .B(n1110), .Z(n1111) );
  NAND U4198 ( .A(n1112), .B(n1111), .Z(n1171) );
  ANDN U4199 ( .B(n1113), .A(n1171), .Z(n1137) );
  IV U4200 ( .A(n1122), .Z(n1128) );
  XOR U4201 ( .A(n1130), .B(n1126), .Z(n1114) );
  NANDN U4202 ( .A(n1128), .B(n1114), .Z(n1117) );
  NANDN U4203 ( .A(n1126), .B(n1128), .Z(n1115) );
  NANDN U4204 ( .A(n1125), .B(n1115), .Z(n1116) );
  NAND U4205 ( .A(n1117), .B(n1116), .Z(n1181) );
  XNOR U4206 ( .A(n1171), .B(n1181), .Z(n1147) );
  AND U4207 ( .A(n1118), .B(n1147), .Z(n1140) );
  OR U4208 ( .A(n1125), .B(n1122), .Z(n1124) );
  ANDN U4209 ( .B(n1125), .A(n1119), .Z(n1120) );
  XNOR U4210 ( .A(n1120), .B(n1130), .Z(n1121) );
  NAND U4211 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U4212 ( .A(n1124), .B(n1123), .Z(n1144) );
  NAND U4213 ( .A(n1126), .B(n1130), .Z(n1132) );
  NAND U4214 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U4215 ( .A(n1128), .B(n1127), .Z(n1129) );
  NANDN U4216 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U4217 ( .A(n1132), .B(n1131), .Z(n1188) );
  NAND U4218 ( .A(n1163), .B(n1133), .Z(n1134) );
  XNOR U4219 ( .A(n1140), .B(n1134), .Z(n1183) );
  XOR U4220 ( .A(n1171), .B(n1188), .Z(n1173) );
  AND U4221 ( .A(n1135), .B(n1173), .Z(n1158) );
  XNOR U4222 ( .A(n1183), .B(n1158), .Z(n1136) );
  XNOR U4223 ( .A(n1137), .B(n1136), .Z(n1191) );
  NAND U4224 ( .A(n1149), .B(n1138), .Z(n1139) );
  XNOR U4225 ( .A(n1140), .B(n1139), .Z(n1166) );
  AND U4226 ( .A(n1141), .B(n1151), .Z(n1182) );
  NANDN U4227 ( .A(n1142), .B(n1144), .Z(n1143) );
  XNOR U4228 ( .A(n1182), .B(n1143), .Z(n1170) );
  XNOR U4229 ( .A(n1166), .B(n1170), .Z(n1155) );
  XOR U4230 ( .A(n1191), .B(n1155), .Z(z[40]) );
  AND U4231 ( .A(n1145), .B(n1144), .Z(n1154) );
  AND U4232 ( .A(n1147), .B(n1146), .Z(n1165) );
  NAND U4233 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U4234 ( .A(n1165), .B(n1150), .Z(n1192) );
  AND U4235 ( .A(n1152), .B(n1151), .Z(n1159) );
  XNOR U4236 ( .A(n1192), .B(n1159), .Z(n1153) );
  XNOR U4237 ( .A(n1154), .B(n1153), .Z(n1179) );
  XNOR U4238 ( .A(n1179), .B(n1155), .Z(n1197) );
  AND U4239 ( .A(n1156), .B(n1181), .Z(n1161) );
  NANDN U4240 ( .A(n1188), .B(n1186), .Z(n1157) );
  XNOR U4241 ( .A(n1158), .B(n1157), .Z(n1169) );
  XNOR U4242 ( .A(n1159), .B(n1169), .Z(n1160) );
  XNOR U4243 ( .A(n1161), .B(n1160), .Z(n1168) );
  NAND U4244 ( .A(n1163), .B(n1162), .Z(n1164) );
  XNOR U4245 ( .A(n1165), .B(n1164), .Z(n1175) );
  XNOR U4246 ( .A(n1166), .B(n1175), .Z(n1167) );
  XNOR U4247 ( .A(n1168), .B(n1167), .Z(n1178) );
  XNOR U4248 ( .A(n1197), .B(n1178), .Z(z[41]) );
  XNOR U4249 ( .A(n1170), .B(n1169), .Z(z[42]) );
  NOR U4250 ( .A(n1172), .B(n1171), .Z(n1177) );
  AND U4251 ( .A(n1174), .B(n1173), .Z(n1190) );
  XNOR U4252 ( .A(n1175), .B(n1190), .Z(n1176) );
  XNOR U4253 ( .A(n1177), .B(n1176), .Z(n1196) );
  XOR U4254 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4255 ( .A(n1196), .B(n1180), .Z(z[43]) );
  XOR U4256 ( .A(n1191), .B(z[42]), .Z(z[44]) );
  AND U4257 ( .A(x[40]), .B(n1181), .Z(n1185) );
  XNOR U4258 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U4259 ( .A(n1185), .B(n1184), .Z(n1198) );
  XOR U4260 ( .A(n1186), .B(x[41]), .Z(n1187) );
  NANDN U4261 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U4262 ( .A(n1190), .B(n1189), .Z(n1194) );
  XNOR U4263 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U4264 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U4265 ( .A(n1198), .B(n1195), .Z(z[45]) );
  XNOR U4266 ( .A(n1197), .B(n1196), .Z(z[46]) );
  XOR U4267 ( .A(n1198), .B(z[41]), .Z(z[47]) );
  XOR U4268 ( .A(x[51]), .B(x[49]), .Z(n1201) );
  XNOR U4269 ( .A(x[48]), .B(x[54]), .Z(n1200) );
  XOR U4270 ( .A(n1200), .B(x[50]), .Z(n1199) );
  XNOR U4271 ( .A(n1201), .B(n1199), .Z(n1236) );
  XNOR U4272 ( .A(x[53]), .B(n1200), .Z(n1309) );
  XOR U4273 ( .A(n1309), .B(x[52]), .Z(n1279) );
  IV U4274 ( .A(n1279), .Z(n1210) );
  XNOR U4275 ( .A(x[55]), .B(x[52]), .Z(n1204) );
  XNOR U4276 ( .A(n1201), .B(n1204), .Z(n1264) );
  NOR U4277 ( .A(n1210), .B(n1264), .Z(n1203) );
  XNOR U4278 ( .A(n1309), .B(x[55]), .Z(n1295) );
  XNOR U4279 ( .A(x[50]), .B(n1295), .Z(n1219) );
  XNOR U4280 ( .A(x[49]), .B(n1219), .Z(n1214) );
  AND U4281 ( .A(x[48]), .B(n1214), .Z(n1202) );
  XNOR U4282 ( .A(n1203), .B(n1202), .Z(n1207) );
  XNOR U4283 ( .A(n1236), .B(n1295), .Z(n1226) );
  IV U4284 ( .A(n1236), .Z(n1221) );
  XNOR U4285 ( .A(x[48]), .B(n1221), .Z(n1241) );
  IV U4286 ( .A(n1204), .Z(n1269) );
  AND U4287 ( .A(n1241), .B(n1269), .Z(n1209) );
  IV U4288 ( .A(n1309), .Z(n1228) );
  XNOR U4289 ( .A(n1236), .B(n1228), .Z(n1258) );
  XOR U4290 ( .A(n1258), .B(n1264), .Z(n1261) );
  XOR U4291 ( .A(x[50]), .B(x[52]), .Z(n1271) );
  NAND U4292 ( .A(n1261), .B(n1271), .Z(n1205) );
  XNOR U4293 ( .A(n1209), .B(n1205), .Z(n1230) );
  XNOR U4294 ( .A(n1226), .B(n1230), .Z(n1206) );
  XNOR U4295 ( .A(n1207), .B(n1206), .Z(n1253) );
  XOR U4296 ( .A(x[50]), .B(x[55]), .Z(n1285) );
  XNOR U4297 ( .A(x[48]), .B(n1264), .Z(n1265) );
  XNOR U4298 ( .A(n1309), .B(n1265), .Z(n1256) );
  NAND U4299 ( .A(n1285), .B(n1256), .Z(n1208) );
  XNOR U4300 ( .A(n1209), .B(n1208), .Z(n1222) );
  IV U4301 ( .A(n1214), .Z(n1268) );
  XNOR U4302 ( .A(n1268), .B(n1210), .Z(n1275) );
  AND U4303 ( .A(n1264), .B(n1275), .Z(n1212) );
  AND U4304 ( .A(x[48]), .B(n1279), .Z(n1211) );
  XNOR U4305 ( .A(n1212), .B(n1211), .Z(n1213) );
  NANDN U4306 ( .A(n1265), .B(n1213), .Z(n1217) );
  NAND U4307 ( .A(x[48]), .B(n1264), .Z(n1215) );
  OR U4308 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4309 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U4310 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U4311 ( .A(n1222), .B(n1220), .Z(n1242) );
  IV U4312 ( .A(n1242), .Z(n1249) );
  AND U4313 ( .A(n1295), .B(n1221), .Z(n1224) );
  XOR U4314 ( .A(x[49]), .B(x[55]), .Z(n1297) );
  AND U4315 ( .A(n1258), .B(n1297), .Z(n1227) );
  XNOR U4316 ( .A(n1227), .B(n1222), .Z(n1223) );
  XNOR U4317 ( .A(n1224), .B(n1223), .Z(n1248) );
  NANDN U4318 ( .A(n1249), .B(n1248), .Z(n1225) );
  NAND U4319 ( .A(n1253), .B(n1225), .Z(n1235) );
  XNOR U4320 ( .A(n1227), .B(n1226), .Z(n1232) );
  ANDN U4321 ( .B(n1228), .A(x[49]), .Z(n1229) );
  XNOR U4322 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U4323 ( .A(n1232), .B(n1231), .Z(n1245) );
  XOR U4324 ( .A(n1248), .B(n1245), .Z(n1233) );
  NAND U4325 ( .A(n1249), .B(n1233), .Z(n1234) );
  NAND U4326 ( .A(n1235), .B(n1234), .Z(n1294) );
  ANDN U4327 ( .B(n1236), .A(n1294), .Z(n1260) );
  IV U4328 ( .A(n1245), .Z(n1251) );
  XOR U4329 ( .A(n1253), .B(n1249), .Z(n1237) );
  NANDN U4330 ( .A(n1251), .B(n1237), .Z(n1240) );
  NANDN U4331 ( .A(n1249), .B(n1251), .Z(n1238) );
  NANDN U4332 ( .A(n1248), .B(n1238), .Z(n1239) );
  NAND U4333 ( .A(n1240), .B(n1239), .Z(n1304) );
  XNOR U4334 ( .A(n1294), .B(n1304), .Z(n1270) );
  AND U4335 ( .A(n1241), .B(n1270), .Z(n1263) );
  OR U4336 ( .A(n1248), .B(n1245), .Z(n1247) );
  ANDN U4337 ( .B(n1248), .A(n1242), .Z(n1243) );
  XNOR U4338 ( .A(n1243), .B(n1253), .Z(n1244) );
  NAND U4339 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U4340 ( .A(n1247), .B(n1246), .Z(n1267) );
  NAND U4341 ( .A(n1249), .B(n1253), .Z(n1255) );
  NAND U4342 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U4343 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U4344 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U4345 ( .A(n1255), .B(n1254), .Z(n1311) );
  NAND U4346 ( .A(n1286), .B(n1256), .Z(n1257) );
  XNOR U4347 ( .A(n1263), .B(n1257), .Z(n1306) );
  XOR U4348 ( .A(n1294), .B(n1311), .Z(n1296) );
  AND U4349 ( .A(n1258), .B(n1296), .Z(n1281) );
  XNOR U4350 ( .A(n1306), .B(n1281), .Z(n1259) );
  XNOR U4351 ( .A(n1260), .B(n1259), .Z(n1314) );
  NAND U4352 ( .A(n1272), .B(n1261), .Z(n1262) );
  XNOR U4353 ( .A(n1263), .B(n1262), .Z(n1289) );
  AND U4354 ( .A(n1264), .B(n1274), .Z(n1305) );
  NANDN U4355 ( .A(n1265), .B(n1267), .Z(n1266) );
  XNOR U4356 ( .A(n1305), .B(n1266), .Z(n1293) );
  XNOR U4357 ( .A(n1289), .B(n1293), .Z(n1278) );
  XOR U4358 ( .A(n1314), .B(n1278), .Z(z[48]) );
  AND U4359 ( .A(n1268), .B(n1267), .Z(n1277) );
  AND U4360 ( .A(n1270), .B(n1269), .Z(n1288) );
  NAND U4361 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U4362 ( .A(n1288), .B(n1273), .Z(n1315) );
  AND U4363 ( .A(n1275), .B(n1274), .Z(n1282) );
  XNOR U4364 ( .A(n1315), .B(n1282), .Z(n1276) );
  XNOR U4365 ( .A(n1277), .B(n1276), .Z(n1302) );
  XNOR U4366 ( .A(n1302), .B(n1278), .Z(n1320) );
  AND U4367 ( .A(n1279), .B(n1304), .Z(n1284) );
  NANDN U4368 ( .A(n1311), .B(n1309), .Z(n1280) );
  XNOR U4369 ( .A(n1281), .B(n1280), .Z(n1292) );
  XNOR U4370 ( .A(n1282), .B(n1292), .Z(n1283) );
  XNOR U4371 ( .A(n1284), .B(n1283), .Z(n1291) );
  NAND U4372 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U4373 ( .A(n1288), .B(n1287), .Z(n1298) );
  XNOR U4374 ( .A(n1289), .B(n1298), .Z(n1290) );
  XNOR U4375 ( .A(n1291), .B(n1290), .Z(n1301) );
  XNOR U4376 ( .A(n1320), .B(n1301), .Z(z[49]) );
  XOR U4377 ( .A(n1437), .B(z[2]), .Z(z[4]) );
  XNOR U4378 ( .A(n1293), .B(n1292), .Z(z[50]) );
  NOR U4379 ( .A(n1295), .B(n1294), .Z(n1300) );
  AND U4380 ( .A(n1297), .B(n1296), .Z(n1313) );
  XNOR U4381 ( .A(n1298), .B(n1313), .Z(n1299) );
  XNOR U4382 ( .A(n1300), .B(n1299), .Z(n1319) );
  XOR U4383 ( .A(n1302), .B(n1301), .Z(n1303) );
  XNOR U4384 ( .A(n1319), .B(n1303), .Z(z[51]) );
  XOR U4385 ( .A(n1314), .B(z[50]), .Z(z[52]) );
  AND U4386 ( .A(x[48]), .B(n1304), .Z(n1308) );
  XNOR U4387 ( .A(n1306), .B(n1305), .Z(n1307) );
  XNOR U4388 ( .A(n1308), .B(n1307), .Z(n1321) );
  XOR U4389 ( .A(n1309), .B(x[49]), .Z(n1310) );
  NANDN U4390 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U4391 ( .A(n1313), .B(n1312), .Z(n1317) );
  XNOR U4392 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U4393 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U4394 ( .A(n1321), .B(n1318), .Z(z[53]) );
  XNOR U4395 ( .A(n1320), .B(n1319), .Z(z[54]) );
  XOR U4396 ( .A(n1321), .B(z[49]), .Z(z[55]) );
  XOR U4397 ( .A(x[59]), .B(x[57]), .Z(n1324) );
  XNOR U4398 ( .A(x[56]), .B(x[62]), .Z(n1323) );
  XOR U4399 ( .A(n1323), .B(x[58]), .Z(n1322) );
  XNOR U4400 ( .A(n1324), .B(n1322), .Z(n1359) );
  XNOR U4401 ( .A(x[61]), .B(n1323), .Z(n1447) );
  XOR U4402 ( .A(n1447), .B(x[60]), .Z(n1402) );
  IV U4403 ( .A(n1402), .Z(n1333) );
  XNOR U4404 ( .A(x[63]), .B(x[60]), .Z(n1327) );
  XNOR U4405 ( .A(n1324), .B(n1327), .Z(n1387) );
  NOR U4406 ( .A(n1333), .B(n1387), .Z(n1326) );
  XNOR U4407 ( .A(n1447), .B(x[63]), .Z(n1418) );
  XNOR U4408 ( .A(x[58]), .B(n1418), .Z(n1342) );
  XNOR U4409 ( .A(x[57]), .B(n1342), .Z(n1337) );
  AND U4410 ( .A(x[56]), .B(n1337), .Z(n1325) );
  XNOR U4411 ( .A(n1326), .B(n1325), .Z(n1330) );
  XNOR U4412 ( .A(n1359), .B(n1418), .Z(n1349) );
  IV U4413 ( .A(n1359), .Z(n1344) );
  XNOR U4414 ( .A(x[56]), .B(n1344), .Z(n1364) );
  IV U4415 ( .A(n1327), .Z(n1392) );
  AND U4416 ( .A(n1364), .B(n1392), .Z(n1332) );
  IV U4417 ( .A(n1447), .Z(n1351) );
  XNOR U4418 ( .A(n1359), .B(n1351), .Z(n1381) );
  XOR U4419 ( .A(n1381), .B(n1387), .Z(n1384) );
  XOR U4420 ( .A(x[58]), .B(x[60]), .Z(n1394) );
  NAND U4421 ( .A(n1384), .B(n1394), .Z(n1328) );
  XNOR U4422 ( .A(n1332), .B(n1328), .Z(n1353) );
  XNOR U4423 ( .A(n1349), .B(n1353), .Z(n1329) );
  XNOR U4424 ( .A(n1330), .B(n1329), .Z(n1376) );
  XOR U4425 ( .A(x[58]), .B(x[63]), .Z(n1408) );
  XNOR U4426 ( .A(x[56]), .B(n1387), .Z(n1388) );
  XNOR U4427 ( .A(n1447), .B(n1388), .Z(n1379) );
  NAND U4428 ( .A(n1408), .B(n1379), .Z(n1331) );
  XNOR U4429 ( .A(n1332), .B(n1331), .Z(n1345) );
  IV U4430 ( .A(n1337), .Z(n1391) );
  XNOR U4431 ( .A(n1391), .B(n1333), .Z(n1398) );
  AND U4432 ( .A(n1387), .B(n1398), .Z(n1335) );
  AND U4433 ( .A(x[56]), .B(n1402), .Z(n1334) );
  XNOR U4434 ( .A(n1335), .B(n1334), .Z(n1336) );
  NANDN U4435 ( .A(n1388), .B(n1336), .Z(n1340) );
  NAND U4436 ( .A(x[56]), .B(n1387), .Z(n1338) );
  OR U4437 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U4438 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4439 ( .A(n1342), .B(n1341), .Z(n1343) );
  XNOR U4440 ( .A(n1345), .B(n1343), .Z(n1365) );
  IV U4441 ( .A(n1365), .Z(n1372) );
  AND U4442 ( .A(n1418), .B(n1344), .Z(n1347) );
  XOR U4443 ( .A(x[57]), .B(x[63]), .Z(n1420) );
  AND U4444 ( .A(n1381), .B(n1420), .Z(n1350) );
  XNOR U4445 ( .A(n1350), .B(n1345), .Z(n1346) );
  XNOR U4446 ( .A(n1347), .B(n1346), .Z(n1371) );
  NANDN U4447 ( .A(n1372), .B(n1371), .Z(n1348) );
  NAND U4448 ( .A(n1376), .B(n1348), .Z(n1358) );
  XNOR U4449 ( .A(n1350), .B(n1349), .Z(n1355) );
  ANDN U4450 ( .B(n1351), .A(x[57]), .Z(n1352) );
  XNOR U4451 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U4452 ( .A(n1355), .B(n1354), .Z(n1368) );
  XOR U4453 ( .A(n1371), .B(n1368), .Z(n1356) );
  NAND U4454 ( .A(n1372), .B(n1356), .Z(n1357) );
  NAND U4455 ( .A(n1358), .B(n1357), .Z(n1417) );
  ANDN U4456 ( .B(n1359), .A(n1417), .Z(n1383) );
  IV U4457 ( .A(n1368), .Z(n1374) );
  XOR U4458 ( .A(n1376), .B(n1372), .Z(n1360) );
  NANDN U4459 ( .A(n1374), .B(n1360), .Z(n1363) );
  NANDN U4460 ( .A(n1372), .B(n1374), .Z(n1361) );
  NANDN U4461 ( .A(n1371), .B(n1361), .Z(n1362) );
  NAND U4462 ( .A(n1363), .B(n1362), .Z(n1442) );
  XNOR U4463 ( .A(n1417), .B(n1442), .Z(n1393) );
  AND U4464 ( .A(n1364), .B(n1393), .Z(n1386) );
  OR U4465 ( .A(n1371), .B(n1368), .Z(n1370) );
  ANDN U4466 ( .B(n1371), .A(n1365), .Z(n1366) );
  XNOR U4467 ( .A(n1366), .B(n1376), .Z(n1367) );
  NAND U4468 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U4469 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U4470 ( .A(n1372), .B(n1376), .Z(n1378) );
  NAND U4471 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4472 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U4473 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U4474 ( .A(n1378), .B(n1377), .Z(n1449) );
  NAND U4475 ( .A(n1409), .B(n1379), .Z(n1380) );
  XNOR U4476 ( .A(n1386), .B(n1380), .Z(n1444) );
  XOR U4477 ( .A(n1417), .B(n1449), .Z(n1419) );
  AND U4478 ( .A(n1381), .B(n1419), .Z(n1404) );
  XNOR U4479 ( .A(n1444), .B(n1404), .Z(n1382) );
  XNOR U4480 ( .A(n1383), .B(n1382), .Z(n1452) );
  NAND U4481 ( .A(n1395), .B(n1384), .Z(n1385) );
  XNOR U4482 ( .A(n1386), .B(n1385), .Z(n1412) );
  AND U4483 ( .A(n1387), .B(n1397), .Z(n1443) );
  NANDN U4484 ( .A(n1388), .B(n1390), .Z(n1389) );
  XNOR U4485 ( .A(n1443), .B(n1389), .Z(n1416) );
  XNOR U4486 ( .A(n1412), .B(n1416), .Z(n1401) );
  XOR U4487 ( .A(n1452), .B(n1401), .Z(z[56]) );
  AND U4488 ( .A(n1391), .B(n1390), .Z(n1400) );
  AND U4489 ( .A(n1393), .B(n1392), .Z(n1411) );
  NAND U4490 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U4491 ( .A(n1411), .B(n1396), .Z(n1453) );
  AND U4492 ( .A(n1398), .B(n1397), .Z(n1405) );
  XNOR U4493 ( .A(n1453), .B(n1405), .Z(n1399) );
  XNOR U4494 ( .A(n1400), .B(n1399), .Z(n1425) );
  XNOR U4495 ( .A(n1425), .B(n1401), .Z(n1458) );
  AND U4496 ( .A(n1402), .B(n1442), .Z(n1407) );
  NANDN U4497 ( .A(n1449), .B(n1447), .Z(n1403) );
  XNOR U4498 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U4499 ( .A(n1405), .B(n1415), .Z(n1406) );
  XNOR U4500 ( .A(n1407), .B(n1406), .Z(n1414) );
  NAND U4501 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U4502 ( .A(n1411), .B(n1410), .Z(n1421) );
  XNOR U4503 ( .A(n1412), .B(n1421), .Z(n1413) );
  XNOR U4504 ( .A(n1414), .B(n1413), .Z(n1424) );
  XNOR U4505 ( .A(n1458), .B(n1424), .Z(z[57]) );
  XNOR U4506 ( .A(n1416), .B(n1415), .Z(z[58]) );
  NOR U4507 ( .A(n1418), .B(n1417), .Z(n1423) );
  AND U4508 ( .A(n1420), .B(n1419), .Z(n1451) );
  XNOR U4509 ( .A(n1421), .B(n1451), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1457) );
  XOR U4511 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U4512 ( .A(n1457), .B(n1426), .Z(z[59]) );
  AND U4513 ( .A(x[0]), .B(n1427), .Z(n1431) );
  XNOR U4514 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U4515 ( .A(n1431), .B(n1430), .Z(n1708) );
  XOR U4516 ( .A(n1432), .B(x[1]), .Z(n1433) );
  NANDN U4517 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U4518 ( .A(n1436), .B(n1435), .Z(n1440) );
  XNOR U4519 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U4520 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U4521 ( .A(n1708), .B(n1441), .Z(z[5]) );
  XOR U4522 ( .A(n1452), .B(z[58]), .Z(z[60]) );
  AND U4523 ( .A(x[56]), .B(n1442), .Z(n1446) );
  XNOR U4524 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U4525 ( .A(n1446), .B(n1445), .Z(n1459) );
  XOR U4526 ( .A(n1447), .B(x[57]), .Z(n1448) );
  NANDN U4527 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U4528 ( .A(n1451), .B(n1450), .Z(n1455) );
  XNOR U4529 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U4530 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U4531 ( .A(n1459), .B(n1456), .Z(z[61]) );
  XNOR U4532 ( .A(n1458), .B(n1457), .Z(z[62]) );
  XOR U4533 ( .A(n1459), .B(z[57]), .Z(z[63]) );
  XOR U4534 ( .A(x[67]), .B(x[65]), .Z(n1462) );
  XNOR U4535 ( .A(x[64]), .B(x[70]), .Z(n1461) );
  XOR U4536 ( .A(n1461), .B(x[66]), .Z(n1460) );
  XNOR U4537 ( .A(n1462), .B(n1460), .Z(n1497) );
  XNOR U4538 ( .A(x[69]), .B(n1461), .Z(n1570) );
  XOR U4539 ( .A(n1570), .B(x[68]), .Z(n1540) );
  IV U4540 ( .A(n1540), .Z(n1471) );
  XNOR U4541 ( .A(x[71]), .B(x[68]), .Z(n1465) );
  XNOR U4542 ( .A(n1462), .B(n1465), .Z(n1525) );
  NOR U4543 ( .A(n1471), .B(n1525), .Z(n1464) );
  XNOR U4544 ( .A(n1570), .B(x[71]), .Z(n1556) );
  XNOR U4545 ( .A(x[66]), .B(n1556), .Z(n1480) );
  XNOR U4546 ( .A(x[65]), .B(n1480), .Z(n1475) );
  AND U4547 ( .A(x[64]), .B(n1475), .Z(n1463) );
  XNOR U4548 ( .A(n1464), .B(n1463), .Z(n1468) );
  XNOR U4549 ( .A(n1497), .B(n1556), .Z(n1487) );
  IV U4550 ( .A(n1497), .Z(n1482) );
  XNOR U4551 ( .A(x[64]), .B(n1482), .Z(n1502) );
  IV U4552 ( .A(n1465), .Z(n1530) );
  AND U4553 ( .A(n1502), .B(n1530), .Z(n1470) );
  IV U4554 ( .A(n1570), .Z(n1489) );
  XNOR U4555 ( .A(n1497), .B(n1489), .Z(n1519) );
  XOR U4556 ( .A(n1519), .B(n1525), .Z(n1522) );
  XOR U4557 ( .A(x[66]), .B(x[68]), .Z(n1532) );
  NAND U4558 ( .A(n1522), .B(n1532), .Z(n1466) );
  XNOR U4559 ( .A(n1470), .B(n1466), .Z(n1491) );
  XNOR U4560 ( .A(n1487), .B(n1491), .Z(n1467) );
  XNOR U4561 ( .A(n1468), .B(n1467), .Z(n1514) );
  XOR U4562 ( .A(x[66]), .B(x[71]), .Z(n1546) );
  XNOR U4563 ( .A(x[64]), .B(n1525), .Z(n1526) );
  XNOR U4564 ( .A(n1570), .B(n1526), .Z(n1517) );
  NAND U4565 ( .A(n1546), .B(n1517), .Z(n1469) );
  XNOR U4566 ( .A(n1470), .B(n1469), .Z(n1483) );
  IV U4567 ( .A(n1475), .Z(n1529) );
  XNOR U4568 ( .A(n1529), .B(n1471), .Z(n1536) );
  AND U4569 ( .A(n1525), .B(n1536), .Z(n1473) );
  AND U4570 ( .A(x[64]), .B(n1540), .Z(n1472) );
  XNOR U4571 ( .A(n1473), .B(n1472), .Z(n1474) );
  NANDN U4572 ( .A(n1526), .B(n1474), .Z(n1478) );
  NAND U4573 ( .A(x[64]), .B(n1525), .Z(n1476) );
  OR U4574 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U4575 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4576 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR U4577 ( .A(n1483), .B(n1481), .Z(n1503) );
  IV U4578 ( .A(n1503), .Z(n1510) );
  AND U4579 ( .A(n1556), .B(n1482), .Z(n1485) );
  XOR U4580 ( .A(x[65]), .B(x[71]), .Z(n1558) );
  AND U4581 ( .A(n1519), .B(n1558), .Z(n1488) );
  XNOR U4582 ( .A(n1488), .B(n1483), .Z(n1484) );
  XNOR U4583 ( .A(n1485), .B(n1484), .Z(n1509) );
  NANDN U4584 ( .A(n1510), .B(n1509), .Z(n1486) );
  NAND U4585 ( .A(n1514), .B(n1486), .Z(n1496) );
  XNOR U4586 ( .A(n1488), .B(n1487), .Z(n1493) );
  ANDN U4587 ( .B(n1489), .A(x[65]), .Z(n1490) );
  XNOR U4588 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U4589 ( .A(n1493), .B(n1492), .Z(n1506) );
  XOR U4590 ( .A(n1509), .B(n1506), .Z(n1494) );
  NAND U4591 ( .A(n1510), .B(n1494), .Z(n1495) );
  NAND U4592 ( .A(n1496), .B(n1495), .Z(n1555) );
  ANDN U4593 ( .B(n1497), .A(n1555), .Z(n1521) );
  IV U4594 ( .A(n1506), .Z(n1512) );
  XOR U4595 ( .A(n1514), .B(n1510), .Z(n1498) );
  NANDN U4596 ( .A(n1512), .B(n1498), .Z(n1501) );
  NANDN U4597 ( .A(n1510), .B(n1512), .Z(n1499) );
  NANDN U4598 ( .A(n1509), .B(n1499), .Z(n1500) );
  NAND U4599 ( .A(n1501), .B(n1500), .Z(n1565) );
  XNOR U4600 ( .A(n1555), .B(n1565), .Z(n1531) );
  AND U4601 ( .A(n1502), .B(n1531), .Z(n1524) );
  OR U4602 ( .A(n1509), .B(n1506), .Z(n1508) );
  ANDN U4603 ( .B(n1509), .A(n1503), .Z(n1504) );
  XNOR U4604 ( .A(n1504), .B(n1514), .Z(n1505) );
  NAND U4605 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U4606 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U4607 ( .A(n1510), .B(n1514), .Z(n1516) );
  NAND U4608 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4609 ( .A(n1512), .B(n1511), .Z(n1513) );
  NANDN U4610 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U4611 ( .A(n1516), .B(n1515), .Z(n1572) );
  NAND U4612 ( .A(n1547), .B(n1517), .Z(n1518) );
  XNOR U4613 ( .A(n1524), .B(n1518), .Z(n1567) );
  XOR U4614 ( .A(n1555), .B(n1572), .Z(n1557) );
  AND U4615 ( .A(n1519), .B(n1557), .Z(n1542) );
  XNOR U4616 ( .A(n1567), .B(n1542), .Z(n1520) );
  XNOR U4617 ( .A(n1521), .B(n1520), .Z(n1575) );
  NAND U4618 ( .A(n1533), .B(n1522), .Z(n1523) );
  XNOR U4619 ( .A(n1524), .B(n1523), .Z(n1550) );
  AND U4620 ( .A(n1525), .B(n1535), .Z(n1566) );
  NANDN U4621 ( .A(n1526), .B(n1528), .Z(n1527) );
  XNOR U4622 ( .A(n1566), .B(n1527), .Z(n1554) );
  XNOR U4623 ( .A(n1550), .B(n1554), .Z(n1539) );
  XOR U4624 ( .A(n1575), .B(n1539), .Z(z[64]) );
  AND U4625 ( .A(n1529), .B(n1528), .Z(n1538) );
  AND U4626 ( .A(n1531), .B(n1530), .Z(n1549) );
  NAND U4627 ( .A(n1533), .B(n1532), .Z(n1534) );
  XNOR U4628 ( .A(n1549), .B(n1534), .Z(n1576) );
  AND U4629 ( .A(n1536), .B(n1535), .Z(n1543) );
  XNOR U4630 ( .A(n1576), .B(n1543), .Z(n1537) );
  XNOR U4631 ( .A(n1538), .B(n1537), .Z(n1563) );
  XNOR U4632 ( .A(n1563), .B(n1539), .Z(n1583) );
  AND U4633 ( .A(n1540), .B(n1565), .Z(n1545) );
  NANDN U4634 ( .A(n1572), .B(n1570), .Z(n1541) );
  XNOR U4635 ( .A(n1542), .B(n1541), .Z(n1553) );
  XNOR U4636 ( .A(n1543), .B(n1553), .Z(n1544) );
  XNOR U4637 ( .A(n1545), .B(n1544), .Z(n1552) );
  NAND U4638 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U4639 ( .A(n1549), .B(n1548), .Z(n1559) );
  XNOR U4640 ( .A(n1550), .B(n1559), .Z(n1551) );
  XNOR U4641 ( .A(n1552), .B(n1551), .Z(n1562) );
  XNOR U4642 ( .A(n1583), .B(n1562), .Z(z[65]) );
  XNOR U4643 ( .A(n1554), .B(n1553), .Z(z[66]) );
  NOR U4644 ( .A(n1556), .B(n1555), .Z(n1561) );
  AND U4645 ( .A(n1558), .B(n1557), .Z(n1574) );
  XNOR U4646 ( .A(n1559), .B(n1574), .Z(n1560) );
  XNOR U4647 ( .A(n1561), .B(n1560), .Z(n1582) );
  XOR U4648 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U4649 ( .A(n1582), .B(n1564), .Z(z[67]) );
  XOR U4650 ( .A(n1575), .B(z[66]), .Z(z[68]) );
  AND U4651 ( .A(x[64]), .B(n1565), .Z(n1569) );
  XNOR U4652 ( .A(n1567), .B(n1566), .Z(n1568) );
  XNOR U4653 ( .A(n1569), .B(n1568), .Z(n1584) );
  XOR U4654 ( .A(n1570), .B(x[65]), .Z(n1571) );
  NANDN U4655 ( .A(n1572), .B(n1571), .Z(n1573) );
  XNOR U4656 ( .A(n1574), .B(n1573), .Z(n1578) );
  XNOR U4657 ( .A(n1576), .B(n1575), .Z(n1577) );
  XNOR U4658 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U4659 ( .A(n1584), .B(n1579), .Z(z[69]) );
  XNOR U4660 ( .A(n1581), .B(n1580), .Z(z[6]) );
  XNOR U4661 ( .A(n1583), .B(n1582), .Z(z[70]) );
  XOR U4662 ( .A(n1584), .B(z[65]), .Z(z[71]) );
  XOR U4663 ( .A(x[75]), .B(x[73]), .Z(n1587) );
  XNOR U4664 ( .A(x[72]), .B(x[78]), .Z(n1586) );
  XOR U4665 ( .A(n1586), .B(x[74]), .Z(n1585) );
  XNOR U4666 ( .A(n1587), .B(n1585), .Z(n1622) );
  XNOR U4667 ( .A(x[77]), .B(n1586), .Z(n1695) );
  XOR U4668 ( .A(n1695), .B(x[76]), .Z(n1665) );
  IV U4669 ( .A(n1665), .Z(n1596) );
  XNOR U4670 ( .A(x[79]), .B(x[76]), .Z(n1590) );
  XNOR U4671 ( .A(n1587), .B(n1590), .Z(n1650) );
  NOR U4672 ( .A(n1596), .B(n1650), .Z(n1589) );
  XNOR U4673 ( .A(n1695), .B(x[79]), .Z(n1681) );
  XNOR U4674 ( .A(x[74]), .B(n1681), .Z(n1605) );
  XNOR U4675 ( .A(x[73]), .B(n1605), .Z(n1600) );
  AND U4676 ( .A(x[72]), .B(n1600), .Z(n1588) );
  XNOR U4677 ( .A(n1589), .B(n1588), .Z(n1593) );
  XNOR U4678 ( .A(n1622), .B(n1681), .Z(n1612) );
  IV U4679 ( .A(n1622), .Z(n1607) );
  XNOR U4680 ( .A(x[72]), .B(n1607), .Z(n1627) );
  IV U4681 ( .A(n1590), .Z(n1655) );
  AND U4682 ( .A(n1627), .B(n1655), .Z(n1595) );
  IV U4683 ( .A(n1695), .Z(n1614) );
  XNOR U4684 ( .A(n1622), .B(n1614), .Z(n1644) );
  XOR U4685 ( .A(n1644), .B(n1650), .Z(n1647) );
  XOR U4686 ( .A(x[74]), .B(x[76]), .Z(n1657) );
  NAND U4687 ( .A(n1647), .B(n1657), .Z(n1591) );
  XNOR U4688 ( .A(n1595), .B(n1591), .Z(n1616) );
  XNOR U4689 ( .A(n1612), .B(n1616), .Z(n1592) );
  XNOR U4690 ( .A(n1593), .B(n1592), .Z(n1639) );
  XOR U4691 ( .A(x[74]), .B(x[79]), .Z(n1671) );
  XNOR U4692 ( .A(x[72]), .B(n1650), .Z(n1651) );
  XNOR U4693 ( .A(n1695), .B(n1651), .Z(n1642) );
  NAND U4694 ( .A(n1671), .B(n1642), .Z(n1594) );
  XNOR U4695 ( .A(n1595), .B(n1594), .Z(n1608) );
  IV U4696 ( .A(n1600), .Z(n1654) );
  XNOR U4697 ( .A(n1654), .B(n1596), .Z(n1661) );
  AND U4698 ( .A(n1650), .B(n1661), .Z(n1598) );
  AND U4699 ( .A(x[72]), .B(n1665), .Z(n1597) );
  XNOR U4700 ( .A(n1598), .B(n1597), .Z(n1599) );
  NANDN U4701 ( .A(n1651), .B(n1599), .Z(n1603) );
  NAND U4702 ( .A(x[72]), .B(n1650), .Z(n1601) );
  OR U4703 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U4704 ( .A(n1603), .B(n1602), .Z(n1604) );
  XNOR U4705 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U4706 ( .A(n1608), .B(n1606), .Z(n1628) );
  IV U4707 ( .A(n1628), .Z(n1635) );
  AND U4708 ( .A(n1681), .B(n1607), .Z(n1610) );
  XOR U4709 ( .A(x[73]), .B(x[79]), .Z(n1683) );
  AND U4710 ( .A(n1644), .B(n1683), .Z(n1613) );
  XNOR U4711 ( .A(n1613), .B(n1608), .Z(n1609) );
  XNOR U4712 ( .A(n1610), .B(n1609), .Z(n1634) );
  NANDN U4713 ( .A(n1635), .B(n1634), .Z(n1611) );
  NAND U4714 ( .A(n1639), .B(n1611), .Z(n1621) );
  XNOR U4715 ( .A(n1613), .B(n1612), .Z(n1618) );
  ANDN U4716 ( .B(n1614), .A(x[73]), .Z(n1615) );
  XNOR U4717 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4718 ( .A(n1618), .B(n1617), .Z(n1631) );
  XOR U4719 ( .A(n1634), .B(n1631), .Z(n1619) );
  NAND U4720 ( .A(n1635), .B(n1619), .Z(n1620) );
  NAND U4721 ( .A(n1621), .B(n1620), .Z(n1680) );
  ANDN U4722 ( .B(n1622), .A(n1680), .Z(n1646) );
  IV U4723 ( .A(n1631), .Z(n1637) );
  XOR U4724 ( .A(n1639), .B(n1635), .Z(n1623) );
  NANDN U4725 ( .A(n1637), .B(n1623), .Z(n1626) );
  NANDN U4726 ( .A(n1635), .B(n1637), .Z(n1624) );
  NANDN U4727 ( .A(n1634), .B(n1624), .Z(n1625) );
  NAND U4728 ( .A(n1626), .B(n1625), .Z(n1690) );
  XNOR U4729 ( .A(n1680), .B(n1690), .Z(n1656) );
  AND U4730 ( .A(n1627), .B(n1656), .Z(n1649) );
  OR U4731 ( .A(n1634), .B(n1631), .Z(n1633) );
  ANDN U4732 ( .B(n1634), .A(n1628), .Z(n1629) );
  XNOR U4733 ( .A(n1629), .B(n1639), .Z(n1630) );
  NAND U4734 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U4735 ( .A(n1633), .B(n1632), .Z(n1653) );
  NAND U4736 ( .A(n1635), .B(n1639), .Z(n1641) );
  NAND U4737 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U4738 ( .A(n1637), .B(n1636), .Z(n1638) );
  NANDN U4739 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U4740 ( .A(n1641), .B(n1640), .Z(n1697) );
  NAND U4741 ( .A(n1672), .B(n1642), .Z(n1643) );
  XNOR U4742 ( .A(n1649), .B(n1643), .Z(n1692) );
  XOR U4743 ( .A(n1680), .B(n1697), .Z(n1682) );
  AND U4744 ( .A(n1644), .B(n1682), .Z(n1667) );
  XNOR U4745 ( .A(n1692), .B(n1667), .Z(n1645) );
  XNOR U4746 ( .A(n1646), .B(n1645), .Z(n1700) );
  NAND U4747 ( .A(n1658), .B(n1647), .Z(n1648) );
  XNOR U4748 ( .A(n1649), .B(n1648), .Z(n1675) );
  AND U4749 ( .A(n1650), .B(n1660), .Z(n1691) );
  NANDN U4750 ( .A(n1651), .B(n1653), .Z(n1652) );
  XNOR U4751 ( .A(n1691), .B(n1652), .Z(n1679) );
  XNOR U4752 ( .A(n1675), .B(n1679), .Z(n1664) );
  XOR U4753 ( .A(n1700), .B(n1664), .Z(z[72]) );
  AND U4754 ( .A(n1654), .B(n1653), .Z(n1663) );
  AND U4755 ( .A(n1656), .B(n1655), .Z(n1674) );
  NAND U4756 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U4757 ( .A(n1674), .B(n1659), .Z(n1701) );
  AND U4758 ( .A(n1661), .B(n1660), .Z(n1668) );
  XNOR U4759 ( .A(n1701), .B(n1668), .Z(n1662) );
  XNOR U4760 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U4761 ( .A(n1688), .B(n1664), .Z(n1706) );
  AND U4762 ( .A(n1665), .B(n1690), .Z(n1670) );
  NANDN U4763 ( .A(n1697), .B(n1695), .Z(n1666) );
  XNOR U4764 ( .A(n1667), .B(n1666), .Z(n1678) );
  XNOR U4765 ( .A(n1668), .B(n1678), .Z(n1669) );
  XNOR U4766 ( .A(n1670), .B(n1669), .Z(n1677) );
  NAND U4767 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR U4768 ( .A(n1674), .B(n1673), .Z(n1684) );
  XNOR U4769 ( .A(n1675), .B(n1684), .Z(n1676) );
  XNOR U4770 ( .A(n1677), .B(n1676), .Z(n1687) );
  XNOR U4771 ( .A(n1706), .B(n1687), .Z(z[73]) );
  XNOR U4772 ( .A(n1679), .B(n1678), .Z(z[74]) );
  NOR U4773 ( .A(n1681), .B(n1680), .Z(n1686) );
  AND U4774 ( .A(n1683), .B(n1682), .Z(n1699) );
  XNOR U4775 ( .A(n1684), .B(n1699), .Z(n1685) );
  XNOR U4776 ( .A(n1686), .B(n1685), .Z(n1705) );
  XOR U4777 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4778 ( .A(n1705), .B(n1689), .Z(z[75]) );
  XOR U4779 ( .A(n1700), .B(z[74]), .Z(z[76]) );
  AND U4780 ( .A(x[72]), .B(n1690), .Z(n1694) );
  XNOR U4781 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4782 ( .A(n1694), .B(n1693), .Z(n1707) );
  XOR U4783 ( .A(n1695), .B(x[73]), .Z(n1696) );
  NANDN U4784 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U4785 ( .A(n1699), .B(n1698), .Z(n1703) );
  XNOR U4786 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U4787 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U4788 ( .A(n1707), .B(n1704), .Z(z[77]) );
  XNOR U4789 ( .A(n1706), .B(n1705), .Z(z[78]) );
  XOR U4790 ( .A(n1707), .B(z[73]), .Z(z[79]) );
  XOR U4791 ( .A(n1708), .B(z[1]), .Z(z[7]) );
  XOR U4792 ( .A(x[83]), .B(x[81]), .Z(n1711) );
  XNOR U4793 ( .A(x[80]), .B(x[86]), .Z(n1710) );
  XOR U4794 ( .A(n1710), .B(x[82]), .Z(n1709) );
  XNOR U4795 ( .A(n1711), .B(n1709), .Z(n1746) );
  XNOR U4796 ( .A(x[85]), .B(n1710), .Z(n1819) );
  XOR U4797 ( .A(n1819), .B(x[84]), .Z(n1789) );
  IV U4798 ( .A(n1789), .Z(n1720) );
  XNOR U4799 ( .A(x[87]), .B(x[84]), .Z(n1714) );
  XNOR U4800 ( .A(n1711), .B(n1714), .Z(n1774) );
  NOR U4801 ( .A(n1720), .B(n1774), .Z(n1713) );
  XNOR U4802 ( .A(n1819), .B(x[87]), .Z(n1805) );
  XNOR U4803 ( .A(x[82]), .B(n1805), .Z(n1729) );
  XNOR U4804 ( .A(x[81]), .B(n1729), .Z(n1724) );
  AND U4805 ( .A(x[80]), .B(n1724), .Z(n1712) );
  XNOR U4806 ( .A(n1713), .B(n1712), .Z(n1717) );
  XNOR U4807 ( .A(n1746), .B(n1805), .Z(n1736) );
  IV U4808 ( .A(n1746), .Z(n1731) );
  XNOR U4809 ( .A(x[80]), .B(n1731), .Z(n1751) );
  IV U4810 ( .A(n1714), .Z(n1779) );
  AND U4811 ( .A(n1751), .B(n1779), .Z(n1719) );
  IV U4812 ( .A(n1819), .Z(n1738) );
  XNOR U4813 ( .A(n1746), .B(n1738), .Z(n1768) );
  XOR U4814 ( .A(n1768), .B(n1774), .Z(n1771) );
  XOR U4815 ( .A(x[82]), .B(x[84]), .Z(n1781) );
  NAND U4816 ( .A(n1771), .B(n1781), .Z(n1715) );
  XNOR U4817 ( .A(n1719), .B(n1715), .Z(n1740) );
  XNOR U4818 ( .A(n1736), .B(n1740), .Z(n1716) );
  XNOR U4819 ( .A(n1717), .B(n1716), .Z(n1763) );
  XOR U4820 ( .A(x[82]), .B(x[87]), .Z(n1795) );
  XNOR U4821 ( .A(x[80]), .B(n1774), .Z(n1775) );
  XNOR U4822 ( .A(n1819), .B(n1775), .Z(n1766) );
  NAND U4823 ( .A(n1795), .B(n1766), .Z(n1718) );
  XNOR U4824 ( .A(n1719), .B(n1718), .Z(n1732) );
  IV U4825 ( .A(n1724), .Z(n1778) );
  XNOR U4826 ( .A(n1778), .B(n1720), .Z(n1785) );
  AND U4827 ( .A(n1774), .B(n1785), .Z(n1722) );
  AND U4828 ( .A(x[80]), .B(n1789), .Z(n1721) );
  XNOR U4829 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U4830 ( .A(n1775), .B(n1723), .Z(n1727) );
  NAND U4831 ( .A(x[80]), .B(n1774), .Z(n1725) );
  OR U4832 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U4833 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U4834 ( .A(n1729), .B(n1728), .Z(n1730) );
  XNOR U4835 ( .A(n1732), .B(n1730), .Z(n1752) );
  IV U4836 ( .A(n1752), .Z(n1759) );
  AND U4837 ( .A(n1805), .B(n1731), .Z(n1734) );
  XOR U4838 ( .A(x[81]), .B(x[87]), .Z(n1807) );
  AND U4839 ( .A(n1768), .B(n1807), .Z(n1737) );
  XNOR U4840 ( .A(n1737), .B(n1732), .Z(n1733) );
  XNOR U4841 ( .A(n1734), .B(n1733), .Z(n1758) );
  NANDN U4842 ( .A(n1759), .B(n1758), .Z(n1735) );
  NAND U4843 ( .A(n1763), .B(n1735), .Z(n1745) );
  XNOR U4844 ( .A(n1737), .B(n1736), .Z(n1742) );
  ANDN U4845 ( .B(n1738), .A(x[81]), .Z(n1739) );
  XNOR U4846 ( .A(n1740), .B(n1739), .Z(n1741) );
  XNOR U4847 ( .A(n1742), .B(n1741), .Z(n1755) );
  XOR U4848 ( .A(n1758), .B(n1755), .Z(n1743) );
  NAND U4849 ( .A(n1759), .B(n1743), .Z(n1744) );
  NAND U4850 ( .A(n1745), .B(n1744), .Z(n1804) );
  ANDN U4851 ( .B(n1746), .A(n1804), .Z(n1770) );
  IV U4852 ( .A(n1755), .Z(n1761) );
  XOR U4853 ( .A(n1763), .B(n1759), .Z(n1747) );
  NANDN U4854 ( .A(n1761), .B(n1747), .Z(n1750) );
  NANDN U4855 ( .A(n1759), .B(n1761), .Z(n1748) );
  NANDN U4856 ( .A(n1758), .B(n1748), .Z(n1749) );
  NAND U4857 ( .A(n1750), .B(n1749), .Z(n1814) );
  XNOR U4858 ( .A(n1804), .B(n1814), .Z(n1780) );
  AND U4859 ( .A(n1751), .B(n1780), .Z(n1773) );
  OR U4860 ( .A(n1758), .B(n1755), .Z(n1757) );
  ANDN U4861 ( .B(n1758), .A(n1752), .Z(n1753) );
  XNOR U4862 ( .A(n1753), .B(n1763), .Z(n1754) );
  NAND U4863 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U4864 ( .A(n1757), .B(n1756), .Z(n1777) );
  NAND U4865 ( .A(n1759), .B(n1763), .Z(n1765) );
  NAND U4866 ( .A(n1759), .B(n1758), .Z(n1760) );
  XNOR U4867 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U4868 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1821) );
  NAND U4870 ( .A(n1796), .B(n1766), .Z(n1767) );
  XNOR U4871 ( .A(n1773), .B(n1767), .Z(n1816) );
  XOR U4872 ( .A(n1804), .B(n1821), .Z(n1806) );
  AND U4873 ( .A(n1768), .B(n1806), .Z(n1791) );
  XNOR U4874 ( .A(n1816), .B(n1791), .Z(n1769) );
  XNOR U4875 ( .A(n1770), .B(n1769), .Z(n1824) );
  NAND U4876 ( .A(n1782), .B(n1771), .Z(n1772) );
  XNOR U4877 ( .A(n1773), .B(n1772), .Z(n1799) );
  AND U4878 ( .A(n1774), .B(n1784), .Z(n1815) );
  NANDN U4879 ( .A(n1775), .B(n1777), .Z(n1776) );
  XNOR U4880 ( .A(n1815), .B(n1776), .Z(n1803) );
  XNOR U4881 ( .A(n1799), .B(n1803), .Z(n1788) );
  XOR U4882 ( .A(n1824), .B(n1788), .Z(z[80]) );
  AND U4883 ( .A(n1778), .B(n1777), .Z(n1787) );
  AND U4884 ( .A(n1780), .B(n1779), .Z(n1798) );
  NAND U4885 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U4886 ( .A(n1798), .B(n1783), .Z(n1825) );
  AND U4887 ( .A(n1785), .B(n1784), .Z(n1792) );
  XNOR U4888 ( .A(n1825), .B(n1792), .Z(n1786) );
  XNOR U4889 ( .A(n1787), .B(n1786), .Z(n1812) );
  XNOR U4890 ( .A(n1812), .B(n1788), .Z(n1830) );
  AND U4891 ( .A(n1789), .B(n1814), .Z(n1794) );
  NANDN U4892 ( .A(n1821), .B(n1819), .Z(n1790) );
  XNOR U4893 ( .A(n1791), .B(n1790), .Z(n1802) );
  XNOR U4894 ( .A(n1792), .B(n1802), .Z(n1793) );
  XNOR U4895 ( .A(n1794), .B(n1793), .Z(n1801) );
  NAND U4896 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U4897 ( .A(n1798), .B(n1797), .Z(n1808) );
  XNOR U4898 ( .A(n1799), .B(n1808), .Z(n1800) );
  XNOR U4899 ( .A(n1801), .B(n1800), .Z(n1811) );
  XNOR U4900 ( .A(n1830), .B(n1811), .Z(z[81]) );
  XNOR U4901 ( .A(n1803), .B(n1802), .Z(z[82]) );
  NOR U4902 ( .A(n1805), .B(n1804), .Z(n1810) );
  AND U4903 ( .A(n1807), .B(n1806), .Z(n1823) );
  XNOR U4904 ( .A(n1808), .B(n1823), .Z(n1809) );
  XNOR U4905 ( .A(n1810), .B(n1809), .Z(n1829) );
  XOR U4906 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U4907 ( .A(n1829), .B(n1813), .Z(z[83]) );
  XOR U4908 ( .A(n1824), .B(z[82]), .Z(z[84]) );
  AND U4909 ( .A(x[80]), .B(n1814), .Z(n1818) );
  XNOR U4910 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U4911 ( .A(n1818), .B(n1817), .Z(n1831) );
  XOR U4912 ( .A(n1819), .B(x[81]), .Z(n1820) );
  NANDN U4913 ( .A(n1821), .B(n1820), .Z(n1822) );
  XNOR U4914 ( .A(n1823), .B(n1822), .Z(n1827) );
  XNOR U4915 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U4916 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U4917 ( .A(n1831), .B(n1828), .Z(z[85]) );
  XNOR U4918 ( .A(n1830), .B(n1829), .Z(z[86]) );
  XOR U4919 ( .A(n1831), .B(z[81]), .Z(z[87]) );
  XOR U4920 ( .A(x[91]), .B(x[89]), .Z(n1834) );
  XNOR U4921 ( .A(x[88]), .B(x[94]), .Z(n1833) );
  XOR U4922 ( .A(n1833), .B(x[90]), .Z(n1832) );
  XNOR U4923 ( .A(n1834), .B(n1832), .Z(n1869) );
  XNOR U4924 ( .A(x[93]), .B(n1833), .Z(n1944) );
  XOR U4925 ( .A(n1944), .B(x[92]), .Z(n1912) );
  IV U4926 ( .A(n1912), .Z(n1843) );
  XNOR U4927 ( .A(x[95]), .B(x[92]), .Z(n1837) );
  XNOR U4928 ( .A(n1834), .B(n1837), .Z(n1897) );
  NOR U4929 ( .A(n1843), .B(n1897), .Z(n1836) );
  XNOR U4930 ( .A(n1944), .B(x[95]), .Z(n1930) );
  XNOR U4931 ( .A(x[90]), .B(n1930), .Z(n1852) );
  XNOR U4932 ( .A(x[89]), .B(n1852), .Z(n1847) );
  AND U4933 ( .A(x[88]), .B(n1847), .Z(n1835) );
  XNOR U4934 ( .A(n1836), .B(n1835), .Z(n1840) );
  XNOR U4935 ( .A(n1869), .B(n1930), .Z(n1859) );
  IV U4936 ( .A(n1869), .Z(n1854) );
  XNOR U4937 ( .A(x[88]), .B(n1854), .Z(n1874) );
  IV U4938 ( .A(n1837), .Z(n1902) );
  AND U4939 ( .A(n1874), .B(n1902), .Z(n1842) );
  IV U4940 ( .A(n1944), .Z(n1861) );
  XNOR U4941 ( .A(n1869), .B(n1861), .Z(n1891) );
  XOR U4942 ( .A(n1891), .B(n1897), .Z(n1894) );
  XOR U4943 ( .A(x[90]), .B(x[92]), .Z(n1904) );
  NAND U4944 ( .A(n1894), .B(n1904), .Z(n1838) );
  XNOR U4945 ( .A(n1842), .B(n1838), .Z(n1863) );
  XNOR U4946 ( .A(n1859), .B(n1863), .Z(n1839) );
  XNOR U4947 ( .A(n1840), .B(n1839), .Z(n1886) );
  XOR U4948 ( .A(x[90]), .B(x[95]), .Z(n1918) );
  XNOR U4949 ( .A(x[88]), .B(n1897), .Z(n1898) );
  XNOR U4950 ( .A(n1944), .B(n1898), .Z(n1889) );
  NAND U4951 ( .A(n1918), .B(n1889), .Z(n1841) );
  XNOR U4952 ( .A(n1842), .B(n1841), .Z(n1855) );
  IV U4953 ( .A(n1847), .Z(n1901) );
  XNOR U4954 ( .A(n1901), .B(n1843), .Z(n1908) );
  AND U4955 ( .A(n1897), .B(n1908), .Z(n1845) );
  AND U4956 ( .A(x[88]), .B(n1912), .Z(n1844) );
  XNOR U4957 ( .A(n1845), .B(n1844), .Z(n1846) );
  NANDN U4958 ( .A(n1898), .B(n1846), .Z(n1850) );
  NAND U4959 ( .A(x[88]), .B(n1897), .Z(n1848) );
  OR U4960 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U4961 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U4962 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U4963 ( .A(n1855), .B(n1853), .Z(n1875) );
  IV U4964 ( .A(n1875), .Z(n1882) );
  AND U4965 ( .A(n1930), .B(n1854), .Z(n1857) );
  XOR U4966 ( .A(x[89]), .B(x[95]), .Z(n1932) );
  AND U4967 ( .A(n1891), .B(n1932), .Z(n1860) );
  XNOR U4968 ( .A(n1860), .B(n1855), .Z(n1856) );
  XNOR U4969 ( .A(n1857), .B(n1856), .Z(n1881) );
  NANDN U4970 ( .A(n1882), .B(n1881), .Z(n1858) );
  NAND U4971 ( .A(n1886), .B(n1858), .Z(n1868) );
  XNOR U4972 ( .A(n1860), .B(n1859), .Z(n1865) );
  ANDN U4973 ( .B(n1861), .A(x[89]), .Z(n1862) );
  XNOR U4974 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U4975 ( .A(n1865), .B(n1864), .Z(n1878) );
  XOR U4976 ( .A(n1881), .B(n1878), .Z(n1866) );
  NAND U4977 ( .A(n1882), .B(n1866), .Z(n1867) );
  NAND U4978 ( .A(n1868), .B(n1867), .Z(n1929) );
  ANDN U4979 ( .B(n1869), .A(n1929), .Z(n1893) );
  IV U4980 ( .A(n1878), .Z(n1884) );
  XOR U4981 ( .A(n1886), .B(n1882), .Z(n1870) );
  NANDN U4982 ( .A(n1884), .B(n1870), .Z(n1873) );
  NANDN U4983 ( .A(n1882), .B(n1884), .Z(n1871) );
  NANDN U4984 ( .A(n1881), .B(n1871), .Z(n1872) );
  NAND U4985 ( .A(n1873), .B(n1872), .Z(n1939) );
  XNOR U4986 ( .A(n1929), .B(n1939), .Z(n1903) );
  AND U4987 ( .A(n1874), .B(n1903), .Z(n1896) );
  OR U4988 ( .A(n1881), .B(n1878), .Z(n1880) );
  ANDN U4989 ( .B(n1881), .A(n1875), .Z(n1876) );
  XNOR U4990 ( .A(n1876), .B(n1886), .Z(n1877) );
  NAND U4991 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U4992 ( .A(n1880), .B(n1879), .Z(n1900) );
  NAND U4993 ( .A(n1882), .B(n1886), .Z(n1888) );
  NAND U4994 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U4995 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U4996 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4997 ( .A(n1888), .B(n1887), .Z(n1946) );
  NAND U4998 ( .A(n1919), .B(n1889), .Z(n1890) );
  XNOR U4999 ( .A(n1896), .B(n1890), .Z(n1941) );
  XOR U5000 ( .A(n1929), .B(n1946), .Z(n1931) );
  AND U5001 ( .A(n1891), .B(n1931), .Z(n1914) );
  XNOR U5002 ( .A(n1941), .B(n1914), .Z(n1892) );
  XNOR U5003 ( .A(n1893), .B(n1892), .Z(n1949) );
  NAND U5004 ( .A(n1905), .B(n1894), .Z(n1895) );
  XNOR U5005 ( .A(n1896), .B(n1895), .Z(n1922) );
  AND U5006 ( .A(n1897), .B(n1907), .Z(n1940) );
  NANDN U5007 ( .A(n1898), .B(n1900), .Z(n1899) );
  XNOR U5008 ( .A(n1940), .B(n1899), .Z(n1928) );
  XNOR U5009 ( .A(n1922), .B(n1928), .Z(n1911) );
  XOR U5010 ( .A(n1949), .B(n1911), .Z(z[88]) );
  AND U5011 ( .A(n1901), .B(n1900), .Z(n1910) );
  AND U5012 ( .A(n1903), .B(n1902), .Z(n1921) );
  NAND U5013 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U5014 ( .A(n1921), .B(n1906), .Z(n1950) );
  AND U5015 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U5016 ( .A(n1950), .B(n1915), .Z(n1909) );
  XNOR U5017 ( .A(n1910), .B(n1909), .Z(n1937) );
  XNOR U5018 ( .A(n1937), .B(n1911), .Z(n1955) );
  AND U5019 ( .A(n1912), .B(n1939), .Z(n1917) );
  NANDN U5020 ( .A(n1946), .B(n1944), .Z(n1913) );
  XNOR U5021 ( .A(n1914), .B(n1913), .Z(n1927) );
  XNOR U5022 ( .A(n1915), .B(n1927), .Z(n1916) );
  XNOR U5023 ( .A(n1917), .B(n1916), .Z(n1924) );
  NAND U5024 ( .A(n1919), .B(n1918), .Z(n1920) );
  XNOR U5025 ( .A(n1921), .B(n1920), .Z(n1933) );
  XNOR U5026 ( .A(n1922), .B(n1933), .Z(n1923) );
  XNOR U5027 ( .A(n1924), .B(n1923), .Z(n1936) );
  XNOR U5028 ( .A(n1955), .B(n1936), .Z(z[89]) );
  XOR U5029 ( .A(n1926), .B(n1925), .Z(z[8]) );
  XNOR U5030 ( .A(n1928), .B(n1927), .Z(z[90]) );
  NOR U5031 ( .A(n1930), .B(n1929), .Z(n1935) );
  AND U5032 ( .A(n1932), .B(n1931), .Z(n1948) );
  XNOR U5033 ( .A(n1933), .B(n1948), .Z(n1934) );
  XNOR U5034 ( .A(n1935), .B(n1934), .Z(n1954) );
  XOR U5035 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U5036 ( .A(n1954), .B(n1938), .Z(z[91]) );
  XOR U5037 ( .A(n1949), .B(z[90]), .Z(z[92]) );
  AND U5038 ( .A(x[88]), .B(n1939), .Z(n1943) );
  XNOR U5039 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5040 ( .A(n1943), .B(n1942), .Z(n1956) );
  XOR U5041 ( .A(n1944), .B(x[89]), .Z(n1945) );
  NANDN U5042 ( .A(n1946), .B(n1945), .Z(n1947) );
  XNOR U5043 ( .A(n1948), .B(n1947), .Z(n1952) );
  XNOR U5044 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U5045 ( .A(n1952), .B(n1951), .Z(n1953) );
  XNOR U5046 ( .A(n1956), .B(n1953), .Z(z[93]) );
  XNOR U5047 ( .A(n1955), .B(n1954), .Z(z[94]) );
  XOR U5048 ( .A(n1956), .B(z[89]), .Z(z[95]) );
  XOR U5049 ( .A(n1958), .B(n1957), .Z(z[96]) );
  XOR U5050 ( .A(n1960), .B(n1959), .Z(n1961) );
  XNOR U5051 ( .A(n1962), .B(n1961), .Z(z[99]) );
endmodule


module aes_2 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [639:0] key;
  output [127:0] out;
  input clk, rst;
  wire   init, \w0[4][127] , \w0[4][126] , \w0[4][125] , \w0[4][124] ,
         \w0[4][123] , \w0[4][122] , \w0[4][121] , \w0[4][120] , \w0[4][119] ,
         \w0[4][118] , \w0[4][117] , \w0[4][116] , \w0[4][115] , \w0[4][114] ,
         \w0[4][113] , \w0[4][112] , \w0[4][111] , \w0[4][110] , \w0[4][109] ,
         \w0[4][108] , \w0[4][107] , \w0[4][106] , \w0[4][105] , \w0[4][104] ,
         \w0[4][103] , \w0[4][102] , \w0[4][101] , \w0[4][100] , \w0[4][99] ,
         \w0[4][98] , \w0[4][97] , \w0[4][96] , \w0[4][95] , \w0[4][94] ,
         \w0[4][93] , \w0[4][92] , \w0[4][91] , \w0[4][90] , \w0[4][89] ,
         \w0[4][88] , \w0[4][87] , \w0[4][86] , \w0[4][85] , \w0[4][84] ,
         \w0[4][83] , \w0[4][82] , \w0[4][81] , \w0[4][80] , \w0[4][79] ,
         \w0[4][78] , \w0[4][77] , \w0[4][76] , \w0[4][75] , \w0[4][74] ,
         \w0[4][73] , \w0[4][72] , \w0[4][71] , \w0[4][70] , \w0[4][69] ,
         \w0[4][68] , \w0[4][67] , \w0[4][66] , \w0[4][65] , \w0[4][64] ,
         \w0[4][63] , \w0[4][62] , \w0[4][61] , \w0[4][60] , \w0[4][59] ,
         \w0[4][58] , \w0[4][57] , \w0[4][56] , \w0[4][55] , \w0[4][54] ,
         \w0[4][53] , \w0[4][52] , \w0[4][51] , \w0[4][50] , \w0[4][49] ,
         \w0[4][48] , \w0[4][47] , \w0[4][46] , \w0[4][45] , \w0[4][44] ,
         \w0[4][43] , \w0[4][42] , \w0[4][41] , \w0[4][40] , \w0[4][39] ,
         \w0[4][38] , \w0[4][37] , \w0[4][36] , \w0[4][35] , \w0[4][34] ,
         \w0[4][33] , \w0[4][32] , \w0[4][31] , \w0[4][30] , \w0[4][29] ,
         \w0[4][28] , \w0[4][27] , \w0[4][26] , \w0[4][25] , \w0[4][24] ,
         \w0[4][23] , \w0[4][22] , \w0[4][21] , \w0[4][20] , \w0[4][19] ,
         \w0[4][18] , \w0[4][17] , \w0[4][16] , \w0[4][15] , \w0[4][14] ,
         \w0[4][13] , \w0[4][12] , \w0[4][11] , \w0[4][10] , \w0[4][9] ,
         \w0[4][8] , \w0[4][7] , \w0[4][6] , \w0[4][5] , \w0[4][4] ,
         \w0[4][3] , \w0[4][2] , \w0[4][1] , \w0[4][0] , \w1[4][127] ,
         \w1[4][126] , \w1[4][125] , \w1[4][124] , \w1[4][123] , \w1[4][122] ,
         \w1[4][121] , \w1[4][120] , \w1[4][119] , \w1[4][118] , \w1[4][117] ,
         \w1[4][116] , \w1[4][115] , \w1[4][114] , \w1[4][113] , \w1[4][112] ,
         \w1[4][111] , \w1[4][110] , \w1[4][109] , \w1[4][108] , \w1[4][107] ,
         \w1[4][106] , \w1[4][105] , \w1[4][104] , \w1[4][103] , \w1[4][102] ,
         \w1[4][101] , \w1[4][100] , \w1[4][99] , \w1[4][98] , \w1[4][97] ,
         \w1[4][96] , \w1[4][95] , \w1[4][94] , \w1[4][93] , \w1[4][92] ,
         \w1[4][91] , \w1[4][90] , \w1[4][89] , \w1[4][88] , \w1[4][87] ,
         \w1[4][86] , \w1[4][85] , \w1[4][84] , \w1[4][83] , \w1[4][82] ,
         \w1[4][81] , \w1[4][80] , \w1[4][79] , \w1[4][78] , \w1[4][77] ,
         \w1[4][76] , \w1[4][75] , \w1[4][74] , \w1[4][73] , \w1[4][72] ,
         \w1[4][71] , \w1[4][70] , \w1[4][69] , \w1[4][68] , \w1[4][67] ,
         \w1[4][66] , \w1[4][65] , \w1[4][64] , \w1[4][63] , \w1[4][62] ,
         \w1[4][61] , \w1[4][60] , \w1[4][59] , \w1[4][58] , \w1[4][57] ,
         \w1[4][56] , \w1[4][55] , \w1[4][54] , \w1[4][53] , \w1[4][52] ,
         \w1[4][51] , \w1[4][50] , \w1[4][49] , \w1[4][48] , \w1[4][47] ,
         \w1[4][46] , \w1[4][45] , \w1[4][44] , \w1[4][43] , \w1[4][42] ,
         \w1[4][41] , \w1[4][40] , \w1[4][39] , \w1[4][38] , \w1[4][37] ,
         \w1[4][36] , \w1[4][35] , \w1[4][34] , \w1[4][33] , \w1[4][32] ,
         \w1[4][31] , \w1[4][30] , \w1[4][29] , \w1[4][28] , \w1[4][27] ,
         \w1[4][26] , \w1[4][25] , \w1[4][24] , \w1[4][23] , \w1[4][22] ,
         \w1[4][21] , \w1[4][20] , \w1[4][19] , \w1[4][18] , \w1[4][17] ,
         \w1[4][16] , \w1[4][15] , \w1[4][14] , \w1[4][13] , \w1[4][12] ,
         \w1[4][11] , \w1[4][10] , \w1[4][9] , \w1[4][8] , \w1[4][7] ,
         \w1[4][6] , \w1[4][5] , \w1[4][4] , \w1[4][3] , \w1[4][2] ,
         \w1[4][1] , \w1[4][0] , \w1[3][127] , \w1[3][126] , \w1[3][125] ,
         \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] , \w1[3][120] ,
         \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] , \w1[3][115] ,
         \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] , \w1[3][110] ,
         \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] , \w1[3][105] ,
         \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] , \w1[3][100] ,
         \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] , \w1[3][95] ,
         \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] , \w1[3][90] ,
         \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] , \w1[3][85] ,
         \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] , \w1[3][80] ,
         \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] , \w1[3][75] ,
         \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] , \w1[3][70] ,
         \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] , \w1[3][65] ,
         \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] , \w1[3][60] ,
         \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] , \w1[3][55] ,
         \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] , \w1[3][50] ,
         \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] , \w1[3][45] ,
         \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] , \w1[3][40] ,
         \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] , \w1[3][35] ,
         \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] , \w1[3][30] ,
         \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] , \w1[3][25] ,
         \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] , \w1[3][20] ,
         \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] , \w1[3][15] ,
         \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] , \w1[3][10] ,
         \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] , \w1[3][5] ,
         \w1[3][4] , \w1[3][3] , \w1[3][2] , \w1[3][1] , \w1[3][0] ,
         \w1[2][127] , \w1[2][126] , \w1[2][125] , \w1[2][124] , \w1[2][123] ,
         \w1[2][122] , \w1[2][121] , \w1[2][120] , \w1[2][119] , \w1[2][118] ,
         \w1[2][117] , \w1[2][116] , \w1[2][115] , \w1[2][114] , \w1[2][113] ,
         \w1[2][112] , \w1[2][111] , \w1[2][110] , \w1[2][109] , \w1[2][108] ,
         \w1[2][107] , \w1[2][106] , \w1[2][105] , \w1[2][104] , \w1[2][103] ,
         \w1[2][102] , \w1[2][101] , \w1[2][100] , \w1[2][99] , \w1[2][98] ,
         \w1[2][97] , \w1[2][96] , \w1[2][95] , \w1[2][94] , \w1[2][93] ,
         \w1[2][92] , \w1[2][91] , \w1[2][90] , \w1[2][89] , \w1[2][88] ,
         \w1[2][87] , \w1[2][86] , \w1[2][85] , \w1[2][84] , \w1[2][83] ,
         \w1[2][82] , \w1[2][81] , \w1[2][80] , \w1[2][79] , \w1[2][78] ,
         \w1[2][77] , \w1[2][76] , \w1[2][75] , \w1[2][74] , \w1[2][73] ,
         \w1[2][72] , \w1[2][71] , \w1[2][70] , \w1[2][69] , \w1[2][68] ,
         \w1[2][67] , \w1[2][66] , \w1[2][65] , \w1[2][64] , \w1[2][63] ,
         \w1[2][62] , \w1[2][61] , \w1[2][60] , \w1[2][59] , \w1[2][58] ,
         \w1[2][57] , \w1[2][56] , \w1[2][55] , \w1[2][54] , \w1[2][53] ,
         \w1[2][52] , \w1[2][51] , \w1[2][50] , \w1[2][49] , \w1[2][48] ,
         \w1[2][47] , \w1[2][46] , \w1[2][45] , \w1[2][44] , \w1[2][43] ,
         \w1[2][42] , \w1[2][41] , \w1[2][40] , \w1[2][39] , \w1[2][38] ,
         \w1[2][37] , \w1[2][36] , \w1[2][35] , \w1[2][34] , \w1[2][33] ,
         \w1[2][32] , \w1[2][31] , \w1[2][30] , \w1[2][29] , \w1[2][28] ,
         \w1[2][27] , \w1[2][26] , \w1[2][25] , \w1[2][24] , \w1[2][23] ,
         \w1[2][22] , \w1[2][21] , \w1[2][20] , \w1[2][19] , \w1[2][18] ,
         \w1[2][17] , \w1[2][16] , \w1[2][15] , \w1[2][14] , \w1[2][13] ,
         \w1[2][12] , \w1[2][11] , \w1[2][10] , \w1[2][9] , \w1[2][8] ,
         \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] , \w1[2][3] ,
         \w1[2][2] , \w1[2][1] , \w1[2][0] , \w1[1][127] , \w1[1][126] ,
         \w1[1][125] , \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] ,
         \w1[1][120] , \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] ,
         \w1[1][115] , \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] ,
         \w1[1][110] , \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] ,
         \w1[1][105] , \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] ,
         \w1[1][100] , \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] ,
         \w1[1][95] , \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] ,
         \w1[1][90] , \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] ,
         \w1[1][85] , \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] ,
         \w1[1][80] , \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] ,
         \w1[1][75] , \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] ,
         \w1[1][70] , \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] ,
         \w1[1][65] , \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] ,
         \w1[1][60] , \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] ,
         \w1[1][55] , \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] ,
         \w1[1][50] , \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] ,
         \w1[1][45] , \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] ,
         \w1[1][40] , \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] ,
         \w1[1][35] , \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] ,
         \w1[1][30] , \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] ,
         \w1[1][25] , \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] ,
         \w1[1][20] , \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] ,
         \w1[1][15] , \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] ,
         \w1[1][10] , \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] ,
         \w1[1][5] , \w1[1][4] , \w1[1][3] , \w1[1][2] , \w1[1][1] ,
         \w1[1][0] , \w1[0][127] , \w1[0][126] , \w1[0][125] , \w1[0][124] ,
         \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , \w1[0][119] ,
         \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , \w1[0][114] ,
         \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , \w1[0][109] ,
         \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , \w1[0][104] ,
         \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , \w1[0][99] ,
         \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , \w1[0][94] ,
         \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , \w1[0][89] ,
         \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , \w1[0][84] ,
         \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , \w1[0][79] ,
         \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , \w1[0][74] ,
         \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , \w1[0][69] ,
         \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , \w1[0][64] ,
         \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , \w1[0][59] ,
         \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , \w1[0][54] ,
         \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , \w1[0][49] ,
         \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , \w1[0][44] ,
         \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , \w1[0][39] ,
         \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , \w1[0][34] ,
         \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , \w1[0][29] ,
         \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , \w1[0][24] ,
         \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , \w1[0][19] ,
         \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , \w1[0][14] ,
         \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , \w1[0][9] ,
         \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] ,
         \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] , \w3[4][127] ,
         \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] , \w3[4][122] ,
         \w3[4][121] , \w3[4][120] , \w3[4][119] , \w3[4][118] , \w3[4][117] ,
         \w3[4][116] , \w3[4][115] , \w3[4][114] , \w3[4][113] , \w3[4][112] ,
         \w3[4][111] , \w3[4][110] , \w3[4][109] , \w3[4][108] , \w3[4][107] ,
         \w3[4][106] , \w3[4][105] , \w3[4][104] , \w3[4][103] , \w3[4][102] ,
         \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] , \w3[4][97] ,
         \w3[4][96] , \w3[4][95] , \w3[4][94] , \w3[4][93] , \w3[4][92] ,
         \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] , \w3[4][87] ,
         \w3[4][86] , \w3[4][85] , \w3[4][84] , \w3[4][83] , \w3[4][82] ,
         \w3[4][81] , \w3[4][80] , \w3[4][79] , \w3[4][78] , \w3[4][77] ,
         \w3[4][76] , \w3[4][75] , \w3[4][74] , \w3[4][73] , \w3[4][72] ,
         \w3[4][71] , \w3[4][70] , \w3[4][69] , \w3[4][68] , \w3[4][67] ,
         \w3[4][66] , \w3[4][65] , \w3[4][64] , \w3[4][63] , \w3[4][62] ,
         \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] , \w3[4][57] ,
         \w3[4][56] , \w3[4][55] , \w3[4][54] , \w3[4][53] , \w3[4][52] ,
         \w3[4][51] , \w3[4][50] , \w3[4][49] , \w3[4][48] , \w3[4][47] ,
         \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] , \w3[4][42] ,
         \w3[4][41] , \w3[4][40] , \w3[4][39] , \w3[4][38] , \w3[4][37] ,
         \w3[4][36] , \w3[4][35] , \w3[4][34] , \w3[4][33] , \w3[4][32] ,
         \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] , \w3[4][27] ,
         \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][23] , \w3[4][22] ,
         \w3[4][21] , \w3[4][20] , \w3[4][19] , \w3[4][18] , \w3[4][17] ,
         \w3[4][16] , \w3[4][15] , \w3[4][14] , \w3[4][13] , \w3[4][12] ,
         \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] , \w3[4][7] ,
         \w3[4][6] , \w3[4][5] , \w3[4][4] , \w3[4][3] , \w3[4][2] ,
         \w3[4][1] , \w3[4][0] , \w3[3][127] , \w3[3][126] , \w3[3][125] ,
         \w3[3][124] , \w3[3][123] , \w3[3][122] , \w3[3][121] , \w3[3][120] ,
         \w3[3][119] , \w3[3][118] , \w3[3][117] , \w3[3][116] , \w3[3][115] ,
         \w3[3][114] , \w3[3][113] , \w3[3][112] , \w3[3][111] , \w3[3][110] ,
         \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] , \w3[3][105] ,
         \w3[3][104] , \w3[3][103] , \w3[3][102] , \w3[3][101] , \w3[3][100] ,
         \w3[3][99] , \w3[3][98] , \w3[3][97] , \w3[3][96] , \w3[3][95] ,
         \w3[3][94] , \w3[3][93] , \w3[3][92] , \w3[3][91] , \w3[3][90] ,
         \w3[3][89] , \w3[3][88] , \w3[3][87] , \w3[3][86] , \w3[3][85] ,
         \w3[3][84] , \w3[3][83] , \w3[3][82] , \w3[3][81] , \w3[3][80] ,
         \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] , \w3[3][75] ,
         \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][71] , \w3[3][70] ,
         \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] , \w3[3][65] ,
         \w3[3][64] , \w3[3][63] , \w3[3][62] , \w3[3][61] , \w3[3][60] ,
         \w3[3][59] , \w3[3][58] , \w3[3][57] , \w3[3][56] , \w3[3][55] ,
         \w3[3][54] , \w3[3][53] , \w3[3][52] , \w3[3][51] , \w3[3][50] ,
         \w3[3][49] , \w3[3][48] , \w3[3][47] , \w3[3][46] , \w3[3][45] ,
         \w3[3][44] , \w3[3][43] , \w3[3][42] , \w3[3][41] , \w3[3][40] ,
         \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] , \w3[3][35] ,
         \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][31] , \w3[3][30] ,
         \w3[3][29] , \w3[3][28] , \w3[3][27] , \w3[3][26] , \w3[3][25] ,
         \w3[3][24] , \w3[3][23] , \w3[3][22] , \w3[3][21] , \w3[3][20] ,
         \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] , \w3[3][15] ,
         \w3[3][14] , \w3[3][13] , \w3[3][12] , \w3[3][11] , \w3[3][10] ,
         \w3[3][9] , \w3[3][8] , \w3[3][7] , \w3[3][6] , \w3[3][5] ,
         \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] , \w3[3][0] ,
         \w3[2][127] , \w3[2][126] , \w3[2][125] , \w3[2][124] , \w3[2][123] ,
         \w3[2][122] , \w3[2][121] , \w3[2][120] , \w3[2][119] , \w3[2][118] ,
         \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] , \w3[2][113] ,
         \w3[2][112] , \w3[2][111] , \w3[2][110] , \w3[2][109] , \w3[2][108] ,
         \w3[2][107] , \w3[2][106] , \w3[2][105] , \w3[2][104] , \w3[2][103] ,
         \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] , \w3[2][98] ,
         \w3[2][97] , \w3[2][96] , \w3[2][95] , \w3[2][94] , \w3[2][93] ,
         \w3[2][92] , \w3[2][91] , \w3[2][90] , \w3[2][89] , \w3[2][88] ,
         \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] , \w3[2][83] ,
         \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][79] , \w3[2][78] ,
         \w3[2][77] , \w3[2][76] , \w3[2][75] , \w3[2][74] , \w3[2][73] ,
         \w3[2][72] , \w3[2][71] , \w3[2][70] , \w3[2][69] , \w3[2][68] ,
         \w3[2][67] , \w3[2][66] , \w3[2][65] , \w3[2][64] , \w3[2][63] ,
         \w3[2][62] , \w3[2][61] , \w3[2][60] , \w3[2][59] , \w3[2][58] ,
         \w3[2][57] , \w3[2][56] , \w3[2][55] , \w3[2][54] , \w3[2][53] ,
         \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] , \w3[2][48] ,
         \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] , \w3[2][43] ,
         \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][39] , \w3[2][38] ,
         \w3[2][37] , \w3[2][36] , \w3[2][35] , \w3[2][34] , \w3[2][33] ,
         \w3[2][32] , \w3[2][31] , \w3[2][30] , \w3[2][29] , \w3[2][28] ,
         \w3[2][27] , \w3[2][26] , \w3[2][25] , \w3[2][24] , \w3[2][23] ,
         \w3[2][22] , \w3[2][21] , \w3[2][20] , \w3[2][19] , \w3[2][18] ,
         \w3[2][17] , \w3[2][16] , \w3[2][15] , \w3[2][14] , \w3[2][13] ,
         \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] , \w3[2][8] ,
         \w3[2][7] , \w3[2][6] , \w3[2][5] , \w3[2][4] , \w3[2][3] ,
         \w3[2][2] , \w3[2][1] , \w3[2][0] , \w3[1][127] , \w3[1][126] ,
         \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , \w3[1][121] ,
         \w3[1][120] , \w3[1][119] , \w3[1][118] , \w3[1][117] , \w3[1][116] ,
         \w3[1][115] , \w3[1][114] , \w3[1][113] , \w3[1][112] , \w3[1][111] ,
         \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] ,
         \w3[1][105] , \w3[1][104] , \w3[1][103] , \w3[1][102] , \w3[1][101] ,
         \w3[1][100] , \w3[1][99] , \w3[1][98] , \w3[1][97] , \w3[1][96] ,
         \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , \w3[1][91] ,
         \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][87] , \w3[1][86] ,
         \w3[1][85] , \w3[1][84] , \w3[1][83] , \w3[1][82] , \w3[1][81] ,
         \w3[1][80] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] ,
         \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][71] ,
         \w3[1][70] , \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] ,
         \w3[1][65] , \w3[1][64] , \w3[1][63] , \w3[1][62] , \w3[1][61] ,
         \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , \w3[1][56] ,
         \w3[1][55] , \w3[1][54] , \w3[1][53] , \w3[1][52] , \w3[1][51] ,
         \w3[1][50] , \w3[1][49] , \w3[1][48] , \w3[1][47] , \w3[1][46] ,
         \w3[1][45] , \w3[1][44] , \w3[1][43] , \w3[1][42] , \w3[1][41] ,
         \w3[1][40] , \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] ,
         \w3[1][35] , \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][31] ,
         \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , \w3[1][26] ,
         \w3[1][25] , \w3[1][24] , \w3[1][23] , \w3[1][22] , \w3[1][21] ,
         \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] ,
         \w3[1][15] , \w3[1][14] , \w3[1][13] , \w3[1][12] , \w3[1][11] ,
         \w3[1][10] , \w3[1][9] , \w3[1][8] , \w3[1][7] , \w3[1][6] ,
         \w3[1][5] , \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] ,
         \w3[1][0] , \w3[0][127] , \w3[0][126] , \w3[0][125] , \w3[0][124] ,
         \w3[0][123] , \w3[0][122] , \w3[0][121] , \w3[0][120] , \w3[0][119] ,
         \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] ,
         \w3[0][113] , \w3[0][112] , \w3[0][111] , \w3[0][110] , \w3[0][109] ,
         \w3[0][108] , \w3[0][107] , \w3[0][106] , \w3[0][105] , \w3[0][104] ,
         \w3[0][103] , \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] ,
         \w3[0][98] , \w3[0][97] , \w3[0][96] , \w3[0][95] , \w3[0][94] ,
         \w3[0][93] , \w3[0][92] , \w3[0][91] , \w3[0][90] , \w3[0][89] ,
         \w3[0][88] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] ,
         \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][79] ,
         \w3[0][78] , \w3[0][77] , \w3[0][76] , \w3[0][75] , \w3[0][74] ,
         \w3[0][73] , \w3[0][72] , \w3[0][71] , \w3[0][70] , \w3[0][69] ,
         \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , \w3[0][64] ,
         \w3[0][63] , \w3[0][62] , \w3[0][61] , \w3[0][60] , \w3[0][59] ,
         \w3[0][58] , \w3[0][57] , \w3[0][56] , \w3[0][55] , \w3[0][54] ,
         \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] ,
         \w3[0][48] , \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] ,
         \w3[0][43] , \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][39] ,
         \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , \w3[0][34] ,
         \w3[0][33] , \w3[0][32] , \w3[0][31] , \w3[0][30] , \w3[0][29] ,
         \w3[0][28] , \w3[0][27] , \w3[0][26] , \w3[0][25] , \w3[0][24] ,
         \w3[0][23] , \w3[0][22] , \w3[0][21] , \w3[0][20] , \w3[0][19] ,
         \w3[0][18] , \w3[0][17] , \w3[0][16] , \w3[0][15] , \w3[0][14] ,
         \w3[0][13] , \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] ,
         \w3[0][8] , \w3[0][7] , \w3[0][6] , \w3[0][5] , \w3[0][4] ,
         \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904;
  wire   [127:0] state;

  SubBytes_0 \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  SubBytes_4 \SUBBYTES[1].a  ( .x({\w1[1][127] , \w1[1][126] , \w1[1][125] , 
        \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] , \w1[1][120] , 
        \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] , \w1[1][115] , 
        \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] , \w1[1][110] , 
        \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] , \w1[1][105] , 
        \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] , \w1[1][100] , 
        \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] , \w1[1][95] , 
        \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] , \w1[1][90] , 
        \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] , \w1[1][85] , 
        \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] , \w1[1][80] , 
        \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] , \w1[1][75] , 
        \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] , \w1[1][70] , 
        \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] , \w1[1][65] , 
        \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] , \w1[1][60] , 
        \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] , \w1[1][55] , 
        \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] , \w1[1][50] , 
        \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] , \w1[1][45] , 
        \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] , \w1[1][40] , 
        \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] , \w1[1][35] , 
        \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] , \w1[1][30] , 
        \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] , \w1[1][25] , 
        \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] , \w1[1][20] , 
        \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] , \w1[1][15] , 
        \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] , \w1[1][10] , 
        \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] , \w1[1][5] , \w1[1][4] , 
        \w1[1][3] , \w1[1][2] , \w1[1][1] , \w1[1][0] }), .z({\w3[1][127] , 
        \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , 
        \w3[1][121] , \w3[1][120] , \w3[1][23] , \w3[1][22] , \w3[1][21] , 
        \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] , 
        \w3[1][47] , \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , 
        \w3[1][42] , \w3[1][41] , \w3[1][40] , \w3[1][71] , \w3[1][70] , 
        \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] , \w3[1][65] , 
        \w3[1][64] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , 
        \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][119] , 
        \w3[1][118] , \w3[1][117] , \w3[1][116] , \w3[1][115] , \w3[1][114] , 
        \w3[1][113] , \w3[1][112] , \w3[1][15] , \w3[1][14] , \w3[1][13] , 
        \w3[1][12] , \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , 
        \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] , \w3[1][35] , 
        \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][63] , \w3[1][62] , 
        \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , 
        \w3[1][56] , \w3[1][87] , \w3[1][86] , \w3[1][85] , \w3[1][84] , 
        \w3[1][83] , \w3[1][82] , \w3[1][81] , \w3[1][80] , \w3[1][111] , 
        \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] , 
        \w3[1][105] , \w3[1][104] , \w3[1][7] , \w3[1][6] , \w3[1][5] , 
        \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] , \w3[1][0] , 
        \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , 
        \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][55] , \w3[1][54] , 
        \w3[1][53] , \w3[1][52] , \w3[1][51] , \w3[1][50] , \w3[1][49] , 
        \w3[1][48] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] , 
        \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][103] , 
        \w3[1][102] , \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , 
        \w3[1][97] , \w3[1][96] }) );
  SubBytes_3 \SUBBYTES[2].a  ( .x({\w1[2][127] , \w1[2][126] , \w1[2][125] , 
        \w1[2][124] , \w1[2][123] , \w1[2][122] , \w1[2][121] , \w1[2][120] , 
        \w1[2][119] , \w1[2][118] , \w1[2][117] , \w1[2][116] , \w1[2][115] , 
        \w1[2][114] , \w1[2][113] , \w1[2][112] , \w1[2][111] , \w1[2][110] , 
        \w1[2][109] , \w1[2][108] , \w1[2][107] , \w1[2][106] , \w1[2][105] , 
        \w1[2][104] , \w1[2][103] , \w1[2][102] , \w1[2][101] , \w1[2][100] , 
        \w1[2][99] , \w1[2][98] , \w1[2][97] , \w1[2][96] , \w1[2][95] , 
        \w1[2][94] , \w1[2][93] , \w1[2][92] , \w1[2][91] , \w1[2][90] , 
        \w1[2][89] , \w1[2][88] , \w1[2][87] , \w1[2][86] , \w1[2][85] , 
        \w1[2][84] , \w1[2][83] , \w1[2][82] , \w1[2][81] , \w1[2][80] , 
        \w1[2][79] , \w1[2][78] , \w1[2][77] , \w1[2][76] , \w1[2][75] , 
        \w1[2][74] , \w1[2][73] , \w1[2][72] , \w1[2][71] , \w1[2][70] , 
        \w1[2][69] , \w1[2][68] , \w1[2][67] , \w1[2][66] , \w1[2][65] , 
        \w1[2][64] , \w1[2][63] , \w1[2][62] , \w1[2][61] , \w1[2][60] , 
        \w1[2][59] , \w1[2][58] , \w1[2][57] , \w1[2][56] , \w1[2][55] , 
        \w1[2][54] , \w1[2][53] , \w1[2][52] , \w1[2][51] , \w1[2][50] , 
        \w1[2][49] , \w1[2][48] , \w1[2][47] , \w1[2][46] , \w1[2][45] , 
        \w1[2][44] , \w1[2][43] , \w1[2][42] , \w1[2][41] , \w1[2][40] , 
        \w1[2][39] , \w1[2][38] , \w1[2][37] , \w1[2][36] , \w1[2][35] , 
        \w1[2][34] , \w1[2][33] , \w1[2][32] , \w1[2][31] , \w1[2][30] , 
        \w1[2][29] , \w1[2][28] , \w1[2][27] , \w1[2][26] , \w1[2][25] , 
        \w1[2][24] , \w1[2][23] , \w1[2][22] , \w1[2][21] , \w1[2][20] , 
        \w1[2][19] , \w1[2][18] , \w1[2][17] , \w1[2][16] , \w1[2][15] , 
        \w1[2][14] , \w1[2][13] , \w1[2][12] , \w1[2][11] , \w1[2][10] , 
        \w1[2][9] , \w1[2][8] , \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] , 
        \w1[2][3] , \w1[2][2] , \w1[2][1] , \w1[2][0] }), .z({\w3[2][127] , 
        \w3[2][126] , \w3[2][125] , \w3[2][124] , \w3[2][123] , \w3[2][122] , 
        \w3[2][121] , \w3[2][120] , \w3[2][23] , \w3[2][22] , \w3[2][21] , 
        \w3[2][20] , \w3[2][19] , \w3[2][18] , \w3[2][17] , \w3[2][16] , 
        \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] , \w3[2][43] , 
        \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][71] , \w3[2][70] , 
        \w3[2][69] , \w3[2][68] , \w3[2][67] , \w3[2][66] , \w3[2][65] , 
        \w3[2][64] , \w3[2][95] , \w3[2][94] , \w3[2][93] , \w3[2][92] , 
        \w3[2][91] , \w3[2][90] , \w3[2][89] , \w3[2][88] , \w3[2][119] , 
        \w3[2][118] , \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] , 
        \w3[2][113] , \w3[2][112] , \w3[2][15] , \w3[2][14] , \w3[2][13] , 
        \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] , \w3[2][8] , 
        \w3[2][39] , \w3[2][38] , \w3[2][37] , \w3[2][36] , \w3[2][35] , 
        \w3[2][34] , \w3[2][33] , \w3[2][32] , \w3[2][63] , \w3[2][62] , 
        \w3[2][61] , \w3[2][60] , \w3[2][59] , \w3[2][58] , \w3[2][57] , 
        \w3[2][56] , \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] , 
        \w3[2][83] , \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][111] , 
        \w3[2][110] , \w3[2][109] , \w3[2][108] , \w3[2][107] , \w3[2][106] , 
        \w3[2][105] , \w3[2][104] , \w3[2][7] , \w3[2][6] , \w3[2][5] , 
        \w3[2][4] , \w3[2][3] , \w3[2][2] , \w3[2][1] , \w3[2][0] , 
        \w3[2][31] , \w3[2][30] , \w3[2][29] , \w3[2][28] , \w3[2][27] , 
        \w3[2][26] , \w3[2][25] , \w3[2][24] , \w3[2][55] , \w3[2][54] , 
        \w3[2][53] , \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] , 
        \w3[2][48] , \w3[2][79] , \w3[2][78] , \w3[2][77] , \w3[2][76] , 
        \w3[2][75] , \w3[2][74] , \w3[2][73] , \w3[2][72] , \w3[2][103] , 
        \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] , \w3[2][98] , 
        \w3[2][97] , \w3[2][96] }) );
  SubBytes_2 \SUBBYTES[3].a  ( .x({\w1[3][127] , \w1[3][126] , \w1[3][125] , 
        \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] , \w1[3][120] , 
        \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] , \w1[3][115] , 
        \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] , \w1[3][110] , 
        \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] , \w1[3][105] , 
        \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] , \w1[3][100] , 
        \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] , \w1[3][95] , 
        \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] , \w1[3][90] , 
        \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] , \w1[3][85] , 
        \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] , \w1[3][80] , 
        \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] , \w1[3][75] , 
        \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] , \w1[3][70] , 
        \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] , \w1[3][65] , 
        \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] , \w1[3][60] , 
        \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] , \w1[3][55] , 
        \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] , \w1[3][50] , 
        \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] , \w1[3][45] , 
        \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] , \w1[3][40] , 
        \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] , \w1[3][35] , 
        \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] , \w1[3][30] , 
        \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] , \w1[3][25] , 
        \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] , \w1[3][20] , 
        \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] , \w1[3][15] , 
        \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] , \w1[3][10] , 
        \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] , \w1[3][5] , \w1[3][4] , 
        \w1[3][3] , \w1[3][2] , \w1[3][1] , \w1[3][0] }), .z({\w3[3][127] , 
        \w3[3][126] , \w3[3][125] , \w3[3][124] , \w3[3][123] , \w3[3][122] , 
        \w3[3][121] , \w3[3][120] , \w3[3][23] , \w3[3][22] , \w3[3][21] , 
        \w3[3][20] , \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] , 
        \w3[3][47] , \w3[3][46] , \w3[3][45] , \w3[3][44] , \w3[3][43] , 
        \w3[3][42] , \w3[3][41] , \w3[3][40] , \w3[3][71] , \w3[3][70] , 
        \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] , \w3[3][65] , 
        \w3[3][64] , \w3[3][95] , \w3[3][94] , \w3[3][93] , \w3[3][92] , 
        \w3[3][91] , \w3[3][90] , \w3[3][89] , \w3[3][88] , \w3[3][119] , 
        \w3[3][118] , \w3[3][117] , \w3[3][116] , \w3[3][115] , \w3[3][114] , 
        \w3[3][113] , \w3[3][112] , \w3[3][15] , \w3[3][14] , \w3[3][13] , 
        \w3[3][12] , \w3[3][11] , \w3[3][10] , \w3[3][9] , \w3[3][8] , 
        \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] , \w3[3][35] , 
        \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][63] , \w3[3][62] , 
        \w3[3][61] , \w3[3][60] , \w3[3][59] , \w3[3][58] , \w3[3][57] , 
        \w3[3][56] , \w3[3][87] , \w3[3][86] , \w3[3][85] , \w3[3][84] , 
        \w3[3][83] , \w3[3][82] , \w3[3][81] , \w3[3][80] , \w3[3][111] , 
        \w3[3][110] , \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] , 
        \w3[3][105] , \w3[3][104] , \w3[3][7] , \w3[3][6] , \w3[3][5] , 
        \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] , \w3[3][0] , 
        \w3[3][31] , \w3[3][30] , \w3[3][29] , \w3[3][28] , \w3[3][27] , 
        \w3[3][26] , \w3[3][25] , \w3[3][24] , \w3[3][55] , \w3[3][54] , 
        \w3[3][53] , \w3[3][52] , \w3[3][51] , \w3[3][50] , \w3[3][49] , 
        \w3[3][48] , \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] , 
        \w3[3][75] , \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][103] , 
        \w3[3][102] , \w3[3][101] , \w3[3][100] , \w3[3][99] , \w3[3][98] , 
        \w3[3][97] , \w3[3][96] }) );
  SubBytes_1 \SUBBYTES[4].a  ( .x({\w1[4][127] , \w1[4][126] , \w1[4][125] , 
        \w1[4][124] , \w1[4][123] , \w1[4][122] , \w1[4][121] , \w1[4][120] , 
        \w1[4][119] , \w1[4][118] , \w1[4][117] , \w1[4][116] , \w1[4][115] , 
        \w1[4][114] , \w1[4][113] , \w1[4][112] , \w1[4][111] , \w1[4][110] , 
        \w1[4][109] , \w1[4][108] , \w1[4][107] , \w1[4][106] , \w1[4][105] , 
        \w1[4][104] , \w1[4][103] , \w1[4][102] , \w1[4][101] , \w1[4][100] , 
        \w1[4][99] , \w1[4][98] , \w1[4][97] , \w1[4][96] , \w1[4][95] , 
        \w1[4][94] , \w1[4][93] , \w1[4][92] , \w1[4][91] , \w1[4][90] , 
        \w1[4][89] , \w1[4][88] , \w1[4][87] , \w1[4][86] , \w1[4][85] , 
        \w1[4][84] , \w1[4][83] , \w1[4][82] , \w1[4][81] , \w1[4][80] , 
        \w1[4][79] , \w1[4][78] , \w1[4][77] , \w1[4][76] , \w1[4][75] , 
        \w1[4][74] , \w1[4][73] , \w1[4][72] , \w1[4][71] , \w1[4][70] , 
        \w1[4][69] , \w1[4][68] , \w1[4][67] , \w1[4][66] , \w1[4][65] , 
        \w1[4][64] , \w1[4][63] , \w1[4][62] , \w1[4][61] , \w1[4][60] , 
        \w1[4][59] , \w1[4][58] , \w1[4][57] , \w1[4][56] , \w1[4][55] , 
        \w1[4][54] , \w1[4][53] , \w1[4][52] , \w1[4][51] , \w1[4][50] , 
        \w1[4][49] , \w1[4][48] , \w1[4][47] , \w1[4][46] , \w1[4][45] , 
        \w1[4][44] , \w1[4][43] , \w1[4][42] , \w1[4][41] , \w1[4][40] , 
        \w1[4][39] , \w1[4][38] , \w1[4][37] , \w1[4][36] , \w1[4][35] , 
        \w1[4][34] , \w1[4][33] , \w1[4][32] , \w1[4][31] , \w1[4][30] , 
        \w1[4][29] , \w1[4][28] , \w1[4][27] , \w1[4][26] , \w1[4][25] , 
        \w1[4][24] , \w1[4][23] , \w1[4][22] , \w1[4][21] , \w1[4][20] , 
        \w1[4][19] , \w1[4][18] , \w1[4][17] , \w1[4][16] , \w1[4][15] , 
        \w1[4][14] , \w1[4][13] , \w1[4][12] , \w1[4][11] , \w1[4][10] , 
        \w1[4][9] , \w1[4][8] , \w1[4][7] , \w1[4][6] , \w1[4][5] , \w1[4][4] , 
        \w1[4][3] , \w1[4][2] , \w1[4][1] , \w1[4][0] }), .z({\w3[4][127] , 
        \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] , \w3[4][122] , 
        \w3[4][121] , \w3[4][120] , \w3[4][23] , \w3[4][22] , \w3[4][21] , 
        \w3[4][20] , \w3[4][19] , \w3[4][18] , \w3[4][17] , \w3[4][16] , 
        \w3[4][47] , \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] , 
        \w3[4][42] , \w3[4][41] , \w3[4][40] , \w3[4][71] , \w3[4][70] , 
        \w3[4][69] , \w3[4][68] , \w3[4][67] , \w3[4][66] , \w3[4][65] , 
        \w3[4][64] , \w3[4][95] , \w3[4][94] , \w3[4][93] , \w3[4][92] , 
        \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] , \w3[4][119] , 
        \w3[4][118] , \w3[4][117] , \w3[4][116] , \w3[4][115] , \w3[4][114] , 
        \w3[4][113] , \w3[4][112] , \w3[4][15] , \w3[4][14] , \w3[4][13] , 
        \w3[4][12] , \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] , 
        \w3[4][39] , \w3[4][38] , \w3[4][37] , \w3[4][36] , \w3[4][35] , 
        \w3[4][34] , \w3[4][33] , \w3[4][32] , \w3[4][63] , \w3[4][62] , 
        \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] , \w3[4][57] , 
        \w3[4][56] , \w3[4][87] , \w3[4][86] , \w3[4][85] , \w3[4][84] , 
        \w3[4][83] , \w3[4][82] , \w3[4][81] , \w3[4][80] , \w3[4][111] , 
        \w3[4][110] , \w3[4][109] , \w3[4][108] , \w3[4][107] , \w3[4][106] , 
        \w3[4][105] , \w3[4][104] , \w3[4][7] , \w3[4][6] , \w3[4][5] , 
        \w3[4][4] , \w3[4][3] , \w3[4][2] , \w3[4][1] , \w3[4][0] , 
        \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] , \w3[4][27] , 
        \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][55] , \w3[4][54] , 
        \w3[4][53] , \w3[4][52] , \w3[4][51] , \w3[4][50] , \w3[4][49] , 
        \w3[4][48] , \w3[4][79] , \w3[4][78] , \w3[4][77] , \w3[4][76] , 
        \w3[4][75] , \w3[4][74] , \w3[4][73] , \w3[4][72] , \w3[4][103] , 
        \w3[4][102] , \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] , 
        \w3[4][97] , \w3[4][96] }) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \state_reg[0]  ( .D(\w0[4][0] ), .CLK(clk), .RST(rst), .Q(state[0]) );
  DFF \state_reg[71]  ( .D(\w0[4][71] ), .CLK(clk), .RST(rst), .Q(state[71])
         );
  DFF \state_reg[88]  ( .D(\w0[4][88] ), .CLK(clk), .RST(rst), .Q(state[88])
         );
  DFF \state_reg[80]  ( .D(\w0[4][80] ), .CLK(clk), .RST(rst), .Q(state[80])
         );
  DFF \state_reg[81]  ( .D(\w0[4][81] ), .CLK(clk), .RST(rst), .Q(state[81])
         );
  DFF \state_reg[64]  ( .D(\w0[4][64] ), .CLK(clk), .RST(rst), .Q(state[64])
         );
  DFF \state_reg[72]  ( .D(\w0[4][72] ), .CLK(clk), .RST(rst), .Q(state[72])
         );
  DFF \state_reg[89]  ( .D(\w0[4][89] ), .CLK(clk), .RST(rst), .Q(state[89])
         );
  DFF \state_reg[82]  ( .D(\w0[4][82] ), .CLK(clk), .RST(rst), .Q(state[82])
         );
  DFF \state_reg[65]  ( .D(\w0[4][65] ), .CLK(clk), .RST(rst), .Q(state[65])
         );
  DFF \state_reg[73]  ( .D(\w0[4][73] ), .CLK(clk), .RST(rst), .Q(state[73])
         );
  DFF \state_reg[90]  ( .D(\w0[4][90] ), .CLK(clk), .RST(rst), .Q(state[90])
         );
  DFF \state_reg[83]  ( .D(\w0[4][83] ), .CLK(clk), .RST(rst), .Q(state[83])
         );
  DFF \state_reg[66]  ( .D(\w0[4][66] ), .CLK(clk), .RST(rst), .Q(state[66])
         );
  DFF \state_reg[74]  ( .D(\w0[4][74] ), .CLK(clk), .RST(rst), .Q(state[74])
         );
  DFF \state_reg[91]  ( .D(\w0[4][91] ), .CLK(clk), .RST(rst), .Q(state[91])
         );
  DFF \state_reg[75]  ( .D(\w0[4][75] ), .CLK(clk), .RST(rst), .Q(state[75])
         );
  DFF \state_reg[67]  ( .D(\w0[4][67] ), .CLK(clk), .RST(rst), .Q(state[67])
         );
  DFF \state_reg[84]  ( .D(\w0[4][84] ), .CLK(clk), .RST(rst), .Q(state[84])
         );
  DFF \state_reg[92]  ( .D(\w0[4][92] ), .CLK(clk), .RST(rst), .Q(state[92])
         );
  DFF \state_reg[76]  ( .D(\w0[4][76] ), .CLK(clk), .RST(rst), .Q(state[76])
         );
  DFF \state_reg[68]  ( .D(\w0[4][68] ), .CLK(clk), .RST(rst), .Q(state[68])
         );
  DFF \state_reg[85]  ( .D(\w0[4][85] ), .CLK(clk), .RST(rst), .Q(state[85])
         );
  DFF \state_reg[93]  ( .D(\w0[4][93] ), .CLK(clk), .RST(rst), .Q(state[93])
         );
  DFF \state_reg[86]  ( .D(\w0[4][86] ), .CLK(clk), .RST(rst), .Q(state[86])
         );
  DFF \state_reg[69]  ( .D(\w0[4][69] ), .CLK(clk), .RST(rst), .Q(state[69])
         );
  DFF \state_reg[77]  ( .D(\w0[4][77] ), .CLK(clk), .RST(rst), .Q(state[77])
         );
  DFF \state_reg[94]  ( .D(\w0[4][94] ), .CLK(clk), .RST(rst), .Q(state[94])
         );
  DFF \state_reg[78]  ( .D(\w0[4][78] ), .CLK(clk), .RST(rst), .Q(state[78])
         );
  DFF \state_reg[70]  ( .D(\w0[4][70] ), .CLK(clk), .RST(rst), .Q(state[70])
         );
  DFF \state_reg[87]  ( .D(\w0[4][87] ), .CLK(clk), .RST(rst), .Q(state[87])
         );
  DFF \state_reg[79]  ( .D(\w0[4][79] ), .CLK(clk), .RST(rst), .Q(state[79])
         );
  DFF \state_reg[95]  ( .D(\w0[4][95] ), .CLK(clk), .RST(rst), .Q(state[95])
         );
  DFF \state_reg[32]  ( .D(\w0[4][32] ), .CLK(clk), .RST(rst), .Q(state[32])
         );
  DFF \state_reg[56]  ( .D(\w0[4][56] ), .CLK(clk), .RST(rst), .Q(state[56])
         );
  DFF \state_reg[47]  ( .D(\w0[4][47] ), .CLK(clk), .RST(rst), .Q(state[47])
         );
  DFF \state_reg[57]  ( .D(\w0[4][57] ), .CLK(clk), .RST(rst), .Q(state[57])
         );
  DFF \state_reg[48]  ( .D(\w0[4][48] ), .CLK(clk), .RST(rst), .Q(state[48])
         );
  DFF \state_reg[33]  ( .D(\w0[4][33] ), .CLK(clk), .RST(rst), .Q(state[33])
         );
  DFF \state_reg[40]  ( .D(\w0[4][40] ), .CLK(clk), .RST(rst), .Q(state[40])
         );
  DFF \state_reg[58]  ( .D(\w0[4][58] ), .CLK(clk), .RST(rst), .Q(state[58])
         );
  DFF \state_reg[49]  ( .D(\w0[4][49] ), .CLK(clk), .RST(rst), .Q(state[49])
         );
  DFF \state_reg[34]  ( .D(\w0[4][34] ), .CLK(clk), .RST(rst), .Q(state[34])
         );
  DFF \state_reg[41]  ( .D(\w0[4][41] ), .CLK(clk), .RST(rst), .Q(state[41])
         );
  DFF \state_reg[50]  ( .D(\w0[4][50] ), .CLK(clk), .RST(rst), .Q(state[50])
         );
  DFF \state_reg[59]  ( .D(\w0[4][59] ), .CLK(clk), .RST(rst), .Q(state[59])
         );
  DFF \state_reg[35]  ( .D(\w0[4][35] ), .CLK(clk), .RST(rst), .Q(state[35])
         );
  DFF \state_reg[42]  ( .D(\w0[4][42] ), .CLK(clk), .RST(rst), .Q(state[42])
         );
  DFF \state_reg[60]  ( .D(\w0[4][60] ), .CLK(clk), .RST(rst), .Q(state[60])
         );
  DFF \state_reg[36]  ( .D(\w0[4][36] ), .CLK(clk), .RST(rst), .Q(state[36])
         );
  DFF \state_reg[51]  ( .D(\w0[4][51] ), .CLK(clk), .RST(rst), .Q(state[51])
         );
  DFF \state_reg[43]  ( .D(\w0[4][43] ), .CLK(clk), .RST(rst), .Q(state[43])
         );
  DFF \state_reg[61]  ( .D(\w0[4][61] ), .CLK(clk), .RST(rst), .Q(state[61])
         );
  DFF \state_reg[37]  ( .D(\w0[4][37] ), .CLK(clk), .RST(rst), .Q(state[37])
         );
  DFF \state_reg[52]  ( .D(\w0[4][52] ), .CLK(clk), .RST(rst), .Q(state[52])
         );
  DFF \state_reg[44]  ( .D(\w0[4][44] ), .CLK(clk), .RST(rst), .Q(state[44])
         );
  DFF \state_reg[53]  ( .D(\w0[4][53] ), .CLK(clk), .RST(rst), .Q(state[53])
         );
  DFF \state_reg[62]  ( .D(\w0[4][62] ), .CLK(clk), .RST(rst), .Q(state[62])
         );
  DFF \state_reg[38]  ( .D(\w0[4][38] ), .CLK(clk), .RST(rst), .Q(state[38])
         );
  DFF \state_reg[45]  ( .D(\w0[4][45] ), .CLK(clk), .RST(rst), .Q(state[45])
         );
  DFF \state_reg[63]  ( .D(\w0[4][63] ), .CLK(clk), .RST(rst), .Q(state[63])
         );
  DFF \state_reg[39]  ( .D(\w0[4][39] ), .CLK(clk), .RST(rst), .Q(state[39])
         );
  DFF \state_reg[55]  ( .D(\w0[4][55] ), .CLK(clk), .RST(rst), .Q(state[55])
         );
  DFF \state_reg[54]  ( .D(\w0[4][54] ), .CLK(clk), .RST(rst), .Q(state[54])
         );
  DFF \state_reg[46]  ( .D(\w0[4][46] ), .CLK(clk), .RST(rst), .Q(state[46])
         );
  DFF \state_reg[8]  ( .D(\w0[4][8] ), .CLK(clk), .RST(rst), .Q(state[8]) );
  DFF \state_reg[23]  ( .D(\w0[4][23] ), .CLK(clk), .RST(rst), .Q(state[23])
         );
  DFF \state_reg[1]  ( .D(\w0[4][1] ), .CLK(clk), .RST(rst), .Q(state[1]) );
  DFF \state_reg[16]  ( .D(\w0[4][16] ), .CLK(clk), .RST(rst), .Q(state[16])
         );
  DFF \state_reg[24]  ( .D(\w0[4][24] ), .CLK(clk), .RST(rst), .Q(state[24])
         );
  DFF \state_reg[9]  ( .D(\w0[4][9] ), .CLK(clk), .RST(rst), .Q(state[9]) );
  DFF \state_reg[10]  ( .D(\w0[4][10] ), .CLK(clk), .RST(rst), .Q(state[10])
         );
  DFF \state_reg[2]  ( .D(\w0[4][2] ), .CLK(clk), .RST(rst), .Q(state[2]) );
  DFF \state_reg[17]  ( .D(\w0[4][17] ), .CLK(clk), .RST(rst), .Q(state[17])
         );
  DFF \state_reg[25]  ( .D(\w0[4][25] ), .CLK(clk), .RST(rst), .Q(state[25])
         );
  DFF \state_reg[11]  ( .D(\w0[4][11] ), .CLK(clk), .RST(rst), .Q(state[11])
         );
  DFF \state_reg[3]  ( .D(\w0[4][3] ), .CLK(clk), .RST(rst), .Q(state[3]) );
  DFF \state_reg[18]  ( .D(\w0[4][18] ), .CLK(clk), .RST(rst), .Q(state[18])
         );
  DFF \state_reg[26]  ( .D(\w0[4][26] ), .CLK(clk), .RST(rst), .Q(state[26])
         );
  DFF \state_reg[12]  ( .D(\w0[4][12] ), .CLK(clk), .RST(rst), .Q(state[12])
         );
  DFF \state_reg[27]  ( .D(\w0[4][27] ), .CLK(clk), .RST(rst), .Q(state[27])
         );
  DFF \state_reg[19]  ( .D(\w0[4][19] ), .CLK(clk), .RST(rst), .Q(state[19])
         );
  DFF \state_reg[4]  ( .D(\w0[4][4] ), .CLK(clk), .RST(rst), .Q(state[4]) );
  DFF \state_reg[13]  ( .D(\w0[4][13] ), .CLK(clk), .RST(rst), .Q(state[13])
         );
  DFF \state_reg[28]  ( .D(\w0[4][28] ), .CLK(clk), .RST(rst), .Q(state[28])
         );
  DFF \state_reg[20]  ( .D(\w0[4][20] ), .CLK(clk), .RST(rst), .Q(state[20])
         );
  DFF \state_reg[5]  ( .D(\w0[4][5] ), .CLK(clk), .RST(rst), .Q(state[5]) );
  DFF \state_reg[14]  ( .D(\w0[4][14] ), .CLK(clk), .RST(rst), .Q(state[14])
         );
  DFF \state_reg[6]  ( .D(\w0[4][6] ), .CLK(clk), .RST(rst), .Q(state[6]) );
  DFF \state_reg[21]  ( .D(\w0[4][21] ), .CLK(clk), .RST(rst), .Q(state[21])
         );
  DFF \state_reg[29]  ( .D(\w0[4][29] ), .CLK(clk), .RST(rst), .Q(state[29])
         );
  DFF \state_reg[15]  ( .D(\w0[4][15] ), .CLK(clk), .RST(rst), .Q(state[15])
         );
  DFF \state_reg[30]  ( .D(\w0[4][30] ), .CLK(clk), .RST(rst), .Q(state[30])
         );
  DFF \state_reg[22]  ( .D(\w0[4][22] ), .CLK(clk), .RST(rst), .Q(state[22])
         );
  DFF \state_reg[7]  ( .D(\w0[4][7] ), .CLK(clk), .RST(rst), .Q(state[7]) );
  DFF \state_reg[31]  ( .D(\w0[4][31] ), .CLK(clk), .RST(rst), .Q(state[31])
         );
  DFF \state_reg[127]  ( .D(\w0[4][127] ), .CLK(clk), .RST(rst), .Q(state[127]) );
  DFF \state_reg[104]  ( .D(\w0[4][104] ), .CLK(clk), .RST(rst), .Q(state[104]) );
  DFF \state_reg[112]  ( .D(\w0[4][112] ), .CLK(clk), .RST(rst), .Q(state[112]) );
  DFF \state_reg[96]  ( .D(\w0[4][96] ), .CLK(clk), .RST(rst), .Q(state[96])
         );
  DFF \state_reg[113]  ( .D(\w0[4][113] ), .CLK(clk), .RST(rst), .Q(state[113]) );
  DFF \state_reg[105]  ( .D(\w0[4][105] ), .CLK(clk), .RST(rst), .Q(state[105]) );
  DFF \state_reg[120]  ( .D(\w0[4][120] ), .CLK(clk), .RST(rst), .Q(state[120]) );
  DFF \state_reg[97]  ( .D(\w0[4][97] ), .CLK(clk), .RST(rst), .Q(state[97])
         );
  DFF \state_reg[114]  ( .D(\w0[4][114] ), .CLK(clk), .RST(rst), .Q(state[114]) );
  DFF \state_reg[106]  ( .D(\w0[4][106] ), .CLK(clk), .RST(rst), .Q(state[106]) );
  DFF \state_reg[121]  ( .D(\w0[4][121] ), .CLK(clk), .RST(rst), .Q(state[121]) );
  DFF \state_reg[98]  ( .D(\w0[4][98] ), .CLK(clk), .RST(rst), .Q(state[98])
         );
  DFF \state_reg[115]  ( .D(\w0[4][115] ), .CLK(clk), .RST(rst), .Q(state[115]) );
  DFF \state_reg[107]  ( .D(\w0[4][107] ), .CLK(clk), .RST(rst), .Q(state[107]) );
  DFF \state_reg[122]  ( .D(\w0[4][122] ), .CLK(clk), .RST(rst), .Q(state[122]) );
  DFF \state_reg[116]  ( .D(\w0[4][116] ), .CLK(clk), .RST(rst), .Q(state[116]) );
  DFF \state_reg[108]  ( .D(\w0[4][108] ), .CLK(clk), .RST(rst), .Q(state[108]) );
  DFF \state_reg[99]  ( .D(\w0[4][99] ), .CLK(clk), .RST(rst), .Q(state[99])
         );
  DFF \state_reg[123]  ( .D(\w0[4][123] ), .CLK(clk), .RST(rst), .Q(state[123]) );
  DFF \state_reg[124]  ( .D(\w0[4][124] ), .CLK(clk), .RST(rst), .Q(state[124]) );
  DFF \state_reg[100]  ( .D(\w0[4][100] ), .CLK(clk), .RST(rst), .Q(state[100]) );
  DFF \state_reg[117]  ( .D(\w0[4][117] ), .CLK(clk), .RST(rst), .Q(state[117]) );
  DFF \state_reg[109]  ( .D(\w0[4][109] ), .CLK(clk), .RST(rst), .Q(state[109]) );
  DFF \state_reg[118]  ( .D(\w0[4][118] ), .CLK(clk), .RST(rst), .Q(state[118]) );
  DFF \state_reg[110]  ( .D(\w0[4][110] ), .CLK(clk), .RST(rst), .Q(state[110]) );
  DFF \state_reg[101]  ( .D(\w0[4][101] ), .CLK(clk), .RST(rst), .Q(state[101]) );
  DFF \state_reg[125]  ( .D(\w0[4][125] ), .CLK(clk), .RST(rst), .Q(state[125]) );
  DFF \state_reg[103]  ( .D(\w0[4][103] ), .CLK(clk), .RST(rst), .Q(state[103]) );
  DFF \state_reg[126]  ( .D(\w0[4][126] ), .CLK(clk), .RST(rst), .Q(state[126]) );
  DFF \state_reg[102]  ( .D(\w0[4][102] ), .CLK(clk), .RST(rst), .Q(state[102]) );
  DFF \state_reg[119]  ( .D(\w0[4][119] ), .CLK(clk), .RST(rst), .Q(state[119]) );
  DFF \state_reg[111]  ( .D(\w0[4][111] ), .CLK(clk), .RST(rst), .Q(state[111]) );
  XOR U2851 ( .A(key[512]), .B(\w3[4][0] ), .Z(out[0]) );
  XOR U2852 ( .A(key[612]), .B(\w3[4][100] ), .Z(out[100]) );
  XOR U2853 ( .A(key[613]), .B(\w3[4][101] ), .Z(out[101]) );
  XOR U2854 ( .A(key[614]), .B(\w3[4][102] ), .Z(out[102]) );
  XOR U2855 ( .A(key[615]), .B(\w3[4][103] ), .Z(out[103]) );
  XOR U2856 ( .A(key[616]), .B(\w3[4][104] ), .Z(out[104]) );
  XOR U2857 ( .A(key[617]), .B(\w3[4][105] ), .Z(out[105]) );
  XOR U2858 ( .A(key[618]), .B(\w3[4][106] ), .Z(out[106]) );
  XOR U2859 ( .A(key[619]), .B(\w3[4][107] ), .Z(out[107]) );
  XOR U2860 ( .A(key[620]), .B(\w3[4][108] ), .Z(out[108]) );
  XOR U2861 ( .A(key[621]), .B(\w3[4][109] ), .Z(out[109]) );
  XOR U2862 ( .A(key[522]), .B(\w3[4][10] ), .Z(out[10]) );
  XOR U2863 ( .A(key[622]), .B(\w3[4][110] ), .Z(out[110]) );
  XOR U2864 ( .A(key[623]), .B(\w3[4][111] ), .Z(out[111]) );
  XOR U2865 ( .A(key[624]), .B(\w3[4][112] ), .Z(out[112]) );
  XOR U2866 ( .A(key[625]), .B(\w3[4][113] ), .Z(out[113]) );
  XOR U2867 ( .A(key[626]), .B(\w3[4][114] ), .Z(out[114]) );
  XOR U2868 ( .A(key[627]), .B(\w3[4][115] ), .Z(out[115]) );
  XOR U2869 ( .A(key[628]), .B(\w3[4][116] ), .Z(out[116]) );
  XOR U2870 ( .A(key[629]), .B(\w3[4][117] ), .Z(out[117]) );
  XOR U2871 ( .A(key[630]), .B(\w3[4][118] ), .Z(out[118]) );
  XOR U2872 ( .A(key[631]), .B(\w3[4][119] ), .Z(out[119]) );
  XOR U2873 ( .A(key[523]), .B(\w3[4][11] ), .Z(out[11]) );
  XOR U2874 ( .A(key[632]), .B(\w3[4][120] ), .Z(out[120]) );
  XOR U2875 ( .A(key[633]), .B(\w3[4][121] ), .Z(out[121]) );
  XOR U2876 ( .A(key[634]), .B(\w3[4][122] ), .Z(out[122]) );
  XOR U2877 ( .A(key[635]), .B(\w3[4][123] ), .Z(out[123]) );
  XOR U2878 ( .A(key[636]), .B(\w3[4][124] ), .Z(out[124]) );
  XOR U2879 ( .A(key[637]), .B(\w3[4][125] ), .Z(out[125]) );
  XOR U2880 ( .A(key[638]), .B(\w3[4][126] ), .Z(out[126]) );
  XOR U2881 ( .A(key[639]), .B(\w3[4][127] ), .Z(out[127]) );
  XOR U2882 ( .A(key[524]), .B(\w3[4][12] ), .Z(out[12]) );
  XOR U2883 ( .A(key[525]), .B(\w3[4][13] ), .Z(out[13]) );
  XOR U2884 ( .A(key[526]), .B(\w3[4][14] ), .Z(out[14]) );
  XOR U2885 ( .A(key[527]), .B(\w3[4][15] ), .Z(out[15]) );
  XOR U2886 ( .A(key[528]), .B(\w3[4][16] ), .Z(out[16]) );
  XOR U2887 ( .A(key[529]), .B(\w3[4][17] ), .Z(out[17]) );
  XOR U2888 ( .A(key[530]), .B(\w3[4][18] ), .Z(out[18]) );
  XOR U2889 ( .A(key[531]), .B(\w3[4][19] ), .Z(out[19]) );
  XOR U2890 ( .A(key[513]), .B(\w3[4][1] ), .Z(out[1]) );
  XOR U2891 ( .A(key[532]), .B(\w3[4][20] ), .Z(out[20]) );
  XOR U2892 ( .A(key[533]), .B(\w3[4][21] ), .Z(out[21]) );
  XOR U2893 ( .A(key[534]), .B(\w3[4][22] ), .Z(out[22]) );
  XOR U2894 ( .A(key[535]), .B(\w3[4][23] ), .Z(out[23]) );
  XOR U2895 ( .A(key[536]), .B(\w3[4][24] ), .Z(out[24]) );
  XOR U2896 ( .A(key[537]), .B(\w3[4][25] ), .Z(out[25]) );
  XOR U2897 ( .A(key[538]), .B(\w3[4][26] ), .Z(out[26]) );
  XOR U2898 ( .A(key[539]), .B(\w3[4][27] ), .Z(out[27]) );
  XOR U2899 ( .A(key[540]), .B(\w3[4][28] ), .Z(out[28]) );
  XOR U2900 ( .A(key[541]), .B(\w3[4][29] ), .Z(out[29]) );
  XOR U2901 ( .A(key[514]), .B(\w3[4][2] ), .Z(out[2]) );
  XOR U2902 ( .A(key[542]), .B(\w3[4][30] ), .Z(out[30]) );
  XOR U2903 ( .A(key[543]), .B(\w3[4][31] ), .Z(out[31]) );
  XOR U2904 ( .A(key[544]), .B(\w3[4][32] ), .Z(out[32]) );
  XOR U2905 ( .A(key[545]), .B(\w3[4][33] ), .Z(out[33]) );
  XOR U2906 ( .A(key[546]), .B(\w3[4][34] ), .Z(out[34]) );
  XOR U2907 ( .A(key[547]), .B(\w3[4][35] ), .Z(out[35]) );
  XOR U2908 ( .A(key[548]), .B(\w3[4][36] ), .Z(out[36]) );
  XOR U2909 ( .A(key[549]), .B(\w3[4][37] ), .Z(out[37]) );
  XOR U2910 ( .A(key[550]), .B(\w3[4][38] ), .Z(out[38]) );
  XOR U2911 ( .A(key[551]), .B(\w3[4][39] ), .Z(out[39]) );
  XOR U2912 ( .A(key[515]), .B(\w3[4][3] ), .Z(out[3]) );
  XOR U2913 ( .A(key[552]), .B(\w3[4][40] ), .Z(out[40]) );
  XOR U2914 ( .A(key[553]), .B(\w3[4][41] ), .Z(out[41]) );
  XOR U2915 ( .A(key[554]), .B(\w3[4][42] ), .Z(out[42]) );
  XOR U2916 ( .A(key[555]), .B(\w3[4][43] ), .Z(out[43]) );
  XOR U2917 ( .A(key[556]), .B(\w3[4][44] ), .Z(out[44]) );
  XOR U2918 ( .A(key[557]), .B(\w3[4][45] ), .Z(out[45]) );
  XOR U2919 ( .A(key[558]), .B(\w3[4][46] ), .Z(out[46]) );
  XOR U2920 ( .A(key[559]), .B(\w3[4][47] ), .Z(out[47]) );
  XOR U2921 ( .A(key[560]), .B(\w3[4][48] ), .Z(out[48]) );
  XOR U2922 ( .A(key[561]), .B(\w3[4][49] ), .Z(out[49]) );
  XOR U2923 ( .A(key[516]), .B(\w3[4][4] ), .Z(out[4]) );
  XOR U2924 ( .A(key[562]), .B(\w3[4][50] ), .Z(out[50]) );
  XOR U2925 ( .A(key[563]), .B(\w3[4][51] ), .Z(out[51]) );
  XOR U2926 ( .A(key[564]), .B(\w3[4][52] ), .Z(out[52]) );
  XOR U2927 ( .A(key[565]), .B(\w3[4][53] ), .Z(out[53]) );
  XOR U2928 ( .A(key[566]), .B(\w3[4][54] ), .Z(out[54]) );
  XOR U2929 ( .A(key[567]), .B(\w3[4][55] ), .Z(out[55]) );
  XOR U2930 ( .A(key[568]), .B(\w3[4][56] ), .Z(out[56]) );
  XOR U2931 ( .A(key[569]), .B(\w3[4][57] ), .Z(out[57]) );
  XOR U2932 ( .A(key[570]), .B(\w3[4][58] ), .Z(out[58]) );
  XOR U2933 ( .A(key[571]), .B(\w3[4][59] ), .Z(out[59]) );
  XOR U2934 ( .A(key[517]), .B(\w3[4][5] ), .Z(out[5]) );
  XOR U2935 ( .A(key[572]), .B(\w3[4][60] ), .Z(out[60]) );
  XOR U2936 ( .A(key[573]), .B(\w3[4][61] ), .Z(out[61]) );
  XOR U2937 ( .A(key[574]), .B(\w3[4][62] ), .Z(out[62]) );
  XOR U2938 ( .A(key[575]), .B(\w3[4][63] ), .Z(out[63]) );
  XOR U2939 ( .A(key[576]), .B(\w3[4][64] ), .Z(out[64]) );
  XOR U2940 ( .A(key[577]), .B(\w3[4][65] ), .Z(out[65]) );
  XOR U2941 ( .A(key[578]), .B(\w3[4][66] ), .Z(out[66]) );
  XOR U2942 ( .A(key[579]), .B(\w3[4][67] ), .Z(out[67]) );
  XOR U2943 ( .A(key[580]), .B(\w3[4][68] ), .Z(out[68]) );
  XOR U2944 ( .A(key[581]), .B(\w3[4][69] ), .Z(out[69]) );
  XOR U2945 ( .A(key[518]), .B(\w3[4][6] ), .Z(out[6]) );
  XOR U2946 ( .A(key[582]), .B(\w3[4][70] ), .Z(out[70]) );
  XOR U2947 ( .A(key[583]), .B(\w3[4][71] ), .Z(out[71]) );
  XOR U2948 ( .A(key[584]), .B(\w3[4][72] ), .Z(out[72]) );
  XOR U2949 ( .A(key[585]), .B(\w3[4][73] ), .Z(out[73]) );
  XOR U2950 ( .A(key[586]), .B(\w3[4][74] ), .Z(out[74]) );
  XOR U2951 ( .A(key[587]), .B(\w3[4][75] ), .Z(out[75]) );
  XOR U2952 ( .A(key[588]), .B(\w3[4][76] ), .Z(out[76]) );
  XOR U2953 ( .A(key[589]), .B(\w3[4][77] ), .Z(out[77]) );
  XOR U2954 ( .A(key[590]), .B(\w3[4][78] ), .Z(out[78]) );
  XOR U2955 ( .A(key[591]), .B(\w3[4][79] ), .Z(out[79]) );
  XOR U2956 ( .A(key[519]), .B(\w3[4][7] ), .Z(out[7]) );
  XOR U2957 ( .A(key[592]), .B(\w3[4][80] ), .Z(out[80]) );
  XOR U2958 ( .A(key[593]), .B(\w3[4][81] ), .Z(out[81]) );
  XOR U2959 ( .A(key[594]), .B(\w3[4][82] ), .Z(out[82]) );
  XOR U2960 ( .A(key[595]), .B(\w3[4][83] ), .Z(out[83]) );
  XOR U2961 ( .A(key[596]), .B(\w3[4][84] ), .Z(out[84]) );
  XOR U2962 ( .A(key[597]), .B(\w3[4][85] ), .Z(out[85]) );
  XOR U2963 ( .A(key[598]), .B(\w3[4][86] ), .Z(out[86]) );
  XOR U2964 ( .A(key[599]), .B(\w3[4][87] ), .Z(out[87]) );
  XOR U2965 ( .A(key[600]), .B(\w3[4][88] ), .Z(out[88]) );
  XOR U2966 ( .A(key[601]), .B(\w3[4][89] ), .Z(out[89]) );
  XOR U2967 ( .A(key[520]), .B(\w3[4][8] ), .Z(out[8]) );
  XOR U2968 ( .A(key[602]), .B(\w3[4][90] ), .Z(out[90]) );
  XOR U2969 ( .A(key[603]), .B(\w3[4][91] ), .Z(out[91]) );
  XOR U2970 ( .A(key[604]), .B(\w3[4][92] ), .Z(out[92]) );
  XOR U2971 ( .A(key[605]), .B(\w3[4][93] ), .Z(out[93]) );
  XOR U2972 ( .A(key[606]), .B(\w3[4][94] ), .Z(out[94]) );
  XOR U2973 ( .A(key[607]), .B(\w3[4][95] ), .Z(out[95]) );
  XOR U2974 ( .A(key[608]), .B(\w3[4][96] ), .Z(out[96]) );
  XOR U2975 ( .A(key[609]), .B(\w3[4][97] ), .Z(out[97]) );
  XOR U2976 ( .A(key[610]), .B(\w3[4][98] ), .Z(out[98]) );
  XOR U2977 ( .A(key[611]), .B(\w3[4][99] ), .Z(out[99]) );
  XOR U2978 ( .A(key[521]), .B(\w3[4][9] ), .Z(out[9]) );
  XOR U2979 ( .A(\w3[3][1] ), .B(\w3[3][25] ), .Z(n2246) );
  XOR U2980 ( .A(\w3[3][16] ), .B(\w3[3][24] ), .Z(n2213) );
  XNOR U2981 ( .A(n2246), .B(n2213), .Z(n1953) );
  XNOR U2982 ( .A(\w3[3][8] ), .B(n1953), .Z(\w0[4][0] ) );
  XOR U2983 ( .A(\w3[3][96] ), .B(\w3[3][101] ), .Z(n1971) );
  XOR U2984 ( .A(\w3[3][108] ), .B(\w3[3][116] ), .Z(n1955) );
  XNOR U2985 ( .A(\w3[3][120] ), .B(\w3[3][125] ), .Z(n1954) );
  XNOR U2986 ( .A(n1955), .B(n1954), .Z(n2009) );
  XNOR U2987 ( .A(\w3[3][124] ), .B(n2009), .Z(n1956) );
  XNOR U2988 ( .A(n1971), .B(n1956), .Z(\w0[4][100] ) );
  XOR U2989 ( .A(\w3[3][102] ), .B(\w3[3][126] ), .Z(n1977) );
  XOR U2990 ( .A(\w3[3][109] ), .B(\w3[3][117] ), .Z(n2012) );
  XNOR U2991 ( .A(\w3[3][125] ), .B(n2012), .Z(n1957) );
  XNOR U2992 ( .A(n1977), .B(n1957), .Z(\w0[4][101] ) );
  XOR U2993 ( .A(\w3[3][96] ), .B(\w3[3][103] ), .Z(n1978) );
  XOR U2994 ( .A(\w3[3][110] ), .B(\w3[3][118] ), .Z(n1988) );
  XNOR U2995 ( .A(\w3[3][120] ), .B(\w3[3][127] ), .Z(n1959) );
  XNOR U2996 ( .A(n1988), .B(n1959), .Z(n2015) );
  XNOR U2997 ( .A(\w3[3][126] ), .B(n2015), .Z(n1958) );
  XNOR U2998 ( .A(n1978), .B(n1958), .Z(\w0[4][102] ) );
  XNOR U2999 ( .A(\w3[3][111] ), .B(\w3[3][119] ), .Z(n2019) );
  XNOR U3000 ( .A(\w3[3][96] ), .B(n1959), .Z(n1960) );
  XNOR U3001 ( .A(n2019), .B(n1960), .Z(\w0[4][103] ) );
  XOR U3002 ( .A(\w3[3][120] ), .B(\w3[3][112] ), .Z(n2235) );
  XOR U3003 ( .A(n2235), .B(\w3[3][97] ), .Z(n1962) );
  XNOR U3004 ( .A(\w3[3][96] ), .B(\w3[3][105] ), .Z(n1961) );
  XNOR U3005 ( .A(n1962), .B(n1961), .Z(\w0[4][104] ) );
  XOR U3006 ( .A(\w3[3][97] ), .B(\w3[3][121] ), .Z(n2234) );
  XOR U3007 ( .A(\w3[3][98] ), .B(n2234), .Z(n1964) );
  XNOR U3008 ( .A(\w3[3][106] ), .B(\w3[3][113] ), .Z(n1963) );
  XNOR U3009 ( .A(n1964), .B(n1963), .Z(\w0[4][105] ) );
  XOR U3010 ( .A(\w3[3][114] ), .B(\w3[3][122] ), .Z(n2240) );
  XOR U3011 ( .A(n2240), .B(\w3[3][99] ), .Z(n1966) );
  XNOR U3012 ( .A(\w3[3][98] ), .B(\w3[3][107] ), .Z(n1965) );
  XNOR U3013 ( .A(n1966), .B(n1965), .Z(\w0[4][106] ) );
  XOR U3014 ( .A(\w3[3][99] ), .B(\w3[3][123] ), .Z(n2242) );
  XNOR U3015 ( .A(\w3[3][108] ), .B(n2242), .Z(n1967) );
  XNOR U3016 ( .A(\w3[3][104] ), .B(n1967), .Z(n1984) );
  XOR U3017 ( .A(\w3[3][96] ), .B(\w3[3][100] ), .Z(n2243) );
  XNOR U3018 ( .A(\w3[3][115] ), .B(n2243), .Z(n1968) );
  XNOR U3019 ( .A(n1984), .B(n1968), .Z(\w0[4][107] ) );
  XOR U3020 ( .A(\w3[3][100] ), .B(\w3[3][104] ), .Z(n1970) );
  XNOR U3021 ( .A(\w3[3][124] ), .B(\w3[3][109] ), .Z(n1969) );
  XNOR U3022 ( .A(n1970), .B(n1969), .Z(n1986) );
  XNOR U3023 ( .A(\w3[3][116] ), .B(n1971), .Z(n1972) );
  XNOR U3024 ( .A(n1986), .B(n1972), .Z(\w0[4][108] ) );
  XOR U3025 ( .A(\w3[3][125] ), .B(\w3[3][101] ), .Z(n1990) );
  XOR U3026 ( .A(\w3[3][110] ), .B(n1990), .Z(n1974) );
  XNOR U3027 ( .A(\w3[3][117] ), .B(\w3[3][102] ), .Z(n1973) );
  XNOR U3028 ( .A(n1974), .B(n1973), .Z(\w0[4][109] ) );
  XOR U3029 ( .A(\w3[3][2] ), .B(\w3[3][26] ), .Z(n2032) );
  XOR U3030 ( .A(\w3[3][3] ), .B(n2032), .Z(n1976) );
  XNOR U3031 ( .A(\w3[3][11] ), .B(\w3[3][18] ), .Z(n1975) );
  XNOR U3032 ( .A(n1976), .B(n1975), .Z(\w0[4][10] ) );
  XNOR U3033 ( .A(\w3[3][111] ), .B(\w3[3][104] ), .Z(n1995) );
  XNOR U3034 ( .A(n1977), .B(n1995), .Z(n1991) );
  XNOR U3035 ( .A(\w3[3][118] ), .B(n1978), .Z(n1979) );
  XNOR U3036 ( .A(n1991), .B(n1979), .Z(\w0[4][110] ) );
  XOR U3037 ( .A(\w3[3][127] ), .B(\w3[3][103] ), .Z(n1993) );
  XOR U3038 ( .A(\w3[3][96] ), .B(\w3[3][104] ), .Z(n1998) );
  XNOR U3039 ( .A(\w3[3][119] ), .B(n1998), .Z(n1980) );
  XNOR U3040 ( .A(n1993), .B(n1980), .Z(\w0[4][111] ) );
  XOR U3041 ( .A(\w3[3][105] ), .B(\w3[3][113] ), .Z(n2001) );
  XNOR U3042 ( .A(\w3[3][120] ), .B(n1998), .Z(n1981) );
  XNOR U3043 ( .A(n2001), .B(n1981), .Z(\w0[4][112] ) );
  XOR U3044 ( .A(\w3[3][106] ), .B(\w3[3][114] ), .Z(n2002) );
  XNOR U3045 ( .A(\w3[3][105] ), .B(n2234), .Z(n1982) );
  XNOR U3046 ( .A(n2002), .B(n1982), .Z(\w0[4][113] ) );
  XOR U3047 ( .A(\w3[3][98] ), .B(\w3[3][122] ), .Z(n2237) );
  XOR U3048 ( .A(\w3[3][107] ), .B(\w3[3][115] ), .Z(n2006) );
  XNOR U3049 ( .A(\w3[3][106] ), .B(n2006), .Z(n1983) );
  XNOR U3050 ( .A(n2237), .B(n1983), .Z(\w0[4][114] ) );
  XOR U3051 ( .A(\w3[3][116] ), .B(\w3[3][112] ), .Z(n2007) );
  XNOR U3052 ( .A(\w3[3][107] ), .B(n1984), .Z(n1985) );
  XNOR U3053 ( .A(n2007), .B(n1985), .Z(\w0[4][115] ) );
  XOR U3054 ( .A(\w3[3][117] ), .B(\w3[3][112] ), .Z(n2011) );
  XNOR U3055 ( .A(\w3[3][108] ), .B(n1986), .Z(n1987) );
  XNOR U3056 ( .A(n2011), .B(n1987), .Z(\w0[4][116] ) );
  XNOR U3057 ( .A(\w3[3][109] ), .B(n1988), .Z(n1989) );
  XNOR U3058 ( .A(n1990), .B(n1989), .Z(\w0[4][117] ) );
  XOR U3059 ( .A(\w3[3][119] ), .B(\w3[3][112] ), .Z(n2017) );
  XNOR U3060 ( .A(\w3[3][110] ), .B(n1991), .Z(n1992) );
  XNOR U3061 ( .A(n2017), .B(n1992), .Z(\w0[4][118] ) );
  XOR U3062 ( .A(\w3[3][112] ), .B(n1993), .Z(n1994) );
  XNOR U3063 ( .A(n1995), .B(n1994), .Z(\w0[4][119] ) );
  XOR U3064 ( .A(\w3[3][3] ), .B(\w3[3][27] ), .Z(n2061) );
  XNOR U3065 ( .A(\w3[3][8] ), .B(\w3[3][12] ), .Z(n1996) );
  XNOR U3066 ( .A(n2061), .B(n1996), .Z(n2030) );
  XOR U3067 ( .A(\w3[3][0] ), .B(\w3[3][4] ), .Z(n2080) );
  XNOR U3068 ( .A(\w3[3][19] ), .B(n2080), .Z(n1997) );
  XNOR U3069 ( .A(n2030), .B(n1997), .Z(\w0[4][11] ) );
  XOR U3070 ( .A(\w3[3][113] ), .B(\w3[3][121] ), .Z(n2239) );
  XNOR U3071 ( .A(\w3[3][112] ), .B(n1998), .Z(n1999) );
  XNOR U3072 ( .A(n2239), .B(n1999), .Z(\w0[4][120] ) );
  XNOR U3073 ( .A(\w3[3][97] ), .B(n2240), .Z(n2000) );
  XNOR U3074 ( .A(n2001), .B(n2000), .Z(\w0[4][121] ) );
  XOR U3075 ( .A(\w3[3][123] ), .B(n2002), .Z(n2004) );
  XNOR U3076 ( .A(\w3[3][98] ), .B(\w3[3][115] ), .Z(n2003) );
  XNOR U3077 ( .A(n2004), .B(n2003), .Z(\w0[4][122] ) );
  XNOR U3078 ( .A(\w3[3][124] ), .B(\w3[3][120] ), .Z(n2005) );
  XNOR U3079 ( .A(n2006), .B(n2005), .Z(n2245) );
  XNOR U3080 ( .A(\w3[3][99] ), .B(n2007), .Z(n2008) );
  XNOR U3081 ( .A(n2245), .B(n2008), .Z(\w0[4][123] ) );
  XNOR U3082 ( .A(n2009), .B(\w3[3][100] ), .Z(n2010) );
  XNOR U3083 ( .A(n2011), .B(n2010), .Z(\w0[4][124] ) );
  XOR U3084 ( .A(\w3[3][126] ), .B(\w3[3][118] ), .Z(n2014) );
  XNOR U3085 ( .A(\w3[3][101] ), .B(n2012), .Z(n2013) );
  XNOR U3086 ( .A(n2014), .B(n2013), .Z(\w0[4][125] ) );
  XNOR U3087 ( .A(\w3[3][102] ), .B(n2015), .Z(n2016) );
  XNOR U3088 ( .A(n2017), .B(n2016), .Z(\w0[4][126] ) );
  XOR U3089 ( .A(\w3[3][103] ), .B(n2235), .Z(n2018) );
  XNOR U3090 ( .A(n2019), .B(n2018), .Z(\w0[4][127] ) );
  XOR U3091 ( .A(\w3[3][13] ), .B(\w3[3][28] ), .Z(n2021) );
  XNOR U3092 ( .A(\w3[3][8] ), .B(\w3[3][4] ), .Z(n2020) );
  XNOR U3093 ( .A(n2021), .B(n2020), .Z(n2034) );
  XOR U3094 ( .A(\w3[3][0] ), .B(\w3[3][5] ), .Z(n2106) );
  XNOR U3095 ( .A(\w3[3][20] ), .B(n2106), .Z(n2022) );
  XNOR U3096 ( .A(n2034), .B(n2022), .Z(\w0[4][12] ) );
  XOR U3097 ( .A(\w3[3][5] ), .B(\w3[3][29] ), .Z(n2036) );
  XOR U3098 ( .A(\w3[3][6] ), .B(n2036), .Z(n2024) );
  XNOR U3099 ( .A(\w3[3][14] ), .B(\w3[3][21] ), .Z(n2023) );
  XNOR U3100 ( .A(n2024), .B(n2023), .Z(\w0[4][13] ) );
  XOR U3101 ( .A(\w3[3][6] ), .B(\w3[3][30] ), .Z(n2136) );
  XNOR U3102 ( .A(\w3[3][8] ), .B(\w3[3][15] ), .Z(n2042) );
  XNOR U3103 ( .A(n2136), .B(n2042), .Z(n2038) );
  XOR U3104 ( .A(\w3[3][0] ), .B(\w3[3][7] ), .Z(n2160) );
  XNOR U3105 ( .A(\w3[3][22] ), .B(n2160), .Z(n2025) );
  XNOR U3106 ( .A(n2038), .B(n2025), .Z(\w0[4][14] ) );
  XOR U3107 ( .A(\w3[3][7] ), .B(\w3[3][31] ), .Z(n2040) );
  XOR U3108 ( .A(\w3[3][8] ), .B(\w3[3][0] ), .Z(n2043) );
  XNOR U3109 ( .A(\w3[3][23] ), .B(n2043), .Z(n2026) );
  XNOR U3110 ( .A(n2040), .B(n2026), .Z(\w0[4][15] ) );
  XOR U3111 ( .A(\w3[3][17] ), .B(\w3[3][9] ), .Z(n2046) );
  XNOR U3112 ( .A(\w3[3][24] ), .B(n2043), .Z(n2027) );
  XNOR U3113 ( .A(n2046), .B(n2027), .Z(\w0[4][16] ) );
  XOR U3114 ( .A(\w3[3][18] ), .B(\w3[3][10] ), .Z(n2063) );
  XNOR U3115 ( .A(n2246), .B(\w3[3][9] ), .Z(n2028) );
  XNOR U3116 ( .A(n2063), .B(n2028), .Z(\w0[4][17] ) );
  XOR U3117 ( .A(\w3[3][11] ), .B(\w3[3][19] ), .Z(n2052) );
  XNOR U3118 ( .A(n2032), .B(\w3[3][10] ), .Z(n2029) );
  XNOR U3119 ( .A(n2052), .B(n2029), .Z(\w0[4][18] ) );
  XOR U3120 ( .A(\w3[3][16] ), .B(\w3[3][20] ), .Z(n2053) );
  XNOR U3121 ( .A(\w3[3][11] ), .B(n2030), .Z(n2031) );
  XNOR U3122 ( .A(n2053), .B(n2031), .Z(\w0[4][19] ) );
  XNOR U3123 ( .A(\w3[3][25] ), .B(n2032), .Z(n2033) );
  XNOR U3124 ( .A(n2046), .B(n2033), .Z(\w0[4][1] ) );
  XOR U3125 ( .A(\w3[3][16] ), .B(\w3[3][21] ), .Z(n2057) );
  XNOR U3126 ( .A(\w3[3][12] ), .B(n2034), .Z(n2035) );
  XNOR U3127 ( .A(n2057), .B(n2035), .Z(\w0[4][20] ) );
  XOR U3128 ( .A(\w3[3][14] ), .B(\w3[3][22] ), .Z(n2064) );
  XNOR U3129 ( .A(\w3[3][13] ), .B(n2036), .Z(n2037) );
  XNOR U3130 ( .A(n2064), .B(n2037), .Z(\w0[4][21] ) );
  XOR U3131 ( .A(\w3[3][16] ), .B(\w3[3][23] ), .Z(n2065) );
  XNOR U3132 ( .A(\w3[3][14] ), .B(n2038), .Z(n2039) );
  XNOR U3133 ( .A(n2065), .B(n2039), .Z(\w0[4][22] ) );
  XOR U3134 ( .A(\w3[3][16] ), .B(n2040), .Z(n2041) );
  XNOR U3135 ( .A(n2042), .B(n2041), .Z(\w0[4][23] ) );
  XOR U3136 ( .A(n2043), .B(\w3[3][17] ), .Z(n2045) );
  XNOR U3137 ( .A(\w3[3][25] ), .B(\w3[3][16] ), .Z(n2044) );
  XNOR U3138 ( .A(n2045), .B(n2044), .Z(\w0[4][24] ) );
  XOR U3139 ( .A(\w3[3][26] ), .B(n2046), .Z(n2048) );
  XNOR U3140 ( .A(\w3[3][1] ), .B(\w3[3][18] ), .Z(n2047) );
  XNOR U3141 ( .A(n2048), .B(n2047), .Z(\w0[4][25] ) );
  XOR U3142 ( .A(\w3[3][27] ), .B(n2063), .Z(n2050) );
  XNOR U3143 ( .A(\w3[3][2] ), .B(\w3[3][19] ), .Z(n2049) );
  XNOR U3144 ( .A(n2050), .B(n2049), .Z(\w0[4][26] ) );
  XNOR U3145 ( .A(\w3[3][24] ), .B(\w3[3][28] ), .Z(n2051) );
  XNOR U3146 ( .A(n2052), .B(n2051), .Z(n2082) );
  XNOR U3147 ( .A(\w3[3][3] ), .B(n2053), .Z(n2054) );
  XNOR U3148 ( .A(n2082), .B(n2054), .Z(\w0[4][27] ) );
  XOR U3149 ( .A(\w3[3][20] ), .B(\w3[3][29] ), .Z(n2056) );
  XNOR U3150 ( .A(\w3[3][24] ), .B(\w3[3][12] ), .Z(n2055) );
  XNOR U3151 ( .A(n2056), .B(n2055), .Z(n2108) );
  XNOR U3152 ( .A(\w3[3][4] ), .B(n2057), .Z(n2058) );
  XNOR U3153 ( .A(n2108), .B(n2058), .Z(\w0[4][28] ) );
  XOR U3154 ( .A(\w3[3][13] ), .B(\w3[3][21] ), .Z(n2138) );
  XOR U3155 ( .A(\w3[3][30] ), .B(n2138), .Z(n2060) );
  XNOR U3156 ( .A(\w3[3][5] ), .B(\w3[3][22] ), .Z(n2059) );
  XNOR U3157 ( .A(n2060), .B(n2059), .Z(\w0[4][29] ) );
  XNOR U3158 ( .A(\w3[3][26] ), .B(n2061), .Z(n2062) );
  XNOR U3159 ( .A(n2063), .B(n2062), .Z(\w0[4][2] ) );
  XNOR U3160 ( .A(\w3[3][24] ), .B(\w3[3][31] ), .Z(n2188) );
  XNOR U3161 ( .A(n2064), .B(n2188), .Z(n2162) );
  XNOR U3162 ( .A(\w3[3][6] ), .B(n2065), .Z(n2066) );
  XNOR U3163 ( .A(n2162), .B(n2066), .Z(\w0[4][30] ) );
  XOR U3164 ( .A(\w3[3][15] ), .B(\w3[3][23] ), .Z(n2186) );
  XNOR U3165 ( .A(n2213), .B(\w3[3][7] ), .Z(n2067) );
  XNOR U3166 ( .A(n2186), .B(n2067), .Z(\w0[4][31] ) );
  XOR U3167 ( .A(\w3[3][33] ), .B(\w3[3][57] ), .Z(n2104) );
  XOR U3168 ( .A(\w3[3][48] ), .B(\w3[3][56] ), .Z(n2148) );
  XNOR U3169 ( .A(n2148), .B(\w3[3][40] ), .Z(n2068) );
  XNOR U3170 ( .A(n2104), .B(n2068), .Z(\w0[4][32] ) );
  XOR U3171 ( .A(\w3[3][34] ), .B(\w3[3][58] ), .Z(n2109) );
  XOR U3172 ( .A(\w3[3][41] ), .B(\w3[3][49] ), .Z(n2127) );
  XNOR U3173 ( .A(\w3[3][57] ), .B(n2127), .Z(n2069) );
  XNOR U3174 ( .A(n2109), .B(n2069), .Z(\w0[4][33] ) );
  XOR U3175 ( .A(\w3[3][35] ), .B(\w3[3][59] ), .Z(n2089) );
  XOR U3176 ( .A(\w3[3][58] ), .B(\w3[3][50] ), .Z(n2129) );
  XNOR U3177 ( .A(\w3[3][42] ), .B(n2129), .Z(n2070) );
  XNOR U3178 ( .A(n2089), .B(n2070), .Z(\w0[4][34] ) );
  XOR U3179 ( .A(\w3[3][36] ), .B(\w3[3][32] ), .Z(n2091) );
  XOR U3180 ( .A(\w3[3][43] ), .B(\w3[3][51] ), .Z(n2111) );
  XNOR U3181 ( .A(\w3[3][56] ), .B(n2111), .Z(n2071) );
  XNOR U3182 ( .A(\w3[3][60] ), .B(n2071), .Z(n2133) );
  XNOR U3183 ( .A(\w3[3][59] ), .B(n2133), .Z(n2072) );
  XNOR U3184 ( .A(n2091), .B(n2072), .Z(\w0[4][35] ) );
  XOR U3185 ( .A(\w3[3][32] ), .B(\w3[3][37] ), .Z(n2095) );
  XOR U3186 ( .A(\w3[3][44] ), .B(\w3[3][52] ), .Z(n2074) );
  XNOR U3187 ( .A(\w3[3][56] ), .B(\w3[3][61] ), .Z(n2073) );
  XNOR U3188 ( .A(n2074), .B(n2073), .Z(n2139) );
  XNOR U3189 ( .A(\w3[3][60] ), .B(n2139), .Z(n2075) );
  XNOR U3190 ( .A(n2095), .B(n2075), .Z(\w0[4][36] ) );
  XOR U3191 ( .A(\w3[3][38] ), .B(\w3[3][62] ), .Z(n2099) );
  XOR U3192 ( .A(\w3[3][45] ), .B(\w3[3][53] ), .Z(n2142) );
  XNOR U3193 ( .A(\w3[3][61] ), .B(n2142), .Z(n2076) );
  XNOR U3194 ( .A(n2099), .B(n2076), .Z(\w0[4][37] ) );
  XOR U3195 ( .A(\w3[3][32] ), .B(\w3[3][39] ), .Z(n2100) );
  XOR U3196 ( .A(\w3[3][46] ), .B(\w3[3][54] ), .Z(n2116) );
  XNOR U3197 ( .A(\w3[3][56] ), .B(\w3[3][63] ), .Z(n2078) );
  XNOR U3198 ( .A(n2116), .B(n2078), .Z(n2145) );
  XNOR U3199 ( .A(\w3[3][62] ), .B(n2145), .Z(n2077) );
  XNOR U3200 ( .A(n2100), .B(n2077), .Z(\w0[4][38] ) );
  XNOR U3201 ( .A(\w3[3][47] ), .B(\w3[3][55] ), .Z(n2150) );
  XNOR U3202 ( .A(\w3[3][32] ), .B(n2078), .Z(n2079) );
  XNOR U3203 ( .A(n2150), .B(n2079), .Z(\w0[4][39] ) );
  XNOR U3204 ( .A(n2080), .B(\w3[3][27] ), .Z(n2081) );
  XNOR U3205 ( .A(n2082), .B(n2081), .Z(\w0[4][3] ) );
  XOR U3206 ( .A(\w3[3][41] ), .B(\w3[3][32] ), .Z(n2084) );
  XNOR U3207 ( .A(n2148), .B(\w3[3][33] ), .Z(n2083) );
  XNOR U3208 ( .A(n2084), .B(n2083), .Z(\w0[4][40] ) );
  XOR U3209 ( .A(\w3[3][34] ), .B(\w3[3][42] ), .Z(n2086) );
  XNOR U3210 ( .A(n2104), .B(\w3[3][49] ), .Z(n2085) );
  XNOR U3211 ( .A(n2086), .B(n2085), .Z(\w0[4][41] ) );
  XOR U3212 ( .A(\w3[3][35] ), .B(\w3[3][43] ), .Z(n2088) );
  XNOR U3213 ( .A(n2109), .B(\w3[3][50] ), .Z(n2087) );
  XNOR U3214 ( .A(n2088), .B(n2087), .Z(\w0[4][42] ) );
  XNOR U3215 ( .A(\w3[3][40] ), .B(n2089), .Z(n2090) );
  XNOR U3216 ( .A(\w3[3][44] ), .B(n2090), .Z(n2112) );
  XNOR U3217 ( .A(\w3[3][51] ), .B(n2091), .Z(n2092) );
  XNOR U3218 ( .A(n2112), .B(n2092), .Z(\w0[4][43] ) );
  XOR U3219 ( .A(\w3[3][36] ), .B(\w3[3][45] ), .Z(n2094) );
  XNOR U3220 ( .A(\w3[3][40] ), .B(\w3[3][60] ), .Z(n2093) );
  XNOR U3221 ( .A(n2094), .B(n2093), .Z(n2114) );
  XNOR U3222 ( .A(\w3[3][52] ), .B(n2095), .Z(n2096) );
  XNOR U3223 ( .A(n2114), .B(n2096), .Z(\w0[4][44] ) );
  XOR U3224 ( .A(\w3[3][61] ), .B(\w3[3][37] ), .Z(n2118) );
  XOR U3225 ( .A(\w3[3][46] ), .B(n2118), .Z(n2098) );
  XNOR U3226 ( .A(\w3[3][53] ), .B(\w3[3][38] ), .Z(n2097) );
  XNOR U3227 ( .A(n2098), .B(n2097), .Z(\w0[4][45] ) );
  XNOR U3228 ( .A(\w3[3][40] ), .B(\w3[3][47] ), .Z(n2123) );
  XNOR U3229 ( .A(n2099), .B(n2123), .Z(n2119) );
  XNOR U3230 ( .A(\w3[3][54] ), .B(n2100), .Z(n2101) );
  XNOR U3231 ( .A(n2119), .B(n2101), .Z(\w0[4][46] ) );
  XOR U3232 ( .A(\w3[3][63] ), .B(\w3[3][39] ), .Z(n2121) );
  XOR U3233 ( .A(\w3[3][40] ), .B(\w3[3][32] ), .Z(n2124) );
  XNOR U3234 ( .A(\w3[3][55] ), .B(n2124), .Z(n2102) );
  XNOR U3235 ( .A(n2121), .B(n2102), .Z(\w0[4][47] ) );
  XNOR U3236 ( .A(\w3[3][56] ), .B(n2127), .Z(n2103) );
  XNOR U3237 ( .A(n2124), .B(n2103), .Z(\w0[4][48] ) );
  XOR U3238 ( .A(\w3[3][42] ), .B(\w3[3][50] ), .Z(n2130) );
  XNOR U3239 ( .A(n2104), .B(\w3[3][41] ), .Z(n2105) );
  XNOR U3240 ( .A(n2130), .B(n2105), .Z(\w0[4][49] ) );
  XNOR U3241 ( .A(n2106), .B(\w3[3][28] ), .Z(n2107) );
  XNOR U3242 ( .A(n2108), .B(n2107), .Z(\w0[4][4] ) );
  XNOR U3243 ( .A(n2109), .B(\w3[3][42] ), .Z(n2110) );
  XNOR U3244 ( .A(n2111), .B(n2110), .Z(\w0[4][50] ) );
  XOR U3245 ( .A(\w3[3][48] ), .B(\w3[3][52] ), .Z(n2135) );
  XNOR U3246 ( .A(\w3[3][43] ), .B(n2112), .Z(n2113) );
  XNOR U3247 ( .A(n2135), .B(n2113), .Z(\w0[4][51] ) );
  XOR U3248 ( .A(\w3[3][48] ), .B(\w3[3][53] ), .Z(n2141) );
  XNOR U3249 ( .A(\w3[3][44] ), .B(n2114), .Z(n2115) );
  XNOR U3250 ( .A(n2141), .B(n2115), .Z(\w0[4][52] ) );
  XNOR U3251 ( .A(\w3[3][45] ), .B(n2116), .Z(n2117) );
  XNOR U3252 ( .A(n2118), .B(n2117), .Z(\w0[4][53] ) );
  XOR U3253 ( .A(\w3[3][48] ), .B(\w3[3][55] ), .Z(n2147) );
  XNOR U3254 ( .A(\w3[3][46] ), .B(n2119), .Z(n2120) );
  XNOR U3255 ( .A(n2147), .B(n2120), .Z(\w0[4][54] ) );
  XOR U3256 ( .A(\w3[3][48] ), .B(n2121), .Z(n2122) );
  XNOR U3257 ( .A(n2123), .B(n2122), .Z(\w0[4][55] ) );
  XOR U3258 ( .A(\w3[3][49] ), .B(n2124), .Z(n2126) );
  XNOR U3259 ( .A(\w3[3][48] ), .B(\w3[3][57] ), .Z(n2125) );
  XNOR U3260 ( .A(n2126), .B(n2125), .Z(\w0[4][56] ) );
  XNOR U3261 ( .A(\w3[3][33] ), .B(n2127), .Z(n2128) );
  XNOR U3262 ( .A(n2129), .B(n2128), .Z(\w0[4][57] ) );
  XOR U3263 ( .A(\w3[3][51] ), .B(n2130), .Z(n2132) );
  XNOR U3264 ( .A(\w3[3][34] ), .B(\w3[3][59] ), .Z(n2131) );
  XNOR U3265 ( .A(n2132), .B(n2131), .Z(\w0[4][58] ) );
  XNOR U3266 ( .A(\w3[3][35] ), .B(n2133), .Z(n2134) );
  XNOR U3267 ( .A(n2135), .B(n2134), .Z(\w0[4][59] ) );
  XNOR U3268 ( .A(\w3[3][29] ), .B(n2136), .Z(n2137) );
  XNOR U3269 ( .A(n2138), .B(n2137), .Z(\w0[4][5] ) );
  XNOR U3270 ( .A(\w3[3][36] ), .B(n2139), .Z(n2140) );
  XNOR U3271 ( .A(n2141), .B(n2140), .Z(\w0[4][60] ) );
  XOR U3272 ( .A(\w3[3][62] ), .B(\w3[3][54] ), .Z(n2144) );
  XNOR U3273 ( .A(\w3[3][37] ), .B(n2142), .Z(n2143) );
  XNOR U3274 ( .A(n2144), .B(n2143), .Z(\w0[4][61] ) );
  XNOR U3275 ( .A(\w3[3][38] ), .B(n2145), .Z(n2146) );
  XNOR U3276 ( .A(n2147), .B(n2146), .Z(\w0[4][62] ) );
  XOR U3277 ( .A(n2148), .B(\w3[3][39] ), .Z(n2149) );
  XNOR U3278 ( .A(n2150), .B(n2149), .Z(\w0[4][63] ) );
  XOR U3279 ( .A(\w3[3][65] ), .B(\w3[3][89] ), .Z(n2190) );
  XOR U3280 ( .A(\w3[3][80] ), .B(\w3[3][88] ), .Z(n2231) );
  XNOR U3281 ( .A(n2231), .B(\w3[3][72] ), .Z(n2151) );
  XNOR U3282 ( .A(n2190), .B(n2151), .Z(\w0[4][64] ) );
  XOR U3283 ( .A(\w3[3][66] ), .B(\w3[3][90] ), .Z(n2192) );
  XOR U3284 ( .A(\w3[3][73] ), .B(\w3[3][81] ), .Z(n2210) );
  XNOR U3285 ( .A(\w3[3][89] ), .B(n2210), .Z(n2152) );
  XNOR U3286 ( .A(n2192), .B(n2152), .Z(\w0[4][65] ) );
  XOR U3287 ( .A(\w3[3][67] ), .B(\w3[3][91] ), .Z(n2172) );
  XOR U3288 ( .A(\w3[3][74] ), .B(\w3[3][82] ), .Z(n2216) );
  XNOR U3289 ( .A(\w3[3][90] ), .B(n2216), .Z(n2153) );
  XNOR U3290 ( .A(n2172), .B(n2153), .Z(\w0[4][66] ) );
  XOR U3291 ( .A(\w3[3][68] ), .B(\w3[3][64] ), .Z(n2174) );
  XOR U3292 ( .A(\w3[3][75] ), .B(\w3[3][83] ), .Z(n2194) );
  XNOR U3293 ( .A(\w3[3][88] ), .B(n2194), .Z(n2154) );
  XNOR U3294 ( .A(\w3[3][92] ), .B(n2154), .Z(n2219) );
  XNOR U3295 ( .A(\w3[3][91] ), .B(n2219), .Z(n2155) );
  XNOR U3296 ( .A(n2174), .B(n2155), .Z(\w0[4][67] ) );
  XOR U3297 ( .A(\w3[3][64] ), .B(\w3[3][69] ), .Z(n2178) );
  XOR U3298 ( .A(\w3[3][76] ), .B(\w3[3][84] ), .Z(n2157) );
  XNOR U3299 ( .A(\w3[3][88] ), .B(\w3[3][93] ), .Z(n2156) );
  XNOR U3300 ( .A(n2157), .B(n2156), .Z(n2222) );
  XNOR U3301 ( .A(\w3[3][92] ), .B(n2222), .Z(n2158) );
  XNOR U3302 ( .A(n2178), .B(n2158), .Z(\w0[4][68] ) );
  XOR U3303 ( .A(\w3[3][70] ), .B(\w3[3][94] ), .Z(n2182) );
  XOR U3304 ( .A(\w3[3][77] ), .B(\w3[3][85] ), .Z(n2225) );
  XNOR U3305 ( .A(\w3[3][93] ), .B(n2225), .Z(n2159) );
  XNOR U3306 ( .A(n2182), .B(n2159), .Z(\w0[4][69] ) );
  XNOR U3307 ( .A(n2160), .B(\w3[3][30] ), .Z(n2161) );
  XNOR U3308 ( .A(n2162), .B(n2161), .Z(\w0[4][6] ) );
  XOR U3309 ( .A(\w3[3][64] ), .B(\w3[3][71] ), .Z(n2183) );
  XOR U3310 ( .A(\w3[3][78] ), .B(\w3[3][86] ), .Z(n2199) );
  XNOR U3311 ( .A(\w3[3][88] ), .B(\w3[3][95] ), .Z(n2164) );
  XNOR U3312 ( .A(n2199), .B(n2164), .Z(n2228) );
  XNOR U3313 ( .A(\w3[3][94] ), .B(n2228), .Z(n2163) );
  XNOR U3314 ( .A(n2183), .B(n2163), .Z(\w0[4][70] ) );
  XNOR U3315 ( .A(\w3[3][79] ), .B(\w3[3][87] ), .Z(n2233) );
  XNOR U3316 ( .A(\w3[3][64] ), .B(n2164), .Z(n2165) );
  XNOR U3317 ( .A(n2233), .B(n2165), .Z(\w0[4][71] ) );
  XOR U3318 ( .A(\w3[3][73] ), .B(\w3[3][64] ), .Z(n2167) );
  XNOR U3319 ( .A(n2231), .B(\w3[3][65] ), .Z(n2166) );
  XNOR U3320 ( .A(n2167), .B(n2166), .Z(\w0[4][72] ) );
  XOR U3321 ( .A(\w3[3][66] ), .B(\w3[3][74] ), .Z(n2169) );
  XNOR U3322 ( .A(n2190), .B(\w3[3][81] ), .Z(n2168) );
  XNOR U3323 ( .A(n2169), .B(n2168), .Z(\w0[4][73] ) );
  XOR U3324 ( .A(\w3[3][67] ), .B(\w3[3][75] ), .Z(n2171) );
  XNOR U3325 ( .A(n2192), .B(\w3[3][82] ), .Z(n2170) );
  XNOR U3326 ( .A(n2171), .B(n2170), .Z(\w0[4][74] ) );
  XNOR U3327 ( .A(\w3[3][72] ), .B(n2172), .Z(n2173) );
  XNOR U3328 ( .A(\w3[3][76] ), .B(n2173), .Z(n2195) );
  XNOR U3329 ( .A(\w3[3][83] ), .B(n2174), .Z(n2175) );
  XNOR U3330 ( .A(n2195), .B(n2175), .Z(\w0[4][75] ) );
  XOR U3331 ( .A(\w3[3][68] ), .B(\w3[3][77] ), .Z(n2177) );
  XNOR U3332 ( .A(\w3[3][72] ), .B(\w3[3][92] ), .Z(n2176) );
  XNOR U3333 ( .A(n2177), .B(n2176), .Z(n2197) );
  XNOR U3334 ( .A(\w3[3][84] ), .B(n2178), .Z(n2179) );
  XNOR U3335 ( .A(n2197), .B(n2179), .Z(\w0[4][76] ) );
  XOR U3336 ( .A(\w3[3][93] ), .B(\w3[3][69] ), .Z(n2201) );
  XOR U3337 ( .A(\w3[3][78] ), .B(n2201), .Z(n2181) );
  XNOR U3338 ( .A(\w3[3][85] ), .B(\w3[3][70] ), .Z(n2180) );
  XNOR U3339 ( .A(n2181), .B(n2180), .Z(\w0[4][77] ) );
  XNOR U3340 ( .A(\w3[3][72] ), .B(\w3[3][79] ), .Z(n2206) );
  XNOR U3341 ( .A(n2182), .B(n2206), .Z(n2202) );
  XNOR U3342 ( .A(\w3[3][86] ), .B(n2183), .Z(n2184) );
  XNOR U3343 ( .A(n2202), .B(n2184), .Z(\w0[4][78] ) );
  XOR U3344 ( .A(\w3[3][95] ), .B(\w3[3][71] ), .Z(n2204) );
  XOR U3345 ( .A(\w3[3][72] ), .B(\w3[3][64] ), .Z(n2207) );
  XNOR U3346 ( .A(\w3[3][87] ), .B(n2207), .Z(n2185) );
  XNOR U3347 ( .A(n2204), .B(n2185), .Z(\w0[4][79] ) );
  XOR U3348 ( .A(\w3[3][0] ), .B(n2186), .Z(n2187) );
  XNOR U3349 ( .A(n2188), .B(n2187), .Z(\w0[4][7] ) );
  XNOR U3350 ( .A(\w3[3][88] ), .B(n2210), .Z(n2189) );
  XNOR U3351 ( .A(n2207), .B(n2189), .Z(\w0[4][80] ) );
  XNOR U3352 ( .A(n2190), .B(\w3[3][73] ), .Z(n2191) );
  XNOR U3353 ( .A(n2216), .B(n2191), .Z(\w0[4][81] ) );
  XNOR U3354 ( .A(n2192), .B(\w3[3][74] ), .Z(n2193) );
  XNOR U3355 ( .A(n2194), .B(n2193), .Z(\w0[4][82] ) );
  XOR U3356 ( .A(\w3[3][80] ), .B(\w3[3][84] ), .Z(n2221) );
  XNOR U3357 ( .A(\w3[3][75] ), .B(n2195), .Z(n2196) );
  XNOR U3358 ( .A(n2221), .B(n2196), .Z(\w0[4][83] ) );
  XOR U3359 ( .A(\w3[3][80] ), .B(\w3[3][85] ), .Z(n2224) );
  XNOR U3360 ( .A(\w3[3][76] ), .B(n2197), .Z(n2198) );
  XNOR U3361 ( .A(n2224), .B(n2198), .Z(\w0[4][84] ) );
  XNOR U3362 ( .A(\w3[3][77] ), .B(n2199), .Z(n2200) );
  XNOR U3363 ( .A(n2201), .B(n2200), .Z(\w0[4][85] ) );
  XOR U3364 ( .A(\w3[3][80] ), .B(\w3[3][87] ), .Z(n2230) );
  XNOR U3365 ( .A(\w3[3][78] ), .B(n2202), .Z(n2203) );
  XNOR U3366 ( .A(n2230), .B(n2203), .Z(\w0[4][86] ) );
  XOR U3367 ( .A(\w3[3][80] ), .B(n2204), .Z(n2205) );
  XNOR U3368 ( .A(n2206), .B(n2205), .Z(\w0[4][87] ) );
  XOR U3369 ( .A(\w3[3][81] ), .B(n2207), .Z(n2209) );
  XNOR U3370 ( .A(\w3[3][80] ), .B(\w3[3][89] ), .Z(n2208) );
  XNOR U3371 ( .A(n2209), .B(n2208), .Z(\w0[4][88] ) );
  XOR U3372 ( .A(\w3[3][90] ), .B(\w3[3][82] ), .Z(n2212) );
  XNOR U3373 ( .A(\w3[3][65] ), .B(n2210), .Z(n2211) );
  XNOR U3374 ( .A(n2212), .B(n2211), .Z(\w0[4][89] ) );
  XOR U3375 ( .A(\w3[3][0] ), .B(\w3[3][9] ), .Z(n2215) );
  XNOR U3376 ( .A(\w3[3][1] ), .B(n2213), .Z(n2214) );
  XNOR U3377 ( .A(n2215), .B(n2214), .Z(\w0[4][8] ) );
  XOR U3378 ( .A(\w3[3][91] ), .B(\w3[3][83] ), .Z(n2218) );
  XNOR U3379 ( .A(\w3[3][66] ), .B(n2216), .Z(n2217) );
  XNOR U3380 ( .A(n2218), .B(n2217), .Z(\w0[4][90] ) );
  XNOR U3381 ( .A(\w3[3][67] ), .B(n2219), .Z(n2220) );
  XNOR U3382 ( .A(n2221), .B(n2220), .Z(\w0[4][91] ) );
  XNOR U3383 ( .A(\w3[3][68] ), .B(n2222), .Z(n2223) );
  XNOR U3384 ( .A(n2224), .B(n2223), .Z(\w0[4][92] ) );
  XOR U3385 ( .A(\w3[3][94] ), .B(\w3[3][86] ), .Z(n2227) );
  XNOR U3386 ( .A(\w3[3][69] ), .B(n2225), .Z(n2226) );
  XNOR U3387 ( .A(n2227), .B(n2226), .Z(\w0[4][93] ) );
  XNOR U3388 ( .A(\w3[3][70] ), .B(n2228), .Z(n2229) );
  XNOR U3389 ( .A(n2230), .B(n2229), .Z(\w0[4][94] ) );
  XOR U3390 ( .A(n2231), .B(\w3[3][71] ), .Z(n2232) );
  XNOR U3391 ( .A(n2233), .B(n2232), .Z(\w0[4][95] ) );
  XNOR U3392 ( .A(n2235), .B(n2234), .Z(n2236) );
  XNOR U3393 ( .A(\w3[3][104] ), .B(n2236), .Z(\w0[4][96] ) );
  XNOR U3394 ( .A(\w3[3][105] ), .B(n2237), .Z(n2238) );
  XNOR U3395 ( .A(n2239), .B(n2238), .Z(\w0[4][97] ) );
  XNOR U3396 ( .A(\w3[3][106] ), .B(n2240), .Z(n2241) );
  XNOR U3397 ( .A(n2242), .B(n2241), .Z(\w0[4][98] ) );
  XNOR U3398 ( .A(n2243), .B(\w3[3][123] ), .Z(n2244) );
  XNOR U3399 ( .A(n2245), .B(n2244), .Z(\w0[4][99] ) );
  XOR U3400 ( .A(\w3[3][17] ), .B(\w3[3][10] ), .Z(n2248) );
  XNOR U3401 ( .A(n2246), .B(\w3[3][2] ), .Z(n2247) );
  XNOR U3402 ( .A(n2248), .B(n2247), .Z(\w0[4][9] ) );
  NANDN U3403 ( .A(state[0]), .B(init), .Z(n2250) );
  OR U3404 ( .A(init), .B(msg[0]), .Z(n2249) );
  NAND U3405 ( .A(n2250), .B(n2249), .Z(n2251) );
  XNOR U3406 ( .A(key[0]), .B(n2251), .Z(\w1[0][0] ) );
  NANDN U3407 ( .A(state[100]), .B(init), .Z(n2253) );
  OR U3408 ( .A(init), .B(msg[100]), .Z(n2252) );
  NAND U3409 ( .A(n2253), .B(n2252), .Z(n2254) );
  XNOR U3410 ( .A(key[100]), .B(n2254), .Z(\w1[0][100] ) );
  NANDN U3411 ( .A(state[101]), .B(init), .Z(n2256) );
  OR U3412 ( .A(init), .B(msg[101]), .Z(n2255) );
  NAND U3413 ( .A(n2256), .B(n2255), .Z(n2257) );
  XNOR U3414 ( .A(key[101]), .B(n2257), .Z(\w1[0][101] ) );
  NANDN U3415 ( .A(state[102]), .B(init), .Z(n2259) );
  OR U3416 ( .A(init), .B(msg[102]), .Z(n2258) );
  NAND U3417 ( .A(n2259), .B(n2258), .Z(n2260) );
  XNOR U3418 ( .A(key[102]), .B(n2260), .Z(\w1[0][102] ) );
  NANDN U3419 ( .A(state[103]), .B(init), .Z(n2262) );
  OR U3420 ( .A(init), .B(msg[103]), .Z(n2261) );
  NAND U3421 ( .A(n2262), .B(n2261), .Z(n2263) );
  XNOR U3422 ( .A(key[103]), .B(n2263), .Z(\w1[0][103] ) );
  NANDN U3423 ( .A(state[104]), .B(init), .Z(n2265) );
  OR U3424 ( .A(init), .B(msg[104]), .Z(n2264) );
  NAND U3425 ( .A(n2265), .B(n2264), .Z(n2266) );
  XNOR U3426 ( .A(key[104]), .B(n2266), .Z(\w1[0][104] ) );
  NANDN U3427 ( .A(state[105]), .B(init), .Z(n2268) );
  OR U3428 ( .A(init), .B(msg[105]), .Z(n2267) );
  NAND U3429 ( .A(n2268), .B(n2267), .Z(n2269) );
  XNOR U3430 ( .A(key[105]), .B(n2269), .Z(\w1[0][105] ) );
  NANDN U3431 ( .A(state[106]), .B(init), .Z(n2271) );
  OR U3432 ( .A(init), .B(msg[106]), .Z(n2270) );
  NAND U3433 ( .A(n2271), .B(n2270), .Z(n2272) );
  XNOR U3434 ( .A(key[106]), .B(n2272), .Z(\w1[0][106] ) );
  NANDN U3435 ( .A(state[107]), .B(init), .Z(n2274) );
  OR U3436 ( .A(init), .B(msg[107]), .Z(n2273) );
  NAND U3437 ( .A(n2274), .B(n2273), .Z(n2275) );
  XNOR U3438 ( .A(key[107]), .B(n2275), .Z(\w1[0][107] ) );
  NANDN U3439 ( .A(state[108]), .B(init), .Z(n2277) );
  OR U3440 ( .A(init), .B(msg[108]), .Z(n2276) );
  NAND U3441 ( .A(n2277), .B(n2276), .Z(n2278) );
  XNOR U3442 ( .A(key[108]), .B(n2278), .Z(\w1[0][108] ) );
  NANDN U3443 ( .A(state[109]), .B(init), .Z(n2280) );
  OR U3444 ( .A(init), .B(msg[109]), .Z(n2279) );
  NAND U3445 ( .A(n2280), .B(n2279), .Z(n2281) );
  XNOR U3446 ( .A(key[109]), .B(n2281), .Z(\w1[0][109] ) );
  NANDN U3447 ( .A(state[10]), .B(init), .Z(n2283) );
  OR U3448 ( .A(init), .B(msg[10]), .Z(n2282) );
  NAND U3449 ( .A(n2283), .B(n2282), .Z(n2284) );
  XNOR U3450 ( .A(key[10]), .B(n2284), .Z(\w1[0][10] ) );
  NANDN U3451 ( .A(state[110]), .B(init), .Z(n2286) );
  OR U3452 ( .A(init), .B(msg[110]), .Z(n2285) );
  NAND U3453 ( .A(n2286), .B(n2285), .Z(n2287) );
  XNOR U3454 ( .A(key[110]), .B(n2287), .Z(\w1[0][110] ) );
  NANDN U3455 ( .A(state[111]), .B(init), .Z(n2289) );
  OR U3456 ( .A(init), .B(msg[111]), .Z(n2288) );
  NAND U3457 ( .A(n2289), .B(n2288), .Z(n2290) );
  XNOR U3458 ( .A(key[111]), .B(n2290), .Z(\w1[0][111] ) );
  NANDN U3459 ( .A(state[112]), .B(init), .Z(n2292) );
  OR U3460 ( .A(init), .B(msg[112]), .Z(n2291) );
  NAND U3461 ( .A(n2292), .B(n2291), .Z(n2293) );
  XNOR U3462 ( .A(key[112]), .B(n2293), .Z(\w1[0][112] ) );
  NANDN U3463 ( .A(state[113]), .B(init), .Z(n2295) );
  OR U3464 ( .A(init), .B(msg[113]), .Z(n2294) );
  NAND U3465 ( .A(n2295), .B(n2294), .Z(n2296) );
  XNOR U3466 ( .A(key[113]), .B(n2296), .Z(\w1[0][113] ) );
  NANDN U3467 ( .A(state[114]), .B(init), .Z(n2298) );
  OR U3468 ( .A(init), .B(msg[114]), .Z(n2297) );
  NAND U3469 ( .A(n2298), .B(n2297), .Z(n2299) );
  XNOR U3470 ( .A(key[114]), .B(n2299), .Z(\w1[0][114] ) );
  NANDN U3471 ( .A(state[115]), .B(init), .Z(n2301) );
  OR U3472 ( .A(init), .B(msg[115]), .Z(n2300) );
  NAND U3473 ( .A(n2301), .B(n2300), .Z(n2302) );
  XNOR U3474 ( .A(key[115]), .B(n2302), .Z(\w1[0][115] ) );
  NANDN U3475 ( .A(state[116]), .B(init), .Z(n2304) );
  OR U3476 ( .A(init), .B(msg[116]), .Z(n2303) );
  NAND U3477 ( .A(n2304), .B(n2303), .Z(n2305) );
  XNOR U3478 ( .A(key[116]), .B(n2305), .Z(\w1[0][116] ) );
  NANDN U3479 ( .A(state[117]), .B(init), .Z(n2307) );
  OR U3480 ( .A(init), .B(msg[117]), .Z(n2306) );
  NAND U3481 ( .A(n2307), .B(n2306), .Z(n2308) );
  XNOR U3482 ( .A(key[117]), .B(n2308), .Z(\w1[0][117] ) );
  NANDN U3483 ( .A(state[118]), .B(init), .Z(n2310) );
  OR U3484 ( .A(init), .B(msg[118]), .Z(n2309) );
  NAND U3485 ( .A(n2310), .B(n2309), .Z(n2311) );
  XNOR U3486 ( .A(key[118]), .B(n2311), .Z(\w1[0][118] ) );
  NANDN U3487 ( .A(state[119]), .B(init), .Z(n2313) );
  OR U3488 ( .A(init), .B(msg[119]), .Z(n2312) );
  NAND U3489 ( .A(n2313), .B(n2312), .Z(n2314) );
  XNOR U3490 ( .A(key[119]), .B(n2314), .Z(\w1[0][119] ) );
  NANDN U3491 ( .A(state[11]), .B(init), .Z(n2316) );
  OR U3492 ( .A(init), .B(msg[11]), .Z(n2315) );
  NAND U3493 ( .A(n2316), .B(n2315), .Z(n2317) );
  XNOR U3494 ( .A(key[11]), .B(n2317), .Z(\w1[0][11] ) );
  NANDN U3495 ( .A(state[120]), .B(init), .Z(n2319) );
  OR U3496 ( .A(init), .B(msg[120]), .Z(n2318) );
  NAND U3497 ( .A(n2319), .B(n2318), .Z(n2320) );
  XNOR U3498 ( .A(key[120]), .B(n2320), .Z(\w1[0][120] ) );
  NANDN U3499 ( .A(state[121]), .B(init), .Z(n2322) );
  OR U3500 ( .A(init), .B(msg[121]), .Z(n2321) );
  NAND U3501 ( .A(n2322), .B(n2321), .Z(n2323) );
  XNOR U3502 ( .A(key[121]), .B(n2323), .Z(\w1[0][121] ) );
  NANDN U3503 ( .A(state[122]), .B(init), .Z(n2325) );
  OR U3504 ( .A(init), .B(msg[122]), .Z(n2324) );
  NAND U3505 ( .A(n2325), .B(n2324), .Z(n2326) );
  XNOR U3506 ( .A(key[122]), .B(n2326), .Z(\w1[0][122] ) );
  NANDN U3507 ( .A(state[123]), .B(init), .Z(n2328) );
  OR U3508 ( .A(init), .B(msg[123]), .Z(n2327) );
  NAND U3509 ( .A(n2328), .B(n2327), .Z(n2329) );
  XNOR U3510 ( .A(key[123]), .B(n2329), .Z(\w1[0][123] ) );
  NANDN U3511 ( .A(state[124]), .B(init), .Z(n2331) );
  OR U3512 ( .A(init), .B(msg[124]), .Z(n2330) );
  NAND U3513 ( .A(n2331), .B(n2330), .Z(n2332) );
  XNOR U3514 ( .A(key[124]), .B(n2332), .Z(\w1[0][124] ) );
  NANDN U3515 ( .A(state[125]), .B(init), .Z(n2334) );
  OR U3516 ( .A(init), .B(msg[125]), .Z(n2333) );
  NAND U3517 ( .A(n2334), .B(n2333), .Z(n2335) );
  XNOR U3518 ( .A(key[125]), .B(n2335), .Z(\w1[0][125] ) );
  NANDN U3519 ( .A(state[126]), .B(init), .Z(n2337) );
  OR U3520 ( .A(init), .B(msg[126]), .Z(n2336) );
  NAND U3521 ( .A(n2337), .B(n2336), .Z(n2338) );
  XNOR U3522 ( .A(key[126]), .B(n2338), .Z(\w1[0][126] ) );
  NANDN U3523 ( .A(state[127]), .B(init), .Z(n2340) );
  OR U3524 ( .A(init), .B(msg[127]), .Z(n2339) );
  NAND U3525 ( .A(n2340), .B(n2339), .Z(n2341) );
  XNOR U3526 ( .A(key[127]), .B(n2341), .Z(\w1[0][127] ) );
  NANDN U3527 ( .A(state[12]), .B(init), .Z(n2343) );
  OR U3528 ( .A(init), .B(msg[12]), .Z(n2342) );
  NAND U3529 ( .A(n2343), .B(n2342), .Z(n2344) );
  XNOR U3530 ( .A(key[12]), .B(n2344), .Z(\w1[0][12] ) );
  NANDN U3531 ( .A(state[13]), .B(init), .Z(n2346) );
  OR U3532 ( .A(init), .B(msg[13]), .Z(n2345) );
  NAND U3533 ( .A(n2346), .B(n2345), .Z(n2347) );
  XNOR U3534 ( .A(key[13]), .B(n2347), .Z(\w1[0][13] ) );
  NANDN U3535 ( .A(state[14]), .B(init), .Z(n2349) );
  OR U3536 ( .A(init), .B(msg[14]), .Z(n2348) );
  NAND U3537 ( .A(n2349), .B(n2348), .Z(n2350) );
  XNOR U3538 ( .A(key[14]), .B(n2350), .Z(\w1[0][14] ) );
  NANDN U3539 ( .A(state[15]), .B(init), .Z(n2352) );
  OR U3540 ( .A(init), .B(msg[15]), .Z(n2351) );
  NAND U3541 ( .A(n2352), .B(n2351), .Z(n2353) );
  XNOR U3542 ( .A(key[15]), .B(n2353), .Z(\w1[0][15] ) );
  NANDN U3543 ( .A(state[16]), .B(init), .Z(n2355) );
  OR U3544 ( .A(init), .B(msg[16]), .Z(n2354) );
  NAND U3545 ( .A(n2355), .B(n2354), .Z(n2356) );
  XNOR U3546 ( .A(key[16]), .B(n2356), .Z(\w1[0][16] ) );
  NANDN U3547 ( .A(state[17]), .B(init), .Z(n2358) );
  OR U3548 ( .A(init), .B(msg[17]), .Z(n2357) );
  NAND U3549 ( .A(n2358), .B(n2357), .Z(n2359) );
  XNOR U3550 ( .A(key[17]), .B(n2359), .Z(\w1[0][17] ) );
  NANDN U3551 ( .A(state[18]), .B(init), .Z(n2361) );
  OR U3552 ( .A(init), .B(msg[18]), .Z(n2360) );
  NAND U3553 ( .A(n2361), .B(n2360), .Z(n2362) );
  XNOR U3554 ( .A(key[18]), .B(n2362), .Z(\w1[0][18] ) );
  NANDN U3555 ( .A(state[19]), .B(init), .Z(n2364) );
  OR U3556 ( .A(init), .B(msg[19]), .Z(n2363) );
  NAND U3557 ( .A(n2364), .B(n2363), .Z(n2365) );
  XNOR U3558 ( .A(key[19]), .B(n2365), .Z(\w1[0][19] ) );
  NANDN U3559 ( .A(state[1]), .B(init), .Z(n2367) );
  OR U3560 ( .A(init), .B(msg[1]), .Z(n2366) );
  NAND U3561 ( .A(n2367), .B(n2366), .Z(n2368) );
  XNOR U3562 ( .A(key[1]), .B(n2368), .Z(\w1[0][1] ) );
  NANDN U3563 ( .A(state[20]), .B(init), .Z(n2370) );
  OR U3564 ( .A(init), .B(msg[20]), .Z(n2369) );
  NAND U3565 ( .A(n2370), .B(n2369), .Z(n2371) );
  XNOR U3566 ( .A(key[20]), .B(n2371), .Z(\w1[0][20] ) );
  NANDN U3567 ( .A(state[21]), .B(init), .Z(n2373) );
  OR U3568 ( .A(init), .B(msg[21]), .Z(n2372) );
  NAND U3569 ( .A(n2373), .B(n2372), .Z(n2374) );
  XNOR U3570 ( .A(key[21]), .B(n2374), .Z(\w1[0][21] ) );
  NANDN U3571 ( .A(state[22]), .B(init), .Z(n2376) );
  OR U3572 ( .A(init), .B(msg[22]), .Z(n2375) );
  NAND U3573 ( .A(n2376), .B(n2375), .Z(n2377) );
  XNOR U3574 ( .A(key[22]), .B(n2377), .Z(\w1[0][22] ) );
  NANDN U3575 ( .A(state[23]), .B(init), .Z(n2379) );
  OR U3576 ( .A(init), .B(msg[23]), .Z(n2378) );
  NAND U3577 ( .A(n2379), .B(n2378), .Z(n2380) );
  XNOR U3578 ( .A(key[23]), .B(n2380), .Z(\w1[0][23] ) );
  NANDN U3579 ( .A(state[24]), .B(init), .Z(n2382) );
  OR U3580 ( .A(init), .B(msg[24]), .Z(n2381) );
  NAND U3581 ( .A(n2382), .B(n2381), .Z(n2383) );
  XNOR U3582 ( .A(key[24]), .B(n2383), .Z(\w1[0][24] ) );
  NANDN U3583 ( .A(state[25]), .B(init), .Z(n2385) );
  OR U3584 ( .A(init), .B(msg[25]), .Z(n2384) );
  NAND U3585 ( .A(n2385), .B(n2384), .Z(n2386) );
  XNOR U3586 ( .A(key[25]), .B(n2386), .Z(\w1[0][25] ) );
  NANDN U3587 ( .A(state[26]), .B(init), .Z(n2388) );
  OR U3588 ( .A(init), .B(msg[26]), .Z(n2387) );
  NAND U3589 ( .A(n2388), .B(n2387), .Z(n2389) );
  XNOR U3590 ( .A(key[26]), .B(n2389), .Z(\w1[0][26] ) );
  NANDN U3591 ( .A(state[27]), .B(init), .Z(n2391) );
  OR U3592 ( .A(init), .B(msg[27]), .Z(n2390) );
  NAND U3593 ( .A(n2391), .B(n2390), .Z(n2392) );
  XNOR U3594 ( .A(key[27]), .B(n2392), .Z(\w1[0][27] ) );
  NANDN U3595 ( .A(state[28]), .B(init), .Z(n2394) );
  OR U3596 ( .A(init), .B(msg[28]), .Z(n2393) );
  NAND U3597 ( .A(n2394), .B(n2393), .Z(n2395) );
  XNOR U3598 ( .A(key[28]), .B(n2395), .Z(\w1[0][28] ) );
  NANDN U3599 ( .A(state[29]), .B(init), .Z(n2397) );
  OR U3600 ( .A(init), .B(msg[29]), .Z(n2396) );
  NAND U3601 ( .A(n2397), .B(n2396), .Z(n2398) );
  XNOR U3602 ( .A(key[29]), .B(n2398), .Z(\w1[0][29] ) );
  NANDN U3603 ( .A(state[2]), .B(init), .Z(n2400) );
  OR U3604 ( .A(init), .B(msg[2]), .Z(n2399) );
  NAND U3605 ( .A(n2400), .B(n2399), .Z(n2401) );
  XNOR U3606 ( .A(key[2]), .B(n2401), .Z(\w1[0][2] ) );
  NANDN U3607 ( .A(state[30]), .B(init), .Z(n2403) );
  OR U3608 ( .A(init), .B(msg[30]), .Z(n2402) );
  NAND U3609 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3610 ( .A(key[30]), .B(n2404), .Z(\w1[0][30] ) );
  NANDN U3611 ( .A(state[31]), .B(init), .Z(n2406) );
  OR U3612 ( .A(init), .B(msg[31]), .Z(n2405) );
  NAND U3613 ( .A(n2406), .B(n2405), .Z(n2407) );
  XNOR U3614 ( .A(key[31]), .B(n2407), .Z(\w1[0][31] ) );
  NANDN U3615 ( .A(state[32]), .B(init), .Z(n2409) );
  OR U3616 ( .A(init), .B(msg[32]), .Z(n2408) );
  NAND U3617 ( .A(n2409), .B(n2408), .Z(n2410) );
  XNOR U3618 ( .A(key[32]), .B(n2410), .Z(\w1[0][32] ) );
  NANDN U3619 ( .A(state[33]), .B(init), .Z(n2412) );
  OR U3620 ( .A(init), .B(msg[33]), .Z(n2411) );
  NAND U3621 ( .A(n2412), .B(n2411), .Z(n2413) );
  XNOR U3622 ( .A(key[33]), .B(n2413), .Z(\w1[0][33] ) );
  NANDN U3623 ( .A(state[34]), .B(init), .Z(n2415) );
  OR U3624 ( .A(init), .B(msg[34]), .Z(n2414) );
  NAND U3625 ( .A(n2415), .B(n2414), .Z(n2416) );
  XNOR U3626 ( .A(key[34]), .B(n2416), .Z(\w1[0][34] ) );
  NANDN U3627 ( .A(state[35]), .B(init), .Z(n2418) );
  OR U3628 ( .A(init), .B(msg[35]), .Z(n2417) );
  NAND U3629 ( .A(n2418), .B(n2417), .Z(n2419) );
  XNOR U3630 ( .A(key[35]), .B(n2419), .Z(\w1[0][35] ) );
  NANDN U3631 ( .A(state[36]), .B(init), .Z(n2421) );
  OR U3632 ( .A(init), .B(msg[36]), .Z(n2420) );
  NAND U3633 ( .A(n2421), .B(n2420), .Z(n2422) );
  XNOR U3634 ( .A(key[36]), .B(n2422), .Z(\w1[0][36] ) );
  NANDN U3635 ( .A(state[37]), .B(init), .Z(n2424) );
  OR U3636 ( .A(init), .B(msg[37]), .Z(n2423) );
  NAND U3637 ( .A(n2424), .B(n2423), .Z(n2425) );
  XNOR U3638 ( .A(key[37]), .B(n2425), .Z(\w1[0][37] ) );
  NANDN U3639 ( .A(state[38]), .B(init), .Z(n2427) );
  OR U3640 ( .A(init), .B(msg[38]), .Z(n2426) );
  NAND U3641 ( .A(n2427), .B(n2426), .Z(n2428) );
  XNOR U3642 ( .A(key[38]), .B(n2428), .Z(\w1[0][38] ) );
  NANDN U3643 ( .A(state[39]), .B(init), .Z(n2430) );
  OR U3644 ( .A(init), .B(msg[39]), .Z(n2429) );
  NAND U3645 ( .A(n2430), .B(n2429), .Z(n2431) );
  XNOR U3646 ( .A(key[39]), .B(n2431), .Z(\w1[0][39] ) );
  NANDN U3647 ( .A(state[3]), .B(init), .Z(n2433) );
  OR U3648 ( .A(init), .B(msg[3]), .Z(n2432) );
  NAND U3649 ( .A(n2433), .B(n2432), .Z(n2434) );
  XNOR U3650 ( .A(key[3]), .B(n2434), .Z(\w1[0][3] ) );
  NANDN U3651 ( .A(state[40]), .B(init), .Z(n2436) );
  OR U3652 ( .A(init), .B(msg[40]), .Z(n2435) );
  NAND U3653 ( .A(n2436), .B(n2435), .Z(n2437) );
  XNOR U3654 ( .A(key[40]), .B(n2437), .Z(\w1[0][40] ) );
  NANDN U3655 ( .A(state[41]), .B(init), .Z(n2439) );
  OR U3656 ( .A(init), .B(msg[41]), .Z(n2438) );
  NAND U3657 ( .A(n2439), .B(n2438), .Z(n2440) );
  XNOR U3658 ( .A(key[41]), .B(n2440), .Z(\w1[0][41] ) );
  NANDN U3659 ( .A(state[42]), .B(init), .Z(n2442) );
  OR U3660 ( .A(init), .B(msg[42]), .Z(n2441) );
  NAND U3661 ( .A(n2442), .B(n2441), .Z(n2443) );
  XNOR U3662 ( .A(key[42]), .B(n2443), .Z(\w1[0][42] ) );
  NANDN U3663 ( .A(state[43]), .B(init), .Z(n2445) );
  OR U3664 ( .A(init), .B(msg[43]), .Z(n2444) );
  NAND U3665 ( .A(n2445), .B(n2444), .Z(n2446) );
  XNOR U3666 ( .A(key[43]), .B(n2446), .Z(\w1[0][43] ) );
  NANDN U3667 ( .A(state[44]), .B(init), .Z(n2448) );
  OR U3668 ( .A(init), .B(msg[44]), .Z(n2447) );
  NAND U3669 ( .A(n2448), .B(n2447), .Z(n2449) );
  XNOR U3670 ( .A(key[44]), .B(n2449), .Z(\w1[0][44] ) );
  NANDN U3671 ( .A(state[45]), .B(init), .Z(n2451) );
  OR U3672 ( .A(init), .B(msg[45]), .Z(n2450) );
  NAND U3673 ( .A(n2451), .B(n2450), .Z(n2452) );
  XNOR U3674 ( .A(key[45]), .B(n2452), .Z(\w1[0][45] ) );
  NANDN U3675 ( .A(state[46]), .B(init), .Z(n2454) );
  OR U3676 ( .A(init), .B(msg[46]), .Z(n2453) );
  NAND U3677 ( .A(n2454), .B(n2453), .Z(n2455) );
  XNOR U3678 ( .A(key[46]), .B(n2455), .Z(\w1[0][46] ) );
  NANDN U3679 ( .A(state[47]), .B(init), .Z(n2457) );
  OR U3680 ( .A(init), .B(msg[47]), .Z(n2456) );
  NAND U3681 ( .A(n2457), .B(n2456), .Z(n2458) );
  XNOR U3682 ( .A(key[47]), .B(n2458), .Z(\w1[0][47] ) );
  NANDN U3683 ( .A(state[48]), .B(init), .Z(n2460) );
  OR U3684 ( .A(init), .B(msg[48]), .Z(n2459) );
  NAND U3685 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3686 ( .A(key[48]), .B(n2461), .Z(\w1[0][48] ) );
  NANDN U3687 ( .A(state[49]), .B(init), .Z(n2463) );
  OR U3688 ( .A(init), .B(msg[49]), .Z(n2462) );
  NAND U3689 ( .A(n2463), .B(n2462), .Z(n2464) );
  XNOR U3690 ( .A(key[49]), .B(n2464), .Z(\w1[0][49] ) );
  NANDN U3691 ( .A(state[4]), .B(init), .Z(n2466) );
  OR U3692 ( .A(init), .B(msg[4]), .Z(n2465) );
  NAND U3693 ( .A(n2466), .B(n2465), .Z(n2467) );
  XNOR U3694 ( .A(key[4]), .B(n2467), .Z(\w1[0][4] ) );
  NANDN U3695 ( .A(state[50]), .B(init), .Z(n2469) );
  OR U3696 ( .A(init), .B(msg[50]), .Z(n2468) );
  NAND U3697 ( .A(n2469), .B(n2468), .Z(n2470) );
  XNOR U3698 ( .A(key[50]), .B(n2470), .Z(\w1[0][50] ) );
  NANDN U3699 ( .A(state[51]), .B(init), .Z(n2472) );
  OR U3700 ( .A(init), .B(msg[51]), .Z(n2471) );
  NAND U3701 ( .A(n2472), .B(n2471), .Z(n2473) );
  XNOR U3702 ( .A(key[51]), .B(n2473), .Z(\w1[0][51] ) );
  NANDN U3703 ( .A(state[52]), .B(init), .Z(n2475) );
  OR U3704 ( .A(init), .B(msg[52]), .Z(n2474) );
  NAND U3705 ( .A(n2475), .B(n2474), .Z(n2476) );
  XNOR U3706 ( .A(key[52]), .B(n2476), .Z(\w1[0][52] ) );
  NANDN U3707 ( .A(state[53]), .B(init), .Z(n2478) );
  OR U3708 ( .A(init), .B(msg[53]), .Z(n2477) );
  NAND U3709 ( .A(n2478), .B(n2477), .Z(n2479) );
  XNOR U3710 ( .A(key[53]), .B(n2479), .Z(\w1[0][53] ) );
  NANDN U3711 ( .A(state[54]), .B(init), .Z(n2481) );
  OR U3712 ( .A(init), .B(msg[54]), .Z(n2480) );
  NAND U3713 ( .A(n2481), .B(n2480), .Z(n2482) );
  XNOR U3714 ( .A(key[54]), .B(n2482), .Z(\w1[0][54] ) );
  NANDN U3715 ( .A(state[55]), .B(init), .Z(n2484) );
  OR U3716 ( .A(init), .B(msg[55]), .Z(n2483) );
  NAND U3717 ( .A(n2484), .B(n2483), .Z(n2485) );
  XNOR U3718 ( .A(key[55]), .B(n2485), .Z(\w1[0][55] ) );
  NANDN U3719 ( .A(state[56]), .B(init), .Z(n2487) );
  OR U3720 ( .A(init), .B(msg[56]), .Z(n2486) );
  NAND U3721 ( .A(n2487), .B(n2486), .Z(n2488) );
  XNOR U3722 ( .A(key[56]), .B(n2488), .Z(\w1[0][56] ) );
  NANDN U3723 ( .A(state[57]), .B(init), .Z(n2490) );
  OR U3724 ( .A(init), .B(msg[57]), .Z(n2489) );
  NAND U3725 ( .A(n2490), .B(n2489), .Z(n2491) );
  XNOR U3726 ( .A(key[57]), .B(n2491), .Z(\w1[0][57] ) );
  NANDN U3727 ( .A(state[58]), .B(init), .Z(n2493) );
  OR U3728 ( .A(init), .B(msg[58]), .Z(n2492) );
  NAND U3729 ( .A(n2493), .B(n2492), .Z(n2494) );
  XNOR U3730 ( .A(key[58]), .B(n2494), .Z(\w1[0][58] ) );
  NANDN U3731 ( .A(state[59]), .B(init), .Z(n2496) );
  OR U3732 ( .A(init), .B(msg[59]), .Z(n2495) );
  NAND U3733 ( .A(n2496), .B(n2495), .Z(n2497) );
  XNOR U3734 ( .A(key[59]), .B(n2497), .Z(\w1[0][59] ) );
  NANDN U3735 ( .A(state[5]), .B(init), .Z(n2499) );
  OR U3736 ( .A(init), .B(msg[5]), .Z(n2498) );
  NAND U3737 ( .A(n2499), .B(n2498), .Z(n2500) );
  XNOR U3738 ( .A(key[5]), .B(n2500), .Z(\w1[0][5] ) );
  NANDN U3739 ( .A(state[60]), .B(init), .Z(n2502) );
  OR U3740 ( .A(init), .B(msg[60]), .Z(n2501) );
  NAND U3741 ( .A(n2502), .B(n2501), .Z(n2503) );
  XNOR U3742 ( .A(key[60]), .B(n2503), .Z(\w1[0][60] ) );
  NANDN U3743 ( .A(state[61]), .B(init), .Z(n2505) );
  OR U3744 ( .A(init), .B(msg[61]), .Z(n2504) );
  NAND U3745 ( .A(n2505), .B(n2504), .Z(n2506) );
  XNOR U3746 ( .A(key[61]), .B(n2506), .Z(\w1[0][61] ) );
  NANDN U3747 ( .A(state[62]), .B(init), .Z(n2508) );
  OR U3748 ( .A(init), .B(msg[62]), .Z(n2507) );
  NAND U3749 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3750 ( .A(key[62]), .B(n2509), .Z(\w1[0][62] ) );
  NANDN U3751 ( .A(state[63]), .B(init), .Z(n2511) );
  OR U3752 ( .A(init), .B(msg[63]), .Z(n2510) );
  NAND U3753 ( .A(n2511), .B(n2510), .Z(n2512) );
  XNOR U3754 ( .A(key[63]), .B(n2512), .Z(\w1[0][63] ) );
  NANDN U3755 ( .A(state[64]), .B(init), .Z(n2514) );
  OR U3756 ( .A(init), .B(msg[64]), .Z(n2513) );
  NAND U3757 ( .A(n2514), .B(n2513), .Z(n2515) );
  XNOR U3758 ( .A(key[64]), .B(n2515), .Z(\w1[0][64] ) );
  NANDN U3759 ( .A(state[65]), .B(init), .Z(n2517) );
  OR U3760 ( .A(init), .B(msg[65]), .Z(n2516) );
  NAND U3761 ( .A(n2517), .B(n2516), .Z(n2518) );
  XNOR U3762 ( .A(key[65]), .B(n2518), .Z(\w1[0][65] ) );
  NANDN U3763 ( .A(state[66]), .B(init), .Z(n2520) );
  OR U3764 ( .A(init), .B(msg[66]), .Z(n2519) );
  NAND U3765 ( .A(n2520), .B(n2519), .Z(n2521) );
  XNOR U3766 ( .A(key[66]), .B(n2521), .Z(\w1[0][66] ) );
  NANDN U3767 ( .A(state[67]), .B(init), .Z(n2523) );
  OR U3768 ( .A(init), .B(msg[67]), .Z(n2522) );
  NAND U3769 ( .A(n2523), .B(n2522), .Z(n2524) );
  XNOR U3770 ( .A(key[67]), .B(n2524), .Z(\w1[0][67] ) );
  NANDN U3771 ( .A(state[68]), .B(init), .Z(n2526) );
  OR U3772 ( .A(init), .B(msg[68]), .Z(n2525) );
  NAND U3773 ( .A(n2526), .B(n2525), .Z(n2527) );
  XNOR U3774 ( .A(key[68]), .B(n2527), .Z(\w1[0][68] ) );
  NANDN U3775 ( .A(state[69]), .B(init), .Z(n2529) );
  OR U3776 ( .A(init), .B(msg[69]), .Z(n2528) );
  NAND U3777 ( .A(n2529), .B(n2528), .Z(n2530) );
  XNOR U3778 ( .A(key[69]), .B(n2530), .Z(\w1[0][69] ) );
  NANDN U3779 ( .A(state[6]), .B(init), .Z(n2532) );
  OR U3780 ( .A(init), .B(msg[6]), .Z(n2531) );
  NAND U3781 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3782 ( .A(key[6]), .B(n2533), .Z(\w1[0][6] ) );
  NANDN U3783 ( .A(state[70]), .B(init), .Z(n2535) );
  OR U3784 ( .A(init), .B(msg[70]), .Z(n2534) );
  NAND U3785 ( .A(n2535), .B(n2534), .Z(n2536) );
  XNOR U3786 ( .A(key[70]), .B(n2536), .Z(\w1[0][70] ) );
  NANDN U3787 ( .A(state[71]), .B(init), .Z(n2538) );
  OR U3788 ( .A(init), .B(msg[71]), .Z(n2537) );
  NAND U3789 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3790 ( .A(key[71]), .B(n2539), .Z(\w1[0][71] ) );
  NANDN U3791 ( .A(state[72]), .B(init), .Z(n2541) );
  OR U3792 ( .A(init), .B(msg[72]), .Z(n2540) );
  NAND U3793 ( .A(n2541), .B(n2540), .Z(n2542) );
  XNOR U3794 ( .A(key[72]), .B(n2542), .Z(\w1[0][72] ) );
  NANDN U3795 ( .A(state[73]), .B(init), .Z(n2544) );
  OR U3796 ( .A(init), .B(msg[73]), .Z(n2543) );
  NAND U3797 ( .A(n2544), .B(n2543), .Z(n2545) );
  XNOR U3798 ( .A(key[73]), .B(n2545), .Z(\w1[0][73] ) );
  NANDN U3799 ( .A(state[74]), .B(init), .Z(n2547) );
  OR U3800 ( .A(init), .B(msg[74]), .Z(n2546) );
  NAND U3801 ( .A(n2547), .B(n2546), .Z(n2548) );
  XNOR U3802 ( .A(key[74]), .B(n2548), .Z(\w1[0][74] ) );
  NANDN U3803 ( .A(state[75]), .B(init), .Z(n2550) );
  OR U3804 ( .A(init), .B(msg[75]), .Z(n2549) );
  NAND U3805 ( .A(n2550), .B(n2549), .Z(n2551) );
  XNOR U3806 ( .A(key[75]), .B(n2551), .Z(\w1[0][75] ) );
  NANDN U3807 ( .A(state[76]), .B(init), .Z(n2553) );
  OR U3808 ( .A(init), .B(msg[76]), .Z(n2552) );
  NAND U3809 ( .A(n2553), .B(n2552), .Z(n2554) );
  XNOR U3810 ( .A(key[76]), .B(n2554), .Z(\w1[0][76] ) );
  NANDN U3811 ( .A(state[77]), .B(init), .Z(n2556) );
  OR U3812 ( .A(init), .B(msg[77]), .Z(n2555) );
  NAND U3813 ( .A(n2556), .B(n2555), .Z(n2557) );
  XNOR U3814 ( .A(key[77]), .B(n2557), .Z(\w1[0][77] ) );
  NANDN U3815 ( .A(state[78]), .B(init), .Z(n2559) );
  OR U3816 ( .A(init), .B(msg[78]), .Z(n2558) );
  NAND U3817 ( .A(n2559), .B(n2558), .Z(n2560) );
  XNOR U3818 ( .A(key[78]), .B(n2560), .Z(\w1[0][78] ) );
  NANDN U3819 ( .A(state[79]), .B(init), .Z(n2562) );
  OR U3820 ( .A(init), .B(msg[79]), .Z(n2561) );
  NAND U3821 ( .A(n2562), .B(n2561), .Z(n2563) );
  XNOR U3822 ( .A(key[79]), .B(n2563), .Z(\w1[0][79] ) );
  NANDN U3823 ( .A(state[7]), .B(init), .Z(n2565) );
  OR U3824 ( .A(init), .B(msg[7]), .Z(n2564) );
  NAND U3825 ( .A(n2565), .B(n2564), .Z(n2566) );
  XNOR U3826 ( .A(key[7]), .B(n2566), .Z(\w1[0][7] ) );
  NANDN U3827 ( .A(state[80]), .B(init), .Z(n2568) );
  OR U3828 ( .A(init), .B(msg[80]), .Z(n2567) );
  NAND U3829 ( .A(n2568), .B(n2567), .Z(n2569) );
  XNOR U3830 ( .A(key[80]), .B(n2569), .Z(\w1[0][80] ) );
  NANDN U3831 ( .A(state[81]), .B(init), .Z(n2571) );
  OR U3832 ( .A(init), .B(msg[81]), .Z(n2570) );
  NAND U3833 ( .A(n2571), .B(n2570), .Z(n2572) );
  XNOR U3834 ( .A(key[81]), .B(n2572), .Z(\w1[0][81] ) );
  NANDN U3835 ( .A(state[82]), .B(init), .Z(n2574) );
  OR U3836 ( .A(init), .B(msg[82]), .Z(n2573) );
  NAND U3837 ( .A(n2574), .B(n2573), .Z(n2575) );
  XNOR U3838 ( .A(key[82]), .B(n2575), .Z(\w1[0][82] ) );
  NANDN U3839 ( .A(state[83]), .B(init), .Z(n2577) );
  OR U3840 ( .A(init), .B(msg[83]), .Z(n2576) );
  NAND U3841 ( .A(n2577), .B(n2576), .Z(n2578) );
  XNOR U3842 ( .A(key[83]), .B(n2578), .Z(\w1[0][83] ) );
  NANDN U3843 ( .A(state[84]), .B(init), .Z(n2580) );
  OR U3844 ( .A(init), .B(msg[84]), .Z(n2579) );
  NAND U3845 ( .A(n2580), .B(n2579), .Z(n2581) );
  XNOR U3846 ( .A(key[84]), .B(n2581), .Z(\w1[0][84] ) );
  NANDN U3847 ( .A(state[85]), .B(init), .Z(n2583) );
  OR U3848 ( .A(init), .B(msg[85]), .Z(n2582) );
  NAND U3849 ( .A(n2583), .B(n2582), .Z(n2584) );
  XNOR U3850 ( .A(key[85]), .B(n2584), .Z(\w1[0][85] ) );
  NANDN U3851 ( .A(state[86]), .B(init), .Z(n2586) );
  OR U3852 ( .A(init), .B(msg[86]), .Z(n2585) );
  NAND U3853 ( .A(n2586), .B(n2585), .Z(n2587) );
  XNOR U3854 ( .A(key[86]), .B(n2587), .Z(\w1[0][86] ) );
  NANDN U3855 ( .A(state[87]), .B(init), .Z(n2589) );
  OR U3856 ( .A(init), .B(msg[87]), .Z(n2588) );
  NAND U3857 ( .A(n2589), .B(n2588), .Z(n2590) );
  XNOR U3858 ( .A(key[87]), .B(n2590), .Z(\w1[0][87] ) );
  NANDN U3859 ( .A(state[88]), .B(init), .Z(n2592) );
  OR U3860 ( .A(init), .B(msg[88]), .Z(n2591) );
  NAND U3861 ( .A(n2592), .B(n2591), .Z(n2593) );
  XNOR U3862 ( .A(key[88]), .B(n2593), .Z(\w1[0][88] ) );
  NANDN U3863 ( .A(state[89]), .B(init), .Z(n2595) );
  OR U3864 ( .A(init), .B(msg[89]), .Z(n2594) );
  NAND U3865 ( .A(n2595), .B(n2594), .Z(n2596) );
  XNOR U3866 ( .A(key[89]), .B(n2596), .Z(\w1[0][89] ) );
  NANDN U3867 ( .A(state[8]), .B(init), .Z(n2598) );
  OR U3868 ( .A(init), .B(msg[8]), .Z(n2597) );
  NAND U3869 ( .A(n2598), .B(n2597), .Z(n2599) );
  XNOR U3870 ( .A(key[8]), .B(n2599), .Z(\w1[0][8] ) );
  NANDN U3871 ( .A(state[90]), .B(init), .Z(n2601) );
  OR U3872 ( .A(init), .B(msg[90]), .Z(n2600) );
  NAND U3873 ( .A(n2601), .B(n2600), .Z(n2602) );
  XNOR U3874 ( .A(key[90]), .B(n2602), .Z(\w1[0][90] ) );
  NANDN U3875 ( .A(state[91]), .B(init), .Z(n2604) );
  OR U3876 ( .A(init), .B(msg[91]), .Z(n2603) );
  NAND U3877 ( .A(n2604), .B(n2603), .Z(n2605) );
  XNOR U3878 ( .A(key[91]), .B(n2605), .Z(\w1[0][91] ) );
  NANDN U3879 ( .A(state[92]), .B(init), .Z(n2607) );
  OR U3880 ( .A(init), .B(msg[92]), .Z(n2606) );
  NAND U3881 ( .A(n2607), .B(n2606), .Z(n2608) );
  XNOR U3882 ( .A(key[92]), .B(n2608), .Z(\w1[0][92] ) );
  NANDN U3883 ( .A(state[93]), .B(init), .Z(n2610) );
  OR U3884 ( .A(init), .B(msg[93]), .Z(n2609) );
  NAND U3885 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3886 ( .A(key[93]), .B(n2611), .Z(\w1[0][93] ) );
  NANDN U3887 ( .A(state[94]), .B(init), .Z(n2613) );
  OR U3888 ( .A(init), .B(msg[94]), .Z(n2612) );
  NAND U3889 ( .A(n2613), .B(n2612), .Z(n2614) );
  XNOR U3890 ( .A(key[94]), .B(n2614), .Z(\w1[0][94] ) );
  NANDN U3891 ( .A(state[95]), .B(init), .Z(n2616) );
  OR U3892 ( .A(init), .B(msg[95]), .Z(n2615) );
  NAND U3893 ( .A(n2616), .B(n2615), .Z(n2617) );
  XNOR U3894 ( .A(key[95]), .B(n2617), .Z(\w1[0][95] ) );
  NANDN U3895 ( .A(state[96]), .B(init), .Z(n2619) );
  OR U3896 ( .A(init), .B(msg[96]), .Z(n2618) );
  NAND U3897 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3898 ( .A(key[96]), .B(n2620), .Z(\w1[0][96] ) );
  NANDN U3899 ( .A(state[97]), .B(init), .Z(n2622) );
  OR U3900 ( .A(init), .B(msg[97]), .Z(n2621) );
  NAND U3901 ( .A(n2622), .B(n2621), .Z(n2623) );
  XNOR U3902 ( .A(key[97]), .B(n2623), .Z(\w1[0][97] ) );
  NANDN U3903 ( .A(state[98]), .B(init), .Z(n2625) );
  OR U3904 ( .A(init), .B(msg[98]), .Z(n2624) );
  NAND U3905 ( .A(n2625), .B(n2624), .Z(n2626) );
  XNOR U3906 ( .A(key[98]), .B(n2626), .Z(\w1[0][98] ) );
  NANDN U3907 ( .A(state[99]), .B(init), .Z(n2628) );
  OR U3908 ( .A(init), .B(msg[99]), .Z(n2627) );
  NAND U3909 ( .A(n2628), .B(n2627), .Z(n2629) );
  XNOR U3910 ( .A(key[99]), .B(n2629), .Z(\w1[0][99] ) );
  NANDN U3911 ( .A(state[9]), .B(init), .Z(n2631) );
  OR U3912 ( .A(init), .B(msg[9]), .Z(n2630) );
  NAND U3913 ( .A(n2631), .B(n2630), .Z(n2632) );
  XNOR U3914 ( .A(key[9]), .B(n2632), .Z(\w1[0][9] ) );
  XOR U3915 ( .A(\w3[0][8] ), .B(key[128]), .Z(n2634) );
  XOR U3916 ( .A(\w3[0][1] ), .B(\w3[0][25] ), .Z(n3056) );
  XOR U3917 ( .A(\w3[0][16] ), .B(\w3[0][24] ), .Z(n3012) );
  XNOR U3918 ( .A(n3056), .B(n3012), .Z(n2633) );
  XNOR U3919 ( .A(n2634), .B(n2633), .Z(\w1[1][0] ) );
  XOR U3920 ( .A(\w3[0][96] ), .B(\w3[0][101] ), .Z(n2660) );
  XOR U3921 ( .A(n2660), .B(key[228]), .Z(n2638) );
  XOR U3922 ( .A(\w3[0][116] ), .B(\w3[0][125] ), .Z(n2636) );
  XNOR U3923 ( .A(\w3[0][120] ), .B(\w3[0][108] ), .Z(n2635) );
  XNOR U3924 ( .A(n2636), .B(n2635), .Z(n2717) );
  XNOR U3925 ( .A(\w3[0][124] ), .B(n2717), .Z(n2637) );
  XNOR U3926 ( .A(n2638), .B(n2637), .Z(\w1[1][100] ) );
  XOR U3927 ( .A(\w3[0][102] ), .B(\w3[0][126] ), .Z(n2669) );
  XOR U3928 ( .A(n2669), .B(key[229]), .Z(n2640) );
  XOR U3929 ( .A(\w3[0][109] ), .B(\w3[0][117] ), .Z(n2720) );
  XNOR U3930 ( .A(\w3[0][125] ), .B(n2720), .Z(n2639) );
  XNOR U3931 ( .A(n2640), .B(n2639), .Z(\w1[1][101] ) );
  XOR U3932 ( .A(\w3[0][96] ), .B(\w3[0][103] ), .Z(n2670) );
  XOR U3933 ( .A(n2670), .B(key[230]), .Z(n2642) );
  XOR U3934 ( .A(\w3[0][110] ), .B(\w3[0][118] ), .Z(n2688) );
  XNOR U3935 ( .A(\w3[0][120] ), .B(\w3[0][127] ), .Z(n2644) );
  XNOR U3936 ( .A(n2688), .B(n2644), .Z(n2725) );
  XNOR U3937 ( .A(\w3[0][126] ), .B(n2725), .Z(n2641) );
  XNOR U3938 ( .A(n2642), .B(n2641), .Z(\w1[1][102] ) );
  XOR U3939 ( .A(\w3[0][111] ), .B(\w3[0][119] ), .Z(n2728) );
  XNOR U3940 ( .A(n2728), .B(key[231]), .Z(n2643) );
  XNOR U3941 ( .A(n2644), .B(n2643), .Z(n2645) );
  XNOR U3942 ( .A(\w3[0][96] ), .B(n2645), .Z(\w1[1][103] ) );
  XOR U3943 ( .A(key[232]), .B(\w3[0][105] ), .Z(n2647) );
  XNOR U3944 ( .A(\w3[0][96] ), .B(\w3[0][97] ), .Z(n2646) );
  XNOR U3945 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3946 ( .A(\w3[0][120] ), .B(\w3[0][112] ), .Z(n3038) );
  XNOR U3947 ( .A(n2648), .B(n3038), .Z(\w1[1][104] ) );
  XOR U3948 ( .A(\w3[0][106] ), .B(\w3[0][98] ), .Z(n2650) );
  XOR U3949 ( .A(\w3[0][97] ), .B(\w3[0][121] ), .Z(n3037) );
  XNOR U3950 ( .A(n3037), .B(key[233]), .Z(n2649) );
  XNOR U3951 ( .A(n2650), .B(n2649), .Z(n2651) );
  XOR U3952 ( .A(\w3[0][113] ), .B(n2651), .Z(\w1[1][105] ) );
  XOR U3953 ( .A(\w3[0][107] ), .B(\w3[0][114] ), .Z(n2653) );
  XOR U3954 ( .A(\w3[0][98] ), .B(\w3[0][122] ), .Z(n3042) );
  XNOR U3955 ( .A(n3042), .B(key[234]), .Z(n2652) );
  XNOR U3956 ( .A(n2653), .B(n2652), .Z(n2654) );
  XOR U3957 ( .A(\w3[0][99] ), .B(n2654), .Z(\w1[1][106] ) );
  XOR U3958 ( .A(\w3[0][99] ), .B(\w3[0][123] ), .Z(n3046) );
  XNOR U3959 ( .A(\w3[0][108] ), .B(n3046), .Z(n2655) );
  XNOR U3960 ( .A(\w3[0][104] ), .B(n2655), .Z(n2681) );
  XOR U3961 ( .A(n2681), .B(key[235]), .Z(n2657) );
  XOR U3962 ( .A(\w3[0][96] ), .B(\w3[0][100] ), .Z(n3050) );
  XNOR U3963 ( .A(\w3[0][115] ), .B(n3050), .Z(n2656) );
  XNOR U3964 ( .A(n2657), .B(n2656), .Z(\w1[1][107] ) );
  XOR U3965 ( .A(\w3[0][100] ), .B(\w3[0][104] ), .Z(n2659) );
  XNOR U3966 ( .A(\w3[0][124] ), .B(\w3[0][109] ), .Z(n2658) );
  XNOR U3967 ( .A(n2659), .B(n2658), .Z(n2684) );
  XOR U3968 ( .A(n2684), .B(key[236]), .Z(n2662) );
  XNOR U3969 ( .A(\w3[0][116] ), .B(n2660), .Z(n2661) );
  XNOR U3970 ( .A(n2662), .B(n2661), .Z(\w1[1][108] ) );
  XOR U3971 ( .A(\w3[0][125] ), .B(\w3[0][101] ), .Z(n2687) );
  XOR U3972 ( .A(n2687), .B(key[237]), .Z(n2664) );
  XNOR U3973 ( .A(\w3[0][102] ), .B(\w3[0][110] ), .Z(n2663) );
  XNOR U3974 ( .A(n2664), .B(n2663), .Z(n2665) );
  XOR U3975 ( .A(\w3[0][117] ), .B(n2665), .Z(\w1[1][109] ) );
  XOR U3976 ( .A(\w3[0][11] ), .B(\w3[0][18] ), .Z(n2667) );
  XOR U3977 ( .A(\w3[0][2] ), .B(\w3[0][26] ), .Z(n2751) );
  XNOR U3978 ( .A(n2751), .B(key[138]), .Z(n2666) );
  XNOR U3979 ( .A(n2667), .B(n2666), .Z(n2668) );
  XOR U3980 ( .A(\w3[0][3] ), .B(n2668), .Z(\w1[1][10] ) );
  XNOR U3981 ( .A(\w3[0][111] ), .B(\w3[0][104] ), .Z(n2696) );
  XNOR U3982 ( .A(n2669), .B(n2696), .Z(n2691) );
  XOR U3983 ( .A(n2691), .B(key[238]), .Z(n2672) );
  XNOR U3984 ( .A(\w3[0][118] ), .B(n2670), .Z(n2671) );
  XNOR U3985 ( .A(n2672), .B(n2671), .Z(\w1[1][110] ) );
  XOR U3986 ( .A(\w3[0][127] ), .B(\w3[0][103] ), .Z(n2694) );
  XOR U3987 ( .A(n2694), .B(key[239]), .Z(n2674) );
  XOR U3988 ( .A(\w3[0][96] ), .B(\w3[0][104] ), .Z(n2701) );
  XNOR U3989 ( .A(\w3[0][119] ), .B(n2701), .Z(n2673) );
  XNOR U3990 ( .A(n2674), .B(n2673), .Z(\w1[1][111] ) );
  XOR U3991 ( .A(\w3[0][105] ), .B(\w3[0][113] ), .Z(n3041) );
  XOR U3992 ( .A(n3041), .B(key[240]), .Z(n2676) );
  XNOR U3993 ( .A(\w3[0][120] ), .B(n2701), .Z(n2675) );
  XNOR U3994 ( .A(n2676), .B(n2675), .Z(\w1[1][112] ) );
  XOR U3995 ( .A(\w3[0][106] ), .B(\w3[0][114] ), .Z(n3045) );
  XOR U3996 ( .A(n3045), .B(key[241]), .Z(n2678) );
  XNOR U3997 ( .A(\w3[0][105] ), .B(n3037), .Z(n2677) );
  XNOR U3998 ( .A(n2678), .B(n2677), .Z(\w1[1][113] ) );
  XOR U3999 ( .A(\w3[0][107] ), .B(\w3[0][115] ), .Z(n2712) );
  XOR U4000 ( .A(n2712), .B(key[242]), .Z(n2680) );
  XNOR U4001 ( .A(\w3[0][106] ), .B(n3042), .Z(n2679) );
  XNOR U4002 ( .A(n2680), .B(n2679), .Z(\w1[1][114] ) );
  XOR U4003 ( .A(\w3[0][116] ), .B(\w3[0][112] ), .Z(n2713) );
  XOR U4004 ( .A(n2713), .B(key[243]), .Z(n2683) );
  XNOR U4005 ( .A(\w3[0][107] ), .B(n2681), .Z(n2682) );
  XNOR U4006 ( .A(n2683), .B(n2682), .Z(\w1[1][115] ) );
  XOR U4007 ( .A(\w3[0][117] ), .B(\w3[0][112] ), .Z(n2716) );
  XOR U4008 ( .A(n2716), .B(key[244]), .Z(n2686) );
  XNOR U4009 ( .A(\w3[0][108] ), .B(n2684), .Z(n2685) );
  XNOR U4010 ( .A(n2686), .B(n2685), .Z(\w1[1][116] ) );
  XOR U4011 ( .A(n2687), .B(key[245]), .Z(n2690) );
  XNOR U4012 ( .A(\w3[0][109] ), .B(n2688), .Z(n2689) );
  XNOR U4013 ( .A(n2690), .B(n2689), .Z(\w1[1][117] ) );
  XOR U4014 ( .A(\w3[0][119] ), .B(\w3[0][112] ), .Z(n2724) );
  XOR U4015 ( .A(n2724), .B(key[246]), .Z(n2693) );
  XNOR U4016 ( .A(\w3[0][110] ), .B(n2691), .Z(n2692) );
  XNOR U4017 ( .A(n2693), .B(n2692), .Z(\w1[1][118] ) );
  XNOR U4018 ( .A(n2694), .B(key[247]), .Z(n2695) );
  XNOR U4019 ( .A(n2696), .B(n2695), .Z(n2697) );
  XNOR U4020 ( .A(\w3[0][112] ), .B(n2697), .Z(\w1[1][119] ) );
  XOR U4021 ( .A(\w3[0][3] ), .B(\w3[0][27] ), .Z(n2792) );
  XNOR U4022 ( .A(\w3[0][8] ), .B(\w3[0][12] ), .Z(n2698) );
  XNOR U4023 ( .A(n2792), .B(n2698), .Z(n2748) );
  XOR U4024 ( .A(n2748), .B(key[139]), .Z(n2700) );
  XOR U4025 ( .A(\w3[0][0] ), .B(\w3[0][4] ), .Z(n2822) );
  XNOR U4026 ( .A(\w3[0][19] ), .B(n2822), .Z(n2699) );
  XNOR U4027 ( .A(n2700), .B(n2699), .Z(\w1[1][11] ) );
  XOR U4028 ( .A(n2701), .B(key[248]), .Z(n2703) );
  XNOR U4029 ( .A(\w3[0][113] ), .B(\w3[0][121] ), .Z(n2702) );
  XNOR U4030 ( .A(n2703), .B(n2702), .Z(n2704) );
  XOR U4031 ( .A(\w3[0][112] ), .B(n2704), .Z(\w1[1][120] ) );
  XOR U4032 ( .A(n3041), .B(key[249]), .Z(n2706) );
  XNOR U4033 ( .A(\w3[0][122] ), .B(\w3[0][114] ), .Z(n2705) );
  XNOR U4034 ( .A(n2706), .B(n2705), .Z(n2707) );
  XOR U4035 ( .A(\w3[0][97] ), .B(n2707), .Z(\w1[1][121] ) );
  XOR U4036 ( .A(n3045), .B(key[250]), .Z(n2709) );
  XNOR U4037 ( .A(\w3[0][115] ), .B(\w3[0][123] ), .Z(n2708) );
  XNOR U4038 ( .A(n2709), .B(n2708), .Z(n2710) );
  XOR U4039 ( .A(\w3[0][98] ), .B(n2710), .Z(\w1[1][122] ) );
  XNOR U4040 ( .A(\w3[0][124] ), .B(\w3[0][120] ), .Z(n2711) );
  XNOR U4041 ( .A(n2712), .B(n2711), .Z(n3049) );
  XOR U4042 ( .A(n3049), .B(key[251]), .Z(n2715) );
  XNOR U4043 ( .A(\w3[0][99] ), .B(n2713), .Z(n2714) );
  XNOR U4044 ( .A(n2715), .B(n2714), .Z(\w1[1][123] ) );
  XOR U4045 ( .A(n2716), .B(key[252]), .Z(n2719) );
  XNOR U4046 ( .A(n2717), .B(\w3[0][100] ), .Z(n2718) );
  XNOR U4047 ( .A(n2719), .B(n2718), .Z(\w1[1][124] ) );
  XOR U4048 ( .A(\w3[0][118] ), .B(key[253]), .Z(n2722) );
  XNOR U4049 ( .A(n2720), .B(\w3[0][126] ), .Z(n2721) );
  XNOR U4050 ( .A(n2722), .B(n2721), .Z(n2723) );
  XOR U4051 ( .A(\w3[0][101] ), .B(n2723), .Z(\w1[1][125] ) );
  XOR U4052 ( .A(n2724), .B(key[254]), .Z(n2727) );
  XNOR U4053 ( .A(\w3[0][102] ), .B(n2725), .Z(n2726) );
  XNOR U4054 ( .A(n2727), .B(n2726), .Z(\w1[1][126] ) );
  XNOR U4055 ( .A(n2728), .B(key[255]), .Z(n2729) );
  XNOR U4056 ( .A(n3038), .B(n2729), .Z(n2730) );
  XNOR U4057 ( .A(\w3[0][103] ), .B(n2730), .Z(\w1[1][127] ) );
  XOR U4058 ( .A(\w3[0][13] ), .B(\w3[0][28] ), .Z(n2732) );
  XNOR U4059 ( .A(\w3[0][8] ), .B(\w3[0][4] ), .Z(n2731) );
  XNOR U4060 ( .A(n2732), .B(n2731), .Z(n2754) );
  XOR U4061 ( .A(n2754), .B(key[140]), .Z(n2734) );
  XOR U4062 ( .A(\w3[0][0] ), .B(\w3[0][5] ), .Z(n2859) );
  XNOR U4063 ( .A(\w3[0][20] ), .B(n2859), .Z(n2733) );
  XNOR U4064 ( .A(n2734), .B(n2733), .Z(\w1[1][12] ) );
  XOR U4065 ( .A(\w3[0][14] ), .B(\w3[0][21] ), .Z(n2736) );
  XOR U4066 ( .A(\w3[0][5] ), .B(\w3[0][29] ), .Z(n2757) );
  XNOR U4067 ( .A(n2757), .B(key[141]), .Z(n2735) );
  XNOR U4068 ( .A(n2736), .B(n2735), .Z(n2737) );
  XOR U4069 ( .A(\w3[0][6] ), .B(n2737), .Z(\w1[1][13] ) );
  XOR U4070 ( .A(\w3[0][6] ), .B(\w3[0][30] ), .Z(n2900) );
  XNOR U4071 ( .A(\w3[0][8] ), .B(\w3[0][15] ), .Z(n2765) );
  XNOR U4072 ( .A(n2900), .B(n2765), .Z(n2760) );
  XOR U4073 ( .A(n2760), .B(key[142]), .Z(n2739) );
  XOR U4074 ( .A(\w3[0][0] ), .B(\w3[0][7] ), .Z(n2935) );
  XNOR U4075 ( .A(\w3[0][22] ), .B(n2935), .Z(n2738) );
  XNOR U4076 ( .A(n2739), .B(n2738), .Z(\w1[1][14] ) );
  XOR U4077 ( .A(\w3[0][7] ), .B(\w3[0][31] ), .Z(n2763) );
  XOR U4078 ( .A(n2763), .B(key[143]), .Z(n2741) );
  XOR U4079 ( .A(\w3[0][8] ), .B(\w3[0][0] ), .Z(n2767) );
  XNOR U4080 ( .A(\w3[0][23] ), .B(n2767), .Z(n2740) );
  XNOR U4081 ( .A(n2741), .B(n2740), .Z(\w1[1][15] ) );
  XOR U4082 ( .A(\w3[0][17] ), .B(\w3[0][9] ), .Z(n2771) );
  XOR U4083 ( .A(n2771), .B(key[144]), .Z(n2743) );
  XNOR U4084 ( .A(\w3[0][24] ), .B(n2767), .Z(n2742) );
  XNOR U4085 ( .A(n2743), .B(n2742), .Z(\w1[1][16] ) );
  XOR U4086 ( .A(\w3[0][18] ), .B(\w3[0][10] ), .Z(n2791) );
  XOR U4087 ( .A(n2791), .B(key[145]), .Z(n2745) );
  XNOR U4088 ( .A(n3056), .B(\w3[0][9] ), .Z(n2744) );
  XNOR U4089 ( .A(n2745), .B(n2744), .Z(\w1[1][17] ) );
  XOR U4090 ( .A(\w3[0][11] ), .B(\w3[0][19] ), .Z(n2779) );
  XOR U4091 ( .A(n2779), .B(key[146]), .Z(n2747) );
  XNOR U4092 ( .A(n2751), .B(\w3[0][10] ), .Z(n2746) );
  XNOR U4093 ( .A(n2747), .B(n2746), .Z(\w1[1][18] ) );
  XOR U4094 ( .A(\w3[0][16] ), .B(\w3[0][20] ), .Z(n2780) );
  XOR U4095 ( .A(n2780), .B(key[147]), .Z(n2750) );
  XNOR U4096 ( .A(\w3[0][11] ), .B(n2748), .Z(n2749) );
  XNOR U4097 ( .A(n2750), .B(n2749), .Z(\w1[1][19] ) );
  XOR U4098 ( .A(n2771), .B(key[129]), .Z(n2753) );
  XNOR U4099 ( .A(\w3[0][25] ), .B(n2751), .Z(n2752) );
  XNOR U4100 ( .A(n2753), .B(n2752), .Z(\w1[1][1] ) );
  XOR U4101 ( .A(\w3[0][16] ), .B(\w3[0][21] ), .Z(n2785) );
  XOR U4102 ( .A(n2785), .B(key[148]), .Z(n2756) );
  XNOR U4103 ( .A(\w3[0][12] ), .B(n2754), .Z(n2755) );
  XNOR U4104 ( .A(n2756), .B(n2755), .Z(\w1[1][20] ) );
  XOR U4105 ( .A(\w3[0][14] ), .B(\w3[0][22] ), .Z(n2795) );
  XOR U4106 ( .A(n2795), .B(key[149]), .Z(n2759) );
  XNOR U4107 ( .A(\w3[0][13] ), .B(n2757), .Z(n2758) );
  XNOR U4108 ( .A(n2759), .B(n2758), .Z(\w1[1][21] ) );
  XOR U4109 ( .A(\w3[0][16] ), .B(\w3[0][23] ), .Z(n2796) );
  XOR U4110 ( .A(n2796), .B(key[150]), .Z(n2762) );
  XNOR U4111 ( .A(\w3[0][14] ), .B(n2760), .Z(n2761) );
  XNOR U4112 ( .A(n2762), .B(n2761), .Z(\w1[1][22] ) );
  XNOR U4113 ( .A(n2763), .B(key[151]), .Z(n2764) );
  XNOR U4114 ( .A(n2765), .B(n2764), .Z(n2766) );
  XNOR U4115 ( .A(\w3[0][16] ), .B(n2766), .Z(\w1[1][23] ) );
  XOR U4116 ( .A(\w3[0][17] ), .B(key[152]), .Z(n2769) );
  XNOR U4117 ( .A(\w3[0][25] ), .B(n2767), .Z(n2768) );
  XNOR U4118 ( .A(n2769), .B(n2768), .Z(n2770) );
  XOR U4119 ( .A(\w3[0][16] ), .B(n2770), .Z(\w1[1][24] ) );
  XOR U4120 ( .A(n2771), .B(key[153]), .Z(n2773) );
  XNOR U4121 ( .A(\w3[0][1] ), .B(\w3[0][26] ), .Z(n2772) );
  XNOR U4122 ( .A(n2773), .B(n2772), .Z(n2774) );
  XOR U4123 ( .A(\w3[0][18] ), .B(n2774), .Z(\w1[1][25] ) );
  XOR U4124 ( .A(n2791), .B(key[154]), .Z(n2776) );
  XNOR U4125 ( .A(\w3[0][2] ), .B(\w3[0][19] ), .Z(n2775) );
  XNOR U4126 ( .A(n2776), .B(n2775), .Z(n2777) );
  XOR U4127 ( .A(\w3[0][27] ), .B(n2777), .Z(\w1[1][26] ) );
  XNOR U4128 ( .A(\w3[0][24] ), .B(\w3[0][28] ), .Z(n2778) );
  XNOR U4129 ( .A(n2779), .B(n2778), .Z(n2821) );
  XOR U4130 ( .A(n2821), .B(key[155]), .Z(n2782) );
  XNOR U4131 ( .A(\w3[0][3] ), .B(n2780), .Z(n2781) );
  XNOR U4132 ( .A(n2782), .B(n2781), .Z(\w1[1][27] ) );
  XOR U4133 ( .A(\w3[0][20] ), .B(\w3[0][29] ), .Z(n2784) );
  XNOR U4134 ( .A(\w3[0][24] ), .B(\w3[0][12] ), .Z(n2783) );
  XNOR U4135 ( .A(n2784), .B(n2783), .Z(n2858) );
  XOR U4136 ( .A(n2858), .B(key[156]), .Z(n2787) );
  XNOR U4137 ( .A(\w3[0][4] ), .B(n2785), .Z(n2786) );
  XNOR U4138 ( .A(n2787), .B(n2786), .Z(\w1[1][28] ) );
  XOR U4139 ( .A(\w3[0][13] ), .B(\w3[0][21] ), .Z(n2899) );
  XOR U4140 ( .A(n2899), .B(key[157]), .Z(n2789) );
  XNOR U4141 ( .A(\w3[0][22] ), .B(\w3[0][30] ), .Z(n2788) );
  XNOR U4142 ( .A(n2789), .B(n2788), .Z(n2790) );
  XOR U4143 ( .A(\w3[0][5] ), .B(n2790), .Z(\w1[1][29] ) );
  XOR U4144 ( .A(n2791), .B(key[130]), .Z(n2794) );
  XNOR U4145 ( .A(\w3[0][26] ), .B(n2792), .Z(n2793) );
  XNOR U4146 ( .A(n2794), .B(n2793), .Z(\w1[1][2] ) );
  XNOR U4147 ( .A(\w3[0][24] ), .B(\w3[0][31] ), .Z(n2973) );
  XNOR U4148 ( .A(n2795), .B(n2973), .Z(n2934) );
  XOR U4149 ( .A(n2934), .B(key[158]), .Z(n2798) );
  XNOR U4150 ( .A(\w3[0][6] ), .B(n2796), .Z(n2797) );
  XNOR U4151 ( .A(n2798), .B(n2797), .Z(\w1[1][30] ) );
  XOR U4152 ( .A(\w3[0][15] ), .B(\w3[0][23] ), .Z(n2971) );
  XOR U4153 ( .A(n2971), .B(key[159]), .Z(n2800) );
  XNOR U4154 ( .A(n3012), .B(\w3[0][7] ), .Z(n2799) );
  XNOR U4155 ( .A(n2800), .B(n2799), .Z(\w1[1][31] ) );
  XOR U4156 ( .A(\w3[0][33] ), .B(\w3[0][57] ), .Z(n2855) );
  XOR U4157 ( .A(n2855), .B(key[160]), .Z(n2802) );
  XOR U4158 ( .A(\w3[0][48] ), .B(\w3[0][56] ), .Z(n2916) );
  XNOR U4159 ( .A(n2916), .B(\w3[0][40] ), .Z(n2801) );
  XNOR U4160 ( .A(n2802), .B(n2801), .Z(\w1[1][32] ) );
  XOR U4161 ( .A(\w3[0][34] ), .B(\w3[0][58] ), .Z(n2863) );
  XOR U4162 ( .A(n2863), .B(key[161]), .Z(n2804) );
  XOR U4163 ( .A(\w3[0][41] ), .B(\w3[0][49] ), .Z(n2887) );
  XNOR U4164 ( .A(\w3[0][57] ), .B(n2887), .Z(n2803) );
  XNOR U4165 ( .A(n2804), .B(n2803), .Z(\w1[1][33] ) );
  XOR U4166 ( .A(\w3[0][35] ), .B(\w3[0][59] ), .Z(n2834) );
  XOR U4167 ( .A(n2834), .B(key[162]), .Z(n2806) );
  XOR U4168 ( .A(\w3[0][42] ), .B(\w3[0][50] ), .Z(n2891) );
  XNOR U4169 ( .A(\w3[0][58] ), .B(n2891), .Z(n2805) );
  XNOR U4170 ( .A(n2806), .B(n2805), .Z(\w1[1][34] ) );
  XOR U4171 ( .A(\w3[0][36] ), .B(\w3[0][32] ), .Z(n2836) );
  XOR U4172 ( .A(n2836), .B(key[163]), .Z(n2809) );
  XOR U4173 ( .A(\w3[0][43] ), .B(\w3[0][51] ), .Z(n2862) );
  XNOR U4174 ( .A(\w3[0][56] ), .B(n2862), .Z(n2807) );
  XNOR U4175 ( .A(\w3[0][60] ), .B(n2807), .Z(n2896) );
  XNOR U4176 ( .A(\w3[0][59] ), .B(n2896), .Z(n2808) );
  XNOR U4177 ( .A(n2809), .B(n2808), .Z(\w1[1][35] ) );
  XOR U4178 ( .A(\w3[0][32] ), .B(\w3[0][37] ), .Z(n2841) );
  XOR U4179 ( .A(n2841), .B(key[164]), .Z(n2813) );
  XOR U4180 ( .A(\w3[0][52] ), .B(\w3[0][61] ), .Z(n2811) );
  XNOR U4181 ( .A(\w3[0][56] ), .B(\w3[0][44] ), .Z(n2810) );
  XNOR U4182 ( .A(n2811), .B(n2810), .Z(n2904) );
  XNOR U4183 ( .A(\w3[0][60] ), .B(n2904), .Z(n2812) );
  XNOR U4184 ( .A(n2813), .B(n2812), .Z(\w1[1][36] ) );
  XOR U4185 ( .A(\w3[0][38] ), .B(\w3[0][62] ), .Z(n2847) );
  XOR U4186 ( .A(n2847), .B(key[165]), .Z(n2815) );
  XOR U4187 ( .A(\w3[0][45] ), .B(\w3[0][53] ), .Z(n2907) );
  XNOR U4188 ( .A(\w3[0][61] ), .B(n2907), .Z(n2814) );
  XNOR U4189 ( .A(n2815), .B(n2814), .Z(\w1[1][37] ) );
  XOR U4190 ( .A(\w3[0][32] ), .B(\w3[0][39] ), .Z(n2848) );
  XOR U4191 ( .A(n2848), .B(key[166]), .Z(n2817) );
  XOR U4192 ( .A(\w3[0][46] ), .B(\w3[0][54] ), .Z(n2873) );
  XNOR U4193 ( .A(\w3[0][56] ), .B(\w3[0][63] ), .Z(n2819) );
  XNOR U4194 ( .A(n2873), .B(n2819), .Z(n2912) );
  XNOR U4195 ( .A(\w3[0][62] ), .B(n2912), .Z(n2816) );
  XNOR U4196 ( .A(n2817), .B(n2816), .Z(\w1[1][38] ) );
  XOR U4197 ( .A(\w3[0][47] ), .B(\w3[0][55] ), .Z(n2915) );
  XNOR U4198 ( .A(n2915), .B(key[167]), .Z(n2818) );
  XNOR U4199 ( .A(n2819), .B(n2818), .Z(n2820) );
  XNOR U4200 ( .A(\w3[0][32] ), .B(n2820), .Z(\w1[1][39] ) );
  XOR U4201 ( .A(n2821), .B(key[131]), .Z(n2824) );
  XNOR U4202 ( .A(n2822), .B(\w3[0][27] ), .Z(n2823) );
  XNOR U4203 ( .A(n2824), .B(n2823), .Z(\w1[1][3] ) );
  XOR U4204 ( .A(\w3[0][32] ), .B(key[168]), .Z(n2826) );
  XNOR U4205 ( .A(\w3[0][33] ), .B(\w3[0][41] ), .Z(n2825) );
  XNOR U4206 ( .A(n2826), .B(n2825), .Z(n2827) );
  XOR U4207 ( .A(n2916), .B(n2827), .Z(\w1[1][40] ) );
  XOR U4208 ( .A(\w3[0][42] ), .B(key[169]), .Z(n2829) );
  XNOR U4209 ( .A(\w3[0][49] ), .B(\w3[0][34] ), .Z(n2828) );
  XNOR U4210 ( .A(n2829), .B(n2828), .Z(n2830) );
  XOR U4211 ( .A(n2855), .B(n2830), .Z(\w1[1][41] ) );
  XOR U4212 ( .A(\w3[0][43] ), .B(key[170]), .Z(n2832) );
  XNOR U4213 ( .A(\w3[0][50] ), .B(\w3[0][35] ), .Z(n2831) );
  XNOR U4214 ( .A(n2832), .B(n2831), .Z(n2833) );
  XOR U4215 ( .A(n2863), .B(n2833), .Z(\w1[1][42] ) );
  XNOR U4216 ( .A(\w3[0][40] ), .B(n2834), .Z(n2835) );
  XNOR U4217 ( .A(\w3[0][44] ), .B(n2835), .Z(n2866) );
  XOR U4218 ( .A(n2866), .B(key[171]), .Z(n2838) );
  XNOR U4219 ( .A(\w3[0][51] ), .B(n2836), .Z(n2837) );
  XNOR U4220 ( .A(n2838), .B(n2837), .Z(\w1[1][43] ) );
  XOR U4221 ( .A(\w3[0][36] ), .B(\w3[0][45] ), .Z(n2840) );
  XNOR U4222 ( .A(\w3[0][40] ), .B(\w3[0][60] ), .Z(n2839) );
  XNOR U4223 ( .A(n2840), .B(n2839), .Z(n2869) );
  XOR U4224 ( .A(n2869), .B(key[172]), .Z(n2843) );
  XNOR U4225 ( .A(\w3[0][52] ), .B(n2841), .Z(n2842) );
  XNOR U4226 ( .A(n2843), .B(n2842), .Z(\w1[1][44] ) );
  XOR U4227 ( .A(\w3[0][61] ), .B(\w3[0][37] ), .Z(n2872) );
  XOR U4228 ( .A(n2872), .B(key[173]), .Z(n2845) );
  XNOR U4229 ( .A(\w3[0][38] ), .B(\w3[0][46] ), .Z(n2844) );
  XNOR U4230 ( .A(n2845), .B(n2844), .Z(n2846) );
  XOR U4231 ( .A(\w3[0][53] ), .B(n2846), .Z(\w1[1][45] ) );
  XNOR U4232 ( .A(\w3[0][40] ), .B(\w3[0][47] ), .Z(n2881) );
  XNOR U4233 ( .A(n2847), .B(n2881), .Z(n2876) );
  XOR U4234 ( .A(n2876), .B(key[174]), .Z(n2850) );
  XNOR U4235 ( .A(\w3[0][54] ), .B(n2848), .Z(n2849) );
  XNOR U4236 ( .A(n2850), .B(n2849), .Z(\w1[1][46] ) );
  XOR U4237 ( .A(\w3[0][63] ), .B(\w3[0][39] ), .Z(n2879) );
  XOR U4238 ( .A(n2879), .B(key[175]), .Z(n2852) );
  XOR U4239 ( .A(\w3[0][40] ), .B(\w3[0][32] ), .Z(n2883) );
  XNOR U4240 ( .A(\w3[0][55] ), .B(n2883), .Z(n2851) );
  XNOR U4241 ( .A(n2852), .B(n2851), .Z(\w1[1][47] ) );
  XOR U4242 ( .A(n2883), .B(key[176]), .Z(n2854) );
  XNOR U4243 ( .A(\w3[0][56] ), .B(n2887), .Z(n2853) );
  XNOR U4244 ( .A(n2854), .B(n2853), .Z(\w1[1][48] ) );
  XOR U4245 ( .A(n2891), .B(key[177]), .Z(n2857) );
  XNOR U4246 ( .A(n2855), .B(\w3[0][41] ), .Z(n2856) );
  XNOR U4247 ( .A(n2857), .B(n2856), .Z(\w1[1][49] ) );
  XOR U4248 ( .A(n2858), .B(key[132]), .Z(n2861) );
  XNOR U4249 ( .A(n2859), .B(\w3[0][28] ), .Z(n2860) );
  XNOR U4250 ( .A(n2861), .B(n2860), .Z(\w1[1][4] ) );
  XOR U4251 ( .A(n2862), .B(key[178]), .Z(n2865) );
  XNOR U4252 ( .A(n2863), .B(\w3[0][42] ), .Z(n2864) );
  XNOR U4253 ( .A(n2865), .B(n2864), .Z(\w1[1][50] ) );
  XOR U4254 ( .A(\w3[0][48] ), .B(\w3[0][52] ), .Z(n2895) );
  XOR U4255 ( .A(n2895), .B(key[179]), .Z(n2868) );
  XNOR U4256 ( .A(\w3[0][43] ), .B(n2866), .Z(n2867) );
  XNOR U4257 ( .A(n2868), .B(n2867), .Z(\w1[1][51] ) );
  XOR U4258 ( .A(\w3[0][48] ), .B(\w3[0][53] ), .Z(n2903) );
  XOR U4259 ( .A(n2903), .B(key[180]), .Z(n2871) );
  XNOR U4260 ( .A(\w3[0][44] ), .B(n2869), .Z(n2870) );
  XNOR U4261 ( .A(n2871), .B(n2870), .Z(\w1[1][52] ) );
  XOR U4262 ( .A(n2872), .B(key[181]), .Z(n2875) );
  XNOR U4263 ( .A(\w3[0][45] ), .B(n2873), .Z(n2874) );
  XNOR U4264 ( .A(n2875), .B(n2874), .Z(\w1[1][53] ) );
  XOR U4265 ( .A(\w3[0][48] ), .B(\w3[0][55] ), .Z(n2911) );
  XOR U4266 ( .A(n2911), .B(key[182]), .Z(n2878) );
  XNOR U4267 ( .A(\w3[0][46] ), .B(n2876), .Z(n2877) );
  XNOR U4268 ( .A(n2878), .B(n2877), .Z(\w1[1][54] ) );
  XNOR U4269 ( .A(n2879), .B(key[183]), .Z(n2880) );
  XNOR U4270 ( .A(n2881), .B(n2880), .Z(n2882) );
  XNOR U4271 ( .A(\w3[0][48] ), .B(n2882), .Z(\w1[1][55] ) );
  XOR U4272 ( .A(n2883), .B(key[184]), .Z(n2885) );
  XNOR U4273 ( .A(\w3[0][48] ), .B(\w3[0][49] ), .Z(n2884) );
  XNOR U4274 ( .A(n2885), .B(n2884), .Z(n2886) );
  XOR U4275 ( .A(\w3[0][57] ), .B(n2886), .Z(\w1[1][56] ) );
  XOR U4276 ( .A(\w3[0][50] ), .B(key[185]), .Z(n2889) );
  XNOR U4277 ( .A(n2887), .B(\w3[0][58] ), .Z(n2888) );
  XNOR U4278 ( .A(n2889), .B(n2888), .Z(n2890) );
  XOR U4279 ( .A(\w3[0][33] ), .B(n2890), .Z(\w1[1][57] ) );
  XOR U4280 ( .A(\w3[0][51] ), .B(key[186]), .Z(n2893) );
  XNOR U4281 ( .A(n2891), .B(\w3[0][59] ), .Z(n2892) );
  XNOR U4282 ( .A(n2893), .B(n2892), .Z(n2894) );
  XOR U4283 ( .A(\w3[0][34] ), .B(n2894), .Z(\w1[1][58] ) );
  XOR U4284 ( .A(n2895), .B(key[187]), .Z(n2898) );
  XNOR U4285 ( .A(\w3[0][35] ), .B(n2896), .Z(n2897) );
  XNOR U4286 ( .A(n2898), .B(n2897), .Z(\w1[1][59] ) );
  XOR U4287 ( .A(n2899), .B(key[133]), .Z(n2902) );
  XNOR U4288 ( .A(\w3[0][29] ), .B(n2900), .Z(n2901) );
  XNOR U4289 ( .A(n2902), .B(n2901), .Z(\w1[1][5] ) );
  XOR U4290 ( .A(n2903), .B(key[188]), .Z(n2906) );
  XNOR U4291 ( .A(\w3[0][36] ), .B(n2904), .Z(n2905) );
  XNOR U4292 ( .A(n2906), .B(n2905), .Z(\w1[1][60] ) );
  XOR U4293 ( .A(\w3[0][54] ), .B(key[189]), .Z(n2909) );
  XNOR U4294 ( .A(n2907), .B(\w3[0][62] ), .Z(n2908) );
  XNOR U4295 ( .A(n2909), .B(n2908), .Z(n2910) );
  XOR U4296 ( .A(\w3[0][37] ), .B(n2910), .Z(\w1[1][61] ) );
  XOR U4297 ( .A(n2911), .B(key[190]), .Z(n2914) );
  XNOR U4298 ( .A(\w3[0][38] ), .B(n2912), .Z(n2913) );
  XNOR U4299 ( .A(n2914), .B(n2913), .Z(\w1[1][62] ) );
  XOR U4300 ( .A(n2915), .B(key[191]), .Z(n2918) );
  XNOR U4301 ( .A(n2916), .B(\w3[0][39] ), .Z(n2917) );
  XNOR U4302 ( .A(n2918), .B(n2917), .Z(\w1[1][63] ) );
  XOR U4303 ( .A(\w3[0][65] ), .B(\w3[0][89] ), .Z(n2977) );
  XOR U4304 ( .A(n2977), .B(key[192]), .Z(n2920) );
  XOR U4305 ( .A(\w3[0][80] ), .B(\w3[0][88] ), .Z(n3034) );
  XNOR U4306 ( .A(n3034), .B(\w3[0][72] ), .Z(n2919) );
  XNOR U4307 ( .A(n2920), .B(n2919), .Z(\w1[1][64] ) );
  XOR U4308 ( .A(\w3[0][66] ), .B(\w3[0][90] ), .Z(n2981) );
  XOR U4309 ( .A(n2981), .B(key[193]), .Z(n2922) );
  XOR U4310 ( .A(\w3[0][73] ), .B(\w3[0][81] ), .Z(n3005) );
  XNOR U4311 ( .A(\w3[0][89] ), .B(n3005), .Z(n2921) );
  XNOR U4312 ( .A(n2922), .B(n2921), .Z(\w1[1][65] ) );
  XOR U4313 ( .A(\w3[0][67] ), .B(\w3[0][91] ), .Z(n2952) );
  XOR U4314 ( .A(n2952), .B(key[194]), .Z(n2924) );
  XOR U4315 ( .A(\w3[0][74] ), .B(\w3[0][82] ), .Z(n3013) );
  XNOR U4316 ( .A(\w3[0][90] ), .B(n3013), .Z(n2923) );
  XNOR U4317 ( .A(n2924), .B(n2923), .Z(\w1[1][66] ) );
  XOR U4318 ( .A(\w3[0][68] ), .B(\w3[0][64] ), .Z(n2954) );
  XOR U4319 ( .A(n2954), .B(key[195]), .Z(n2927) );
  XOR U4320 ( .A(\w3[0][75] ), .B(\w3[0][83] ), .Z(n2980) );
  XNOR U4321 ( .A(\w3[0][88] ), .B(n2980), .Z(n2925) );
  XNOR U4322 ( .A(\w3[0][92] ), .B(n2925), .Z(n3018) );
  XNOR U4323 ( .A(\w3[0][91] ), .B(n3018), .Z(n2926) );
  XNOR U4324 ( .A(n2927), .B(n2926), .Z(\w1[1][67] ) );
  XOR U4325 ( .A(\w3[0][64] ), .B(\w3[0][69] ), .Z(n2959) );
  XOR U4326 ( .A(n2959), .B(key[196]), .Z(n2931) );
  XOR U4327 ( .A(\w3[0][84] ), .B(\w3[0][93] ), .Z(n2929) );
  XNOR U4328 ( .A(\w3[0][88] ), .B(\w3[0][76] ), .Z(n2928) );
  XNOR U4329 ( .A(n2929), .B(n2928), .Z(n3022) );
  XNOR U4330 ( .A(\w3[0][92] ), .B(n3022), .Z(n2930) );
  XNOR U4331 ( .A(n2931), .B(n2930), .Z(\w1[1][68] ) );
  XOR U4332 ( .A(\w3[0][70] ), .B(\w3[0][94] ), .Z(n2965) );
  XOR U4333 ( .A(n2965), .B(key[197]), .Z(n2933) );
  XOR U4334 ( .A(\w3[0][77] ), .B(\w3[0][85] ), .Z(n3025) );
  XNOR U4335 ( .A(\w3[0][93] ), .B(n3025), .Z(n2932) );
  XNOR U4336 ( .A(n2933), .B(n2932), .Z(\w1[1][69] ) );
  XOR U4337 ( .A(n2934), .B(key[134]), .Z(n2937) );
  XNOR U4338 ( .A(n2935), .B(\w3[0][30] ), .Z(n2936) );
  XNOR U4339 ( .A(n2937), .B(n2936), .Z(\w1[1][6] ) );
  XOR U4340 ( .A(\w3[0][64] ), .B(\w3[0][71] ), .Z(n2966) );
  XOR U4341 ( .A(n2966), .B(key[198]), .Z(n2939) );
  XOR U4342 ( .A(\w3[0][78] ), .B(\w3[0][86] ), .Z(n2991) );
  XNOR U4343 ( .A(\w3[0][88] ), .B(\w3[0][95] ), .Z(n2941) );
  XNOR U4344 ( .A(n2991), .B(n2941), .Z(n3030) );
  XNOR U4345 ( .A(\w3[0][94] ), .B(n3030), .Z(n2938) );
  XNOR U4346 ( .A(n2939), .B(n2938), .Z(\w1[1][70] ) );
  XOR U4347 ( .A(\w3[0][79] ), .B(\w3[0][87] ), .Z(n3033) );
  XNOR U4348 ( .A(n3033), .B(key[199]), .Z(n2940) );
  XNOR U4349 ( .A(n2941), .B(n2940), .Z(n2942) );
  XNOR U4350 ( .A(\w3[0][64] ), .B(n2942), .Z(\w1[1][71] ) );
  XOR U4351 ( .A(\w3[0][64] ), .B(key[200]), .Z(n2944) );
  XNOR U4352 ( .A(\w3[0][65] ), .B(\w3[0][73] ), .Z(n2943) );
  XNOR U4353 ( .A(n2944), .B(n2943), .Z(n2945) );
  XOR U4354 ( .A(n3034), .B(n2945), .Z(\w1[1][72] ) );
  XOR U4355 ( .A(\w3[0][74] ), .B(key[201]), .Z(n2947) );
  XNOR U4356 ( .A(\w3[0][81] ), .B(\w3[0][66] ), .Z(n2946) );
  XNOR U4357 ( .A(n2947), .B(n2946), .Z(n2948) );
  XOR U4358 ( .A(n2977), .B(n2948), .Z(\w1[1][73] ) );
  XOR U4359 ( .A(\w3[0][75] ), .B(key[202]), .Z(n2950) );
  XNOR U4360 ( .A(\w3[0][82] ), .B(\w3[0][67] ), .Z(n2949) );
  XNOR U4361 ( .A(n2950), .B(n2949), .Z(n2951) );
  XOR U4362 ( .A(n2981), .B(n2951), .Z(\w1[1][74] ) );
  XNOR U4363 ( .A(\w3[0][72] ), .B(n2952), .Z(n2953) );
  XNOR U4364 ( .A(\w3[0][76] ), .B(n2953), .Z(n2984) );
  XOR U4365 ( .A(n2984), .B(key[203]), .Z(n2956) );
  XNOR U4366 ( .A(\w3[0][83] ), .B(n2954), .Z(n2955) );
  XNOR U4367 ( .A(n2956), .B(n2955), .Z(\w1[1][75] ) );
  XOR U4368 ( .A(\w3[0][68] ), .B(\w3[0][77] ), .Z(n2958) );
  XNOR U4369 ( .A(\w3[0][72] ), .B(\w3[0][92] ), .Z(n2957) );
  XNOR U4370 ( .A(n2958), .B(n2957), .Z(n2987) );
  XOR U4371 ( .A(n2987), .B(key[204]), .Z(n2961) );
  XNOR U4372 ( .A(\w3[0][84] ), .B(n2959), .Z(n2960) );
  XNOR U4373 ( .A(n2961), .B(n2960), .Z(\w1[1][76] ) );
  XOR U4374 ( .A(\w3[0][93] ), .B(\w3[0][69] ), .Z(n2990) );
  XOR U4375 ( .A(n2990), .B(key[205]), .Z(n2963) );
  XNOR U4376 ( .A(\w3[0][70] ), .B(\w3[0][78] ), .Z(n2962) );
  XNOR U4377 ( .A(n2963), .B(n2962), .Z(n2964) );
  XOR U4378 ( .A(\w3[0][85] ), .B(n2964), .Z(\w1[1][77] ) );
  XNOR U4379 ( .A(\w3[0][72] ), .B(\w3[0][79] ), .Z(n2999) );
  XNOR U4380 ( .A(n2965), .B(n2999), .Z(n2994) );
  XOR U4381 ( .A(n2994), .B(key[206]), .Z(n2968) );
  XNOR U4382 ( .A(\w3[0][86] ), .B(n2966), .Z(n2967) );
  XNOR U4383 ( .A(n2968), .B(n2967), .Z(\w1[1][78] ) );
  XOR U4384 ( .A(\w3[0][95] ), .B(\w3[0][71] ), .Z(n2997) );
  XOR U4385 ( .A(n2997), .B(key[207]), .Z(n2970) );
  XOR U4386 ( .A(\w3[0][72] ), .B(\w3[0][64] ), .Z(n3001) );
  XNOR U4387 ( .A(\w3[0][87] ), .B(n3001), .Z(n2969) );
  XNOR U4388 ( .A(n2970), .B(n2969), .Z(\w1[1][79] ) );
  XNOR U4389 ( .A(n2971), .B(key[135]), .Z(n2972) );
  XNOR U4390 ( .A(n2973), .B(n2972), .Z(n2974) );
  XNOR U4391 ( .A(\w3[0][0] ), .B(n2974), .Z(\w1[1][7] ) );
  XOR U4392 ( .A(n3001), .B(key[208]), .Z(n2976) );
  XNOR U4393 ( .A(\w3[0][88] ), .B(n3005), .Z(n2975) );
  XNOR U4394 ( .A(n2976), .B(n2975), .Z(\w1[1][80] ) );
  XOR U4395 ( .A(n3013), .B(key[209]), .Z(n2979) );
  XNOR U4396 ( .A(n2977), .B(\w3[0][73] ), .Z(n2978) );
  XNOR U4397 ( .A(n2979), .B(n2978), .Z(\w1[1][81] ) );
  XOR U4398 ( .A(n2980), .B(key[210]), .Z(n2983) );
  XNOR U4399 ( .A(n2981), .B(\w3[0][74] ), .Z(n2982) );
  XNOR U4400 ( .A(n2983), .B(n2982), .Z(\w1[1][82] ) );
  XOR U4401 ( .A(\w3[0][80] ), .B(\w3[0][84] ), .Z(n3017) );
  XOR U4402 ( .A(n3017), .B(key[211]), .Z(n2986) );
  XNOR U4403 ( .A(\w3[0][75] ), .B(n2984), .Z(n2985) );
  XNOR U4404 ( .A(n2986), .B(n2985), .Z(\w1[1][83] ) );
  XOR U4405 ( .A(\w3[0][80] ), .B(\w3[0][85] ), .Z(n3021) );
  XOR U4406 ( .A(n3021), .B(key[212]), .Z(n2989) );
  XNOR U4407 ( .A(\w3[0][76] ), .B(n2987), .Z(n2988) );
  XNOR U4408 ( .A(n2989), .B(n2988), .Z(\w1[1][84] ) );
  XOR U4409 ( .A(n2990), .B(key[213]), .Z(n2993) );
  XNOR U4410 ( .A(\w3[0][77] ), .B(n2991), .Z(n2992) );
  XNOR U4411 ( .A(n2993), .B(n2992), .Z(\w1[1][85] ) );
  XOR U4412 ( .A(\w3[0][80] ), .B(\w3[0][87] ), .Z(n3029) );
  XOR U4413 ( .A(n3029), .B(key[214]), .Z(n2996) );
  XNOR U4414 ( .A(\w3[0][78] ), .B(n2994), .Z(n2995) );
  XNOR U4415 ( .A(n2996), .B(n2995), .Z(\w1[1][86] ) );
  XNOR U4416 ( .A(n2997), .B(key[215]), .Z(n2998) );
  XNOR U4417 ( .A(n2999), .B(n2998), .Z(n3000) );
  XNOR U4418 ( .A(\w3[0][80] ), .B(n3000), .Z(\w1[1][87] ) );
  XOR U4419 ( .A(n3001), .B(key[216]), .Z(n3003) );
  XNOR U4420 ( .A(\w3[0][80] ), .B(\w3[0][81] ), .Z(n3002) );
  XNOR U4421 ( .A(n3003), .B(n3002), .Z(n3004) );
  XOR U4422 ( .A(\w3[0][89] ), .B(n3004), .Z(\w1[1][88] ) );
  XOR U4423 ( .A(\w3[0][82] ), .B(key[217]), .Z(n3007) );
  XNOR U4424 ( .A(n3005), .B(\w3[0][90] ), .Z(n3006) );
  XNOR U4425 ( .A(n3007), .B(n3006), .Z(n3008) );
  XOR U4426 ( .A(\w3[0][65] ), .B(n3008), .Z(\w1[1][89] ) );
  XOR U4427 ( .A(\w3[0][9] ), .B(key[136]), .Z(n3010) );
  XNOR U4428 ( .A(\w3[0][1] ), .B(\w3[0][0] ), .Z(n3009) );
  XNOR U4429 ( .A(n3010), .B(n3009), .Z(n3011) );
  XOR U4430 ( .A(n3012), .B(n3011), .Z(\w1[1][8] ) );
  XOR U4431 ( .A(\w3[0][83] ), .B(key[218]), .Z(n3015) );
  XNOR U4432 ( .A(n3013), .B(\w3[0][91] ), .Z(n3014) );
  XNOR U4433 ( .A(n3015), .B(n3014), .Z(n3016) );
  XOR U4434 ( .A(\w3[0][66] ), .B(n3016), .Z(\w1[1][90] ) );
  XOR U4435 ( .A(n3017), .B(key[219]), .Z(n3020) );
  XNOR U4436 ( .A(\w3[0][67] ), .B(n3018), .Z(n3019) );
  XNOR U4437 ( .A(n3020), .B(n3019), .Z(\w1[1][91] ) );
  XOR U4438 ( .A(n3021), .B(key[220]), .Z(n3024) );
  XNOR U4439 ( .A(\w3[0][68] ), .B(n3022), .Z(n3023) );
  XNOR U4440 ( .A(n3024), .B(n3023), .Z(\w1[1][92] ) );
  XOR U4441 ( .A(\w3[0][86] ), .B(key[221]), .Z(n3027) );
  XNOR U4442 ( .A(n3025), .B(\w3[0][94] ), .Z(n3026) );
  XNOR U4443 ( .A(n3027), .B(n3026), .Z(n3028) );
  XOR U4444 ( .A(\w3[0][69] ), .B(n3028), .Z(\w1[1][93] ) );
  XOR U4445 ( .A(n3029), .B(key[222]), .Z(n3032) );
  XNOR U4446 ( .A(\w3[0][70] ), .B(n3030), .Z(n3031) );
  XNOR U4447 ( .A(n3032), .B(n3031), .Z(\w1[1][94] ) );
  XOR U4448 ( .A(n3033), .B(key[223]), .Z(n3036) );
  XNOR U4449 ( .A(n3034), .B(\w3[0][71] ), .Z(n3035) );
  XNOR U4450 ( .A(n3036), .B(n3035), .Z(\w1[1][95] ) );
  XOR U4451 ( .A(\w3[0][104] ), .B(key[224]), .Z(n3040) );
  XOR U4452 ( .A(n3038), .B(n3037), .Z(n3039) );
  XNOR U4453 ( .A(n3040), .B(n3039), .Z(\w1[1][96] ) );
  XOR U4454 ( .A(n3041), .B(key[225]), .Z(n3044) );
  XNOR U4455 ( .A(\w3[0][121] ), .B(n3042), .Z(n3043) );
  XNOR U4456 ( .A(n3044), .B(n3043), .Z(\w1[1][97] ) );
  XOR U4457 ( .A(n3045), .B(key[226]), .Z(n3048) );
  XNOR U4458 ( .A(\w3[0][122] ), .B(n3046), .Z(n3047) );
  XNOR U4459 ( .A(n3048), .B(n3047), .Z(\w1[1][98] ) );
  XOR U4460 ( .A(n3049), .B(key[227]), .Z(n3052) );
  XNOR U4461 ( .A(n3050), .B(\w3[0][123] ), .Z(n3051) );
  XNOR U4462 ( .A(n3052), .B(n3051), .Z(\w1[1][99] ) );
  XOR U4463 ( .A(\w3[0][10] ), .B(key[137]), .Z(n3054) );
  XNOR U4464 ( .A(\w3[0][2] ), .B(\w3[0][17] ), .Z(n3053) );
  XNOR U4465 ( .A(n3054), .B(n3053), .Z(n3055) );
  XOR U4466 ( .A(n3056), .B(n3055), .Z(\w1[1][9] ) );
  XOR U4467 ( .A(\w3[1][8] ), .B(key[256]), .Z(n3058) );
  XOR U4468 ( .A(\w3[1][1] ), .B(\w3[1][25] ), .Z(n3480) );
  XOR U4469 ( .A(\w3[1][16] ), .B(\w3[1][24] ), .Z(n3436) );
  XNOR U4470 ( .A(n3480), .B(n3436), .Z(n3057) );
  XNOR U4471 ( .A(n3058), .B(n3057), .Z(\w1[2][0] ) );
  XOR U4472 ( .A(\w3[1][96] ), .B(\w3[1][101] ), .Z(n3083) );
  XOR U4473 ( .A(n3083), .B(key[356]), .Z(n3062) );
  XOR U4474 ( .A(\w3[1][116] ), .B(\w3[1][125] ), .Z(n3060) );
  XNOR U4475 ( .A(\w3[1][120] ), .B(\w3[1][108] ), .Z(n3059) );
  XNOR U4476 ( .A(n3060), .B(n3059), .Z(n3141) );
  XNOR U4477 ( .A(\w3[1][124] ), .B(n3141), .Z(n3061) );
  XNOR U4478 ( .A(n3062), .B(n3061), .Z(\w1[2][100] ) );
  XOR U4479 ( .A(\w3[1][102] ), .B(\w3[1][126] ), .Z(n3092) );
  XOR U4480 ( .A(n3092), .B(key[357]), .Z(n3064) );
  XOR U4481 ( .A(\w3[1][109] ), .B(\w3[1][117] ), .Z(n3144) );
  XNOR U4482 ( .A(\w3[1][125] ), .B(n3144), .Z(n3063) );
  XNOR U4483 ( .A(n3064), .B(n3063), .Z(\w1[2][101] ) );
  XOR U4484 ( .A(\w3[1][96] ), .B(\w3[1][103] ), .Z(n3093) );
  XOR U4485 ( .A(n3093), .B(key[358]), .Z(n3066) );
  XOR U4486 ( .A(\w3[1][110] ), .B(\w3[1][118] ), .Z(n3112) );
  XNOR U4487 ( .A(\w3[1][120] ), .B(\w3[1][127] ), .Z(n3068) );
  XNOR U4488 ( .A(n3112), .B(n3068), .Z(n3149) );
  XNOR U4489 ( .A(\w3[1][126] ), .B(n3149), .Z(n3065) );
  XNOR U4490 ( .A(n3066), .B(n3065), .Z(\w1[2][102] ) );
  XOR U4491 ( .A(\w3[1][111] ), .B(\w3[1][119] ), .Z(n3152) );
  XNOR U4492 ( .A(n3152), .B(key[359]), .Z(n3067) );
  XNOR U4493 ( .A(n3068), .B(n3067), .Z(n3069) );
  XNOR U4494 ( .A(\w3[1][96] ), .B(n3069), .Z(\w1[2][103] ) );
  XOR U4495 ( .A(\w3[1][105] ), .B(\w3[1][97] ), .Z(n3100) );
  XOR U4496 ( .A(n3100), .B(key[360]), .Z(n3071) );
  XOR U4497 ( .A(\w3[1][120] ), .B(\w3[1][112] ), .Z(n3462) );
  XNOR U4498 ( .A(\w3[1][96] ), .B(n3462), .Z(n3070) );
  XNOR U4499 ( .A(n3071), .B(n3070), .Z(\w1[2][104] ) );
  XOR U4500 ( .A(\w3[1][106] ), .B(\w3[1][98] ), .Z(n3073) );
  XOR U4501 ( .A(\w3[1][97] ), .B(\w3[1][121] ), .Z(n3461) );
  XNOR U4502 ( .A(n3461), .B(key[361]), .Z(n3072) );
  XNOR U4503 ( .A(n3073), .B(n3072), .Z(n3074) );
  XOR U4504 ( .A(\w3[1][113] ), .B(n3074), .Z(\w1[2][105] ) );
  XOR U4505 ( .A(\w3[1][107] ), .B(\w3[1][99] ), .Z(n3076) );
  XOR U4506 ( .A(\w3[1][98] ), .B(\w3[1][122] ), .Z(n3466) );
  XNOR U4507 ( .A(n3466), .B(key[362]), .Z(n3075) );
  XNOR U4508 ( .A(n3076), .B(n3075), .Z(n3077) );
  XOR U4509 ( .A(\w3[1][114] ), .B(n3077), .Z(\w1[2][106] ) );
  XOR U4510 ( .A(\w3[1][99] ), .B(\w3[1][123] ), .Z(n3470) );
  XNOR U4511 ( .A(\w3[1][108] ), .B(n3470), .Z(n3078) );
  XNOR U4512 ( .A(\w3[1][104] ), .B(n3078), .Z(n3105) );
  XOR U4513 ( .A(n3105), .B(key[363]), .Z(n3080) );
  XOR U4514 ( .A(\w3[1][96] ), .B(\w3[1][100] ), .Z(n3474) );
  XNOR U4515 ( .A(\w3[1][115] ), .B(n3474), .Z(n3079) );
  XNOR U4516 ( .A(n3080), .B(n3079), .Z(\w1[2][107] ) );
  XOR U4517 ( .A(\w3[1][100] ), .B(\w3[1][104] ), .Z(n3082) );
  XNOR U4518 ( .A(\w3[1][124] ), .B(\w3[1][109] ), .Z(n3081) );
  XNOR U4519 ( .A(n3082), .B(n3081), .Z(n3108) );
  XOR U4520 ( .A(n3108), .B(key[364]), .Z(n3085) );
  XNOR U4521 ( .A(\w3[1][116] ), .B(n3083), .Z(n3084) );
  XNOR U4522 ( .A(n3085), .B(n3084), .Z(\w1[2][108] ) );
  XOR U4523 ( .A(\w3[1][125] ), .B(\w3[1][101] ), .Z(n3111) );
  XOR U4524 ( .A(n3111), .B(key[365]), .Z(n3087) );
  XNOR U4525 ( .A(\w3[1][102] ), .B(\w3[1][110] ), .Z(n3086) );
  XNOR U4526 ( .A(n3087), .B(n3086), .Z(n3088) );
  XOR U4527 ( .A(\w3[1][117] ), .B(n3088), .Z(\w1[2][109] ) );
  XOR U4528 ( .A(\w3[1][11] ), .B(\w3[1][18] ), .Z(n3090) );
  XOR U4529 ( .A(\w3[1][2] ), .B(\w3[1][26] ), .Z(n3175) );
  XNOR U4530 ( .A(n3175), .B(key[266]), .Z(n3089) );
  XNOR U4531 ( .A(n3090), .B(n3089), .Z(n3091) );
  XOR U4532 ( .A(\w3[1][3] ), .B(n3091), .Z(\w1[2][10] ) );
  XNOR U4533 ( .A(\w3[1][111] ), .B(\w3[1][104] ), .Z(n3120) );
  XNOR U4534 ( .A(n3092), .B(n3120), .Z(n3115) );
  XOR U4535 ( .A(n3115), .B(key[366]), .Z(n3095) );
  XNOR U4536 ( .A(\w3[1][118] ), .B(n3093), .Z(n3094) );
  XNOR U4537 ( .A(n3095), .B(n3094), .Z(\w1[2][110] ) );
  XOR U4538 ( .A(\w3[1][127] ), .B(\w3[1][103] ), .Z(n3118) );
  XOR U4539 ( .A(n3118), .B(key[367]), .Z(n3097) );
  XOR U4540 ( .A(\w3[1][96] ), .B(\w3[1][104] ), .Z(n3125) );
  XNOR U4541 ( .A(\w3[1][119] ), .B(n3125), .Z(n3096) );
  XNOR U4542 ( .A(n3097), .B(n3096), .Z(\w1[2][111] ) );
  XOR U4543 ( .A(\w3[1][105] ), .B(\w3[1][113] ), .Z(n3465) );
  XOR U4544 ( .A(n3465), .B(key[368]), .Z(n3099) );
  XNOR U4545 ( .A(\w3[1][120] ), .B(n3125), .Z(n3098) );
  XNOR U4546 ( .A(n3099), .B(n3098), .Z(\w1[2][112] ) );
  XOR U4547 ( .A(\w3[1][106] ), .B(\w3[1][114] ), .Z(n3469) );
  XOR U4548 ( .A(n3469), .B(key[369]), .Z(n3102) );
  XNOR U4549 ( .A(n3100), .B(\w3[1][121] ), .Z(n3101) );
  XNOR U4550 ( .A(n3102), .B(n3101), .Z(\w1[2][113] ) );
  XOR U4551 ( .A(\w3[1][107] ), .B(\w3[1][115] ), .Z(n3136) );
  XOR U4552 ( .A(n3136), .B(key[370]), .Z(n3104) );
  XNOR U4553 ( .A(\w3[1][106] ), .B(n3466), .Z(n3103) );
  XNOR U4554 ( .A(n3104), .B(n3103), .Z(\w1[2][114] ) );
  XOR U4555 ( .A(\w3[1][116] ), .B(\w3[1][112] ), .Z(n3137) );
  XOR U4556 ( .A(n3137), .B(key[371]), .Z(n3107) );
  XNOR U4557 ( .A(\w3[1][107] ), .B(n3105), .Z(n3106) );
  XNOR U4558 ( .A(n3107), .B(n3106), .Z(\w1[2][115] ) );
  XOR U4559 ( .A(\w3[1][117] ), .B(\w3[1][112] ), .Z(n3140) );
  XOR U4560 ( .A(n3140), .B(key[372]), .Z(n3110) );
  XNOR U4561 ( .A(\w3[1][108] ), .B(n3108), .Z(n3109) );
  XNOR U4562 ( .A(n3110), .B(n3109), .Z(\w1[2][116] ) );
  XOR U4563 ( .A(n3111), .B(key[373]), .Z(n3114) );
  XNOR U4564 ( .A(\w3[1][109] ), .B(n3112), .Z(n3113) );
  XNOR U4565 ( .A(n3114), .B(n3113), .Z(\w1[2][117] ) );
  XOR U4566 ( .A(\w3[1][119] ), .B(\w3[1][112] ), .Z(n3148) );
  XOR U4567 ( .A(n3148), .B(key[374]), .Z(n3117) );
  XNOR U4568 ( .A(\w3[1][110] ), .B(n3115), .Z(n3116) );
  XNOR U4569 ( .A(n3117), .B(n3116), .Z(\w1[2][118] ) );
  XNOR U4570 ( .A(n3118), .B(key[375]), .Z(n3119) );
  XNOR U4571 ( .A(n3120), .B(n3119), .Z(n3121) );
  XNOR U4572 ( .A(\w3[1][112] ), .B(n3121), .Z(\w1[2][119] ) );
  XOR U4573 ( .A(\w3[1][3] ), .B(\w3[1][27] ), .Z(n3216) );
  XNOR U4574 ( .A(\w3[1][8] ), .B(\w3[1][12] ), .Z(n3122) );
  XNOR U4575 ( .A(n3216), .B(n3122), .Z(n3172) );
  XOR U4576 ( .A(n3172), .B(key[267]), .Z(n3124) );
  XOR U4577 ( .A(\w3[1][0] ), .B(\w3[1][4] ), .Z(n3246) );
  XNOR U4578 ( .A(\w3[1][19] ), .B(n3246), .Z(n3123) );
  XNOR U4579 ( .A(n3124), .B(n3123), .Z(\w1[2][11] ) );
  XOR U4580 ( .A(n3125), .B(key[376]), .Z(n3127) );
  XNOR U4581 ( .A(\w3[1][113] ), .B(\w3[1][121] ), .Z(n3126) );
  XNOR U4582 ( .A(n3127), .B(n3126), .Z(n3128) );
  XOR U4583 ( .A(\w3[1][112] ), .B(n3128), .Z(\w1[2][120] ) );
  XOR U4584 ( .A(n3465), .B(key[377]), .Z(n3130) );
  XNOR U4585 ( .A(\w3[1][114] ), .B(\w3[1][122] ), .Z(n3129) );
  XNOR U4586 ( .A(n3130), .B(n3129), .Z(n3131) );
  XOR U4587 ( .A(\w3[1][97] ), .B(n3131), .Z(\w1[2][121] ) );
  XOR U4588 ( .A(n3469), .B(key[378]), .Z(n3133) );
  XNOR U4589 ( .A(\w3[1][115] ), .B(\w3[1][123] ), .Z(n3132) );
  XNOR U4590 ( .A(n3133), .B(n3132), .Z(n3134) );
  XOR U4591 ( .A(\w3[1][98] ), .B(n3134), .Z(\w1[2][122] ) );
  XNOR U4592 ( .A(\w3[1][124] ), .B(\w3[1][120] ), .Z(n3135) );
  XNOR U4593 ( .A(n3136), .B(n3135), .Z(n3473) );
  XOR U4594 ( .A(n3473), .B(key[379]), .Z(n3139) );
  XNOR U4595 ( .A(\w3[1][99] ), .B(n3137), .Z(n3138) );
  XNOR U4596 ( .A(n3139), .B(n3138), .Z(\w1[2][123] ) );
  XOR U4597 ( .A(n3140), .B(key[380]), .Z(n3143) );
  XNOR U4598 ( .A(n3141), .B(\w3[1][100] ), .Z(n3142) );
  XNOR U4599 ( .A(n3143), .B(n3142), .Z(\w1[2][124] ) );
  XOR U4600 ( .A(\w3[1][118] ), .B(key[381]), .Z(n3146) );
  XNOR U4601 ( .A(n3144), .B(\w3[1][126] ), .Z(n3145) );
  XNOR U4602 ( .A(n3146), .B(n3145), .Z(n3147) );
  XOR U4603 ( .A(\w3[1][101] ), .B(n3147), .Z(\w1[2][125] ) );
  XOR U4604 ( .A(n3148), .B(key[382]), .Z(n3151) );
  XNOR U4605 ( .A(\w3[1][102] ), .B(n3149), .Z(n3150) );
  XNOR U4606 ( .A(n3151), .B(n3150), .Z(\w1[2][126] ) );
  XOR U4607 ( .A(n3462), .B(key[383]), .Z(n3154) );
  XNOR U4608 ( .A(\w3[1][103] ), .B(n3152), .Z(n3153) );
  XNOR U4609 ( .A(n3154), .B(n3153), .Z(\w1[2][127] ) );
  XOR U4610 ( .A(\w3[1][13] ), .B(\w3[1][28] ), .Z(n3156) );
  XNOR U4611 ( .A(\w3[1][8] ), .B(\w3[1][4] ), .Z(n3155) );
  XNOR U4612 ( .A(n3156), .B(n3155), .Z(n3178) );
  XOR U4613 ( .A(n3178), .B(key[268]), .Z(n3158) );
  XOR U4614 ( .A(\w3[1][0] ), .B(\w3[1][5] ), .Z(n3283) );
  XNOR U4615 ( .A(\w3[1][20] ), .B(n3283), .Z(n3157) );
  XNOR U4616 ( .A(n3158), .B(n3157), .Z(\w1[2][12] ) );
  XOR U4617 ( .A(\w3[1][14] ), .B(\w3[1][21] ), .Z(n3160) );
  XOR U4618 ( .A(\w3[1][5] ), .B(\w3[1][29] ), .Z(n3181) );
  XNOR U4619 ( .A(n3181), .B(key[269]), .Z(n3159) );
  XNOR U4620 ( .A(n3160), .B(n3159), .Z(n3161) );
  XOR U4621 ( .A(\w3[1][6] ), .B(n3161), .Z(\w1[2][13] ) );
  XOR U4622 ( .A(\w3[1][6] ), .B(\w3[1][30] ), .Z(n3324) );
  XNOR U4623 ( .A(\w3[1][8] ), .B(\w3[1][15] ), .Z(n3189) );
  XNOR U4624 ( .A(n3324), .B(n3189), .Z(n3184) );
  XOR U4625 ( .A(n3184), .B(key[270]), .Z(n3163) );
  XOR U4626 ( .A(\w3[1][0] ), .B(\w3[1][7] ), .Z(n3359) );
  XNOR U4627 ( .A(\w3[1][22] ), .B(n3359), .Z(n3162) );
  XNOR U4628 ( .A(n3163), .B(n3162), .Z(\w1[2][14] ) );
  XOR U4629 ( .A(\w3[1][7] ), .B(\w3[1][31] ), .Z(n3187) );
  XOR U4630 ( .A(n3187), .B(key[271]), .Z(n3165) );
  XOR U4631 ( .A(\w3[1][8] ), .B(\w3[1][0] ), .Z(n3191) );
  XNOR U4632 ( .A(\w3[1][23] ), .B(n3191), .Z(n3164) );
  XNOR U4633 ( .A(n3165), .B(n3164), .Z(\w1[2][15] ) );
  XOR U4634 ( .A(\w3[1][17] ), .B(\w3[1][9] ), .Z(n3195) );
  XOR U4635 ( .A(n3195), .B(key[272]), .Z(n3167) );
  XNOR U4636 ( .A(\w3[1][24] ), .B(n3191), .Z(n3166) );
  XNOR U4637 ( .A(n3167), .B(n3166), .Z(\w1[2][16] ) );
  XOR U4638 ( .A(\w3[1][18] ), .B(\w3[1][10] ), .Z(n3215) );
  XOR U4639 ( .A(n3215), .B(key[273]), .Z(n3169) );
  XNOR U4640 ( .A(n3480), .B(\w3[1][9] ), .Z(n3168) );
  XNOR U4641 ( .A(n3169), .B(n3168), .Z(\w1[2][17] ) );
  XOR U4642 ( .A(\w3[1][11] ), .B(\w3[1][19] ), .Z(n3203) );
  XOR U4643 ( .A(n3203), .B(key[274]), .Z(n3171) );
  XNOR U4644 ( .A(n3175), .B(\w3[1][10] ), .Z(n3170) );
  XNOR U4645 ( .A(n3171), .B(n3170), .Z(\w1[2][18] ) );
  XOR U4646 ( .A(\w3[1][16] ), .B(\w3[1][20] ), .Z(n3204) );
  XOR U4647 ( .A(n3204), .B(key[275]), .Z(n3174) );
  XNOR U4648 ( .A(\w3[1][11] ), .B(n3172), .Z(n3173) );
  XNOR U4649 ( .A(n3174), .B(n3173), .Z(\w1[2][19] ) );
  XOR U4650 ( .A(n3195), .B(key[257]), .Z(n3177) );
  XNOR U4651 ( .A(\w3[1][25] ), .B(n3175), .Z(n3176) );
  XNOR U4652 ( .A(n3177), .B(n3176), .Z(\w1[2][1] ) );
  XOR U4653 ( .A(\w3[1][16] ), .B(\w3[1][21] ), .Z(n3209) );
  XOR U4654 ( .A(n3209), .B(key[276]), .Z(n3180) );
  XNOR U4655 ( .A(\w3[1][12] ), .B(n3178), .Z(n3179) );
  XNOR U4656 ( .A(n3180), .B(n3179), .Z(\w1[2][20] ) );
  XOR U4657 ( .A(\w3[1][14] ), .B(\w3[1][22] ), .Z(n3219) );
  XOR U4658 ( .A(n3219), .B(key[277]), .Z(n3183) );
  XNOR U4659 ( .A(\w3[1][13] ), .B(n3181), .Z(n3182) );
  XNOR U4660 ( .A(n3183), .B(n3182), .Z(\w1[2][21] ) );
  XOR U4661 ( .A(\w3[1][16] ), .B(\w3[1][23] ), .Z(n3220) );
  XOR U4662 ( .A(n3220), .B(key[278]), .Z(n3186) );
  XNOR U4663 ( .A(\w3[1][14] ), .B(n3184), .Z(n3185) );
  XNOR U4664 ( .A(n3186), .B(n3185), .Z(\w1[2][22] ) );
  XNOR U4665 ( .A(n3187), .B(key[279]), .Z(n3188) );
  XNOR U4666 ( .A(n3189), .B(n3188), .Z(n3190) );
  XNOR U4667 ( .A(\w3[1][16] ), .B(n3190), .Z(\w1[2][23] ) );
  XOR U4668 ( .A(\w3[1][17] ), .B(key[280]), .Z(n3193) );
  XNOR U4669 ( .A(\w3[1][25] ), .B(n3191), .Z(n3192) );
  XNOR U4670 ( .A(n3193), .B(n3192), .Z(n3194) );
  XOR U4671 ( .A(\w3[1][16] ), .B(n3194), .Z(\w1[2][24] ) );
  XOR U4672 ( .A(n3195), .B(key[281]), .Z(n3197) );
  XNOR U4673 ( .A(\w3[1][1] ), .B(\w3[1][26] ), .Z(n3196) );
  XNOR U4674 ( .A(n3197), .B(n3196), .Z(n3198) );
  XOR U4675 ( .A(\w3[1][18] ), .B(n3198), .Z(\w1[2][25] ) );
  XOR U4676 ( .A(n3215), .B(key[282]), .Z(n3200) );
  XNOR U4677 ( .A(\w3[1][2] ), .B(\w3[1][19] ), .Z(n3199) );
  XNOR U4678 ( .A(n3200), .B(n3199), .Z(n3201) );
  XOR U4679 ( .A(\w3[1][27] ), .B(n3201), .Z(\w1[2][26] ) );
  XNOR U4680 ( .A(\w3[1][24] ), .B(\w3[1][28] ), .Z(n3202) );
  XNOR U4681 ( .A(n3203), .B(n3202), .Z(n3245) );
  XOR U4682 ( .A(n3245), .B(key[283]), .Z(n3206) );
  XNOR U4683 ( .A(\w3[1][3] ), .B(n3204), .Z(n3205) );
  XNOR U4684 ( .A(n3206), .B(n3205), .Z(\w1[2][27] ) );
  XOR U4685 ( .A(\w3[1][20] ), .B(\w3[1][29] ), .Z(n3208) );
  XNOR U4686 ( .A(\w3[1][24] ), .B(\w3[1][12] ), .Z(n3207) );
  XNOR U4687 ( .A(n3208), .B(n3207), .Z(n3282) );
  XOR U4688 ( .A(n3282), .B(key[284]), .Z(n3211) );
  XNOR U4689 ( .A(\w3[1][4] ), .B(n3209), .Z(n3210) );
  XNOR U4690 ( .A(n3211), .B(n3210), .Z(\w1[2][28] ) );
  XOR U4691 ( .A(\w3[1][13] ), .B(\w3[1][21] ), .Z(n3323) );
  XOR U4692 ( .A(n3323), .B(key[285]), .Z(n3213) );
  XNOR U4693 ( .A(\w3[1][22] ), .B(\w3[1][30] ), .Z(n3212) );
  XNOR U4694 ( .A(n3213), .B(n3212), .Z(n3214) );
  XOR U4695 ( .A(\w3[1][5] ), .B(n3214), .Z(\w1[2][29] ) );
  XOR U4696 ( .A(n3215), .B(key[258]), .Z(n3218) );
  XNOR U4697 ( .A(\w3[1][26] ), .B(n3216), .Z(n3217) );
  XNOR U4698 ( .A(n3218), .B(n3217), .Z(\w1[2][2] ) );
  XNOR U4699 ( .A(\w3[1][24] ), .B(\w3[1][31] ), .Z(n3397) );
  XNOR U4700 ( .A(n3219), .B(n3397), .Z(n3358) );
  XOR U4701 ( .A(n3358), .B(key[286]), .Z(n3222) );
  XNOR U4702 ( .A(\w3[1][6] ), .B(n3220), .Z(n3221) );
  XNOR U4703 ( .A(n3222), .B(n3221), .Z(\w1[2][30] ) );
  XOR U4704 ( .A(\w3[1][15] ), .B(\w3[1][23] ), .Z(n3395) );
  XOR U4705 ( .A(n3395), .B(key[287]), .Z(n3224) );
  XNOR U4706 ( .A(n3436), .B(\w3[1][7] ), .Z(n3223) );
  XNOR U4707 ( .A(n3224), .B(n3223), .Z(\w1[2][31] ) );
  XOR U4708 ( .A(\w3[1][33] ), .B(\w3[1][57] ), .Z(n3279) );
  XOR U4709 ( .A(n3279), .B(key[288]), .Z(n3226) );
  XOR U4710 ( .A(\w3[1][48] ), .B(\w3[1][56] ), .Z(n3340) );
  XNOR U4711 ( .A(n3340), .B(\w3[1][40] ), .Z(n3225) );
  XNOR U4712 ( .A(n3226), .B(n3225), .Z(\w1[2][32] ) );
  XOR U4713 ( .A(\w3[1][34] ), .B(\w3[1][58] ), .Z(n3287) );
  XOR U4714 ( .A(n3287), .B(key[289]), .Z(n3228) );
  XOR U4715 ( .A(\w3[1][41] ), .B(\w3[1][49] ), .Z(n3311) );
  XNOR U4716 ( .A(\w3[1][57] ), .B(n3311), .Z(n3227) );
  XNOR U4717 ( .A(n3228), .B(n3227), .Z(\w1[2][33] ) );
  XOR U4718 ( .A(\w3[1][35] ), .B(\w3[1][59] ), .Z(n3258) );
  XOR U4719 ( .A(n3258), .B(key[290]), .Z(n3230) );
  XOR U4720 ( .A(\w3[1][42] ), .B(\w3[1][50] ), .Z(n3315) );
  XNOR U4721 ( .A(\w3[1][58] ), .B(n3315), .Z(n3229) );
  XNOR U4722 ( .A(n3230), .B(n3229), .Z(\w1[2][34] ) );
  XOR U4723 ( .A(\w3[1][36] ), .B(\w3[1][32] ), .Z(n3260) );
  XOR U4724 ( .A(n3260), .B(key[291]), .Z(n3233) );
  XOR U4725 ( .A(\w3[1][43] ), .B(\w3[1][51] ), .Z(n3286) );
  XNOR U4726 ( .A(\w3[1][56] ), .B(n3286), .Z(n3231) );
  XNOR U4727 ( .A(\w3[1][60] ), .B(n3231), .Z(n3320) );
  XNOR U4728 ( .A(\w3[1][59] ), .B(n3320), .Z(n3232) );
  XNOR U4729 ( .A(n3233), .B(n3232), .Z(\w1[2][35] ) );
  XOR U4730 ( .A(\w3[1][32] ), .B(\w3[1][37] ), .Z(n3265) );
  XOR U4731 ( .A(n3265), .B(key[292]), .Z(n3237) );
  XOR U4732 ( .A(\w3[1][52] ), .B(\w3[1][61] ), .Z(n3235) );
  XNOR U4733 ( .A(\w3[1][56] ), .B(\w3[1][44] ), .Z(n3234) );
  XNOR U4734 ( .A(n3235), .B(n3234), .Z(n3328) );
  XNOR U4735 ( .A(\w3[1][60] ), .B(n3328), .Z(n3236) );
  XNOR U4736 ( .A(n3237), .B(n3236), .Z(\w1[2][36] ) );
  XOR U4737 ( .A(\w3[1][38] ), .B(\w3[1][62] ), .Z(n3271) );
  XOR U4738 ( .A(n3271), .B(key[293]), .Z(n3239) );
  XOR U4739 ( .A(\w3[1][45] ), .B(\w3[1][53] ), .Z(n3331) );
  XNOR U4740 ( .A(\w3[1][61] ), .B(n3331), .Z(n3238) );
  XNOR U4741 ( .A(n3239), .B(n3238), .Z(\w1[2][37] ) );
  XOR U4742 ( .A(\w3[1][32] ), .B(\w3[1][39] ), .Z(n3272) );
  XOR U4743 ( .A(n3272), .B(key[294]), .Z(n3241) );
  XOR U4744 ( .A(\w3[1][46] ), .B(\w3[1][54] ), .Z(n3297) );
  XNOR U4745 ( .A(\w3[1][56] ), .B(\w3[1][63] ), .Z(n3243) );
  XNOR U4746 ( .A(n3297), .B(n3243), .Z(n3336) );
  XNOR U4747 ( .A(\w3[1][62] ), .B(n3336), .Z(n3240) );
  XNOR U4748 ( .A(n3241), .B(n3240), .Z(\w1[2][38] ) );
  XOR U4749 ( .A(\w3[1][47] ), .B(\w3[1][55] ), .Z(n3339) );
  XNOR U4750 ( .A(n3339), .B(key[295]), .Z(n3242) );
  XNOR U4751 ( .A(n3243), .B(n3242), .Z(n3244) );
  XNOR U4752 ( .A(\w3[1][32] ), .B(n3244), .Z(\w1[2][39] ) );
  XOR U4753 ( .A(n3245), .B(key[259]), .Z(n3248) );
  XNOR U4754 ( .A(n3246), .B(\w3[1][27] ), .Z(n3247) );
  XNOR U4755 ( .A(n3248), .B(n3247), .Z(\w1[2][3] ) );
  XOR U4756 ( .A(\w3[1][32] ), .B(key[296]), .Z(n3250) );
  XNOR U4757 ( .A(\w3[1][33] ), .B(\w3[1][41] ), .Z(n3249) );
  XNOR U4758 ( .A(n3250), .B(n3249), .Z(n3251) );
  XOR U4759 ( .A(n3340), .B(n3251), .Z(\w1[2][40] ) );
  XOR U4760 ( .A(\w3[1][42] ), .B(key[297]), .Z(n3253) );
  XNOR U4761 ( .A(\w3[1][49] ), .B(\w3[1][34] ), .Z(n3252) );
  XNOR U4762 ( .A(n3253), .B(n3252), .Z(n3254) );
  XOR U4763 ( .A(n3279), .B(n3254), .Z(\w1[2][41] ) );
  XOR U4764 ( .A(\w3[1][43] ), .B(key[298]), .Z(n3256) );
  XNOR U4765 ( .A(\w3[1][50] ), .B(\w3[1][35] ), .Z(n3255) );
  XNOR U4766 ( .A(n3256), .B(n3255), .Z(n3257) );
  XOR U4767 ( .A(n3287), .B(n3257), .Z(\w1[2][42] ) );
  XNOR U4768 ( .A(\w3[1][40] ), .B(n3258), .Z(n3259) );
  XNOR U4769 ( .A(\w3[1][44] ), .B(n3259), .Z(n3290) );
  XOR U4770 ( .A(n3290), .B(key[299]), .Z(n3262) );
  XNOR U4771 ( .A(\w3[1][51] ), .B(n3260), .Z(n3261) );
  XNOR U4772 ( .A(n3262), .B(n3261), .Z(\w1[2][43] ) );
  XOR U4773 ( .A(\w3[1][36] ), .B(\w3[1][45] ), .Z(n3264) );
  XNOR U4774 ( .A(\w3[1][40] ), .B(\w3[1][60] ), .Z(n3263) );
  XNOR U4775 ( .A(n3264), .B(n3263), .Z(n3293) );
  XOR U4776 ( .A(n3293), .B(key[300]), .Z(n3267) );
  XNOR U4777 ( .A(\w3[1][52] ), .B(n3265), .Z(n3266) );
  XNOR U4778 ( .A(n3267), .B(n3266), .Z(\w1[2][44] ) );
  XOR U4779 ( .A(\w3[1][61] ), .B(\w3[1][37] ), .Z(n3296) );
  XOR U4780 ( .A(n3296), .B(key[301]), .Z(n3269) );
  XNOR U4781 ( .A(\w3[1][38] ), .B(\w3[1][46] ), .Z(n3268) );
  XNOR U4782 ( .A(n3269), .B(n3268), .Z(n3270) );
  XOR U4783 ( .A(\w3[1][53] ), .B(n3270), .Z(\w1[2][45] ) );
  XNOR U4784 ( .A(\w3[1][40] ), .B(\w3[1][47] ), .Z(n3305) );
  XNOR U4785 ( .A(n3271), .B(n3305), .Z(n3300) );
  XOR U4786 ( .A(n3300), .B(key[302]), .Z(n3274) );
  XNOR U4787 ( .A(\w3[1][54] ), .B(n3272), .Z(n3273) );
  XNOR U4788 ( .A(n3274), .B(n3273), .Z(\w1[2][46] ) );
  XOR U4789 ( .A(\w3[1][63] ), .B(\w3[1][39] ), .Z(n3303) );
  XOR U4790 ( .A(n3303), .B(key[303]), .Z(n3276) );
  XOR U4791 ( .A(\w3[1][40] ), .B(\w3[1][32] ), .Z(n3307) );
  XNOR U4792 ( .A(\w3[1][55] ), .B(n3307), .Z(n3275) );
  XNOR U4793 ( .A(n3276), .B(n3275), .Z(\w1[2][47] ) );
  XOR U4794 ( .A(n3307), .B(key[304]), .Z(n3278) );
  XNOR U4795 ( .A(\w3[1][56] ), .B(n3311), .Z(n3277) );
  XNOR U4796 ( .A(n3278), .B(n3277), .Z(\w1[2][48] ) );
  XOR U4797 ( .A(n3315), .B(key[305]), .Z(n3281) );
  XNOR U4798 ( .A(n3279), .B(\w3[1][41] ), .Z(n3280) );
  XNOR U4799 ( .A(n3281), .B(n3280), .Z(\w1[2][49] ) );
  XOR U4800 ( .A(n3282), .B(key[260]), .Z(n3285) );
  XNOR U4801 ( .A(n3283), .B(\w3[1][28] ), .Z(n3284) );
  XNOR U4802 ( .A(n3285), .B(n3284), .Z(\w1[2][4] ) );
  XOR U4803 ( .A(n3286), .B(key[306]), .Z(n3289) );
  XNOR U4804 ( .A(n3287), .B(\w3[1][42] ), .Z(n3288) );
  XNOR U4805 ( .A(n3289), .B(n3288), .Z(\w1[2][50] ) );
  XOR U4806 ( .A(\w3[1][48] ), .B(\w3[1][52] ), .Z(n3319) );
  XOR U4807 ( .A(n3319), .B(key[307]), .Z(n3292) );
  XNOR U4808 ( .A(\w3[1][43] ), .B(n3290), .Z(n3291) );
  XNOR U4809 ( .A(n3292), .B(n3291), .Z(\w1[2][51] ) );
  XOR U4810 ( .A(\w3[1][48] ), .B(\w3[1][53] ), .Z(n3327) );
  XOR U4811 ( .A(n3327), .B(key[308]), .Z(n3295) );
  XNOR U4812 ( .A(\w3[1][44] ), .B(n3293), .Z(n3294) );
  XNOR U4813 ( .A(n3295), .B(n3294), .Z(\w1[2][52] ) );
  XOR U4814 ( .A(n3296), .B(key[309]), .Z(n3299) );
  XNOR U4815 ( .A(\w3[1][45] ), .B(n3297), .Z(n3298) );
  XNOR U4816 ( .A(n3299), .B(n3298), .Z(\w1[2][53] ) );
  XOR U4817 ( .A(\w3[1][48] ), .B(\w3[1][55] ), .Z(n3335) );
  XOR U4818 ( .A(n3335), .B(key[310]), .Z(n3302) );
  XNOR U4819 ( .A(\w3[1][46] ), .B(n3300), .Z(n3301) );
  XNOR U4820 ( .A(n3302), .B(n3301), .Z(\w1[2][54] ) );
  XNOR U4821 ( .A(n3303), .B(key[311]), .Z(n3304) );
  XNOR U4822 ( .A(n3305), .B(n3304), .Z(n3306) );
  XNOR U4823 ( .A(\w3[1][48] ), .B(n3306), .Z(\w1[2][55] ) );
  XOR U4824 ( .A(n3307), .B(key[312]), .Z(n3309) );
  XNOR U4825 ( .A(\w3[1][48] ), .B(\w3[1][49] ), .Z(n3308) );
  XNOR U4826 ( .A(n3309), .B(n3308), .Z(n3310) );
  XOR U4827 ( .A(\w3[1][57] ), .B(n3310), .Z(\w1[2][56] ) );
  XOR U4828 ( .A(\w3[1][50] ), .B(key[313]), .Z(n3313) );
  XNOR U4829 ( .A(n3311), .B(\w3[1][58] ), .Z(n3312) );
  XNOR U4830 ( .A(n3313), .B(n3312), .Z(n3314) );
  XOR U4831 ( .A(\w3[1][33] ), .B(n3314), .Z(\w1[2][57] ) );
  XOR U4832 ( .A(\w3[1][51] ), .B(key[314]), .Z(n3317) );
  XNOR U4833 ( .A(n3315), .B(\w3[1][59] ), .Z(n3316) );
  XNOR U4834 ( .A(n3317), .B(n3316), .Z(n3318) );
  XOR U4835 ( .A(\w3[1][34] ), .B(n3318), .Z(\w1[2][58] ) );
  XOR U4836 ( .A(n3319), .B(key[315]), .Z(n3322) );
  XNOR U4837 ( .A(\w3[1][35] ), .B(n3320), .Z(n3321) );
  XNOR U4838 ( .A(n3322), .B(n3321), .Z(\w1[2][59] ) );
  XOR U4839 ( .A(n3323), .B(key[261]), .Z(n3326) );
  XNOR U4840 ( .A(\w3[1][29] ), .B(n3324), .Z(n3325) );
  XNOR U4841 ( .A(n3326), .B(n3325), .Z(\w1[2][5] ) );
  XOR U4842 ( .A(n3327), .B(key[316]), .Z(n3330) );
  XNOR U4843 ( .A(\w3[1][36] ), .B(n3328), .Z(n3329) );
  XNOR U4844 ( .A(n3330), .B(n3329), .Z(\w1[2][60] ) );
  XOR U4845 ( .A(\w3[1][54] ), .B(key[317]), .Z(n3333) );
  XNOR U4846 ( .A(n3331), .B(\w3[1][62] ), .Z(n3332) );
  XNOR U4847 ( .A(n3333), .B(n3332), .Z(n3334) );
  XOR U4848 ( .A(\w3[1][37] ), .B(n3334), .Z(\w1[2][61] ) );
  XOR U4849 ( .A(n3335), .B(key[318]), .Z(n3338) );
  XNOR U4850 ( .A(\w3[1][38] ), .B(n3336), .Z(n3337) );
  XNOR U4851 ( .A(n3338), .B(n3337), .Z(\w1[2][62] ) );
  XOR U4852 ( .A(n3339), .B(key[319]), .Z(n3342) );
  XNOR U4853 ( .A(n3340), .B(\w3[1][39] ), .Z(n3341) );
  XNOR U4854 ( .A(n3342), .B(n3341), .Z(\w1[2][63] ) );
  XOR U4855 ( .A(\w3[1][65] ), .B(\w3[1][89] ), .Z(n3401) );
  XOR U4856 ( .A(n3401), .B(key[320]), .Z(n3344) );
  XOR U4857 ( .A(\w3[1][80] ), .B(\w3[1][88] ), .Z(n3458) );
  XNOR U4858 ( .A(n3458), .B(\w3[1][72] ), .Z(n3343) );
  XNOR U4859 ( .A(n3344), .B(n3343), .Z(\w1[2][64] ) );
  XOR U4860 ( .A(\w3[1][66] ), .B(\w3[1][90] ), .Z(n3405) );
  XOR U4861 ( .A(n3405), .B(key[321]), .Z(n3346) );
  XOR U4862 ( .A(\w3[1][73] ), .B(\w3[1][81] ), .Z(n3429) );
  XNOR U4863 ( .A(\w3[1][89] ), .B(n3429), .Z(n3345) );
  XNOR U4864 ( .A(n3346), .B(n3345), .Z(\w1[2][65] ) );
  XOR U4865 ( .A(\w3[1][67] ), .B(\w3[1][91] ), .Z(n3376) );
  XOR U4866 ( .A(n3376), .B(key[322]), .Z(n3348) );
  XOR U4867 ( .A(\w3[1][74] ), .B(\w3[1][82] ), .Z(n3437) );
  XNOR U4868 ( .A(\w3[1][90] ), .B(n3437), .Z(n3347) );
  XNOR U4869 ( .A(n3348), .B(n3347), .Z(\w1[2][66] ) );
  XOR U4870 ( .A(\w3[1][68] ), .B(\w3[1][64] ), .Z(n3378) );
  XOR U4871 ( .A(n3378), .B(key[323]), .Z(n3351) );
  XOR U4872 ( .A(\w3[1][75] ), .B(\w3[1][83] ), .Z(n3404) );
  XNOR U4873 ( .A(\w3[1][88] ), .B(n3404), .Z(n3349) );
  XNOR U4874 ( .A(\w3[1][92] ), .B(n3349), .Z(n3442) );
  XNOR U4875 ( .A(\w3[1][91] ), .B(n3442), .Z(n3350) );
  XNOR U4876 ( .A(n3351), .B(n3350), .Z(\w1[2][67] ) );
  XOR U4877 ( .A(\w3[1][64] ), .B(\w3[1][69] ), .Z(n3383) );
  XOR U4878 ( .A(n3383), .B(key[324]), .Z(n3355) );
  XOR U4879 ( .A(\w3[1][84] ), .B(\w3[1][93] ), .Z(n3353) );
  XNOR U4880 ( .A(\w3[1][88] ), .B(\w3[1][76] ), .Z(n3352) );
  XNOR U4881 ( .A(n3353), .B(n3352), .Z(n3446) );
  XNOR U4882 ( .A(\w3[1][92] ), .B(n3446), .Z(n3354) );
  XNOR U4883 ( .A(n3355), .B(n3354), .Z(\w1[2][68] ) );
  XOR U4884 ( .A(\w3[1][70] ), .B(\w3[1][94] ), .Z(n3389) );
  XOR U4885 ( .A(n3389), .B(key[325]), .Z(n3357) );
  XOR U4886 ( .A(\w3[1][77] ), .B(\w3[1][85] ), .Z(n3449) );
  XNOR U4887 ( .A(\w3[1][93] ), .B(n3449), .Z(n3356) );
  XNOR U4888 ( .A(n3357), .B(n3356), .Z(\w1[2][69] ) );
  XOR U4889 ( .A(n3358), .B(key[262]), .Z(n3361) );
  XNOR U4890 ( .A(n3359), .B(\w3[1][30] ), .Z(n3360) );
  XNOR U4891 ( .A(n3361), .B(n3360), .Z(\w1[2][6] ) );
  XOR U4892 ( .A(\w3[1][64] ), .B(\w3[1][71] ), .Z(n3390) );
  XOR U4893 ( .A(n3390), .B(key[326]), .Z(n3363) );
  XOR U4894 ( .A(\w3[1][78] ), .B(\w3[1][86] ), .Z(n3415) );
  XNOR U4895 ( .A(\w3[1][88] ), .B(\w3[1][95] ), .Z(n3365) );
  XNOR U4896 ( .A(n3415), .B(n3365), .Z(n3454) );
  XNOR U4897 ( .A(\w3[1][94] ), .B(n3454), .Z(n3362) );
  XNOR U4898 ( .A(n3363), .B(n3362), .Z(\w1[2][70] ) );
  XOR U4899 ( .A(\w3[1][79] ), .B(\w3[1][87] ), .Z(n3457) );
  XNOR U4900 ( .A(n3457), .B(key[327]), .Z(n3364) );
  XNOR U4901 ( .A(n3365), .B(n3364), .Z(n3366) );
  XNOR U4902 ( .A(\w3[1][64] ), .B(n3366), .Z(\w1[2][71] ) );
  XOR U4903 ( .A(\w3[1][64] ), .B(key[328]), .Z(n3368) );
  XNOR U4904 ( .A(\w3[1][65] ), .B(\w3[1][73] ), .Z(n3367) );
  XNOR U4905 ( .A(n3368), .B(n3367), .Z(n3369) );
  XOR U4906 ( .A(n3458), .B(n3369), .Z(\w1[2][72] ) );
  XOR U4907 ( .A(\w3[1][74] ), .B(key[329]), .Z(n3371) );
  XNOR U4908 ( .A(\w3[1][81] ), .B(\w3[1][66] ), .Z(n3370) );
  XNOR U4909 ( .A(n3371), .B(n3370), .Z(n3372) );
  XOR U4910 ( .A(n3401), .B(n3372), .Z(\w1[2][73] ) );
  XOR U4911 ( .A(\w3[1][75] ), .B(key[330]), .Z(n3374) );
  XNOR U4912 ( .A(\w3[1][82] ), .B(\w3[1][67] ), .Z(n3373) );
  XNOR U4913 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4914 ( .A(n3405), .B(n3375), .Z(\w1[2][74] ) );
  XNOR U4915 ( .A(\w3[1][72] ), .B(n3376), .Z(n3377) );
  XNOR U4916 ( .A(\w3[1][76] ), .B(n3377), .Z(n3408) );
  XOR U4917 ( .A(n3408), .B(key[331]), .Z(n3380) );
  XNOR U4918 ( .A(\w3[1][83] ), .B(n3378), .Z(n3379) );
  XNOR U4919 ( .A(n3380), .B(n3379), .Z(\w1[2][75] ) );
  XOR U4920 ( .A(\w3[1][68] ), .B(\w3[1][77] ), .Z(n3382) );
  XNOR U4921 ( .A(\w3[1][72] ), .B(\w3[1][92] ), .Z(n3381) );
  XNOR U4922 ( .A(n3382), .B(n3381), .Z(n3411) );
  XOR U4923 ( .A(n3411), .B(key[332]), .Z(n3385) );
  XNOR U4924 ( .A(\w3[1][84] ), .B(n3383), .Z(n3384) );
  XNOR U4925 ( .A(n3385), .B(n3384), .Z(\w1[2][76] ) );
  XOR U4926 ( .A(\w3[1][93] ), .B(\w3[1][69] ), .Z(n3414) );
  XOR U4927 ( .A(n3414), .B(key[333]), .Z(n3387) );
  XNOR U4928 ( .A(\w3[1][70] ), .B(\w3[1][78] ), .Z(n3386) );
  XNOR U4929 ( .A(n3387), .B(n3386), .Z(n3388) );
  XOR U4930 ( .A(\w3[1][85] ), .B(n3388), .Z(\w1[2][77] ) );
  XNOR U4931 ( .A(\w3[1][72] ), .B(\w3[1][79] ), .Z(n3423) );
  XNOR U4932 ( .A(n3389), .B(n3423), .Z(n3418) );
  XOR U4933 ( .A(n3418), .B(key[334]), .Z(n3392) );
  XNOR U4934 ( .A(\w3[1][86] ), .B(n3390), .Z(n3391) );
  XNOR U4935 ( .A(n3392), .B(n3391), .Z(\w1[2][78] ) );
  XOR U4936 ( .A(\w3[1][95] ), .B(\w3[1][71] ), .Z(n3421) );
  XOR U4937 ( .A(n3421), .B(key[335]), .Z(n3394) );
  XOR U4938 ( .A(\w3[1][72] ), .B(\w3[1][64] ), .Z(n3425) );
  XNOR U4939 ( .A(\w3[1][87] ), .B(n3425), .Z(n3393) );
  XNOR U4940 ( .A(n3394), .B(n3393), .Z(\w1[2][79] ) );
  XNOR U4941 ( .A(n3395), .B(key[263]), .Z(n3396) );
  XNOR U4942 ( .A(n3397), .B(n3396), .Z(n3398) );
  XNOR U4943 ( .A(\w3[1][0] ), .B(n3398), .Z(\w1[2][7] ) );
  XOR U4944 ( .A(n3425), .B(key[336]), .Z(n3400) );
  XNOR U4945 ( .A(\w3[1][88] ), .B(n3429), .Z(n3399) );
  XNOR U4946 ( .A(n3400), .B(n3399), .Z(\w1[2][80] ) );
  XOR U4947 ( .A(n3437), .B(key[337]), .Z(n3403) );
  XNOR U4948 ( .A(n3401), .B(\w3[1][73] ), .Z(n3402) );
  XNOR U4949 ( .A(n3403), .B(n3402), .Z(\w1[2][81] ) );
  XOR U4950 ( .A(n3404), .B(key[338]), .Z(n3407) );
  XNOR U4951 ( .A(n3405), .B(\w3[1][74] ), .Z(n3406) );
  XNOR U4952 ( .A(n3407), .B(n3406), .Z(\w1[2][82] ) );
  XOR U4953 ( .A(\w3[1][80] ), .B(\w3[1][84] ), .Z(n3441) );
  XOR U4954 ( .A(n3441), .B(key[339]), .Z(n3410) );
  XNOR U4955 ( .A(\w3[1][75] ), .B(n3408), .Z(n3409) );
  XNOR U4956 ( .A(n3410), .B(n3409), .Z(\w1[2][83] ) );
  XOR U4957 ( .A(\w3[1][80] ), .B(\w3[1][85] ), .Z(n3445) );
  XOR U4958 ( .A(n3445), .B(key[340]), .Z(n3413) );
  XNOR U4959 ( .A(\w3[1][76] ), .B(n3411), .Z(n3412) );
  XNOR U4960 ( .A(n3413), .B(n3412), .Z(\w1[2][84] ) );
  XOR U4961 ( .A(n3414), .B(key[341]), .Z(n3417) );
  XNOR U4962 ( .A(\w3[1][77] ), .B(n3415), .Z(n3416) );
  XNOR U4963 ( .A(n3417), .B(n3416), .Z(\w1[2][85] ) );
  XOR U4964 ( .A(\w3[1][80] ), .B(\w3[1][87] ), .Z(n3453) );
  XOR U4965 ( .A(n3453), .B(key[342]), .Z(n3420) );
  XNOR U4966 ( .A(\w3[1][78] ), .B(n3418), .Z(n3419) );
  XNOR U4967 ( .A(n3420), .B(n3419), .Z(\w1[2][86] ) );
  XNOR U4968 ( .A(n3421), .B(key[343]), .Z(n3422) );
  XNOR U4969 ( .A(n3423), .B(n3422), .Z(n3424) );
  XNOR U4970 ( .A(\w3[1][80] ), .B(n3424), .Z(\w1[2][87] ) );
  XOR U4971 ( .A(n3425), .B(key[344]), .Z(n3427) );
  XNOR U4972 ( .A(\w3[1][80] ), .B(\w3[1][81] ), .Z(n3426) );
  XNOR U4973 ( .A(n3427), .B(n3426), .Z(n3428) );
  XOR U4974 ( .A(\w3[1][89] ), .B(n3428), .Z(\w1[2][88] ) );
  XOR U4975 ( .A(\w3[1][82] ), .B(key[345]), .Z(n3431) );
  XNOR U4976 ( .A(n3429), .B(\w3[1][90] ), .Z(n3430) );
  XNOR U4977 ( .A(n3431), .B(n3430), .Z(n3432) );
  XOR U4978 ( .A(\w3[1][65] ), .B(n3432), .Z(\w1[2][89] ) );
  XOR U4979 ( .A(\w3[1][9] ), .B(key[264]), .Z(n3434) );
  XNOR U4980 ( .A(\w3[1][1] ), .B(\w3[1][0] ), .Z(n3433) );
  XNOR U4981 ( .A(n3434), .B(n3433), .Z(n3435) );
  XOR U4982 ( .A(n3436), .B(n3435), .Z(\w1[2][8] ) );
  XOR U4983 ( .A(\w3[1][83] ), .B(key[346]), .Z(n3439) );
  XNOR U4984 ( .A(n3437), .B(\w3[1][91] ), .Z(n3438) );
  XNOR U4985 ( .A(n3439), .B(n3438), .Z(n3440) );
  XOR U4986 ( .A(\w3[1][66] ), .B(n3440), .Z(\w1[2][90] ) );
  XOR U4987 ( .A(n3441), .B(key[347]), .Z(n3444) );
  XNOR U4988 ( .A(\w3[1][67] ), .B(n3442), .Z(n3443) );
  XNOR U4989 ( .A(n3444), .B(n3443), .Z(\w1[2][91] ) );
  XOR U4990 ( .A(n3445), .B(key[348]), .Z(n3448) );
  XNOR U4991 ( .A(\w3[1][68] ), .B(n3446), .Z(n3447) );
  XNOR U4992 ( .A(n3448), .B(n3447), .Z(\w1[2][92] ) );
  XOR U4993 ( .A(\w3[1][86] ), .B(key[349]), .Z(n3451) );
  XNOR U4994 ( .A(n3449), .B(\w3[1][94] ), .Z(n3450) );
  XNOR U4995 ( .A(n3451), .B(n3450), .Z(n3452) );
  XOR U4996 ( .A(\w3[1][69] ), .B(n3452), .Z(\w1[2][93] ) );
  XOR U4997 ( .A(n3453), .B(key[350]), .Z(n3456) );
  XNOR U4998 ( .A(\w3[1][70] ), .B(n3454), .Z(n3455) );
  XNOR U4999 ( .A(n3456), .B(n3455), .Z(\w1[2][94] ) );
  XOR U5000 ( .A(n3457), .B(key[351]), .Z(n3460) );
  XNOR U5001 ( .A(n3458), .B(\w3[1][71] ), .Z(n3459) );
  XNOR U5002 ( .A(n3460), .B(n3459), .Z(\w1[2][95] ) );
  XOR U5003 ( .A(\w3[1][104] ), .B(key[352]), .Z(n3464) );
  XNOR U5004 ( .A(n3462), .B(n3461), .Z(n3463) );
  XNOR U5005 ( .A(n3464), .B(n3463), .Z(\w1[2][96] ) );
  XOR U5006 ( .A(n3465), .B(key[353]), .Z(n3468) );
  XNOR U5007 ( .A(\w3[1][121] ), .B(n3466), .Z(n3467) );
  XNOR U5008 ( .A(n3468), .B(n3467), .Z(\w1[2][97] ) );
  XOR U5009 ( .A(n3469), .B(key[354]), .Z(n3472) );
  XNOR U5010 ( .A(\w3[1][122] ), .B(n3470), .Z(n3471) );
  XNOR U5011 ( .A(n3472), .B(n3471), .Z(\w1[2][98] ) );
  XOR U5012 ( .A(n3473), .B(key[355]), .Z(n3476) );
  XNOR U5013 ( .A(n3474), .B(\w3[1][123] ), .Z(n3475) );
  XNOR U5014 ( .A(n3476), .B(n3475), .Z(\w1[2][99] ) );
  XOR U5015 ( .A(\w3[1][10] ), .B(key[265]), .Z(n3478) );
  XNOR U5016 ( .A(\w3[1][2] ), .B(\w3[1][17] ), .Z(n3477) );
  XNOR U5017 ( .A(n3478), .B(n3477), .Z(n3479) );
  XOR U5018 ( .A(n3480), .B(n3479), .Z(\w1[2][9] ) );
  XOR U5019 ( .A(\w3[2][8] ), .B(key[384]), .Z(n3482) );
  XOR U5020 ( .A(\w3[2][1] ), .B(\w3[2][25] ), .Z(n3904) );
  XOR U5021 ( .A(\w3[2][16] ), .B(\w3[2][24] ), .Z(n3860) );
  XNOR U5022 ( .A(n3904), .B(n3860), .Z(n3481) );
  XNOR U5023 ( .A(n3482), .B(n3481), .Z(\w1[3][0] ) );
  XOR U5024 ( .A(\w3[2][96] ), .B(\w3[2][101] ), .Z(n3508) );
  XOR U5025 ( .A(n3508), .B(key[484]), .Z(n3486) );
  XOR U5026 ( .A(\w3[2][116] ), .B(\w3[2][125] ), .Z(n3484) );
  XNOR U5027 ( .A(\w3[2][120] ), .B(\w3[2][108] ), .Z(n3483) );
  XNOR U5028 ( .A(n3484), .B(n3483), .Z(n3565) );
  XNOR U5029 ( .A(\w3[2][124] ), .B(n3565), .Z(n3485) );
  XNOR U5030 ( .A(n3486), .B(n3485), .Z(\w1[3][100] ) );
  XOR U5031 ( .A(\w3[2][102] ), .B(\w3[2][126] ), .Z(n3517) );
  XOR U5032 ( .A(n3517), .B(key[485]), .Z(n3488) );
  XOR U5033 ( .A(\w3[2][109] ), .B(\w3[2][117] ), .Z(n3568) );
  XNOR U5034 ( .A(\w3[2][125] ), .B(n3568), .Z(n3487) );
  XNOR U5035 ( .A(n3488), .B(n3487), .Z(\w1[3][101] ) );
  XOR U5036 ( .A(\w3[2][96] ), .B(\w3[2][103] ), .Z(n3518) );
  XOR U5037 ( .A(n3518), .B(key[486]), .Z(n3490) );
  XOR U5038 ( .A(\w3[2][110] ), .B(\w3[2][118] ), .Z(n3536) );
  XNOR U5039 ( .A(\w3[2][120] ), .B(\w3[2][127] ), .Z(n3492) );
  XNOR U5040 ( .A(n3536), .B(n3492), .Z(n3573) );
  XNOR U5041 ( .A(\w3[2][126] ), .B(n3573), .Z(n3489) );
  XNOR U5042 ( .A(n3490), .B(n3489), .Z(\w1[3][102] ) );
  XOR U5043 ( .A(\w3[2][111] ), .B(\w3[2][119] ), .Z(n3576) );
  XNOR U5044 ( .A(n3576), .B(key[487]), .Z(n3491) );
  XNOR U5045 ( .A(n3492), .B(n3491), .Z(n3493) );
  XNOR U5046 ( .A(\w3[2][96] ), .B(n3493), .Z(\w1[3][103] ) );
  XOR U5047 ( .A(key[488]), .B(\w3[2][105] ), .Z(n3495) );
  XNOR U5048 ( .A(\w3[2][96] ), .B(\w3[2][97] ), .Z(n3494) );
  XNOR U5049 ( .A(n3495), .B(n3494), .Z(n3496) );
  XNOR U5050 ( .A(\w3[2][120] ), .B(\w3[2][112] ), .Z(n3886) );
  XNOR U5051 ( .A(n3496), .B(n3886), .Z(\w1[3][104] ) );
  XOR U5052 ( .A(\w3[2][106] ), .B(\w3[2][98] ), .Z(n3498) );
  XOR U5053 ( .A(\w3[2][97] ), .B(\w3[2][121] ), .Z(n3885) );
  XNOR U5054 ( .A(n3885), .B(key[489]), .Z(n3497) );
  XNOR U5055 ( .A(n3498), .B(n3497), .Z(n3499) );
  XOR U5056 ( .A(\w3[2][113] ), .B(n3499), .Z(\w1[3][105] ) );
  XOR U5057 ( .A(\w3[2][107] ), .B(\w3[2][99] ), .Z(n3501) );
  XOR U5058 ( .A(\w3[2][98] ), .B(\w3[2][122] ), .Z(n3890) );
  XNOR U5059 ( .A(n3890), .B(key[490]), .Z(n3500) );
  XNOR U5060 ( .A(n3501), .B(n3500), .Z(n3502) );
  XOR U5061 ( .A(\w3[2][114] ), .B(n3502), .Z(\w1[3][106] ) );
  XOR U5062 ( .A(\w3[2][99] ), .B(\w3[2][123] ), .Z(n3894) );
  XNOR U5063 ( .A(\w3[2][108] ), .B(n3894), .Z(n3503) );
  XNOR U5064 ( .A(\w3[2][104] ), .B(n3503), .Z(n3529) );
  XOR U5065 ( .A(n3529), .B(key[491]), .Z(n3505) );
  XOR U5066 ( .A(\w3[2][96] ), .B(\w3[2][100] ), .Z(n3898) );
  XNOR U5067 ( .A(\w3[2][115] ), .B(n3898), .Z(n3504) );
  XNOR U5068 ( .A(n3505), .B(n3504), .Z(\w1[3][107] ) );
  XOR U5069 ( .A(\w3[2][100] ), .B(\w3[2][104] ), .Z(n3507) );
  XNOR U5070 ( .A(\w3[2][124] ), .B(\w3[2][109] ), .Z(n3506) );
  XNOR U5071 ( .A(n3507), .B(n3506), .Z(n3532) );
  XOR U5072 ( .A(n3532), .B(key[492]), .Z(n3510) );
  XNOR U5073 ( .A(\w3[2][116] ), .B(n3508), .Z(n3509) );
  XNOR U5074 ( .A(n3510), .B(n3509), .Z(\w1[3][108] ) );
  XOR U5075 ( .A(\w3[2][125] ), .B(\w3[2][101] ), .Z(n3535) );
  XOR U5076 ( .A(n3535), .B(key[493]), .Z(n3512) );
  XNOR U5077 ( .A(\w3[2][102] ), .B(\w3[2][110] ), .Z(n3511) );
  XNOR U5078 ( .A(n3512), .B(n3511), .Z(n3513) );
  XOR U5079 ( .A(\w3[2][117] ), .B(n3513), .Z(\w1[3][109] ) );
  XOR U5080 ( .A(\w3[2][11] ), .B(\w3[2][3] ), .Z(n3515) );
  XOR U5081 ( .A(\w3[2][2] ), .B(\w3[2][26] ), .Z(n3599) );
  XNOR U5082 ( .A(n3599), .B(key[394]), .Z(n3514) );
  XNOR U5083 ( .A(n3515), .B(n3514), .Z(n3516) );
  XOR U5084 ( .A(\w3[2][18] ), .B(n3516), .Z(\w1[3][10] ) );
  XNOR U5085 ( .A(\w3[2][111] ), .B(\w3[2][104] ), .Z(n3544) );
  XNOR U5086 ( .A(n3517), .B(n3544), .Z(n3539) );
  XOR U5087 ( .A(n3539), .B(key[494]), .Z(n3520) );
  XNOR U5088 ( .A(\w3[2][118] ), .B(n3518), .Z(n3519) );
  XNOR U5089 ( .A(n3520), .B(n3519), .Z(\w1[3][110] ) );
  XOR U5090 ( .A(\w3[2][127] ), .B(\w3[2][103] ), .Z(n3542) );
  XOR U5091 ( .A(n3542), .B(key[495]), .Z(n3522) );
  XOR U5092 ( .A(\w3[2][96] ), .B(\w3[2][104] ), .Z(n3549) );
  XNOR U5093 ( .A(\w3[2][119] ), .B(n3549), .Z(n3521) );
  XNOR U5094 ( .A(n3522), .B(n3521), .Z(\w1[3][111] ) );
  XOR U5095 ( .A(\w3[2][105] ), .B(\w3[2][113] ), .Z(n3889) );
  XOR U5096 ( .A(n3889), .B(key[496]), .Z(n3524) );
  XNOR U5097 ( .A(\w3[2][120] ), .B(n3549), .Z(n3523) );
  XNOR U5098 ( .A(n3524), .B(n3523), .Z(\w1[3][112] ) );
  XOR U5099 ( .A(\w3[2][106] ), .B(\w3[2][114] ), .Z(n3893) );
  XOR U5100 ( .A(n3893), .B(key[497]), .Z(n3526) );
  XNOR U5101 ( .A(\w3[2][105] ), .B(n3885), .Z(n3525) );
  XNOR U5102 ( .A(n3526), .B(n3525), .Z(\w1[3][113] ) );
  XOR U5103 ( .A(\w3[2][107] ), .B(\w3[2][115] ), .Z(n3560) );
  XOR U5104 ( .A(n3560), .B(key[498]), .Z(n3528) );
  XNOR U5105 ( .A(\w3[2][106] ), .B(n3890), .Z(n3527) );
  XNOR U5106 ( .A(n3528), .B(n3527), .Z(\w1[3][114] ) );
  XOR U5107 ( .A(\w3[2][116] ), .B(\w3[2][112] ), .Z(n3561) );
  XOR U5108 ( .A(n3561), .B(key[499]), .Z(n3531) );
  XNOR U5109 ( .A(\w3[2][107] ), .B(n3529), .Z(n3530) );
  XNOR U5110 ( .A(n3531), .B(n3530), .Z(\w1[3][115] ) );
  XOR U5111 ( .A(\w3[2][117] ), .B(\w3[2][112] ), .Z(n3564) );
  XOR U5112 ( .A(n3564), .B(key[500]), .Z(n3534) );
  XNOR U5113 ( .A(\w3[2][108] ), .B(n3532), .Z(n3533) );
  XNOR U5114 ( .A(n3534), .B(n3533), .Z(\w1[3][116] ) );
  XOR U5115 ( .A(n3535), .B(key[501]), .Z(n3538) );
  XNOR U5116 ( .A(\w3[2][109] ), .B(n3536), .Z(n3537) );
  XNOR U5117 ( .A(n3538), .B(n3537), .Z(\w1[3][117] ) );
  XOR U5118 ( .A(\w3[2][119] ), .B(\w3[2][112] ), .Z(n3572) );
  XOR U5119 ( .A(n3572), .B(key[502]), .Z(n3541) );
  XNOR U5120 ( .A(\w3[2][110] ), .B(n3539), .Z(n3540) );
  XNOR U5121 ( .A(n3541), .B(n3540), .Z(\w1[3][118] ) );
  XNOR U5122 ( .A(n3542), .B(key[503]), .Z(n3543) );
  XNOR U5123 ( .A(n3544), .B(n3543), .Z(n3545) );
  XNOR U5124 ( .A(\w3[2][112] ), .B(n3545), .Z(\w1[3][119] ) );
  XOR U5125 ( .A(\w3[2][3] ), .B(\w3[2][27] ), .Z(n3640) );
  XNOR U5126 ( .A(\w3[2][8] ), .B(\w3[2][12] ), .Z(n3546) );
  XNOR U5127 ( .A(n3640), .B(n3546), .Z(n3596) );
  XOR U5128 ( .A(n3596), .B(key[395]), .Z(n3548) );
  XOR U5129 ( .A(\w3[2][0] ), .B(\w3[2][4] ), .Z(n3670) );
  XNOR U5130 ( .A(\w3[2][19] ), .B(n3670), .Z(n3547) );
  XNOR U5131 ( .A(n3548), .B(n3547), .Z(\w1[3][11] ) );
  XOR U5132 ( .A(n3549), .B(key[504]), .Z(n3551) );
  XNOR U5133 ( .A(\w3[2][113] ), .B(\w3[2][121] ), .Z(n3550) );
  XNOR U5134 ( .A(n3551), .B(n3550), .Z(n3552) );
  XOR U5135 ( .A(\w3[2][112] ), .B(n3552), .Z(\w1[3][120] ) );
  XOR U5136 ( .A(n3889), .B(key[505]), .Z(n3554) );
  XNOR U5137 ( .A(\w3[2][114] ), .B(\w3[2][122] ), .Z(n3553) );
  XNOR U5138 ( .A(n3554), .B(n3553), .Z(n3555) );
  XOR U5139 ( .A(\w3[2][97] ), .B(n3555), .Z(\w1[3][121] ) );
  XOR U5140 ( .A(n3893), .B(key[506]), .Z(n3557) );
  XNOR U5141 ( .A(\w3[2][115] ), .B(\w3[2][123] ), .Z(n3556) );
  XNOR U5142 ( .A(n3557), .B(n3556), .Z(n3558) );
  XOR U5143 ( .A(\w3[2][98] ), .B(n3558), .Z(\w1[3][122] ) );
  XNOR U5144 ( .A(\w3[2][124] ), .B(\w3[2][120] ), .Z(n3559) );
  XNOR U5145 ( .A(n3560), .B(n3559), .Z(n3897) );
  XOR U5146 ( .A(n3897), .B(key[507]), .Z(n3563) );
  XNOR U5147 ( .A(\w3[2][99] ), .B(n3561), .Z(n3562) );
  XNOR U5148 ( .A(n3563), .B(n3562), .Z(\w1[3][123] ) );
  XOR U5149 ( .A(n3564), .B(key[508]), .Z(n3567) );
  XNOR U5150 ( .A(n3565), .B(\w3[2][100] ), .Z(n3566) );
  XNOR U5151 ( .A(n3567), .B(n3566), .Z(\w1[3][124] ) );
  XOR U5152 ( .A(\w3[2][118] ), .B(key[509]), .Z(n3570) );
  XNOR U5153 ( .A(n3568), .B(\w3[2][126] ), .Z(n3569) );
  XNOR U5154 ( .A(n3570), .B(n3569), .Z(n3571) );
  XOR U5155 ( .A(\w3[2][101] ), .B(n3571), .Z(\w1[3][125] ) );
  XOR U5156 ( .A(n3572), .B(key[510]), .Z(n3575) );
  XNOR U5157 ( .A(\w3[2][102] ), .B(n3573), .Z(n3574) );
  XNOR U5158 ( .A(n3575), .B(n3574), .Z(\w1[3][126] ) );
  XNOR U5159 ( .A(n3576), .B(key[511]), .Z(n3577) );
  XNOR U5160 ( .A(n3886), .B(n3577), .Z(n3578) );
  XNOR U5161 ( .A(\w3[2][103] ), .B(n3578), .Z(\w1[3][127] ) );
  XOR U5162 ( .A(\w3[2][13] ), .B(\w3[2][28] ), .Z(n3580) );
  XNOR U5163 ( .A(\w3[2][8] ), .B(\w3[2][4] ), .Z(n3579) );
  XNOR U5164 ( .A(n3580), .B(n3579), .Z(n3602) );
  XOR U5165 ( .A(n3602), .B(key[396]), .Z(n3582) );
  XOR U5166 ( .A(\w3[2][0] ), .B(\w3[2][5] ), .Z(n3707) );
  XNOR U5167 ( .A(\w3[2][20] ), .B(n3707), .Z(n3581) );
  XNOR U5168 ( .A(n3582), .B(n3581), .Z(\w1[3][12] ) );
  XOR U5169 ( .A(\w3[2][14] ), .B(\w3[2][6] ), .Z(n3584) );
  XOR U5170 ( .A(\w3[2][5] ), .B(\w3[2][29] ), .Z(n3605) );
  XNOR U5171 ( .A(n3605), .B(key[397]), .Z(n3583) );
  XNOR U5172 ( .A(n3584), .B(n3583), .Z(n3585) );
  XOR U5173 ( .A(\w3[2][21] ), .B(n3585), .Z(\w1[3][13] ) );
  XOR U5174 ( .A(\w3[2][6] ), .B(\w3[2][30] ), .Z(n3748) );
  XNOR U5175 ( .A(\w3[2][8] ), .B(\w3[2][15] ), .Z(n3613) );
  XNOR U5176 ( .A(n3748), .B(n3613), .Z(n3608) );
  XOR U5177 ( .A(n3608), .B(key[398]), .Z(n3587) );
  XOR U5178 ( .A(\w3[2][0] ), .B(\w3[2][7] ), .Z(n3783) );
  XNOR U5179 ( .A(\w3[2][22] ), .B(n3783), .Z(n3586) );
  XNOR U5180 ( .A(n3587), .B(n3586), .Z(\w1[3][14] ) );
  XOR U5181 ( .A(\w3[2][7] ), .B(\w3[2][31] ), .Z(n3611) );
  XOR U5182 ( .A(n3611), .B(key[399]), .Z(n3589) );
  XOR U5183 ( .A(\w3[2][8] ), .B(\w3[2][0] ), .Z(n3615) );
  XNOR U5184 ( .A(\w3[2][23] ), .B(n3615), .Z(n3588) );
  XNOR U5185 ( .A(n3589), .B(n3588), .Z(\w1[3][15] ) );
  XOR U5186 ( .A(\w3[2][17] ), .B(\w3[2][9] ), .Z(n3619) );
  XOR U5187 ( .A(n3619), .B(key[400]), .Z(n3591) );
  XNOR U5188 ( .A(\w3[2][24] ), .B(n3615), .Z(n3590) );
  XNOR U5189 ( .A(n3591), .B(n3590), .Z(\w1[3][16] ) );
  XOR U5190 ( .A(\w3[2][18] ), .B(\w3[2][10] ), .Z(n3639) );
  XOR U5191 ( .A(n3639), .B(key[401]), .Z(n3593) );
  XNOR U5192 ( .A(n3904), .B(\w3[2][9] ), .Z(n3592) );
  XNOR U5193 ( .A(n3593), .B(n3592), .Z(\w1[3][17] ) );
  XOR U5194 ( .A(\w3[2][11] ), .B(\w3[2][19] ), .Z(n3627) );
  XOR U5195 ( .A(n3627), .B(key[402]), .Z(n3595) );
  XNOR U5196 ( .A(n3599), .B(\w3[2][10] ), .Z(n3594) );
  XNOR U5197 ( .A(n3595), .B(n3594), .Z(\w1[3][18] ) );
  XOR U5198 ( .A(\w3[2][16] ), .B(\w3[2][20] ), .Z(n3628) );
  XOR U5199 ( .A(n3628), .B(key[403]), .Z(n3598) );
  XNOR U5200 ( .A(\w3[2][11] ), .B(n3596), .Z(n3597) );
  XNOR U5201 ( .A(n3598), .B(n3597), .Z(\w1[3][19] ) );
  XOR U5202 ( .A(n3619), .B(key[385]), .Z(n3601) );
  XNOR U5203 ( .A(\w3[2][25] ), .B(n3599), .Z(n3600) );
  XNOR U5204 ( .A(n3601), .B(n3600), .Z(\w1[3][1] ) );
  XOR U5205 ( .A(\w3[2][16] ), .B(\w3[2][21] ), .Z(n3633) );
  XOR U5206 ( .A(n3633), .B(key[404]), .Z(n3604) );
  XNOR U5207 ( .A(\w3[2][12] ), .B(n3602), .Z(n3603) );
  XNOR U5208 ( .A(n3604), .B(n3603), .Z(\w1[3][20] ) );
  XOR U5209 ( .A(\w3[2][14] ), .B(\w3[2][22] ), .Z(n3643) );
  XOR U5210 ( .A(n3643), .B(key[405]), .Z(n3607) );
  XNOR U5211 ( .A(\w3[2][13] ), .B(n3605), .Z(n3606) );
  XNOR U5212 ( .A(n3607), .B(n3606), .Z(\w1[3][21] ) );
  XOR U5213 ( .A(\w3[2][16] ), .B(\w3[2][23] ), .Z(n3644) );
  XOR U5214 ( .A(n3644), .B(key[406]), .Z(n3610) );
  XNOR U5215 ( .A(\w3[2][14] ), .B(n3608), .Z(n3609) );
  XNOR U5216 ( .A(n3610), .B(n3609), .Z(\w1[3][22] ) );
  XNOR U5217 ( .A(n3611), .B(key[407]), .Z(n3612) );
  XNOR U5218 ( .A(n3613), .B(n3612), .Z(n3614) );
  XNOR U5219 ( .A(\w3[2][16] ), .B(n3614), .Z(\w1[3][23] ) );
  XOR U5220 ( .A(\w3[2][17] ), .B(key[408]), .Z(n3617) );
  XNOR U5221 ( .A(\w3[2][25] ), .B(n3615), .Z(n3616) );
  XNOR U5222 ( .A(n3617), .B(n3616), .Z(n3618) );
  XOR U5223 ( .A(\w3[2][16] ), .B(n3618), .Z(\w1[3][24] ) );
  XOR U5224 ( .A(n3619), .B(key[409]), .Z(n3621) );
  XNOR U5225 ( .A(\w3[2][1] ), .B(\w3[2][26] ), .Z(n3620) );
  XNOR U5226 ( .A(n3621), .B(n3620), .Z(n3622) );
  XOR U5227 ( .A(\w3[2][18] ), .B(n3622), .Z(\w1[3][25] ) );
  XOR U5228 ( .A(n3639), .B(key[410]), .Z(n3624) );
  XNOR U5229 ( .A(\w3[2][2] ), .B(\w3[2][19] ), .Z(n3623) );
  XNOR U5230 ( .A(n3624), .B(n3623), .Z(n3625) );
  XOR U5231 ( .A(\w3[2][27] ), .B(n3625), .Z(\w1[3][26] ) );
  XNOR U5232 ( .A(\w3[2][24] ), .B(\w3[2][28] ), .Z(n3626) );
  XNOR U5233 ( .A(n3627), .B(n3626), .Z(n3669) );
  XOR U5234 ( .A(n3669), .B(key[411]), .Z(n3630) );
  XNOR U5235 ( .A(\w3[2][3] ), .B(n3628), .Z(n3629) );
  XNOR U5236 ( .A(n3630), .B(n3629), .Z(\w1[3][27] ) );
  XOR U5237 ( .A(\w3[2][20] ), .B(\w3[2][29] ), .Z(n3632) );
  XNOR U5238 ( .A(\w3[2][24] ), .B(\w3[2][12] ), .Z(n3631) );
  XNOR U5239 ( .A(n3632), .B(n3631), .Z(n3706) );
  XOR U5240 ( .A(n3706), .B(key[412]), .Z(n3635) );
  XNOR U5241 ( .A(\w3[2][4] ), .B(n3633), .Z(n3634) );
  XNOR U5242 ( .A(n3635), .B(n3634), .Z(\w1[3][28] ) );
  XOR U5243 ( .A(\w3[2][13] ), .B(\w3[2][21] ), .Z(n3747) );
  XOR U5244 ( .A(n3747), .B(key[413]), .Z(n3637) );
  XNOR U5245 ( .A(\w3[2][22] ), .B(\w3[2][30] ), .Z(n3636) );
  XNOR U5246 ( .A(n3637), .B(n3636), .Z(n3638) );
  XOR U5247 ( .A(\w3[2][5] ), .B(n3638), .Z(\w1[3][29] ) );
  XOR U5248 ( .A(n3639), .B(key[386]), .Z(n3642) );
  XNOR U5249 ( .A(\w3[2][26] ), .B(n3640), .Z(n3641) );
  XNOR U5250 ( .A(n3642), .B(n3641), .Z(\w1[3][2] ) );
  XNOR U5251 ( .A(\w3[2][24] ), .B(\w3[2][31] ), .Z(n3821) );
  XNOR U5252 ( .A(n3643), .B(n3821), .Z(n3782) );
  XOR U5253 ( .A(n3782), .B(key[414]), .Z(n3646) );
  XNOR U5254 ( .A(\w3[2][6] ), .B(n3644), .Z(n3645) );
  XNOR U5255 ( .A(n3646), .B(n3645), .Z(\w1[3][30] ) );
  XOR U5256 ( .A(\w3[2][15] ), .B(\w3[2][23] ), .Z(n3819) );
  XOR U5257 ( .A(n3819), .B(key[415]), .Z(n3648) );
  XNOR U5258 ( .A(n3860), .B(\w3[2][7] ), .Z(n3647) );
  XNOR U5259 ( .A(n3648), .B(n3647), .Z(\w1[3][31] ) );
  XOR U5260 ( .A(\w3[2][33] ), .B(\w3[2][57] ), .Z(n3703) );
  XOR U5261 ( .A(n3703), .B(key[416]), .Z(n3650) );
  XOR U5262 ( .A(\w3[2][48] ), .B(\w3[2][56] ), .Z(n3764) );
  XNOR U5263 ( .A(n3764), .B(\w3[2][40] ), .Z(n3649) );
  XNOR U5264 ( .A(n3650), .B(n3649), .Z(\w1[3][32] ) );
  XOR U5265 ( .A(\w3[2][34] ), .B(\w3[2][58] ), .Z(n3711) );
  XOR U5266 ( .A(n3711), .B(key[417]), .Z(n3652) );
  XOR U5267 ( .A(\w3[2][41] ), .B(\w3[2][49] ), .Z(n3735) );
  XNOR U5268 ( .A(\w3[2][57] ), .B(n3735), .Z(n3651) );
  XNOR U5269 ( .A(n3652), .B(n3651), .Z(\w1[3][33] ) );
  XOR U5270 ( .A(\w3[2][35] ), .B(\w3[2][59] ), .Z(n3682) );
  XOR U5271 ( .A(n3682), .B(key[418]), .Z(n3654) );
  XOR U5272 ( .A(\w3[2][42] ), .B(\w3[2][50] ), .Z(n3739) );
  XNOR U5273 ( .A(\w3[2][58] ), .B(n3739), .Z(n3653) );
  XNOR U5274 ( .A(n3654), .B(n3653), .Z(\w1[3][34] ) );
  XOR U5275 ( .A(\w3[2][36] ), .B(\w3[2][32] ), .Z(n3684) );
  XOR U5276 ( .A(n3684), .B(key[419]), .Z(n3657) );
  XOR U5277 ( .A(\w3[2][43] ), .B(\w3[2][51] ), .Z(n3710) );
  XNOR U5278 ( .A(\w3[2][56] ), .B(n3710), .Z(n3655) );
  XNOR U5279 ( .A(\w3[2][60] ), .B(n3655), .Z(n3744) );
  XNOR U5280 ( .A(\w3[2][59] ), .B(n3744), .Z(n3656) );
  XNOR U5281 ( .A(n3657), .B(n3656), .Z(\w1[3][35] ) );
  XOR U5282 ( .A(\w3[2][32] ), .B(\w3[2][37] ), .Z(n3689) );
  XOR U5283 ( .A(n3689), .B(key[420]), .Z(n3661) );
  XOR U5284 ( .A(\w3[2][52] ), .B(\w3[2][61] ), .Z(n3659) );
  XNOR U5285 ( .A(\w3[2][56] ), .B(\w3[2][44] ), .Z(n3658) );
  XNOR U5286 ( .A(n3659), .B(n3658), .Z(n3752) );
  XNOR U5287 ( .A(\w3[2][60] ), .B(n3752), .Z(n3660) );
  XNOR U5288 ( .A(n3661), .B(n3660), .Z(\w1[3][36] ) );
  XOR U5289 ( .A(\w3[2][38] ), .B(\w3[2][62] ), .Z(n3695) );
  XOR U5290 ( .A(n3695), .B(key[421]), .Z(n3663) );
  XOR U5291 ( .A(\w3[2][45] ), .B(\w3[2][53] ), .Z(n3755) );
  XNOR U5292 ( .A(\w3[2][61] ), .B(n3755), .Z(n3662) );
  XNOR U5293 ( .A(n3663), .B(n3662), .Z(\w1[3][37] ) );
  XOR U5294 ( .A(\w3[2][32] ), .B(\w3[2][39] ), .Z(n3696) );
  XOR U5295 ( .A(n3696), .B(key[422]), .Z(n3665) );
  XOR U5296 ( .A(\w3[2][46] ), .B(\w3[2][54] ), .Z(n3721) );
  XNOR U5297 ( .A(\w3[2][56] ), .B(\w3[2][63] ), .Z(n3667) );
  XNOR U5298 ( .A(n3721), .B(n3667), .Z(n3760) );
  XNOR U5299 ( .A(\w3[2][62] ), .B(n3760), .Z(n3664) );
  XNOR U5300 ( .A(n3665), .B(n3664), .Z(\w1[3][38] ) );
  XOR U5301 ( .A(\w3[2][47] ), .B(\w3[2][55] ), .Z(n3763) );
  XNOR U5302 ( .A(n3763), .B(key[423]), .Z(n3666) );
  XNOR U5303 ( .A(n3667), .B(n3666), .Z(n3668) );
  XNOR U5304 ( .A(\w3[2][32] ), .B(n3668), .Z(\w1[3][39] ) );
  XOR U5305 ( .A(n3669), .B(key[387]), .Z(n3672) );
  XNOR U5306 ( .A(n3670), .B(\w3[2][27] ), .Z(n3671) );
  XNOR U5307 ( .A(n3672), .B(n3671), .Z(\w1[3][3] ) );
  XOR U5308 ( .A(\w3[2][32] ), .B(key[424]), .Z(n3674) );
  XNOR U5309 ( .A(\w3[2][33] ), .B(\w3[2][41] ), .Z(n3673) );
  XNOR U5310 ( .A(n3674), .B(n3673), .Z(n3675) );
  XOR U5311 ( .A(n3764), .B(n3675), .Z(\w1[3][40] ) );
  XOR U5312 ( .A(\w3[2][42] ), .B(key[425]), .Z(n3677) );
  XNOR U5313 ( .A(\w3[2][49] ), .B(\w3[2][34] ), .Z(n3676) );
  XNOR U5314 ( .A(n3677), .B(n3676), .Z(n3678) );
  XOR U5315 ( .A(n3703), .B(n3678), .Z(\w1[3][41] ) );
  XOR U5316 ( .A(\w3[2][43] ), .B(key[426]), .Z(n3680) );
  XNOR U5317 ( .A(\w3[2][50] ), .B(\w3[2][35] ), .Z(n3679) );
  XNOR U5318 ( .A(n3680), .B(n3679), .Z(n3681) );
  XOR U5319 ( .A(n3711), .B(n3681), .Z(\w1[3][42] ) );
  XNOR U5320 ( .A(\w3[2][40] ), .B(n3682), .Z(n3683) );
  XNOR U5321 ( .A(\w3[2][44] ), .B(n3683), .Z(n3714) );
  XOR U5322 ( .A(n3714), .B(key[427]), .Z(n3686) );
  XNOR U5323 ( .A(\w3[2][51] ), .B(n3684), .Z(n3685) );
  XNOR U5324 ( .A(n3686), .B(n3685), .Z(\w1[3][43] ) );
  XOR U5325 ( .A(\w3[2][36] ), .B(\w3[2][45] ), .Z(n3688) );
  XNOR U5326 ( .A(\w3[2][40] ), .B(\w3[2][60] ), .Z(n3687) );
  XNOR U5327 ( .A(n3688), .B(n3687), .Z(n3717) );
  XOR U5328 ( .A(n3717), .B(key[428]), .Z(n3691) );
  XNOR U5329 ( .A(\w3[2][52] ), .B(n3689), .Z(n3690) );
  XNOR U5330 ( .A(n3691), .B(n3690), .Z(\w1[3][44] ) );
  XOR U5331 ( .A(\w3[2][61] ), .B(\w3[2][37] ), .Z(n3720) );
  XOR U5332 ( .A(n3720), .B(key[429]), .Z(n3693) );
  XNOR U5333 ( .A(\w3[2][38] ), .B(\w3[2][46] ), .Z(n3692) );
  XNOR U5334 ( .A(n3693), .B(n3692), .Z(n3694) );
  XOR U5335 ( .A(\w3[2][53] ), .B(n3694), .Z(\w1[3][45] ) );
  XNOR U5336 ( .A(\w3[2][40] ), .B(\w3[2][47] ), .Z(n3729) );
  XNOR U5337 ( .A(n3695), .B(n3729), .Z(n3724) );
  XOR U5338 ( .A(n3724), .B(key[430]), .Z(n3698) );
  XNOR U5339 ( .A(\w3[2][54] ), .B(n3696), .Z(n3697) );
  XNOR U5340 ( .A(n3698), .B(n3697), .Z(\w1[3][46] ) );
  XOR U5341 ( .A(\w3[2][63] ), .B(\w3[2][39] ), .Z(n3727) );
  XOR U5342 ( .A(n3727), .B(key[431]), .Z(n3700) );
  XOR U5343 ( .A(\w3[2][40] ), .B(\w3[2][32] ), .Z(n3731) );
  XNOR U5344 ( .A(\w3[2][55] ), .B(n3731), .Z(n3699) );
  XNOR U5345 ( .A(n3700), .B(n3699), .Z(\w1[3][47] ) );
  XOR U5346 ( .A(n3731), .B(key[432]), .Z(n3702) );
  XNOR U5347 ( .A(\w3[2][56] ), .B(n3735), .Z(n3701) );
  XNOR U5348 ( .A(n3702), .B(n3701), .Z(\w1[3][48] ) );
  XOR U5349 ( .A(n3739), .B(key[433]), .Z(n3705) );
  XNOR U5350 ( .A(n3703), .B(\w3[2][41] ), .Z(n3704) );
  XNOR U5351 ( .A(n3705), .B(n3704), .Z(\w1[3][49] ) );
  XOR U5352 ( .A(n3706), .B(key[388]), .Z(n3709) );
  XNOR U5353 ( .A(n3707), .B(\w3[2][28] ), .Z(n3708) );
  XNOR U5354 ( .A(n3709), .B(n3708), .Z(\w1[3][4] ) );
  XOR U5355 ( .A(n3710), .B(key[434]), .Z(n3713) );
  XNOR U5356 ( .A(n3711), .B(\w3[2][42] ), .Z(n3712) );
  XNOR U5357 ( .A(n3713), .B(n3712), .Z(\w1[3][50] ) );
  XOR U5358 ( .A(\w3[2][48] ), .B(\w3[2][52] ), .Z(n3743) );
  XOR U5359 ( .A(n3743), .B(key[435]), .Z(n3716) );
  XNOR U5360 ( .A(\w3[2][43] ), .B(n3714), .Z(n3715) );
  XNOR U5361 ( .A(n3716), .B(n3715), .Z(\w1[3][51] ) );
  XOR U5362 ( .A(\w3[2][48] ), .B(\w3[2][53] ), .Z(n3751) );
  XOR U5363 ( .A(n3751), .B(key[436]), .Z(n3719) );
  XNOR U5364 ( .A(\w3[2][44] ), .B(n3717), .Z(n3718) );
  XNOR U5365 ( .A(n3719), .B(n3718), .Z(\w1[3][52] ) );
  XOR U5366 ( .A(n3720), .B(key[437]), .Z(n3723) );
  XNOR U5367 ( .A(\w3[2][45] ), .B(n3721), .Z(n3722) );
  XNOR U5368 ( .A(n3723), .B(n3722), .Z(\w1[3][53] ) );
  XOR U5369 ( .A(\w3[2][48] ), .B(\w3[2][55] ), .Z(n3759) );
  XOR U5370 ( .A(n3759), .B(key[438]), .Z(n3726) );
  XNOR U5371 ( .A(\w3[2][46] ), .B(n3724), .Z(n3725) );
  XNOR U5372 ( .A(n3726), .B(n3725), .Z(\w1[3][54] ) );
  XNOR U5373 ( .A(n3727), .B(key[439]), .Z(n3728) );
  XNOR U5374 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U5375 ( .A(\w3[2][48] ), .B(n3730), .Z(\w1[3][55] ) );
  XOR U5376 ( .A(n3731), .B(key[440]), .Z(n3733) );
  XNOR U5377 ( .A(\w3[2][48] ), .B(\w3[2][49] ), .Z(n3732) );
  XNOR U5378 ( .A(n3733), .B(n3732), .Z(n3734) );
  XOR U5379 ( .A(\w3[2][57] ), .B(n3734), .Z(\w1[3][56] ) );
  XOR U5380 ( .A(\w3[2][50] ), .B(key[441]), .Z(n3737) );
  XNOR U5381 ( .A(n3735), .B(\w3[2][58] ), .Z(n3736) );
  XNOR U5382 ( .A(n3737), .B(n3736), .Z(n3738) );
  XOR U5383 ( .A(\w3[2][33] ), .B(n3738), .Z(\w1[3][57] ) );
  XOR U5384 ( .A(\w3[2][51] ), .B(key[442]), .Z(n3741) );
  XNOR U5385 ( .A(n3739), .B(\w3[2][59] ), .Z(n3740) );
  XNOR U5386 ( .A(n3741), .B(n3740), .Z(n3742) );
  XOR U5387 ( .A(\w3[2][34] ), .B(n3742), .Z(\w1[3][58] ) );
  XOR U5388 ( .A(n3743), .B(key[443]), .Z(n3746) );
  XNOR U5389 ( .A(\w3[2][35] ), .B(n3744), .Z(n3745) );
  XNOR U5390 ( .A(n3746), .B(n3745), .Z(\w1[3][59] ) );
  XOR U5391 ( .A(n3747), .B(key[389]), .Z(n3750) );
  XNOR U5392 ( .A(\w3[2][29] ), .B(n3748), .Z(n3749) );
  XNOR U5393 ( .A(n3750), .B(n3749), .Z(\w1[3][5] ) );
  XOR U5394 ( .A(n3751), .B(key[444]), .Z(n3754) );
  XNOR U5395 ( .A(\w3[2][36] ), .B(n3752), .Z(n3753) );
  XNOR U5396 ( .A(n3754), .B(n3753), .Z(\w1[3][60] ) );
  XOR U5397 ( .A(\w3[2][54] ), .B(key[445]), .Z(n3757) );
  XNOR U5398 ( .A(n3755), .B(\w3[2][62] ), .Z(n3756) );
  XNOR U5399 ( .A(n3757), .B(n3756), .Z(n3758) );
  XOR U5400 ( .A(\w3[2][37] ), .B(n3758), .Z(\w1[3][61] ) );
  XOR U5401 ( .A(n3759), .B(key[446]), .Z(n3762) );
  XNOR U5402 ( .A(\w3[2][38] ), .B(n3760), .Z(n3761) );
  XNOR U5403 ( .A(n3762), .B(n3761), .Z(\w1[3][62] ) );
  XOR U5404 ( .A(n3763), .B(key[447]), .Z(n3766) );
  XNOR U5405 ( .A(n3764), .B(\w3[2][39] ), .Z(n3765) );
  XNOR U5406 ( .A(n3766), .B(n3765), .Z(\w1[3][63] ) );
  XOR U5407 ( .A(\w3[2][65] ), .B(\w3[2][89] ), .Z(n3825) );
  XOR U5408 ( .A(n3825), .B(key[448]), .Z(n3768) );
  XOR U5409 ( .A(\w3[2][80] ), .B(\w3[2][88] ), .Z(n3882) );
  XNOR U5410 ( .A(n3882), .B(\w3[2][72] ), .Z(n3767) );
  XNOR U5411 ( .A(n3768), .B(n3767), .Z(\w1[3][64] ) );
  XOR U5412 ( .A(\w3[2][66] ), .B(\w3[2][90] ), .Z(n3829) );
  XOR U5413 ( .A(n3829), .B(key[449]), .Z(n3770) );
  XOR U5414 ( .A(\w3[2][73] ), .B(\w3[2][81] ), .Z(n3853) );
  XNOR U5415 ( .A(\w3[2][89] ), .B(n3853), .Z(n3769) );
  XNOR U5416 ( .A(n3770), .B(n3769), .Z(\w1[3][65] ) );
  XOR U5417 ( .A(\w3[2][67] ), .B(\w3[2][91] ), .Z(n3800) );
  XOR U5418 ( .A(n3800), .B(key[450]), .Z(n3772) );
  XOR U5419 ( .A(\w3[2][74] ), .B(\w3[2][82] ), .Z(n3861) );
  XNOR U5420 ( .A(\w3[2][90] ), .B(n3861), .Z(n3771) );
  XNOR U5421 ( .A(n3772), .B(n3771), .Z(\w1[3][66] ) );
  XOR U5422 ( .A(\w3[2][68] ), .B(\w3[2][64] ), .Z(n3802) );
  XOR U5423 ( .A(n3802), .B(key[451]), .Z(n3775) );
  XOR U5424 ( .A(\w3[2][75] ), .B(\w3[2][83] ), .Z(n3828) );
  XNOR U5425 ( .A(\w3[2][88] ), .B(n3828), .Z(n3773) );
  XNOR U5426 ( .A(\w3[2][92] ), .B(n3773), .Z(n3866) );
  XNOR U5427 ( .A(\w3[2][91] ), .B(n3866), .Z(n3774) );
  XNOR U5428 ( .A(n3775), .B(n3774), .Z(\w1[3][67] ) );
  XOR U5429 ( .A(\w3[2][64] ), .B(\w3[2][69] ), .Z(n3807) );
  XOR U5430 ( .A(n3807), .B(key[452]), .Z(n3779) );
  XOR U5431 ( .A(\w3[2][84] ), .B(\w3[2][93] ), .Z(n3777) );
  XNOR U5432 ( .A(\w3[2][88] ), .B(\w3[2][76] ), .Z(n3776) );
  XNOR U5433 ( .A(n3777), .B(n3776), .Z(n3870) );
  XNOR U5434 ( .A(\w3[2][92] ), .B(n3870), .Z(n3778) );
  XNOR U5435 ( .A(n3779), .B(n3778), .Z(\w1[3][68] ) );
  XOR U5436 ( .A(\w3[2][70] ), .B(\w3[2][94] ), .Z(n3813) );
  XOR U5437 ( .A(n3813), .B(key[453]), .Z(n3781) );
  XOR U5438 ( .A(\w3[2][77] ), .B(\w3[2][85] ), .Z(n3873) );
  XNOR U5439 ( .A(\w3[2][93] ), .B(n3873), .Z(n3780) );
  XNOR U5440 ( .A(n3781), .B(n3780), .Z(\w1[3][69] ) );
  XOR U5441 ( .A(n3782), .B(key[390]), .Z(n3785) );
  XNOR U5442 ( .A(n3783), .B(\w3[2][30] ), .Z(n3784) );
  XNOR U5443 ( .A(n3785), .B(n3784), .Z(\w1[3][6] ) );
  XOR U5444 ( .A(\w3[2][64] ), .B(\w3[2][71] ), .Z(n3814) );
  XOR U5445 ( .A(n3814), .B(key[454]), .Z(n3787) );
  XOR U5446 ( .A(\w3[2][78] ), .B(\w3[2][86] ), .Z(n3839) );
  XNOR U5447 ( .A(\w3[2][88] ), .B(\w3[2][95] ), .Z(n3789) );
  XNOR U5448 ( .A(n3839), .B(n3789), .Z(n3878) );
  XNOR U5449 ( .A(\w3[2][94] ), .B(n3878), .Z(n3786) );
  XNOR U5450 ( .A(n3787), .B(n3786), .Z(\w1[3][70] ) );
  XOR U5451 ( .A(\w3[2][79] ), .B(\w3[2][87] ), .Z(n3881) );
  XNOR U5452 ( .A(n3881), .B(key[455]), .Z(n3788) );
  XNOR U5453 ( .A(n3789), .B(n3788), .Z(n3790) );
  XNOR U5454 ( .A(\w3[2][64] ), .B(n3790), .Z(\w1[3][71] ) );
  XOR U5455 ( .A(\w3[2][64] ), .B(key[456]), .Z(n3792) );
  XNOR U5456 ( .A(\w3[2][65] ), .B(\w3[2][73] ), .Z(n3791) );
  XNOR U5457 ( .A(n3792), .B(n3791), .Z(n3793) );
  XOR U5458 ( .A(n3882), .B(n3793), .Z(\w1[3][72] ) );
  XOR U5459 ( .A(\w3[2][74] ), .B(key[457]), .Z(n3795) );
  XNOR U5460 ( .A(\w3[2][81] ), .B(\w3[2][66] ), .Z(n3794) );
  XNOR U5461 ( .A(n3795), .B(n3794), .Z(n3796) );
  XOR U5462 ( .A(n3825), .B(n3796), .Z(\w1[3][73] ) );
  XOR U5463 ( .A(\w3[2][75] ), .B(key[458]), .Z(n3798) );
  XNOR U5464 ( .A(\w3[2][82] ), .B(\w3[2][67] ), .Z(n3797) );
  XNOR U5465 ( .A(n3798), .B(n3797), .Z(n3799) );
  XOR U5466 ( .A(n3829), .B(n3799), .Z(\w1[3][74] ) );
  XNOR U5467 ( .A(\w3[2][72] ), .B(n3800), .Z(n3801) );
  XNOR U5468 ( .A(\w3[2][76] ), .B(n3801), .Z(n3832) );
  XOR U5469 ( .A(n3832), .B(key[459]), .Z(n3804) );
  XNOR U5470 ( .A(\w3[2][83] ), .B(n3802), .Z(n3803) );
  XNOR U5471 ( .A(n3804), .B(n3803), .Z(\w1[3][75] ) );
  XOR U5472 ( .A(\w3[2][68] ), .B(\w3[2][77] ), .Z(n3806) );
  XNOR U5473 ( .A(\w3[2][72] ), .B(\w3[2][92] ), .Z(n3805) );
  XNOR U5474 ( .A(n3806), .B(n3805), .Z(n3835) );
  XOR U5475 ( .A(n3835), .B(key[460]), .Z(n3809) );
  XNOR U5476 ( .A(\w3[2][84] ), .B(n3807), .Z(n3808) );
  XNOR U5477 ( .A(n3809), .B(n3808), .Z(\w1[3][76] ) );
  XOR U5478 ( .A(\w3[2][93] ), .B(\w3[2][69] ), .Z(n3838) );
  XOR U5479 ( .A(n3838), .B(key[461]), .Z(n3811) );
  XNOR U5480 ( .A(\w3[2][70] ), .B(\w3[2][78] ), .Z(n3810) );
  XNOR U5481 ( .A(n3811), .B(n3810), .Z(n3812) );
  XOR U5482 ( .A(\w3[2][85] ), .B(n3812), .Z(\w1[3][77] ) );
  XNOR U5483 ( .A(\w3[2][72] ), .B(\w3[2][79] ), .Z(n3847) );
  XNOR U5484 ( .A(n3813), .B(n3847), .Z(n3842) );
  XOR U5485 ( .A(n3842), .B(key[462]), .Z(n3816) );
  XNOR U5486 ( .A(\w3[2][86] ), .B(n3814), .Z(n3815) );
  XNOR U5487 ( .A(n3816), .B(n3815), .Z(\w1[3][78] ) );
  XOR U5488 ( .A(\w3[2][95] ), .B(\w3[2][71] ), .Z(n3845) );
  XOR U5489 ( .A(n3845), .B(key[463]), .Z(n3818) );
  XOR U5490 ( .A(\w3[2][72] ), .B(\w3[2][64] ), .Z(n3849) );
  XNOR U5491 ( .A(\w3[2][87] ), .B(n3849), .Z(n3817) );
  XNOR U5492 ( .A(n3818), .B(n3817), .Z(\w1[3][79] ) );
  XNOR U5493 ( .A(n3819), .B(key[391]), .Z(n3820) );
  XNOR U5494 ( .A(n3821), .B(n3820), .Z(n3822) );
  XNOR U5495 ( .A(\w3[2][0] ), .B(n3822), .Z(\w1[3][7] ) );
  XOR U5496 ( .A(n3849), .B(key[464]), .Z(n3824) );
  XNOR U5497 ( .A(\w3[2][88] ), .B(n3853), .Z(n3823) );
  XNOR U5498 ( .A(n3824), .B(n3823), .Z(\w1[3][80] ) );
  XOR U5499 ( .A(n3861), .B(key[465]), .Z(n3827) );
  XNOR U5500 ( .A(n3825), .B(\w3[2][73] ), .Z(n3826) );
  XNOR U5501 ( .A(n3827), .B(n3826), .Z(\w1[3][81] ) );
  XOR U5502 ( .A(n3828), .B(key[466]), .Z(n3831) );
  XNOR U5503 ( .A(n3829), .B(\w3[2][74] ), .Z(n3830) );
  XNOR U5504 ( .A(n3831), .B(n3830), .Z(\w1[3][82] ) );
  XOR U5505 ( .A(\w3[2][80] ), .B(\w3[2][84] ), .Z(n3865) );
  XOR U5506 ( .A(n3865), .B(key[467]), .Z(n3834) );
  XNOR U5507 ( .A(\w3[2][75] ), .B(n3832), .Z(n3833) );
  XNOR U5508 ( .A(n3834), .B(n3833), .Z(\w1[3][83] ) );
  XOR U5509 ( .A(\w3[2][80] ), .B(\w3[2][85] ), .Z(n3869) );
  XOR U5510 ( .A(n3869), .B(key[468]), .Z(n3837) );
  XNOR U5511 ( .A(\w3[2][76] ), .B(n3835), .Z(n3836) );
  XNOR U5512 ( .A(n3837), .B(n3836), .Z(\w1[3][84] ) );
  XOR U5513 ( .A(n3838), .B(key[469]), .Z(n3841) );
  XNOR U5514 ( .A(\w3[2][77] ), .B(n3839), .Z(n3840) );
  XNOR U5515 ( .A(n3841), .B(n3840), .Z(\w1[3][85] ) );
  XOR U5516 ( .A(\w3[2][80] ), .B(\w3[2][87] ), .Z(n3877) );
  XOR U5517 ( .A(n3877), .B(key[470]), .Z(n3844) );
  XNOR U5518 ( .A(\w3[2][78] ), .B(n3842), .Z(n3843) );
  XNOR U5519 ( .A(n3844), .B(n3843), .Z(\w1[3][86] ) );
  XNOR U5520 ( .A(n3845), .B(key[471]), .Z(n3846) );
  XNOR U5521 ( .A(n3847), .B(n3846), .Z(n3848) );
  XNOR U5522 ( .A(\w3[2][80] ), .B(n3848), .Z(\w1[3][87] ) );
  XOR U5523 ( .A(n3849), .B(key[472]), .Z(n3851) );
  XNOR U5524 ( .A(\w3[2][80] ), .B(\w3[2][81] ), .Z(n3850) );
  XNOR U5525 ( .A(n3851), .B(n3850), .Z(n3852) );
  XOR U5526 ( .A(\w3[2][89] ), .B(n3852), .Z(\w1[3][88] ) );
  XOR U5527 ( .A(\w3[2][82] ), .B(key[473]), .Z(n3855) );
  XNOR U5528 ( .A(n3853), .B(\w3[2][90] ), .Z(n3854) );
  XNOR U5529 ( .A(n3855), .B(n3854), .Z(n3856) );
  XOR U5530 ( .A(\w3[2][65] ), .B(n3856), .Z(\w1[3][89] ) );
  XOR U5531 ( .A(\w3[2][9] ), .B(key[392]), .Z(n3858) );
  XNOR U5532 ( .A(\w3[2][1] ), .B(\w3[2][0] ), .Z(n3857) );
  XNOR U5533 ( .A(n3858), .B(n3857), .Z(n3859) );
  XOR U5534 ( .A(n3860), .B(n3859), .Z(\w1[3][8] ) );
  XOR U5535 ( .A(\w3[2][83] ), .B(key[474]), .Z(n3863) );
  XNOR U5536 ( .A(n3861), .B(\w3[2][91] ), .Z(n3862) );
  XNOR U5537 ( .A(n3863), .B(n3862), .Z(n3864) );
  XOR U5538 ( .A(\w3[2][66] ), .B(n3864), .Z(\w1[3][90] ) );
  XOR U5539 ( .A(n3865), .B(key[475]), .Z(n3868) );
  XNOR U5540 ( .A(\w3[2][67] ), .B(n3866), .Z(n3867) );
  XNOR U5541 ( .A(n3868), .B(n3867), .Z(\w1[3][91] ) );
  XOR U5542 ( .A(n3869), .B(key[476]), .Z(n3872) );
  XNOR U5543 ( .A(\w3[2][68] ), .B(n3870), .Z(n3871) );
  XNOR U5544 ( .A(n3872), .B(n3871), .Z(\w1[3][92] ) );
  XOR U5545 ( .A(\w3[2][86] ), .B(key[477]), .Z(n3875) );
  XNOR U5546 ( .A(n3873), .B(\w3[2][94] ), .Z(n3874) );
  XNOR U5547 ( .A(n3875), .B(n3874), .Z(n3876) );
  XOR U5548 ( .A(\w3[2][69] ), .B(n3876), .Z(\w1[3][93] ) );
  XOR U5549 ( .A(n3877), .B(key[478]), .Z(n3880) );
  XNOR U5550 ( .A(\w3[2][70] ), .B(n3878), .Z(n3879) );
  XNOR U5551 ( .A(n3880), .B(n3879), .Z(\w1[3][94] ) );
  XOR U5552 ( .A(n3881), .B(key[479]), .Z(n3884) );
  XNOR U5553 ( .A(n3882), .B(\w3[2][71] ), .Z(n3883) );
  XNOR U5554 ( .A(n3884), .B(n3883), .Z(\w1[3][95] ) );
  XOR U5555 ( .A(\w3[2][104] ), .B(key[480]), .Z(n3888) );
  XOR U5556 ( .A(n3886), .B(n3885), .Z(n3887) );
  XNOR U5557 ( .A(n3888), .B(n3887), .Z(\w1[3][96] ) );
  XOR U5558 ( .A(n3889), .B(key[481]), .Z(n3892) );
  XNOR U5559 ( .A(\w3[2][121] ), .B(n3890), .Z(n3891) );
  XNOR U5560 ( .A(n3892), .B(n3891), .Z(\w1[3][97] ) );
  XOR U5561 ( .A(n3893), .B(key[482]), .Z(n3896) );
  XNOR U5562 ( .A(\w3[2][122] ), .B(n3894), .Z(n3895) );
  XNOR U5563 ( .A(n3896), .B(n3895), .Z(\w1[3][98] ) );
  XOR U5564 ( .A(n3897), .B(key[483]), .Z(n3900) );
  XNOR U5565 ( .A(n3898), .B(\w3[2][123] ), .Z(n3899) );
  XNOR U5566 ( .A(n3900), .B(n3899), .Z(\w1[3][99] ) );
  XOR U5567 ( .A(\w3[2][10] ), .B(key[393]), .Z(n3902) );
  XNOR U5568 ( .A(\w3[2][2] ), .B(\w3[2][17] ), .Z(n3901) );
  XNOR U5569 ( .A(n3902), .B(n3901), .Z(n3903) );
  XOR U5570 ( .A(n3904), .B(n3903), .Z(\w1[3][9] ) );
  XOR U5571 ( .A(key[512]), .B(\w0[4][0] ), .Z(\w1[4][0] ) );
  XOR U5572 ( .A(key[612]), .B(\w0[4][100] ), .Z(\w1[4][100] ) );
  XOR U5573 ( .A(key[613]), .B(\w0[4][101] ), .Z(\w1[4][101] ) );
  XOR U5574 ( .A(key[614]), .B(\w0[4][102] ), .Z(\w1[4][102] ) );
  XOR U5575 ( .A(key[615]), .B(\w0[4][103] ), .Z(\w1[4][103] ) );
  XOR U5576 ( .A(key[616]), .B(\w0[4][104] ), .Z(\w1[4][104] ) );
  XOR U5577 ( .A(key[617]), .B(\w0[4][105] ), .Z(\w1[4][105] ) );
  XOR U5578 ( .A(key[618]), .B(\w0[4][106] ), .Z(\w1[4][106] ) );
  XOR U5579 ( .A(key[619]), .B(\w0[4][107] ), .Z(\w1[4][107] ) );
  XOR U5580 ( .A(key[620]), .B(\w0[4][108] ), .Z(\w1[4][108] ) );
  XOR U5581 ( .A(key[621]), .B(\w0[4][109] ), .Z(\w1[4][109] ) );
  XOR U5582 ( .A(key[522]), .B(\w0[4][10] ), .Z(\w1[4][10] ) );
  XOR U5583 ( .A(key[622]), .B(\w0[4][110] ), .Z(\w1[4][110] ) );
  XOR U5584 ( .A(key[623]), .B(\w0[4][111] ), .Z(\w1[4][111] ) );
  XOR U5585 ( .A(key[624]), .B(\w0[4][112] ), .Z(\w1[4][112] ) );
  XOR U5586 ( .A(key[625]), .B(\w0[4][113] ), .Z(\w1[4][113] ) );
  XOR U5587 ( .A(key[626]), .B(\w0[4][114] ), .Z(\w1[4][114] ) );
  XOR U5588 ( .A(key[627]), .B(\w0[4][115] ), .Z(\w1[4][115] ) );
  XOR U5589 ( .A(key[628]), .B(\w0[4][116] ), .Z(\w1[4][116] ) );
  XOR U5590 ( .A(key[629]), .B(\w0[4][117] ), .Z(\w1[4][117] ) );
  XOR U5591 ( .A(key[630]), .B(\w0[4][118] ), .Z(\w1[4][118] ) );
  XOR U5592 ( .A(key[631]), .B(\w0[4][119] ), .Z(\w1[4][119] ) );
  XOR U5593 ( .A(key[523]), .B(\w0[4][11] ), .Z(\w1[4][11] ) );
  XOR U5594 ( .A(key[632]), .B(\w0[4][120] ), .Z(\w1[4][120] ) );
  XOR U5595 ( .A(key[633]), .B(\w0[4][121] ), .Z(\w1[4][121] ) );
  XOR U5596 ( .A(key[634]), .B(\w0[4][122] ), .Z(\w1[4][122] ) );
  XOR U5597 ( .A(key[635]), .B(\w0[4][123] ), .Z(\w1[4][123] ) );
  XOR U5598 ( .A(key[636]), .B(\w0[4][124] ), .Z(\w1[4][124] ) );
  XOR U5599 ( .A(key[637]), .B(\w0[4][125] ), .Z(\w1[4][125] ) );
  XOR U5600 ( .A(key[638]), .B(\w0[4][126] ), .Z(\w1[4][126] ) );
  XOR U5601 ( .A(key[639]), .B(\w0[4][127] ), .Z(\w1[4][127] ) );
  XOR U5602 ( .A(key[524]), .B(\w0[4][12] ), .Z(\w1[4][12] ) );
  XOR U5603 ( .A(key[525]), .B(\w0[4][13] ), .Z(\w1[4][13] ) );
  XOR U5604 ( .A(key[526]), .B(\w0[4][14] ), .Z(\w1[4][14] ) );
  XOR U5605 ( .A(key[527]), .B(\w0[4][15] ), .Z(\w1[4][15] ) );
  XOR U5606 ( .A(key[528]), .B(\w0[4][16] ), .Z(\w1[4][16] ) );
  XOR U5607 ( .A(key[529]), .B(\w0[4][17] ), .Z(\w1[4][17] ) );
  XOR U5608 ( .A(key[530]), .B(\w0[4][18] ), .Z(\w1[4][18] ) );
  XOR U5609 ( .A(key[531]), .B(\w0[4][19] ), .Z(\w1[4][19] ) );
  XOR U5610 ( .A(key[513]), .B(\w0[4][1] ), .Z(\w1[4][1] ) );
  XOR U5611 ( .A(key[532]), .B(\w0[4][20] ), .Z(\w1[4][20] ) );
  XOR U5612 ( .A(key[533]), .B(\w0[4][21] ), .Z(\w1[4][21] ) );
  XOR U5613 ( .A(key[534]), .B(\w0[4][22] ), .Z(\w1[4][22] ) );
  XOR U5614 ( .A(key[535]), .B(\w0[4][23] ), .Z(\w1[4][23] ) );
  XOR U5615 ( .A(key[536]), .B(\w0[4][24] ), .Z(\w1[4][24] ) );
  XOR U5616 ( .A(key[537]), .B(\w0[4][25] ), .Z(\w1[4][25] ) );
  XOR U5617 ( .A(key[538]), .B(\w0[4][26] ), .Z(\w1[4][26] ) );
  XOR U5618 ( .A(key[539]), .B(\w0[4][27] ), .Z(\w1[4][27] ) );
  XOR U5619 ( .A(key[540]), .B(\w0[4][28] ), .Z(\w1[4][28] ) );
  XOR U5620 ( .A(key[541]), .B(\w0[4][29] ), .Z(\w1[4][29] ) );
  XOR U5621 ( .A(key[514]), .B(\w0[4][2] ), .Z(\w1[4][2] ) );
  XOR U5622 ( .A(key[542]), .B(\w0[4][30] ), .Z(\w1[4][30] ) );
  XOR U5623 ( .A(key[543]), .B(\w0[4][31] ), .Z(\w1[4][31] ) );
  XOR U5624 ( .A(key[544]), .B(\w0[4][32] ), .Z(\w1[4][32] ) );
  XOR U5625 ( .A(key[545]), .B(\w0[4][33] ), .Z(\w1[4][33] ) );
  XOR U5626 ( .A(key[546]), .B(\w0[4][34] ), .Z(\w1[4][34] ) );
  XOR U5627 ( .A(key[547]), .B(\w0[4][35] ), .Z(\w1[4][35] ) );
  XOR U5628 ( .A(key[548]), .B(\w0[4][36] ), .Z(\w1[4][36] ) );
  XOR U5629 ( .A(key[549]), .B(\w0[4][37] ), .Z(\w1[4][37] ) );
  XOR U5630 ( .A(key[550]), .B(\w0[4][38] ), .Z(\w1[4][38] ) );
  XOR U5631 ( .A(key[551]), .B(\w0[4][39] ), .Z(\w1[4][39] ) );
  XOR U5632 ( .A(key[515]), .B(\w0[4][3] ), .Z(\w1[4][3] ) );
  XOR U5633 ( .A(key[552]), .B(\w0[4][40] ), .Z(\w1[4][40] ) );
  XOR U5634 ( .A(key[553]), .B(\w0[4][41] ), .Z(\w1[4][41] ) );
  XOR U5635 ( .A(key[554]), .B(\w0[4][42] ), .Z(\w1[4][42] ) );
  XOR U5636 ( .A(key[555]), .B(\w0[4][43] ), .Z(\w1[4][43] ) );
  XOR U5637 ( .A(key[556]), .B(\w0[4][44] ), .Z(\w1[4][44] ) );
  XOR U5638 ( .A(key[557]), .B(\w0[4][45] ), .Z(\w1[4][45] ) );
  XOR U5639 ( .A(key[558]), .B(\w0[4][46] ), .Z(\w1[4][46] ) );
  XOR U5640 ( .A(key[559]), .B(\w0[4][47] ), .Z(\w1[4][47] ) );
  XOR U5641 ( .A(key[560]), .B(\w0[4][48] ), .Z(\w1[4][48] ) );
  XOR U5642 ( .A(key[561]), .B(\w0[4][49] ), .Z(\w1[4][49] ) );
  XOR U5643 ( .A(key[516]), .B(\w0[4][4] ), .Z(\w1[4][4] ) );
  XOR U5644 ( .A(key[562]), .B(\w0[4][50] ), .Z(\w1[4][50] ) );
  XOR U5645 ( .A(key[563]), .B(\w0[4][51] ), .Z(\w1[4][51] ) );
  XOR U5646 ( .A(key[564]), .B(\w0[4][52] ), .Z(\w1[4][52] ) );
  XOR U5647 ( .A(key[565]), .B(\w0[4][53] ), .Z(\w1[4][53] ) );
  XOR U5648 ( .A(key[566]), .B(\w0[4][54] ), .Z(\w1[4][54] ) );
  XOR U5649 ( .A(key[567]), .B(\w0[4][55] ), .Z(\w1[4][55] ) );
  XOR U5650 ( .A(key[568]), .B(\w0[4][56] ), .Z(\w1[4][56] ) );
  XOR U5651 ( .A(key[569]), .B(\w0[4][57] ), .Z(\w1[4][57] ) );
  XOR U5652 ( .A(key[570]), .B(\w0[4][58] ), .Z(\w1[4][58] ) );
  XOR U5653 ( .A(key[571]), .B(\w0[4][59] ), .Z(\w1[4][59] ) );
  XOR U5654 ( .A(key[517]), .B(\w0[4][5] ), .Z(\w1[4][5] ) );
  XOR U5655 ( .A(key[572]), .B(\w0[4][60] ), .Z(\w1[4][60] ) );
  XOR U5656 ( .A(key[573]), .B(\w0[4][61] ), .Z(\w1[4][61] ) );
  XOR U5657 ( .A(key[574]), .B(\w0[4][62] ), .Z(\w1[4][62] ) );
  XOR U5658 ( .A(key[575]), .B(\w0[4][63] ), .Z(\w1[4][63] ) );
  XOR U5659 ( .A(key[576]), .B(\w0[4][64] ), .Z(\w1[4][64] ) );
  XOR U5660 ( .A(key[577]), .B(\w0[4][65] ), .Z(\w1[4][65] ) );
  XOR U5661 ( .A(key[578]), .B(\w0[4][66] ), .Z(\w1[4][66] ) );
  XOR U5662 ( .A(key[579]), .B(\w0[4][67] ), .Z(\w1[4][67] ) );
  XOR U5663 ( .A(key[580]), .B(\w0[4][68] ), .Z(\w1[4][68] ) );
  XOR U5664 ( .A(key[581]), .B(\w0[4][69] ), .Z(\w1[4][69] ) );
  XOR U5665 ( .A(key[518]), .B(\w0[4][6] ), .Z(\w1[4][6] ) );
  XOR U5666 ( .A(key[582]), .B(\w0[4][70] ), .Z(\w1[4][70] ) );
  XOR U5667 ( .A(key[583]), .B(\w0[4][71] ), .Z(\w1[4][71] ) );
  XOR U5668 ( .A(key[584]), .B(\w0[4][72] ), .Z(\w1[4][72] ) );
  XOR U5669 ( .A(key[585]), .B(\w0[4][73] ), .Z(\w1[4][73] ) );
  XOR U5670 ( .A(key[586]), .B(\w0[4][74] ), .Z(\w1[4][74] ) );
  XOR U5671 ( .A(key[587]), .B(\w0[4][75] ), .Z(\w1[4][75] ) );
  XOR U5672 ( .A(key[588]), .B(\w0[4][76] ), .Z(\w1[4][76] ) );
  XOR U5673 ( .A(key[589]), .B(\w0[4][77] ), .Z(\w1[4][77] ) );
  XOR U5674 ( .A(key[590]), .B(\w0[4][78] ), .Z(\w1[4][78] ) );
  XOR U5675 ( .A(key[591]), .B(\w0[4][79] ), .Z(\w1[4][79] ) );
  XOR U5676 ( .A(key[519]), .B(\w0[4][7] ), .Z(\w1[4][7] ) );
  XOR U5677 ( .A(key[592]), .B(\w0[4][80] ), .Z(\w1[4][80] ) );
  XOR U5678 ( .A(key[593]), .B(\w0[4][81] ), .Z(\w1[4][81] ) );
  XOR U5679 ( .A(key[594]), .B(\w0[4][82] ), .Z(\w1[4][82] ) );
  XOR U5680 ( .A(key[595]), .B(\w0[4][83] ), .Z(\w1[4][83] ) );
  XOR U5681 ( .A(key[596]), .B(\w0[4][84] ), .Z(\w1[4][84] ) );
  XOR U5682 ( .A(key[597]), .B(\w0[4][85] ), .Z(\w1[4][85] ) );
  XOR U5683 ( .A(key[598]), .B(\w0[4][86] ), .Z(\w1[4][86] ) );
  XOR U5684 ( .A(key[599]), .B(\w0[4][87] ), .Z(\w1[4][87] ) );
  XOR U5685 ( .A(key[600]), .B(\w0[4][88] ), .Z(\w1[4][88] ) );
  XOR U5686 ( .A(key[601]), .B(\w0[4][89] ), .Z(\w1[4][89] ) );
  XOR U5687 ( .A(key[520]), .B(\w0[4][8] ), .Z(\w1[4][8] ) );
  XOR U5688 ( .A(key[602]), .B(\w0[4][90] ), .Z(\w1[4][90] ) );
  XOR U5689 ( .A(key[603]), .B(\w0[4][91] ), .Z(\w1[4][91] ) );
  XOR U5690 ( .A(key[604]), .B(\w0[4][92] ), .Z(\w1[4][92] ) );
  XOR U5691 ( .A(key[605]), .B(\w0[4][93] ), .Z(\w1[4][93] ) );
  XOR U5692 ( .A(key[606]), .B(\w0[4][94] ), .Z(\w1[4][94] ) );
  XOR U5693 ( .A(key[607]), .B(\w0[4][95] ), .Z(\w1[4][95] ) );
  XOR U5694 ( .A(key[608]), .B(\w0[4][96] ), .Z(\w1[4][96] ) );
  XOR U5695 ( .A(key[609]), .B(\w0[4][97] ), .Z(\w1[4][97] ) );
  XOR U5696 ( .A(key[610]), .B(\w0[4][98] ), .Z(\w1[4][98] ) );
  XOR U5697 ( .A(key[611]), .B(\w0[4][99] ), .Z(\w1[4][99] ) );
  XOR U5698 ( .A(key[521]), .B(\w0[4][9] ), .Z(\w1[4][9] ) );
endmodule

