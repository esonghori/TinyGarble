
module aes_seq_CC10 ( clk, rst, e_init, g_input, o );
  input [127:0] e_init;
  input [127:0] g_input;
  output [127:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
  wire   [127:0] state;

  DFF \state_reg[127]  ( .D(state[127]), .CLK(clk), .RST(rst), .I(e_init[127]), 
        .Q(state[127]) );
  DFF \state_reg[126]  ( .D(state[126]), .CLK(clk), .RST(rst), .I(e_init[126]), 
        .Q(state[126]) );
  DFF \state_reg[125]  ( .D(state[125]), .CLK(clk), .RST(rst), .I(e_init[125]), 
        .Q(state[125]) );
  DFF \state_reg[124]  ( .D(state[124]), .CLK(clk), .RST(rst), .I(e_init[124]), 
        .Q(state[124]) );
  DFF \state_reg[123]  ( .D(state[123]), .CLK(clk), .RST(rst), .I(e_init[123]), 
        .Q(state[123]) );
  DFF \state_reg[122]  ( .D(state[122]), .CLK(clk), .RST(rst), .I(e_init[122]), 
        .Q(state[122]) );
  DFF \state_reg[121]  ( .D(state[121]), .CLK(clk), .RST(rst), .I(e_init[121]), 
        .Q(state[121]) );
  DFF \state_reg[120]  ( .D(state[120]), .CLK(clk), .RST(rst), .I(e_init[120]), 
        .Q(state[120]) );
  DFF \state_reg[119]  ( .D(state[119]), .CLK(clk), .RST(rst), .I(e_init[119]), 
        .Q(state[119]) );
  DFF \state_reg[118]  ( .D(state[118]), .CLK(clk), .RST(rst), .I(e_init[118]), 
        .Q(state[118]) );
  DFF \state_reg[117]  ( .D(state[117]), .CLK(clk), .RST(rst), .I(e_init[117]), 
        .Q(state[117]) );
  DFF \state_reg[116]  ( .D(state[116]), .CLK(clk), .RST(rst), .I(e_init[116]), 
        .Q(state[116]) );
  DFF \state_reg[115]  ( .D(state[115]), .CLK(clk), .RST(rst), .I(e_init[115]), 
        .Q(state[115]) );
  DFF \state_reg[114]  ( .D(state[114]), .CLK(clk), .RST(rst), .I(e_init[114]), 
        .Q(state[114]) );
  DFF \state_reg[113]  ( .D(state[113]), .CLK(clk), .RST(rst), .I(e_init[113]), 
        .Q(state[113]) );
  DFF \state_reg[112]  ( .D(state[112]), .CLK(clk), .RST(rst), .I(e_init[112]), 
        .Q(state[112]) );
  DFF \state_reg[111]  ( .D(state[111]), .CLK(clk), .RST(rst), .I(e_init[111]), 
        .Q(state[111]) );
  DFF \state_reg[110]  ( .D(state[110]), .CLK(clk), .RST(rst), .I(e_init[110]), 
        .Q(state[110]) );
  DFF \state_reg[109]  ( .D(state[109]), .CLK(clk), .RST(rst), .I(e_init[109]), 
        .Q(state[109]) );
  DFF \state_reg[108]  ( .D(state[108]), .CLK(clk), .RST(rst), .I(e_init[108]), 
        .Q(state[108]) );
  DFF \state_reg[107]  ( .D(state[107]), .CLK(clk), .RST(rst), .I(e_init[107]), 
        .Q(state[107]) );
  DFF \state_reg[106]  ( .D(state[106]), .CLK(clk), .RST(rst), .I(e_init[106]), 
        .Q(state[106]) );
  DFF \state_reg[105]  ( .D(state[105]), .CLK(clk), .RST(rst), .I(e_init[105]), 
        .Q(state[105]) );
  DFF \state_reg[104]  ( .D(state[104]), .CLK(clk), .RST(rst), .I(e_init[104]), 
        .Q(state[104]) );
  DFF \state_reg[103]  ( .D(state[103]), .CLK(clk), .RST(rst), .I(e_init[103]), 
        .Q(state[103]) );
  DFF \state_reg[102]  ( .D(state[102]), .CLK(clk), .RST(rst), .I(e_init[102]), 
        .Q(state[102]) );
  DFF \state_reg[101]  ( .D(state[101]), .CLK(clk), .RST(rst), .I(e_init[101]), 
        .Q(state[101]) );
  DFF \state_reg[100]  ( .D(state[100]), .CLK(clk), .RST(rst), .I(e_init[100]), 
        .Q(state[100]) );
  DFF \state_reg[99]  ( .D(state[99]), .CLK(clk), .RST(rst), .I(e_init[99]), 
        .Q(state[99]) );
  DFF \state_reg[98]  ( .D(state[98]), .CLK(clk), .RST(rst), .I(e_init[98]), 
        .Q(state[98]) );
  DFF \state_reg[97]  ( .D(state[97]), .CLK(clk), .RST(rst), .I(e_init[97]), 
        .Q(state[97]) );
  DFF \state_reg[96]  ( .D(state[96]), .CLK(clk), .RST(rst), .I(e_init[96]), 
        .Q(state[96]) );
  DFF \state_reg[95]  ( .D(state[95]), .CLK(clk), .RST(rst), .I(e_init[95]), 
        .Q(state[95]) );
  DFF \state_reg[94]  ( .D(state[94]), .CLK(clk), .RST(rst), .I(e_init[94]), 
        .Q(state[94]) );
  DFF \state_reg[93]  ( .D(state[93]), .CLK(clk), .RST(rst), .I(e_init[93]), 
        .Q(state[93]) );
  DFF \state_reg[92]  ( .D(state[92]), .CLK(clk), .RST(rst), .I(e_init[92]), 
        .Q(state[92]) );
  DFF \state_reg[91]  ( .D(state[91]), .CLK(clk), .RST(rst), .I(e_init[91]), 
        .Q(state[91]) );
  DFF \state_reg[90]  ( .D(state[90]), .CLK(clk), .RST(rst), .I(e_init[90]), 
        .Q(state[90]) );
  DFF \state_reg[89]  ( .D(state[89]), .CLK(clk), .RST(rst), .I(e_init[89]), 
        .Q(state[89]) );
  DFF \state_reg[88]  ( .D(state[88]), .CLK(clk), .RST(rst), .I(e_init[88]), 
        .Q(state[88]) );
  DFF \state_reg[87]  ( .D(state[87]), .CLK(clk), .RST(rst), .I(e_init[87]), 
        .Q(state[87]) );
  DFF \state_reg[86]  ( .D(state[86]), .CLK(clk), .RST(rst), .I(e_init[86]), 
        .Q(state[86]) );
  DFF \state_reg[85]  ( .D(state[85]), .CLK(clk), .RST(rst), .I(e_init[85]), 
        .Q(state[85]) );
  DFF \state_reg[84]  ( .D(state[84]), .CLK(clk), .RST(rst), .I(e_init[84]), 
        .Q(state[84]) );
  DFF \state_reg[83]  ( .D(state[83]), .CLK(clk), .RST(rst), .I(e_init[83]), 
        .Q(state[83]) );
  DFF \state_reg[82]  ( .D(state[82]), .CLK(clk), .RST(rst), .I(e_init[82]), 
        .Q(state[82]) );
  DFF \state_reg[81]  ( .D(state[81]), .CLK(clk), .RST(rst), .I(e_init[81]), 
        .Q(state[81]) );
  DFF \state_reg[80]  ( .D(state[80]), .CLK(clk), .RST(rst), .I(e_init[80]), 
        .Q(state[80]) );
  DFF \state_reg[79]  ( .D(state[79]), .CLK(clk), .RST(rst), .I(e_init[79]), 
        .Q(state[79]) );
  DFF \state_reg[78]  ( .D(state[78]), .CLK(clk), .RST(rst), .I(e_init[78]), 
        .Q(state[78]) );
  DFF \state_reg[77]  ( .D(state[77]), .CLK(clk), .RST(rst), .I(e_init[77]), 
        .Q(state[77]) );
  DFF \state_reg[76]  ( .D(state[76]), .CLK(clk), .RST(rst), .I(e_init[76]), 
        .Q(state[76]) );
  DFF \state_reg[75]  ( .D(state[75]), .CLK(clk), .RST(rst), .I(e_init[75]), 
        .Q(state[75]) );
  DFF \state_reg[74]  ( .D(state[74]), .CLK(clk), .RST(rst), .I(e_init[74]), 
        .Q(state[74]) );
  DFF \state_reg[73]  ( .D(state[73]), .CLK(clk), .RST(rst), .I(e_init[73]), 
        .Q(state[73]) );
  DFF \state_reg[72]  ( .D(state[72]), .CLK(clk), .RST(rst), .I(e_init[72]), 
        .Q(state[72]) );
  DFF \state_reg[71]  ( .D(state[71]), .CLK(clk), .RST(rst), .I(e_init[71]), 
        .Q(state[71]) );
  DFF \state_reg[70]  ( .D(state[70]), .CLK(clk), .RST(rst), .I(e_init[70]), 
        .Q(state[70]) );
  DFF \state_reg[69]  ( .D(state[69]), .CLK(clk), .RST(rst), .I(e_init[69]), 
        .Q(state[69]) );
  DFF \state_reg[68]  ( .D(state[68]), .CLK(clk), .RST(rst), .I(e_init[68]), 
        .Q(state[68]) );
  DFF \state_reg[67]  ( .D(state[67]), .CLK(clk), .RST(rst), .I(e_init[67]), 
        .Q(state[67]) );
  DFF \state_reg[66]  ( .D(state[66]), .CLK(clk), .RST(rst), .I(e_init[66]), 
        .Q(state[66]) );
  DFF \state_reg[65]  ( .D(state[65]), .CLK(clk), .RST(rst), .I(e_init[65]), 
        .Q(state[65]) );
  DFF \state_reg[64]  ( .D(state[64]), .CLK(clk), .RST(rst), .I(e_init[64]), 
        .Q(state[64]) );
  DFF \state_reg[63]  ( .D(state[63]), .CLK(clk), .RST(rst), .I(e_init[63]), 
        .Q(state[63]) );
  DFF \state_reg[62]  ( .D(state[62]), .CLK(clk), .RST(rst), .I(e_init[62]), 
        .Q(state[62]) );
  DFF \state_reg[61]  ( .D(state[61]), .CLK(clk), .RST(rst), .I(e_init[61]), 
        .Q(state[61]) );
  DFF \state_reg[60]  ( .D(state[60]), .CLK(clk), .RST(rst), .I(e_init[60]), 
        .Q(state[60]) );
  DFF \state_reg[59]  ( .D(state[59]), .CLK(clk), .RST(rst), .I(e_init[59]), 
        .Q(state[59]) );
  DFF \state_reg[58]  ( .D(state[58]), .CLK(clk), .RST(rst), .I(e_init[58]), 
        .Q(state[58]) );
  DFF \state_reg[57]  ( .D(state[57]), .CLK(clk), .RST(rst), .I(e_init[57]), 
        .Q(state[57]) );
  DFF \state_reg[56]  ( .D(state[56]), .CLK(clk), .RST(rst), .I(e_init[56]), 
        .Q(state[56]) );
  DFF \state_reg[55]  ( .D(state[55]), .CLK(clk), .RST(rst), .I(e_init[55]), 
        .Q(state[55]) );
  DFF \state_reg[54]  ( .D(state[54]), .CLK(clk), .RST(rst), .I(e_init[54]), 
        .Q(state[54]) );
  DFF \state_reg[53]  ( .D(state[53]), .CLK(clk), .RST(rst), .I(e_init[53]), 
        .Q(state[53]) );
  DFF \state_reg[52]  ( .D(state[52]), .CLK(clk), .RST(rst), .I(e_init[52]), 
        .Q(state[52]) );
  DFF \state_reg[51]  ( .D(state[51]), .CLK(clk), .RST(rst), .I(e_init[51]), 
        .Q(state[51]) );
  DFF \state_reg[50]  ( .D(state[50]), .CLK(clk), .RST(rst), .I(e_init[50]), 
        .Q(state[50]) );
  DFF \state_reg[49]  ( .D(state[49]), .CLK(clk), .RST(rst), .I(e_init[49]), 
        .Q(state[49]) );
  DFF \state_reg[48]  ( .D(state[48]), .CLK(clk), .RST(rst), .I(e_init[48]), 
        .Q(state[48]) );
  DFF \state_reg[47]  ( .D(state[47]), .CLK(clk), .RST(rst), .I(e_init[47]), 
        .Q(state[47]) );
  DFF \state_reg[46]  ( .D(state[46]), .CLK(clk), .RST(rst), .I(e_init[46]), 
        .Q(state[46]) );
  DFF \state_reg[45]  ( .D(state[45]), .CLK(clk), .RST(rst), .I(e_init[45]), 
        .Q(state[45]) );
  DFF \state_reg[44]  ( .D(state[44]), .CLK(clk), .RST(rst), .I(e_init[44]), 
        .Q(state[44]) );
  DFF \state_reg[43]  ( .D(state[43]), .CLK(clk), .RST(rst), .I(e_init[43]), 
        .Q(state[43]) );
  DFF \state_reg[42]  ( .D(state[42]), .CLK(clk), .RST(rst), .I(e_init[42]), 
        .Q(state[42]) );
  DFF \state_reg[41]  ( .D(state[41]), .CLK(clk), .RST(rst), .I(e_init[41]), 
        .Q(state[41]) );
  DFF \state_reg[40]  ( .D(state[40]), .CLK(clk), .RST(rst), .I(e_init[40]), 
        .Q(state[40]) );
  DFF \state_reg[39]  ( .D(state[39]), .CLK(clk), .RST(rst), .I(e_init[39]), 
        .Q(state[39]) );
  DFF \state_reg[38]  ( .D(state[38]), .CLK(clk), .RST(rst), .I(e_init[38]), 
        .Q(state[38]) );
  DFF \state_reg[37]  ( .D(state[37]), .CLK(clk), .RST(rst), .I(e_init[37]), 
        .Q(state[37]) );
  DFF \state_reg[36]  ( .D(state[36]), .CLK(clk), .RST(rst), .I(e_init[36]), 
        .Q(state[36]) );
  DFF \state_reg[35]  ( .D(state[35]), .CLK(clk), .RST(rst), .I(e_init[35]), 
        .Q(state[35]) );
  DFF \state_reg[34]  ( .D(state[34]), .CLK(clk), .RST(rst), .I(e_init[34]), 
        .Q(state[34]) );
  DFF \state_reg[33]  ( .D(state[33]), .CLK(clk), .RST(rst), .I(e_init[33]), 
        .Q(state[33]) );
  DFF \state_reg[32]  ( .D(state[32]), .CLK(clk), .RST(rst), .I(e_init[32]), 
        .Q(state[32]) );
  DFF \state_reg[31]  ( .D(state[31]), .CLK(clk), .RST(rst), .I(e_init[31]), 
        .Q(state[31]) );
  DFF \state_reg[30]  ( .D(state[30]), .CLK(clk), .RST(rst), .I(e_init[30]), 
        .Q(state[30]) );
  DFF \state_reg[29]  ( .D(state[29]), .CLK(clk), .RST(rst), .I(e_init[29]), 
        .Q(state[29]) );
  DFF \state_reg[28]  ( .D(state[28]), .CLK(clk), .RST(rst), .I(e_init[28]), 
        .Q(state[28]) );
  DFF \state_reg[27]  ( .D(state[27]), .CLK(clk), .RST(rst), .I(e_init[27]), 
        .Q(state[27]) );
  DFF \state_reg[26]  ( .D(state[26]), .CLK(clk), .RST(rst), .I(e_init[26]), 
        .Q(state[26]) );
  DFF \state_reg[25]  ( .D(state[25]), .CLK(clk), .RST(rst), .I(e_init[25]), 
        .Q(state[25]) );
  DFF \state_reg[24]  ( .D(state[24]), .CLK(clk), .RST(rst), .I(e_init[24]), 
        .Q(state[24]) );
  DFF \state_reg[23]  ( .D(state[23]), .CLK(clk), .RST(rst), .I(e_init[23]), 
        .Q(state[23]) );
  DFF \state_reg[22]  ( .D(state[22]), .CLK(clk), .RST(rst), .I(e_init[22]), 
        .Q(state[22]) );
  DFF \state_reg[21]  ( .D(state[21]), .CLK(clk), .RST(rst), .I(e_init[21]), 
        .Q(state[21]) );
  DFF \state_reg[20]  ( .D(state[20]), .CLK(clk), .RST(rst), .I(e_init[20]), 
        .Q(state[20]) );
  DFF \state_reg[19]  ( .D(state[19]), .CLK(clk), .RST(rst), .I(e_init[19]), 
        .Q(state[19]) );
  DFF \state_reg[18]  ( .D(state[18]), .CLK(clk), .RST(rst), .I(e_init[18]), 
        .Q(state[18]) );
  DFF \state_reg[17]  ( .D(state[17]), .CLK(clk), .RST(rst), .I(e_init[17]), 
        .Q(state[17]) );
  DFF \state_reg[16]  ( .D(state[16]), .CLK(clk), .RST(rst), .I(e_init[16]), 
        .Q(state[16]) );
  DFF \state_reg[15]  ( .D(state[15]), .CLK(clk), .RST(rst), .I(e_init[15]), 
        .Q(state[15]) );
  DFF \state_reg[14]  ( .D(state[14]), .CLK(clk), .RST(rst), .I(e_init[14]), 
        .Q(state[14]) );
  DFF \state_reg[13]  ( .D(state[13]), .CLK(clk), .RST(rst), .I(e_init[13]), 
        .Q(state[13]) );
  DFF \state_reg[12]  ( .D(state[12]), .CLK(clk), .RST(rst), .I(e_init[12]), 
        .Q(state[12]) );
  DFF \state_reg[11]  ( .D(state[11]), .CLK(clk), .RST(rst), .I(e_init[11]), 
        .Q(state[11]) );
  DFF \state_reg[10]  ( .D(state[10]), .CLK(clk), .RST(rst), .I(e_init[10]), 
        .Q(state[10]) );
  DFF \state_reg[9]  ( .D(state[9]), .CLK(clk), .RST(rst), .I(e_init[9]), .Q(
        state[9]) );
  DFF \state_reg[8]  ( .D(state[8]), .CLK(clk), .RST(rst), .I(e_init[8]), .Q(
        state[8]) );
  DFF \state_reg[7]  ( .D(state[7]), .CLK(clk), .RST(rst), .I(e_init[7]), .Q(
        state[7]) );
  DFF \state_reg[6]  ( .D(state[6]), .CLK(clk), .RST(rst), .I(e_init[6]), .Q(
        state[6]) );
  DFF \state_reg[5]  ( .D(state[5]), .CLK(clk), .RST(rst), .I(e_init[5]), .Q(
        state[5]) );
  DFF \state_reg[4]  ( .D(state[4]), .CLK(clk), .RST(rst), .I(e_init[4]), .Q(
        state[4]) );
  DFF \state_reg[3]  ( .D(state[3]), .CLK(clk), .RST(rst), .I(e_init[3]), .Q(
        state[3]) );
  DFF \state_reg[2]  ( .D(state[2]), .CLK(clk), .RST(rst), .I(e_init[2]), .Q(
        state[2]) );
  DFF \state_reg[1]  ( .D(state[1]), .CLK(clk), .RST(rst), .I(e_init[1]), .Q(
        state[1]) );
  DFF \state_reg[0]  ( .D(state[0]), .CLK(clk), .RST(rst), .I(e_init[0]), .Q(
        state[0]) );
  ANDN U4 ( .A(n566), .B(n584), .Z(n575) );
  NOR U5 ( .A(n2301), .B(n2331), .Z(n2378) );
  ANDN U6 ( .A(n2434), .B(n2443), .Z(n2438) );
  XOR U7 ( .A(n2102), .B(n2083), .Z(n2097) );
  ANDN U8 ( .A(n1588), .B(n1597), .Z(n1592) );
  ANDN U9 ( .A(n1405), .B(n1414), .Z(n1409) );
  ANDN U10 ( .A(n1246), .B(n1255), .Z(n1250) );
  ANDN U11 ( .A(n1079), .B(n1088), .Z(n1083) );
  ANDN U12 ( .A(n923), .B(n932), .Z(n927) );
  ANDN U13 ( .A(n765), .B(n774), .Z(n769) );
  XOR U14 ( .A(n520), .B(n570), .Z(n551) );
  ANDN U15 ( .A(n267), .B(n276), .Z(n271) );
  ANDN U16 ( .A(n111), .B(n120), .Z(n115) );
  XNOR U17 ( .A(n2298), .B(n2319), .Z(n2321) );
  ANDN U18 ( .A(n2205), .B(n2214), .Z(n2209) );
  ANDN U19 ( .A(n1964), .B(n1973), .Z(n1968) );
  ANDN U20 ( .A(n1780), .B(n1789), .Z(n1784) );
  XNOR U21 ( .A(n1512), .B(n1516), .Z(n1514) );
  XOR U22 ( .A(n2441), .B(n703), .Z(n2437) );
  XNOR U23 ( .A(n1043), .B(n1047), .Z(n1045) );
  XOR U24 ( .A(n1086), .B(n1015), .Z(n1082) );
  XNOR U25 ( .A(n655), .B(n656), .Z(n642) );
  XNOR U26 ( .A(n231), .B(n235), .Z(n233) );
  XOR U27 ( .A(n274), .B(n203), .Z(n270) );
  ANDN U28 ( .A(n2345), .B(n2344), .Z(n2339) );
  XNOR U29 ( .A(n1859), .B(n1875), .Z(n1867) );
  XOR U30 ( .A(n1536), .B(n1584), .Z(n1552) );
  XNOR U31 ( .A(n1644), .B(n1646), .Z(n1566) );
  XOR U32 ( .A(n1353), .B(n1401), .Z(n1369) );
  XNOR U33 ( .A(n1461), .B(n1463), .Z(n1383) );
  XOR U34 ( .A(n1194), .B(n1242), .Z(n1210) );
  XOR U35 ( .A(n869), .B(n919), .Z(n887) );
  XNOR U36 ( .A(n979), .B(n981), .Z(n901) );
  XOR U37 ( .A(n713), .B(n761), .Z(n729) );
  XNOR U38 ( .A(n821), .B(n823), .Z(n743) );
  XNOR U39 ( .A(n600), .B(n597), .Z(n570) );
  XOR U40 ( .A(n56), .B(n107), .Z(n75) );
  XNOR U41 ( .A(n167), .B(n169), .Z(n89) );
  XOR U42 ( .A(n2153), .B(n2201), .Z(n2169) );
  XOR U43 ( .A(n1912), .B(n1960), .Z(n1928) );
  XOR U44 ( .A(n1728), .B(n1776), .Z(n1744) );
  XNOR U45 ( .A(n1836), .B(n1838), .Z(n1758) );
  XOR U46 ( .A(n2071), .B(n2075), .Z(n2066) );
  XOR U47 ( .A(n447), .B(n439), .Z(n442) );
  XOR U48 ( .A(n1670), .B(n1690), .Z(n1873) );
  XNOR U49 ( .A(n1854), .B(n1859), .Z(n1860) );
  XNOR U50 ( .A(n1552), .B(n1556), .Z(n1554) );
  XOR U51 ( .A(n1595), .B(n1497), .Z(n1591) );
  XNOR U52 ( .A(n1369), .B(n1373), .Z(n1371) );
  XOR U53 ( .A(n1412), .B(n1341), .Z(n1408) );
  XNOR U54 ( .A(n1210), .B(n1214), .Z(n1212) );
  XOR U55 ( .A(n1253), .B(n1182), .Z(n1249) );
  XNOR U56 ( .A(n887), .B(n891), .Z(n889) );
  XOR U57 ( .A(n930), .B(n857), .Z(n926) );
  XNOR U58 ( .A(n729), .B(n733), .Z(n731) );
  XOR U59 ( .A(n772), .B(n685), .Z(n768) );
  XNOR U60 ( .A(n75), .B(n79), .Z(n77) );
  XOR U61 ( .A(n118), .B(n44), .Z(n114) );
  XNOR U62 ( .A(n2309), .B(n2301), .Z(n2307) );
  XNOR U63 ( .A(n2290), .B(n2310), .Z(n2298) );
  XNOR U64 ( .A(n2169), .B(n2173), .Z(n2171) );
  XOR U65 ( .A(n2212), .B(n2141), .Z(n2208) );
  XNOR U66 ( .A(n1928), .B(n1932), .Z(n1930) );
  XOR U67 ( .A(n1971), .B(n1900), .Z(n1967) );
  XNOR U68 ( .A(n1744), .B(n1748), .Z(n1746) );
  XOR U69 ( .A(n1787), .B(n1716), .Z(n1783) );
  XOR U70 ( .A(n1156), .B(n2430), .Z(n1512) );
  XNOR U71 ( .A(n2490), .B(n2492), .Z(n1526) );
  XNOR U72 ( .A(n2111), .B(n2113), .Z(n2044) );
  XOR U73 ( .A(n1027), .B(n1075), .Z(n1043) );
  XNOR U74 ( .A(n1135), .B(n1137), .Z(n1057) );
  XNOR U75 ( .A(n521), .B(n542), .Z(n544) );
  ANDN U76 ( .A(n543), .B(n580), .Z(n558) );
  XNOR U77 ( .A(n491), .B(n493), .Z(n410) );
  XOR U78 ( .A(n215), .B(n263), .Z(n231) );
  XNOR U79 ( .A(n323), .B(n325), .Z(n245) );
  ANDN U80 ( .A(n632), .B(n530), .Z(n528) );
  XOR U81 ( .A(g_input[23]), .B(n1477), .Z(n1476) );
  XOR U82 ( .A(g_input[31]), .B(n1319), .Z(n1318) );
  XOR U83 ( .A(g_input[39]), .B(n1162), .Z(n1161) );
  XOR U84 ( .A(g_input[55]), .B(n837), .Z(n836) );
  XOR U85 ( .A(g_input[63]), .B(n665), .Z(n664) );
  XOR U86 ( .A(g_input[95]), .B(n24), .Z(n23) );
  XOR U87 ( .A(g_input[111]), .B(n2037), .Z(n2036) );
  XOR U88 ( .A(g_input[119]), .B(n1880), .Z(n1879) );
  XOR U89 ( .A(g_input[127]), .B(n1696), .Z(n1695) );
  XOR U90 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U91 ( .A(g_input[9]), .B(n3), .Z(n2) );
  XOR U92 ( .A(n4), .B(n5), .Z(n1) );
  XOR U93 ( .A(n6), .B(n7), .Z(o[99]) );
  XNOR U94 ( .A(n8), .B(n9), .Z(n7) );
  XNOR U95 ( .A(g_input[99]), .B(n10), .Z(n9) );
  XNOR U96 ( .A(n11), .B(n12), .Z(n6) );
  XNOR U97 ( .A(n13), .B(g_input[98]), .Z(o[98]) );
  XOR U98 ( .A(n14), .B(n15), .Z(o[97]) );
  XNOR U99 ( .A(g_input[97]), .B(n8), .Z(n15) );
  XOR U100 ( .A(n16), .B(n12), .Z(n14) );
  XOR U101 ( .A(n17), .B(n18), .Z(o[96]) );
  XNOR U102 ( .A(n19), .B(g_input[96]), .Z(n17) );
  XOR U103 ( .A(n20), .B(n21), .Z(o[95]) );
  XOR U104 ( .A(n22), .B(n23), .Z(n21) );
  XOR U105 ( .A(n25), .B(n26), .Z(n20) );
  XNOR U106 ( .A(n27), .B(n28), .Z(o[94]) );
  XNOR U107 ( .A(n24), .B(g_input[94]), .Z(n27) );
  XOR U108 ( .A(n29), .B(n30), .Z(o[93]) );
  XOR U109 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U110 ( .A(g_input[93]), .B(n33), .Z(n32) );
  NOR U111 ( .A(n34), .B(n35), .Z(n31) );
  XNOR U112 ( .A(n36), .B(n37), .Z(n29) );
  XOR U113 ( .A(n25), .B(n38), .Z(n36) );
  XNOR U114 ( .A(n39), .B(n40), .Z(n25) );
  XNOR U115 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U116 ( .B(n43), .A(n44), .Z(n41) );
  XNOR U117 ( .A(n45), .B(n46), .Z(o[92]) );
  XOR U118 ( .A(n37), .B(g_input[92]), .Z(n45) );
  XOR U119 ( .A(n47), .B(n48), .Z(o[91]) );
  XOR U120 ( .A(n22), .B(n49), .Z(n48) );
  XNOR U121 ( .A(g_input[91]), .B(n50), .Z(n49) );
  XNOR U122 ( .A(n28), .B(n26), .Z(n47) );
  XNOR U123 ( .A(n51), .B(n52), .Z(n28) );
  XNOR U124 ( .A(n53), .B(n33), .Z(n51) );
  NANDN U125 ( .B(n54), .A(n55), .Z(n33) );
  NANDN U126 ( .B(n56), .A(n57), .Z(n53) );
  XOR U127 ( .A(n46), .B(g_input[90]), .Z(o[90]) );
  XOR U128 ( .A(n58), .B(n59), .Z(n46) );
  XNOR U129 ( .A(n60), .B(n61), .Z(o[8]) );
  XOR U130 ( .A(n62), .B(g_input[8]), .Z(n60) );
  XOR U131 ( .A(n63), .B(n64), .Z(o[89]) );
  XOR U132 ( .A(g_input[89]), .B(n24), .Z(n64) );
  XOR U133 ( .A(n50), .B(n59), .Z(n24) );
  XNOR U134 ( .A(n65), .B(n38), .Z(n50) );
  XOR U135 ( .A(n66), .B(n67), .Z(n65) );
  ANDN U136 ( .A(n68), .B(n69), .Z(n67) );
  XNOR U137 ( .A(n58), .B(n22), .Z(n63) );
  XOR U138 ( .A(n70), .B(n52), .Z(n22) );
  XNOR U139 ( .A(n71), .B(n38), .Z(n52) );
  XNOR U140 ( .A(n72), .B(n73), .Z(n38) );
  NOR U141 ( .A(n74), .B(n75), .Z(n73) );
  XOR U142 ( .A(n76), .B(n72), .Z(n71) );
  NOR U143 ( .A(n77), .B(n78), .Z(n72) );
  NANDN U144 ( .B(n79), .A(n80), .Z(n76) );
  XOR U145 ( .A(n66), .B(n81), .Z(n70) );
  ANDN U146 ( .A(n82), .B(n43), .Z(n81) );
  OR U147 ( .A(n83), .B(n84), .Z(n66) );
  IV U148 ( .A(n26), .Z(n58) );
  XNOR U149 ( .A(n85), .B(n86), .Z(n26) );
  XNOR U150 ( .A(n87), .B(n88), .Z(n85) );
  NOR U151 ( .A(n89), .B(n35), .Z(n88) );
  XNOR U152 ( .A(n90), .B(n37), .Z(o[88]) );
  XOR U153 ( .A(n91), .B(n40), .Z(n37) );
  XOR U154 ( .A(n92), .B(n86), .Z(n40) );
  XNOR U155 ( .A(n93), .B(n94), .Z(n92) );
  NOR U156 ( .A(n79), .B(n95), .Z(n94) );
  XNOR U157 ( .A(n87), .B(n96), .Z(n91) );
  NOR U158 ( .A(n56), .B(n97), .Z(n96) );
  ANDN U159 ( .A(n55), .B(n98), .Z(n87) );
  XOR U160 ( .A(n56), .B(n35), .Z(n55) );
  XOR U161 ( .A(n59), .B(g_input[88]), .Z(n90) );
  XNOR U162 ( .A(n99), .B(n86), .Z(n59) );
  XNOR U163 ( .A(n93), .B(n100), .Z(n86) );
  NOR U164 ( .A(n101), .B(n75), .Z(n100) );
  NOR U165 ( .A(n77), .B(n102), .Z(n93) );
  XNOR U166 ( .A(n69), .B(n35), .Z(n79) );
  XNOR U167 ( .A(n103), .B(n104), .Z(n35) );
  ANDN U168 ( .A(n105), .B(n106), .Z(n104) );
  IV U169 ( .A(n107), .Z(n43) );
  XNOR U170 ( .A(n103), .B(n108), .Z(n56) );
  NOR U171 ( .A(n109), .B(n110), .Z(n108) );
  ANDN U172 ( .A(n111), .B(n112), .Z(n103) );
  XNOR U173 ( .A(n113), .B(n42), .Z(n99) );
  OR U174 ( .A(n83), .B(n114), .Z(n42) );
  XOR U175 ( .A(n107), .B(n69), .Z(n83) );
  XOR U176 ( .A(n115), .B(n116), .Z(n107) );
  ANDN U177 ( .A(n117), .B(n110), .Z(n116) );
  OR U178 ( .A(n69), .B(n118), .Z(n113) );
  XOR U179 ( .A(n119), .B(n115), .Z(n69) );
  XOR U180 ( .A(n110), .B(n106), .Z(n111) );
  XNOR U181 ( .A(n121), .B(n122), .Z(n110) );
  XNOR U182 ( .A(n123), .B(n124), .Z(n121) );
  NANDN U183 ( .B(n125), .A(n105), .Z(n123) );
  OR U184 ( .A(n106), .B(n125), .Z(n119) );
  XOR U185 ( .A(n126), .B(n127), .Z(n106) );
  XOR U186 ( .A(n128), .B(n129), .Z(n127) );
  XNOR U187 ( .A(n124), .B(n130), .Z(n129) );
  ANDN U188 ( .A(n117), .B(n109), .Z(n130) );
  OR U189 ( .A(n112), .B(n120), .Z(n124) );
  XNOR U190 ( .A(n131), .B(n117), .Z(n120) );
  XOR U191 ( .A(n105), .B(n109), .Z(n112) );
  IV U192 ( .A(n128), .Z(n109) );
  XNOR U193 ( .A(n132), .B(n133), .Z(n128) );
  XNOR U194 ( .A(n118), .B(n134), .Z(n133) );
  XNOR U195 ( .A(n135), .B(n136), .Z(n134) );
  ANDN U196 ( .A(n44), .B(n137), .Z(n135) );
  XNOR U197 ( .A(n138), .B(n139), .Z(n132) );
  XOR U198 ( .A(n140), .B(n68), .Z(n138) );
  XOR U199 ( .A(n122), .B(n117), .Z(n126) );
  XNOR U200 ( .A(n141), .B(n142), .Z(n117) );
  XNOR U201 ( .A(n143), .B(n144), .Z(n142) );
  ANDN U202 ( .A(n57), .B(n97), .Z(n143) );
  XNOR U203 ( .A(n145), .B(n140), .Z(n141) );
  XOR U204 ( .A(n146), .B(n147), .Z(n140) );
  XNOR U205 ( .A(n148), .B(n149), .Z(n146) );
  NANDN U206 ( .B(n95), .A(n80), .Z(n148) );
  XNOR U207 ( .A(n131), .B(n105), .Z(n122) );
  XNOR U208 ( .A(n150), .B(n151), .Z(n105) );
  XOR U209 ( .A(n44), .B(n152), .Z(n151) );
  XNOR U210 ( .A(n153), .B(n136), .Z(n152) );
  OR U211 ( .A(n84), .B(n114), .Z(n136) );
  XNOR U212 ( .A(n82), .B(n68), .Z(n84) );
  IV U213 ( .A(n137), .Z(n82) );
  ANDN U214 ( .A(n68), .B(n118), .Z(n153) );
  XNOR U215 ( .A(n154), .B(n145), .Z(n150) );
  XOR U216 ( .A(n147), .B(n137), .Z(n154) );
  IV U217 ( .A(n125), .Z(n131) );
  XOR U218 ( .A(n155), .B(n156), .Z(n125) );
  XOR U219 ( .A(n147), .B(n157), .Z(n156) );
  XNOR U220 ( .A(n158), .B(n144), .Z(n157) );
  OR U221 ( .A(n54), .B(n98), .Z(n144) );
  XNOR U222 ( .A(n97), .B(n89), .Z(n98) );
  XNOR U223 ( .A(n159), .B(n57), .Z(n54) );
  ANDN U224 ( .A(n160), .B(n34), .Z(n158) );
  XNOR U225 ( .A(n149), .B(n161), .Z(n147) );
  ANDN U226 ( .A(n162), .B(n74), .Z(n161) );
  OR U227 ( .A(n102), .B(n78), .Z(n149) );
  XOR U228 ( .A(n74), .B(n80), .Z(n78) );
  XNOR U229 ( .A(n34), .B(n68), .Z(n80) );
  XNOR U230 ( .A(n163), .B(n57), .Z(n68) );
  XNOR U231 ( .A(n164), .B(n165), .Z(n163) );
  XOR U232 ( .A(n137), .B(n57), .Z(n74) );
  XOR U233 ( .A(n166), .B(n167), .Z(n137) );
  XNOR U234 ( .A(n168), .B(n169), .Z(n166) );
  XOR U235 ( .A(n162), .B(n95), .Z(n102) );
  XOR U236 ( .A(n160), .B(n118), .Z(n95) );
  XOR U237 ( .A(n170), .B(n171), .Z(n118) );
  XNOR U238 ( .A(n172), .B(n44), .Z(n171) );
  XNOR U239 ( .A(n173), .B(n168), .Z(n170) );
  XOR U240 ( .A(g_input[92]), .B(state[92]), .Z(n168) );
  IV U241 ( .A(n101), .Z(n162) );
  XOR U242 ( .A(n97), .B(n44), .Z(n101) );
  XNOR U243 ( .A(n145), .B(n139), .Z(n155) );
  XNOR U244 ( .A(n159), .B(n160), .Z(n139) );
  IV U245 ( .A(n89), .Z(n160) );
  IV U246 ( .A(n34), .Z(n159) );
  XOR U247 ( .A(n174), .B(n167), .Z(n34) );
  XNOR U248 ( .A(n165), .B(n169), .Z(n174) );
  XOR U249 ( .A(n57), .B(n97), .Z(n145) );
  XNOR U250 ( .A(n164), .B(n175), .Z(n97) );
  XNOR U251 ( .A(n172), .B(n169), .Z(n175) );
  XOR U252 ( .A(n176), .B(n165), .Z(n172) );
  XOR U253 ( .A(g_input[89]), .B(state[89]), .Z(n165) );
  XNOR U254 ( .A(g_input[91]), .B(state[91]), .Z(n176) );
  XOR U255 ( .A(g_input[90]), .B(state[90]), .Z(n164) );
  XNOR U256 ( .A(n177), .B(n167), .Z(n57) );
  XOR U257 ( .A(g_input[93]), .B(state[93]), .Z(n167) );
  XNOR U258 ( .A(n173), .B(n169), .Z(n177) );
  XNOR U259 ( .A(n178), .B(n44), .Z(n169) );
  XOR U260 ( .A(g_input[88]), .B(state[88]), .Z(n44) );
  XNOR U261 ( .A(g_input[94]), .B(state[94]), .Z(n178) );
  XOR U262 ( .A(g_input[95]), .B(state[95]), .Z(n173) );
  XOR U263 ( .A(n179), .B(n180), .Z(o[87]) );
  XOR U264 ( .A(n181), .B(n182), .Z(n180) );
  XOR U265 ( .A(g_input[87]), .B(n183), .Z(n182) );
  XOR U266 ( .A(n184), .B(n185), .Z(n179) );
  XNOR U267 ( .A(n186), .B(n187), .Z(o[86]) );
  XNOR U268 ( .A(n183), .B(g_input[86]), .Z(n186) );
  XOR U269 ( .A(n188), .B(n189), .Z(o[85]) );
  XOR U270 ( .A(n190), .B(n191), .Z(n189) );
  XNOR U271 ( .A(g_input[85]), .B(n192), .Z(n191) );
  NOR U272 ( .A(n193), .B(n194), .Z(n190) );
  XNOR U273 ( .A(n195), .B(n196), .Z(n188) );
  XOR U274 ( .A(n184), .B(n197), .Z(n195) );
  XNOR U275 ( .A(n198), .B(n199), .Z(n184) );
  XNOR U276 ( .A(n200), .B(n201), .Z(n198) );
  NANDN U277 ( .B(n202), .A(n203), .Z(n200) );
  XNOR U278 ( .A(n204), .B(n205), .Z(o[84]) );
  XOR U279 ( .A(n196), .B(g_input[84]), .Z(n204) );
  XOR U280 ( .A(n206), .B(n207), .Z(o[83]) );
  XOR U281 ( .A(n181), .B(n208), .Z(n207) );
  XNOR U282 ( .A(g_input[83]), .B(n209), .Z(n208) );
  XNOR U283 ( .A(n187), .B(n185), .Z(n206) );
  XNOR U284 ( .A(n210), .B(n211), .Z(n187) );
  XNOR U285 ( .A(n212), .B(n192), .Z(n210) );
  NANDN U286 ( .B(n213), .A(n214), .Z(n192) );
  NANDN U287 ( .B(n215), .A(n216), .Z(n212) );
  XOR U288 ( .A(n205), .B(g_input[82]), .Z(o[82]) );
  XOR U289 ( .A(n217), .B(n218), .Z(n205) );
  XOR U290 ( .A(n219), .B(n220), .Z(o[81]) );
  XOR U291 ( .A(g_input[81]), .B(n183), .Z(n220) );
  XOR U292 ( .A(n209), .B(n218), .Z(n183) );
  XNOR U293 ( .A(n221), .B(n197), .Z(n209) );
  XOR U294 ( .A(n222), .B(n223), .Z(n221) );
  ANDN U295 ( .A(n224), .B(n225), .Z(n223) );
  XNOR U296 ( .A(n217), .B(n181), .Z(n219) );
  XOR U297 ( .A(n226), .B(n211), .Z(n181) );
  XNOR U298 ( .A(n227), .B(n197), .Z(n211) );
  XNOR U299 ( .A(n228), .B(n229), .Z(n197) );
  NOR U300 ( .A(n230), .B(n231), .Z(n229) );
  XOR U301 ( .A(n232), .B(n228), .Z(n227) );
  NOR U302 ( .A(n233), .B(n234), .Z(n228) );
  NANDN U303 ( .B(n235), .A(n236), .Z(n232) );
  XOR U304 ( .A(n222), .B(n237), .Z(n226) );
  ANDN U305 ( .A(n238), .B(n202), .Z(n237) );
  OR U306 ( .A(n239), .B(n240), .Z(n222) );
  IV U307 ( .A(n185), .Z(n217) );
  XNOR U308 ( .A(n241), .B(n242), .Z(n185) );
  XNOR U309 ( .A(n243), .B(n244), .Z(n241) );
  NOR U310 ( .A(n245), .B(n194), .Z(n244) );
  XNOR U311 ( .A(n246), .B(n196), .Z(o[80]) );
  XOR U312 ( .A(n247), .B(n199), .Z(n196) );
  XOR U313 ( .A(n248), .B(n242), .Z(n199) );
  XNOR U314 ( .A(n249), .B(n250), .Z(n248) );
  NOR U315 ( .A(n235), .B(n251), .Z(n250) );
  XNOR U316 ( .A(n243), .B(n252), .Z(n247) );
  NOR U317 ( .A(n215), .B(n253), .Z(n252) );
  ANDN U318 ( .A(n214), .B(n254), .Z(n243) );
  XOR U319 ( .A(n215), .B(n194), .Z(n214) );
  XOR U320 ( .A(n218), .B(g_input[80]), .Z(n246) );
  XNOR U321 ( .A(n255), .B(n242), .Z(n218) );
  XNOR U322 ( .A(n249), .B(n256), .Z(n242) );
  NOR U323 ( .A(n257), .B(n231), .Z(n256) );
  NOR U324 ( .A(n233), .B(n258), .Z(n249) );
  XNOR U325 ( .A(n225), .B(n194), .Z(n235) );
  XNOR U326 ( .A(n259), .B(n260), .Z(n194) );
  ANDN U327 ( .A(n261), .B(n262), .Z(n260) );
  IV U328 ( .A(n263), .Z(n202) );
  XNOR U329 ( .A(n259), .B(n264), .Z(n215) );
  NOR U330 ( .A(n265), .B(n266), .Z(n264) );
  ANDN U331 ( .A(n267), .B(n268), .Z(n259) );
  XNOR U332 ( .A(n269), .B(n201), .Z(n255) );
  OR U333 ( .A(n239), .B(n270), .Z(n201) );
  XOR U334 ( .A(n263), .B(n225), .Z(n239) );
  XOR U335 ( .A(n271), .B(n272), .Z(n263) );
  ANDN U336 ( .A(n273), .B(n266), .Z(n272) );
  OR U337 ( .A(n225), .B(n274), .Z(n269) );
  XOR U338 ( .A(n275), .B(n271), .Z(n225) );
  XOR U339 ( .A(n266), .B(n262), .Z(n267) );
  XNOR U340 ( .A(n277), .B(n278), .Z(n266) );
  XNOR U341 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U342 ( .B(n281), .A(n261), .Z(n279) );
  OR U343 ( .A(n262), .B(n281), .Z(n275) );
  XOR U344 ( .A(n282), .B(n283), .Z(n262) );
  XOR U345 ( .A(n284), .B(n285), .Z(n283) );
  XNOR U346 ( .A(n280), .B(n286), .Z(n285) );
  ANDN U347 ( .A(n273), .B(n265), .Z(n286) );
  OR U348 ( .A(n268), .B(n276), .Z(n280) );
  XNOR U349 ( .A(n287), .B(n273), .Z(n276) );
  XOR U350 ( .A(n261), .B(n265), .Z(n268) );
  IV U351 ( .A(n284), .Z(n265) );
  XNOR U352 ( .A(n288), .B(n289), .Z(n284) );
  XNOR U353 ( .A(n274), .B(n290), .Z(n289) );
  XNOR U354 ( .A(n291), .B(n292), .Z(n290) );
  ANDN U355 ( .A(n203), .B(n293), .Z(n291) );
  XNOR U356 ( .A(n294), .B(n295), .Z(n288) );
  XOR U357 ( .A(n296), .B(n224), .Z(n294) );
  XOR U358 ( .A(n278), .B(n273), .Z(n282) );
  XNOR U359 ( .A(n297), .B(n298), .Z(n273) );
  XNOR U360 ( .A(n299), .B(n300), .Z(n298) );
  ANDN U361 ( .A(n216), .B(n253), .Z(n299) );
  XNOR U362 ( .A(n301), .B(n296), .Z(n297) );
  XOR U363 ( .A(n302), .B(n303), .Z(n296) );
  XNOR U364 ( .A(n304), .B(n305), .Z(n302) );
  NANDN U365 ( .B(n251), .A(n236), .Z(n304) );
  XNOR U366 ( .A(n287), .B(n261), .Z(n278) );
  XNOR U367 ( .A(n306), .B(n307), .Z(n261) );
  XOR U368 ( .A(n203), .B(n308), .Z(n307) );
  XNOR U369 ( .A(n309), .B(n292), .Z(n308) );
  OR U370 ( .A(n240), .B(n270), .Z(n292) );
  XNOR U371 ( .A(n238), .B(n224), .Z(n240) );
  IV U372 ( .A(n293), .Z(n238) );
  ANDN U373 ( .A(n224), .B(n274), .Z(n309) );
  XNOR U374 ( .A(n310), .B(n301), .Z(n306) );
  XOR U375 ( .A(n303), .B(n293), .Z(n310) );
  IV U376 ( .A(n281), .Z(n287) );
  XOR U377 ( .A(n311), .B(n312), .Z(n281) );
  XOR U378 ( .A(n303), .B(n313), .Z(n312) );
  XNOR U379 ( .A(n314), .B(n300), .Z(n313) );
  OR U380 ( .A(n213), .B(n254), .Z(n300) );
  XNOR U381 ( .A(n253), .B(n245), .Z(n254) );
  XNOR U382 ( .A(n315), .B(n216), .Z(n213) );
  ANDN U383 ( .A(n316), .B(n193), .Z(n314) );
  XNOR U384 ( .A(n305), .B(n317), .Z(n303) );
  ANDN U385 ( .A(n318), .B(n230), .Z(n317) );
  OR U386 ( .A(n258), .B(n234), .Z(n305) );
  XOR U387 ( .A(n230), .B(n236), .Z(n234) );
  XNOR U388 ( .A(n193), .B(n224), .Z(n236) );
  XNOR U389 ( .A(n319), .B(n216), .Z(n224) );
  XNOR U390 ( .A(n320), .B(n321), .Z(n319) );
  XOR U391 ( .A(n293), .B(n216), .Z(n230) );
  XOR U392 ( .A(n322), .B(n323), .Z(n293) );
  XNOR U393 ( .A(n324), .B(n325), .Z(n322) );
  XOR U394 ( .A(n318), .B(n251), .Z(n258) );
  XOR U395 ( .A(n316), .B(n274), .Z(n251) );
  XOR U396 ( .A(n326), .B(n327), .Z(n274) );
  XNOR U397 ( .A(n328), .B(n203), .Z(n327) );
  XNOR U398 ( .A(n329), .B(n324), .Z(n326) );
  XOR U399 ( .A(g_input[52]), .B(state[52]), .Z(n324) );
  IV U400 ( .A(n257), .Z(n318) );
  XOR U401 ( .A(n253), .B(n203), .Z(n257) );
  XNOR U402 ( .A(n301), .B(n295), .Z(n311) );
  XNOR U403 ( .A(n315), .B(n316), .Z(n295) );
  IV U404 ( .A(n245), .Z(n316) );
  IV U405 ( .A(n193), .Z(n315) );
  XOR U406 ( .A(n330), .B(n323), .Z(n193) );
  XNOR U407 ( .A(n321), .B(n325), .Z(n330) );
  XOR U408 ( .A(n216), .B(n253), .Z(n301) );
  XNOR U409 ( .A(n320), .B(n331), .Z(n253) );
  XNOR U410 ( .A(n328), .B(n325), .Z(n331) );
  XOR U411 ( .A(n332), .B(n321), .Z(n328) );
  XOR U412 ( .A(g_input[49]), .B(state[49]), .Z(n321) );
  XNOR U413 ( .A(g_input[51]), .B(state[51]), .Z(n332) );
  XOR U414 ( .A(g_input[50]), .B(state[50]), .Z(n320) );
  XNOR U415 ( .A(n333), .B(n323), .Z(n216) );
  XOR U416 ( .A(g_input[53]), .B(state[53]), .Z(n323) );
  XNOR U417 ( .A(n329), .B(n325), .Z(n333) );
  XNOR U418 ( .A(n334), .B(n203), .Z(n325) );
  XOR U419 ( .A(g_input[48]), .B(state[48]), .Z(n203) );
  XNOR U420 ( .A(g_input[54]), .B(state[54]), .Z(n334) );
  XOR U421 ( .A(g_input[55]), .B(state[55]), .Z(n329) );
  XOR U422 ( .A(n335), .B(n336), .Z(o[7]) );
  XOR U423 ( .A(n337), .B(n338), .Z(n336) );
  XOR U424 ( .A(g_input[7]), .B(n339), .Z(n338) );
  XOR U425 ( .A(n340), .B(n341), .Z(n335) );
  XOR U426 ( .A(n342), .B(n343), .Z(o[79]) );
  XNOR U427 ( .A(n344), .B(n345), .Z(n343) );
  XNOR U428 ( .A(g_input[79]), .B(n346), .Z(n345) );
  XOR U429 ( .A(n347), .B(n348), .Z(n342) );
  XOR U430 ( .A(n349), .B(n350), .Z(o[78]) );
  XOR U431 ( .A(g_input[78]), .B(n351), .Z(n350) );
  XOR U432 ( .A(n352), .B(n353), .Z(n349) );
  XOR U433 ( .A(n354), .B(n355), .Z(o[77]) );
  XOR U434 ( .A(n356), .B(n357), .Z(n355) );
  XNOR U435 ( .A(g_input[77]), .B(n358), .Z(n357) );
  ANDN U436 ( .A(n359), .B(n360), .Z(n356) );
  XNOR U437 ( .A(n361), .B(n362), .Z(n354) );
  XOR U438 ( .A(n347), .B(n363), .Z(n361) );
  XNOR U439 ( .A(n364), .B(n365), .Z(n347) );
  XNOR U440 ( .A(n366), .B(n367), .Z(n364) );
  NANDN U441 ( .B(n368), .A(n369), .Z(n366) );
  XNOR U442 ( .A(n370), .B(n371), .Z(o[76]) );
  XOR U443 ( .A(n362), .B(g_input[76]), .Z(n370) );
  XOR U444 ( .A(n372), .B(n373), .Z(o[75]) );
  XOR U445 ( .A(n351), .B(n374), .Z(n373) );
  XNOR U446 ( .A(g_input[75]), .B(n346), .Z(n374) );
  XNOR U447 ( .A(n352), .B(n348), .Z(n372) );
  XNOR U448 ( .A(n375), .B(n376), .Z(n352) );
  XNOR U449 ( .A(n377), .B(n358), .Z(n375) );
  OR U450 ( .A(n378), .B(n379), .Z(n358) );
  OR U451 ( .A(n380), .B(n381), .Z(n377) );
  XOR U452 ( .A(n371), .B(g_input[74]), .Z(o[74]) );
  XNOR U453 ( .A(n382), .B(n353), .Z(n371) );
  XOR U454 ( .A(n383), .B(n384), .Z(o[73]) );
  XNOR U455 ( .A(g_input[73]), .B(n346), .Z(n384) );
  XNOR U456 ( .A(n385), .B(n376), .Z(n346) );
  XNOR U457 ( .A(n386), .B(n363), .Z(n376) );
  XNOR U458 ( .A(n387), .B(n388), .Z(n386) );
  AND U459 ( .A(n389), .B(n390), .Z(n388) );
  XOR U460 ( .A(n391), .B(n392), .Z(n385) );
  ANDN U461 ( .A(n393), .B(n394), .Z(n392) );
  XOR U462 ( .A(n382), .B(n344), .Z(n383) );
  XNOR U463 ( .A(n353), .B(n351), .Z(n344) );
  XOR U464 ( .A(n395), .B(n363), .Z(n351) );
  XNOR U465 ( .A(n387), .B(n396), .Z(n363) );
  ANDN U466 ( .A(n397), .B(n398), .Z(n396) );
  ANDN U467 ( .A(n399), .B(n400), .Z(n387) );
  XNOR U468 ( .A(n401), .B(n391), .Z(n395) );
  NANDN U469 ( .B(n402), .A(n403), .Z(n391) );
  OR U470 ( .A(n404), .B(n405), .Z(n401) );
  IV U471 ( .A(n348), .Z(n382) );
  XNOR U472 ( .A(n406), .B(n407), .Z(n348) );
  XNOR U473 ( .A(n408), .B(n409), .Z(n406) );
  NANDN U474 ( .B(n410), .A(n411), .Z(n408) );
  XNOR U475 ( .A(n412), .B(n362), .Z(o[72]) );
  XOR U476 ( .A(n413), .B(n365), .Z(n362) );
  XOR U477 ( .A(n414), .B(n407), .Z(n365) );
  XNOR U478 ( .A(n415), .B(n416), .Z(n414) );
  AND U479 ( .A(n417), .B(n389), .Z(n416) );
  XNOR U480 ( .A(n418), .B(n409), .Z(n413) );
  OR U481 ( .A(n378), .B(n419), .Z(n409) );
  XOR U482 ( .A(n411), .B(n380), .Z(n378) );
  NANDN U483 ( .B(n380), .A(n420), .Z(n418) );
  XNOR U484 ( .A(n353), .B(g_input[72]), .Z(n412) );
  XOR U485 ( .A(n421), .B(n407), .Z(n353) );
  XNOR U486 ( .A(n415), .B(n422), .Z(n407) );
  NOR U487 ( .A(n398), .B(n423), .Z(n422) );
  ANDN U488 ( .A(n399), .B(n424), .Z(n415) );
  XNOR U489 ( .A(n389), .B(n398), .Z(n399) );
  XOR U490 ( .A(n380), .B(n369), .Z(n398) );
  XNOR U491 ( .A(n425), .B(n426), .Z(n380) );
  NANDN U492 ( .B(n427), .A(n428), .Z(n425) );
  XOR U493 ( .A(n360), .B(n404), .Z(n389) );
  IV U494 ( .A(n411), .Z(n360) );
  XNOR U495 ( .A(n426), .B(n429), .Z(n411) );
  AND U496 ( .A(n430), .B(n431), .Z(n429) );
  NAND U497 ( .A(n432), .B(n433), .Z(n426) );
  XOR U498 ( .A(n430), .B(n434), .Z(n432) );
  XNOR U499 ( .A(n435), .B(n367), .Z(n421) );
  NANDN U500 ( .B(n436), .A(n403), .Z(n367) );
  XOR U501 ( .A(n404), .B(n394), .Z(n403) );
  IV U502 ( .A(n369), .Z(n394) );
  XNOR U503 ( .A(n437), .B(n438), .Z(n369) );
  AND U504 ( .A(n428), .B(n439), .Z(n438) );
  NANDN U505 ( .B(n404), .A(n440), .Z(n435) );
  XNOR U506 ( .A(n441), .B(n437), .Z(n404) );
  NANDN U507 ( .B(n442), .A(n433), .Z(n437) );
  XOR U508 ( .A(n431), .B(n428), .Z(n433) );
  XOR U509 ( .A(n443), .B(n444), .Z(n428) );
  XNOR U510 ( .A(n445), .B(n446), .Z(n443) );
  NANDN U511 ( .B(n447), .A(n430), .Z(n445) );
  NANDN U512 ( .B(n447), .A(n431), .Z(n441) );
  XNOR U513 ( .A(n448), .B(n449), .Z(n431) );
  XOR U514 ( .A(n439), .B(n450), .Z(n449) );
  XNOR U515 ( .A(n451), .B(n446), .Z(n450) );
  NANDN U516 ( .B(n442), .A(n452), .Z(n446) );
  XNOR U517 ( .A(n430), .B(n427), .Z(n452) );
  ANDN U518 ( .A(n439), .B(n427), .Z(n451) );
  XNOR U519 ( .A(n453), .B(n454), .Z(n439) );
  XNOR U520 ( .A(n455), .B(n456), .Z(n454) );
  ANDN U521 ( .A(n420), .B(n381), .Z(n455) );
  XOR U522 ( .A(n457), .B(n458), .Z(n453) );
  XNOR U523 ( .A(n444), .B(n427), .Z(n448) );
  IV U524 ( .A(n434), .Z(n427) );
  XNOR U525 ( .A(n459), .B(n460), .Z(n434) );
  XNOR U526 ( .A(n405), .B(n461), .Z(n460) );
  XNOR U527 ( .A(n462), .B(n463), .Z(n461) );
  ANDN U528 ( .A(n393), .B(n368), .Z(n462) );
  XOR U529 ( .A(n464), .B(n465), .Z(n459) );
  XOR U530 ( .A(n457), .B(n440), .Z(n464) );
  XNOR U531 ( .A(n466), .B(n467), .Z(n457) );
  XNOR U532 ( .A(n468), .B(n469), .Z(n466) );
  NAND U533 ( .A(n417), .B(n390), .Z(n468) );
  XOR U534 ( .A(n430), .B(n447), .Z(n444) );
  XNOR U535 ( .A(n470), .B(n471), .Z(n430) );
  XNOR U536 ( .A(n368), .B(n472), .Z(n471) );
  XNOR U537 ( .A(n473), .B(n463), .Z(n472) );
  OR U538 ( .A(n402), .B(n436), .Z(n463) );
  XOR U539 ( .A(n440), .B(n368), .Z(n436) );
  XNOR U540 ( .A(n474), .B(n393), .Z(n402) );
  ANDN U541 ( .A(n440), .B(n405), .Z(n473) );
  IV U542 ( .A(n474), .Z(n405) );
  XNOR U543 ( .A(n475), .B(n467), .Z(n470) );
  XOR U544 ( .A(n476), .B(n393), .Z(n475) );
  XOR U545 ( .A(n477), .B(n478), .Z(n447) );
  XNOR U546 ( .A(n476), .B(n479), .Z(n478) );
  XNOR U547 ( .A(n480), .B(n456), .Z(n479) );
  OR U548 ( .A(n379), .B(n419), .Z(n456) );
  XNOR U549 ( .A(n481), .B(n420), .Z(n419) );
  XNOR U550 ( .A(n359), .B(n482), .Z(n379) );
  IV U551 ( .A(n483), .Z(n359) );
  ANDN U552 ( .A(n481), .B(n483), .Z(n480) );
  IV U553 ( .A(n458), .Z(n476) );
  XOR U554 ( .A(n420), .B(n482), .Z(n458) );
  XOR U555 ( .A(n465), .B(n467), .Z(n477) );
  XOR U556 ( .A(n469), .B(n484), .Z(n467) );
  ANDN U557 ( .A(n397), .B(n423), .Z(n484) );
  OR U558 ( .A(n424), .B(n400), .Z(n469) );
  XNOR U559 ( .A(n390), .B(n397), .Z(n400) );
  XOR U560 ( .A(n393), .B(n482), .Z(n397) );
  IV U561 ( .A(n381), .Z(n482) );
  XOR U562 ( .A(n485), .B(n486), .Z(n393) );
  XNOR U563 ( .A(n483), .B(n474), .Z(n390) );
  XNOR U564 ( .A(n487), .B(n488), .Z(n474) );
  XNOR U565 ( .A(n489), .B(n381), .Z(n487) );
  XOR U566 ( .A(n490), .B(n491), .Z(n381) );
  XNOR U567 ( .A(n492), .B(n493), .Z(n490) );
  XOR U568 ( .A(n417), .B(n423), .Z(n424) );
  XNOR U569 ( .A(n420), .B(n494), .Z(n423) );
  XNOR U570 ( .A(n495), .B(n496), .Z(n420) );
  XNOR U571 ( .A(n488), .B(n493), .Z(n495) );
  XOR U572 ( .A(g_input[10]), .B(state[10]), .Z(n488) );
  XOR U573 ( .A(n440), .B(n481), .Z(n417) );
  IV U574 ( .A(n410), .Z(n481) );
  XNOR U575 ( .A(n497), .B(n498), .Z(n440) );
  XNOR U576 ( .A(n492), .B(n368), .Z(n498) );
  IV U577 ( .A(n494), .Z(n368) );
  XOR U578 ( .A(g_input[15]), .B(state[15]), .Z(n492) );
  XOR U579 ( .A(n486), .B(n496), .Z(n497) );
  XOR U580 ( .A(n499), .B(n489), .Z(n496) );
  XNOR U581 ( .A(g_input[11]), .B(state[11]), .Z(n499) );
  XNOR U582 ( .A(g_input[12]), .B(state[12]), .Z(n486) );
  XOR U583 ( .A(n410), .B(n483), .Z(n465) );
  XNOR U584 ( .A(n485), .B(n489), .Z(n483) );
  XNOR U585 ( .A(g_input[9]), .B(state[9]), .Z(n489) );
  XNOR U586 ( .A(n491), .B(n493), .Z(n485) );
  XNOR U587 ( .A(n500), .B(n494), .Z(n493) );
  XOR U588 ( .A(g_input[8]), .B(state[8]), .Z(n494) );
  XNOR U589 ( .A(g_input[14]), .B(state[14]), .Z(n500) );
  XOR U590 ( .A(g_input[13]), .B(state[13]), .Z(n491) );
  XOR U591 ( .A(n501), .B(n502), .Z(o[71]) );
  XNOR U592 ( .A(n503), .B(n504), .Z(n502) );
  XNOR U593 ( .A(g_input[71]), .B(n505), .Z(n504) );
  XOR U594 ( .A(n506), .B(n507), .Z(n501) );
  XOR U595 ( .A(n508), .B(n509), .Z(o[70]) );
  XNOR U596 ( .A(g_input[70]), .B(n510), .Z(n509) );
  XNOR U597 ( .A(n511), .B(n512), .Z(n508) );
  XNOR U598 ( .A(n513), .B(n514), .Z(o[6]) );
  XNOR U599 ( .A(n339), .B(g_input[6]), .Z(n513) );
  XOR U600 ( .A(n515), .B(n516), .Z(o[69]) );
  XOR U601 ( .A(n517), .B(n518), .Z(n516) );
  XOR U602 ( .A(g_input[69]), .B(n519), .Z(n518) );
  ANDN U603 ( .A(n520), .B(n521), .Z(n519) );
  XNOR U604 ( .A(n522), .B(n523), .Z(n515) );
  XOR U605 ( .A(n506), .B(n524), .Z(n522) );
  XNOR U606 ( .A(n525), .B(n526), .Z(n506) );
  XNOR U607 ( .A(n527), .B(n528), .Z(n525) );
  XNOR U608 ( .A(n531), .B(n532), .Z(o[68]) );
  XOR U609 ( .A(n523), .B(g_input[68]), .Z(n531) );
  XOR U610 ( .A(n533), .B(n534), .Z(o[67]) );
  XOR U611 ( .A(n535), .B(n536), .Z(n534) );
  XNOR U612 ( .A(g_input[67]), .B(n505), .Z(n536) );
  XOR U613 ( .A(n511), .B(n537), .Z(n533) );
  XNOR U614 ( .A(n538), .B(n539), .Z(n511) );
  XNOR U615 ( .A(n517), .B(n540), .Z(n538) );
  ANDN U616 ( .A(n541), .B(n542), .Z(n540) );
  ANDN U617 ( .A(n543), .B(n544), .Z(n517) );
  XOR U618 ( .A(n532), .B(g_input[66]), .Z(o[66]) );
  XNOR U619 ( .A(n510), .B(n503), .Z(n532) );
  IV U620 ( .A(n535), .Z(n503) );
  XOR U621 ( .A(n545), .B(n546), .Z(o[65]) );
  XNOR U622 ( .A(g_input[65]), .B(n505), .Z(n546) );
  XNOR U623 ( .A(n547), .B(n539), .Z(n505) );
  XNOR U624 ( .A(n548), .B(n524), .Z(n539) );
  XNOR U625 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U626 ( .B(n551), .A(n552), .Z(n549) );
  XNOR U627 ( .A(n553), .B(n554), .Z(n547) );
  NANDN U628 ( .B(n530), .A(n555), .Z(n553) );
  XOR U629 ( .A(n507), .B(n535), .Z(n545) );
  XOR U630 ( .A(n556), .B(n557), .Z(n535) );
  XNOR U631 ( .A(n558), .B(n559), .Z(n556) );
  ANDN U632 ( .A(n520), .B(n560), .Z(n559) );
  XOR U633 ( .A(n537), .B(n510), .Z(n507) );
  IV U634 ( .A(n512), .Z(n537) );
  XNOR U635 ( .A(n561), .B(n524), .Z(n512) );
  XOR U636 ( .A(n550), .B(n562), .Z(n524) );
  ANDN U637 ( .A(n563), .B(n564), .Z(n562) );
  NANDN U638 ( .B(n565), .A(n566), .Z(n550) );
  XNOR U639 ( .A(n567), .B(n554), .Z(n561) );
  NANDN U640 ( .B(n568), .A(n569), .Z(n554) );
  NANDN U641 ( .B(n570), .A(n571), .Z(n567) );
  XNOR U642 ( .A(n572), .B(n523), .Z(o[64]) );
  XOR U643 ( .A(n573), .B(n526), .Z(n523) );
  XOR U644 ( .A(n574), .B(n557), .Z(n526) );
  XNOR U645 ( .A(n575), .B(n576), .Z(n574) );
  ANDN U646 ( .A(n577), .B(n551), .Z(n576) );
  XNOR U647 ( .A(n558), .B(n578), .Z(n573) );
  AND U648 ( .A(n579), .B(n541), .Z(n578) );
  XOR U649 ( .A(n520), .B(n541), .Z(n543) );
  XOR U650 ( .A(n510), .B(g_input[64]), .Z(n572) );
  XNOR U651 ( .A(n581), .B(n557), .Z(n510) );
  XNOR U652 ( .A(n575), .B(n582), .Z(n557) );
  ANDN U653 ( .A(n583), .B(n564), .Z(n582) );
  XOR U654 ( .A(n551), .B(n564), .Z(n566) );
  XOR U655 ( .A(n541), .B(n530), .Z(n564) );
  XOR U656 ( .A(n585), .B(n586), .Z(n541) );
  ANDN U657 ( .A(n587), .B(n588), .Z(n586) );
  XOR U658 ( .A(n585), .B(n589), .Z(n520) );
  ANDN U659 ( .A(n590), .B(n591), .Z(n589) );
  AND U660 ( .A(n592), .B(n593), .Z(n585) );
  XNOR U661 ( .A(n527), .B(n594), .Z(n581) );
  ANDN U662 ( .A(n595), .B(n570), .Z(n594) );
  ANDN U663 ( .A(n569), .B(n596), .Z(n527) );
  XOR U664 ( .A(n570), .B(n530), .Z(n569) );
  XOR U665 ( .A(n597), .B(n598), .Z(n530) );
  AND U666 ( .A(n587), .B(n599), .Z(n598) );
  NAND U667 ( .A(n601), .B(n592), .Z(n597) );
  XOR U668 ( .A(n587), .B(n590), .Z(n592) );
  XOR U669 ( .A(n602), .B(n603), .Z(n587) );
  XNOR U670 ( .A(n604), .B(n605), .Z(n602) );
  OR U671 ( .A(n591), .B(n606), .Z(n604) );
  XOR U672 ( .A(n607), .B(n599), .Z(n601) );
  NANDN U673 ( .B(n606), .A(n590), .Z(n600) );
  XNOR U674 ( .A(n608), .B(n609), .Z(n590) );
  XNOR U675 ( .A(n603), .B(n610), .Z(n609) );
  XNOR U676 ( .A(n605), .B(n611), .Z(n610) );
  ANDN U677 ( .A(n599), .B(n588), .Z(n611) );
  NAND U678 ( .A(n612), .B(n593), .Z(n605) );
  XOR U679 ( .A(n588), .B(n591), .Z(n593) );
  XNOR U680 ( .A(n606), .B(n599), .Z(n612) );
  XOR U681 ( .A(n591), .B(n607), .Z(n603) );
  XOR U682 ( .A(n613), .B(n614), .Z(n591) );
  XNOR U683 ( .A(n529), .B(n615), .Z(n614) );
  XNOR U684 ( .A(n616), .B(n617), .Z(n615) );
  ANDN U685 ( .A(n571), .B(n618), .Z(n616) );
  XNOR U686 ( .A(n619), .B(n620), .Z(n613) );
  XNOR U687 ( .A(n621), .B(n622), .Z(n619) );
  XOR U688 ( .A(n588), .B(n599), .Z(n608) );
  XNOR U689 ( .A(n623), .B(n624), .Z(n599) );
  XNOR U690 ( .A(n625), .B(n626), .Z(n624) );
  ANDN U691 ( .A(n579), .B(n542), .Z(n625) );
  XOR U692 ( .A(n627), .B(n620), .Z(n623) );
  XOR U693 ( .A(n628), .B(n629), .Z(n588) );
  XOR U694 ( .A(n571), .B(n630), .Z(n629) );
  XNOR U695 ( .A(n631), .B(n617), .Z(n630) );
  OR U696 ( .A(n568), .B(n596), .Z(n617) );
  XNOR U697 ( .A(n595), .B(n632), .Z(n596) );
  IV U698 ( .A(n618), .Z(n595) );
  XNOR U699 ( .A(n555), .B(n571), .Z(n568) );
  ANDN U700 ( .A(n632), .B(n622), .Z(n631) );
  XOR U701 ( .A(n633), .B(n627), .Z(n628) );
  XOR U702 ( .A(n634), .B(n621), .Z(n627) );
  XNOR U703 ( .A(n635), .B(n636), .Z(n634) );
  NAND U704 ( .A(n577), .B(n552), .Z(n635) );
  XOR U705 ( .A(n637), .B(n618), .Z(n633) );
  IV U706 ( .A(n607), .Z(n606) );
  XNOR U707 ( .A(n638), .B(n639), .Z(n607) );
  XNOR U708 ( .A(n621), .B(n640), .Z(n639) );
  XNOR U709 ( .A(n641), .B(n626), .Z(n640) );
  OR U710 ( .A(n544), .B(n580), .Z(n626) );
  XNOR U711 ( .A(n642), .B(n579), .Z(n580) );
  ANDN U712 ( .A(n642), .B(n521), .Z(n641) );
  XOR U713 ( .A(n636), .B(n644), .Z(n621) );
  AND U714 ( .A(n583), .B(n563), .Z(n644) );
  OR U715 ( .A(n565), .B(n584), .Z(n636) );
  XNOR U716 ( .A(n577), .B(n583), .Z(n584) );
  XOR U717 ( .A(n579), .B(n632), .Z(n583) );
  XNOR U718 ( .A(n618), .B(n642), .Z(n577) );
  XOR U719 ( .A(n645), .B(n646), .Z(n618) );
  XNOR U720 ( .A(n647), .B(n529), .Z(n646) );
  IV U721 ( .A(n632), .Z(n529) );
  XOR U722 ( .A(n648), .B(n649), .Z(n645) );
  XNOR U723 ( .A(n563), .B(n552), .Z(n565) );
  XNOR U724 ( .A(n521), .B(n571), .Z(n552) );
  XOR U725 ( .A(n650), .B(n651), .Z(n571) );
  XNOR U726 ( .A(n652), .B(n542), .Z(n650) );
  XNOR U727 ( .A(n622), .B(n643), .Z(n563) );
  IV U728 ( .A(n555), .Z(n622) );
  XNOR U729 ( .A(n653), .B(n648), .Z(n555) );
  XOR U730 ( .A(g_input[100]), .B(state[100]), .Z(n648) );
  XOR U731 ( .A(n637), .B(n620), .Z(n638) );
  XNOR U732 ( .A(n579), .B(n643), .Z(n620) );
  IV U733 ( .A(n542), .Z(n643) );
  XOR U734 ( .A(n654), .B(n655), .Z(n542) );
  XOR U735 ( .A(n647), .B(n656), .Z(n654) );
  XOR U736 ( .A(g_input[103]), .B(state[103]), .Z(n647) );
  XOR U737 ( .A(n657), .B(n649), .Z(n579) );
  XNOR U738 ( .A(n658), .B(n652), .Z(n649) );
  XNOR U739 ( .A(g_input[99]), .B(state[99]), .Z(n658) );
  XOR U740 ( .A(n651), .B(n659), .Z(n657) );
  XNOR U741 ( .A(g_input[98]), .B(state[98]), .Z(n651) );
  XOR U742 ( .A(n560), .B(n521), .Z(n637) );
  XNOR U743 ( .A(n653), .B(n652), .Z(n521) );
  XNOR U744 ( .A(g_input[97]), .B(state[97]), .Z(n652) );
  XNOR U745 ( .A(n655), .B(n659), .Z(n653) );
  IV U746 ( .A(n642), .Z(n560) );
  IV U747 ( .A(n656), .Z(n659) );
  XOR U748 ( .A(n660), .B(n632), .Z(n656) );
  XOR U749 ( .A(g_input[96]), .B(state[96]), .Z(n632) );
  XNOR U750 ( .A(g_input[102]), .B(state[102]), .Z(n660) );
  XOR U751 ( .A(g_input[101]), .B(state[101]), .Z(n655) );
  XOR U752 ( .A(n661), .B(n662), .Z(o[63]) );
  XOR U753 ( .A(n663), .B(n664), .Z(n662) );
  XOR U754 ( .A(n666), .B(n667), .Z(n661) );
  XNOR U755 ( .A(n668), .B(n669), .Z(o[62]) );
  XNOR U756 ( .A(n665), .B(g_input[62]), .Z(n668) );
  XOR U757 ( .A(n670), .B(n671), .Z(o[61]) );
  XOR U758 ( .A(n672), .B(n673), .Z(n671) );
  XNOR U759 ( .A(g_input[61]), .B(n674), .Z(n673) );
  NOR U760 ( .A(n675), .B(n676), .Z(n672) );
  XNOR U761 ( .A(n677), .B(n678), .Z(n670) );
  XOR U762 ( .A(n666), .B(n679), .Z(n677) );
  XNOR U763 ( .A(n680), .B(n681), .Z(n666) );
  XNOR U764 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U765 ( .B(n684), .A(n685), .Z(n682) );
  XNOR U766 ( .A(n686), .B(n687), .Z(o[60]) );
  XOR U767 ( .A(n678), .B(g_input[60]), .Z(n686) );
  XOR U768 ( .A(n688), .B(n689), .Z(o[5]) );
  XOR U769 ( .A(n690), .B(n691), .Z(n689) );
  XNOR U770 ( .A(g_input[5]), .B(n692), .Z(n691) );
  NOR U771 ( .A(n693), .B(n694), .Z(n690) );
  XNOR U772 ( .A(n695), .B(n696), .Z(n688) );
  XOR U773 ( .A(n340), .B(n697), .Z(n695) );
  XNOR U774 ( .A(n698), .B(n699), .Z(n340) );
  XNOR U775 ( .A(n700), .B(n701), .Z(n698) );
  NANDN U776 ( .B(n702), .A(n703), .Z(n700) );
  XOR U777 ( .A(n704), .B(n705), .Z(o[59]) );
  XOR U778 ( .A(n663), .B(n706), .Z(n705) );
  XNOR U779 ( .A(g_input[59]), .B(n707), .Z(n706) );
  XNOR U780 ( .A(n669), .B(n667), .Z(n704) );
  XNOR U781 ( .A(n708), .B(n709), .Z(n669) );
  XNOR U782 ( .A(n710), .B(n674), .Z(n708) );
  NANDN U783 ( .B(n711), .A(n712), .Z(n674) );
  NANDN U784 ( .B(n713), .A(n714), .Z(n710) );
  XOR U785 ( .A(n687), .B(g_input[58]), .Z(o[58]) );
  XOR U786 ( .A(n715), .B(n716), .Z(n687) );
  XOR U787 ( .A(n717), .B(n718), .Z(o[57]) );
  XOR U788 ( .A(g_input[57]), .B(n665), .Z(n718) );
  XOR U789 ( .A(n707), .B(n716), .Z(n665) );
  XNOR U790 ( .A(n719), .B(n679), .Z(n707) );
  XOR U791 ( .A(n720), .B(n721), .Z(n719) );
  ANDN U792 ( .A(n722), .B(n723), .Z(n721) );
  XNOR U793 ( .A(n715), .B(n663), .Z(n717) );
  XOR U794 ( .A(n724), .B(n709), .Z(n663) );
  XNOR U795 ( .A(n725), .B(n679), .Z(n709) );
  XNOR U796 ( .A(n726), .B(n727), .Z(n679) );
  NOR U797 ( .A(n728), .B(n729), .Z(n727) );
  XOR U798 ( .A(n730), .B(n726), .Z(n725) );
  NOR U799 ( .A(n731), .B(n732), .Z(n726) );
  NANDN U800 ( .B(n733), .A(n734), .Z(n730) );
  XOR U801 ( .A(n720), .B(n735), .Z(n724) );
  ANDN U802 ( .A(n736), .B(n684), .Z(n735) );
  OR U803 ( .A(n737), .B(n738), .Z(n720) );
  IV U804 ( .A(n667), .Z(n715) );
  XNOR U805 ( .A(n739), .B(n740), .Z(n667) );
  XNOR U806 ( .A(n741), .B(n742), .Z(n739) );
  NOR U807 ( .A(n743), .B(n676), .Z(n742) );
  XNOR U808 ( .A(n744), .B(n678), .Z(o[56]) );
  XOR U809 ( .A(n745), .B(n681), .Z(n678) );
  XOR U810 ( .A(n746), .B(n740), .Z(n681) );
  XNOR U811 ( .A(n747), .B(n748), .Z(n746) );
  NOR U812 ( .A(n733), .B(n749), .Z(n748) );
  XNOR U813 ( .A(n741), .B(n750), .Z(n745) );
  NOR U814 ( .A(n713), .B(n751), .Z(n750) );
  ANDN U815 ( .A(n712), .B(n752), .Z(n741) );
  XOR U816 ( .A(n713), .B(n676), .Z(n712) );
  XOR U817 ( .A(n716), .B(g_input[56]), .Z(n744) );
  XNOR U818 ( .A(n753), .B(n740), .Z(n716) );
  XNOR U819 ( .A(n747), .B(n754), .Z(n740) );
  NOR U820 ( .A(n755), .B(n729), .Z(n754) );
  NOR U821 ( .A(n731), .B(n756), .Z(n747) );
  XNOR U822 ( .A(n723), .B(n676), .Z(n733) );
  XNOR U823 ( .A(n757), .B(n758), .Z(n676) );
  ANDN U824 ( .A(n759), .B(n760), .Z(n758) );
  IV U825 ( .A(n761), .Z(n684) );
  XNOR U826 ( .A(n757), .B(n762), .Z(n713) );
  NOR U827 ( .A(n763), .B(n764), .Z(n762) );
  ANDN U828 ( .A(n765), .B(n766), .Z(n757) );
  XNOR U829 ( .A(n767), .B(n683), .Z(n753) );
  OR U830 ( .A(n737), .B(n768), .Z(n683) );
  XOR U831 ( .A(n761), .B(n723), .Z(n737) );
  XOR U832 ( .A(n769), .B(n770), .Z(n761) );
  ANDN U833 ( .A(n771), .B(n764), .Z(n770) );
  OR U834 ( .A(n723), .B(n772), .Z(n767) );
  XOR U835 ( .A(n773), .B(n769), .Z(n723) );
  XOR U836 ( .A(n764), .B(n760), .Z(n765) );
  XNOR U837 ( .A(n775), .B(n776), .Z(n764) );
  XNOR U838 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U839 ( .B(n779), .A(n759), .Z(n777) );
  OR U840 ( .A(n760), .B(n779), .Z(n773) );
  XOR U841 ( .A(n780), .B(n781), .Z(n760) );
  XOR U842 ( .A(n782), .B(n783), .Z(n781) );
  XNOR U843 ( .A(n778), .B(n784), .Z(n783) );
  ANDN U844 ( .A(n771), .B(n763), .Z(n784) );
  OR U845 ( .A(n766), .B(n774), .Z(n778) );
  XNOR U846 ( .A(n785), .B(n771), .Z(n774) );
  XOR U847 ( .A(n759), .B(n763), .Z(n766) );
  IV U848 ( .A(n782), .Z(n763) );
  XNOR U849 ( .A(n786), .B(n787), .Z(n782) );
  XNOR U850 ( .A(n772), .B(n788), .Z(n787) );
  XNOR U851 ( .A(n789), .B(n790), .Z(n788) );
  ANDN U852 ( .A(n685), .B(n791), .Z(n789) );
  XNOR U853 ( .A(n792), .B(n793), .Z(n786) );
  XOR U854 ( .A(n794), .B(n722), .Z(n792) );
  XOR U855 ( .A(n776), .B(n771), .Z(n780) );
  XNOR U856 ( .A(n795), .B(n796), .Z(n771) );
  XNOR U857 ( .A(n797), .B(n798), .Z(n796) );
  ANDN U858 ( .A(n714), .B(n751), .Z(n797) );
  XNOR U859 ( .A(n799), .B(n794), .Z(n795) );
  XOR U860 ( .A(n800), .B(n801), .Z(n794) );
  XNOR U861 ( .A(n802), .B(n803), .Z(n800) );
  NANDN U862 ( .B(n749), .A(n734), .Z(n802) );
  XNOR U863 ( .A(n785), .B(n759), .Z(n776) );
  XNOR U864 ( .A(n804), .B(n805), .Z(n759) );
  XOR U865 ( .A(n685), .B(n806), .Z(n805) );
  XNOR U866 ( .A(n807), .B(n790), .Z(n806) );
  OR U867 ( .A(n738), .B(n768), .Z(n790) );
  XNOR U868 ( .A(n736), .B(n722), .Z(n738) );
  IV U869 ( .A(n791), .Z(n736) );
  ANDN U870 ( .A(n722), .B(n772), .Z(n807) );
  XNOR U871 ( .A(n808), .B(n799), .Z(n804) );
  XOR U872 ( .A(n801), .B(n791), .Z(n808) );
  IV U873 ( .A(n779), .Z(n785) );
  XOR U874 ( .A(n809), .B(n810), .Z(n779) );
  XOR U875 ( .A(n801), .B(n811), .Z(n810) );
  XNOR U876 ( .A(n812), .B(n798), .Z(n811) );
  OR U877 ( .A(n711), .B(n752), .Z(n798) );
  XNOR U878 ( .A(n751), .B(n743), .Z(n752) );
  XNOR U879 ( .A(n813), .B(n714), .Z(n711) );
  ANDN U880 ( .A(n814), .B(n675), .Z(n812) );
  XNOR U881 ( .A(n803), .B(n815), .Z(n801) );
  ANDN U882 ( .A(n816), .B(n728), .Z(n815) );
  OR U883 ( .A(n756), .B(n732), .Z(n803) );
  XOR U884 ( .A(n728), .B(n734), .Z(n732) );
  XNOR U885 ( .A(n675), .B(n722), .Z(n734) );
  XNOR U886 ( .A(n817), .B(n714), .Z(n722) );
  XNOR U887 ( .A(n818), .B(n819), .Z(n817) );
  XOR U888 ( .A(n791), .B(n714), .Z(n728) );
  XOR U889 ( .A(n820), .B(n821), .Z(n791) );
  XNOR U890 ( .A(n822), .B(n823), .Z(n820) );
  XOR U891 ( .A(n816), .B(n749), .Z(n756) );
  XOR U892 ( .A(n814), .B(n772), .Z(n749) );
  XOR U893 ( .A(n824), .B(n825), .Z(n772) );
  XNOR U894 ( .A(n826), .B(n685), .Z(n825) );
  XNOR U895 ( .A(n827), .B(n822), .Z(n824) );
  XOR U896 ( .A(g_input[60]), .B(state[60]), .Z(n822) );
  IV U897 ( .A(n755), .Z(n816) );
  XOR U898 ( .A(n751), .B(n685), .Z(n755) );
  XNOR U899 ( .A(n799), .B(n793), .Z(n809) );
  XNOR U900 ( .A(n813), .B(n814), .Z(n793) );
  IV U901 ( .A(n743), .Z(n814) );
  IV U902 ( .A(n675), .Z(n813) );
  XOR U903 ( .A(n828), .B(n821), .Z(n675) );
  XNOR U904 ( .A(n819), .B(n823), .Z(n828) );
  XOR U905 ( .A(n714), .B(n751), .Z(n799) );
  XNOR U906 ( .A(n818), .B(n829), .Z(n751) );
  XNOR U907 ( .A(n826), .B(n823), .Z(n829) );
  XOR U908 ( .A(n830), .B(n819), .Z(n826) );
  XOR U909 ( .A(g_input[57]), .B(state[57]), .Z(n819) );
  XNOR U910 ( .A(g_input[59]), .B(state[59]), .Z(n830) );
  XOR U911 ( .A(g_input[58]), .B(state[58]), .Z(n818) );
  XNOR U912 ( .A(n831), .B(n821), .Z(n714) );
  XOR U913 ( .A(g_input[61]), .B(state[61]), .Z(n821) );
  XNOR U914 ( .A(n827), .B(n823), .Z(n831) );
  XNOR U915 ( .A(n832), .B(n685), .Z(n823) );
  XOR U916 ( .A(g_input[56]), .B(state[56]), .Z(n685) );
  XNOR U917 ( .A(g_input[62]), .B(state[62]), .Z(n832) );
  XOR U918 ( .A(g_input[63]), .B(state[63]), .Z(n827) );
  XOR U919 ( .A(n833), .B(n834), .Z(o[55]) );
  XOR U920 ( .A(n835), .B(n836), .Z(n834) );
  XOR U921 ( .A(n838), .B(n839), .Z(n833) );
  XNOR U922 ( .A(n840), .B(n841), .Z(o[54]) );
  XNOR U923 ( .A(n837), .B(g_input[54]), .Z(n840) );
  XOR U924 ( .A(n842), .B(n843), .Z(o[53]) );
  XOR U925 ( .A(n844), .B(n845), .Z(n843) );
  XNOR U926 ( .A(g_input[53]), .B(n846), .Z(n845) );
  NOR U927 ( .A(n847), .B(n848), .Z(n844) );
  XNOR U928 ( .A(n849), .B(n850), .Z(n842) );
  XOR U929 ( .A(n838), .B(n851), .Z(n849) );
  XNOR U930 ( .A(n852), .B(n853), .Z(n838) );
  XNOR U931 ( .A(n854), .B(n855), .Z(n852) );
  NANDN U932 ( .B(n856), .A(n857), .Z(n854) );
  XNOR U933 ( .A(n858), .B(n859), .Z(o[52]) );
  XOR U934 ( .A(n850), .B(g_input[52]), .Z(n858) );
  XOR U935 ( .A(n860), .B(n861), .Z(o[51]) );
  XOR U936 ( .A(n835), .B(n862), .Z(n861) );
  XNOR U937 ( .A(g_input[51]), .B(n863), .Z(n862) );
  XNOR U938 ( .A(n841), .B(n839), .Z(n860) );
  XNOR U939 ( .A(n864), .B(n865), .Z(n841) );
  XNOR U940 ( .A(n866), .B(n846), .Z(n864) );
  NANDN U941 ( .B(n867), .A(n868), .Z(n846) );
  NANDN U942 ( .B(n869), .A(n870), .Z(n866) );
  XOR U943 ( .A(n859), .B(g_input[50]), .Z(o[50]) );
  XOR U944 ( .A(n871), .B(n872), .Z(n859) );
  XNOR U945 ( .A(n873), .B(n874), .Z(o[4]) );
  XOR U946 ( .A(n696), .B(g_input[4]), .Z(n873) );
  XOR U947 ( .A(n875), .B(n876), .Z(o[49]) );
  XOR U948 ( .A(g_input[49]), .B(n837), .Z(n876) );
  XOR U949 ( .A(n863), .B(n872), .Z(n837) );
  XNOR U950 ( .A(n877), .B(n851), .Z(n863) );
  XOR U951 ( .A(n878), .B(n879), .Z(n877) );
  ANDN U952 ( .A(n880), .B(n881), .Z(n879) );
  XNOR U953 ( .A(n871), .B(n835), .Z(n875) );
  XOR U954 ( .A(n882), .B(n865), .Z(n835) );
  XNOR U955 ( .A(n883), .B(n851), .Z(n865) );
  XNOR U956 ( .A(n884), .B(n885), .Z(n851) );
  NOR U957 ( .A(n886), .B(n887), .Z(n885) );
  XOR U958 ( .A(n888), .B(n884), .Z(n883) );
  NOR U959 ( .A(n889), .B(n890), .Z(n884) );
  NANDN U960 ( .B(n891), .A(n892), .Z(n888) );
  XOR U961 ( .A(n878), .B(n893), .Z(n882) );
  ANDN U962 ( .A(n894), .B(n856), .Z(n893) );
  OR U963 ( .A(n895), .B(n896), .Z(n878) );
  IV U964 ( .A(n839), .Z(n871) );
  XNOR U965 ( .A(n897), .B(n898), .Z(n839) );
  XNOR U966 ( .A(n899), .B(n900), .Z(n897) );
  NOR U967 ( .A(n901), .B(n848), .Z(n900) );
  XNOR U968 ( .A(n902), .B(n850), .Z(o[48]) );
  XOR U969 ( .A(n903), .B(n853), .Z(n850) );
  XOR U970 ( .A(n904), .B(n898), .Z(n853) );
  XNOR U971 ( .A(n905), .B(n906), .Z(n904) );
  NOR U972 ( .A(n891), .B(n907), .Z(n906) );
  XNOR U973 ( .A(n899), .B(n908), .Z(n903) );
  NOR U974 ( .A(n869), .B(n909), .Z(n908) );
  ANDN U975 ( .A(n868), .B(n910), .Z(n899) );
  XOR U976 ( .A(n869), .B(n848), .Z(n868) );
  XOR U977 ( .A(n872), .B(g_input[48]), .Z(n902) );
  XNOR U978 ( .A(n911), .B(n898), .Z(n872) );
  XNOR U979 ( .A(n905), .B(n912), .Z(n898) );
  NOR U980 ( .A(n913), .B(n887), .Z(n912) );
  NOR U981 ( .A(n889), .B(n914), .Z(n905) );
  XNOR U982 ( .A(n881), .B(n848), .Z(n891) );
  XNOR U983 ( .A(n915), .B(n916), .Z(n848) );
  ANDN U984 ( .A(n917), .B(n918), .Z(n916) );
  IV U985 ( .A(n919), .Z(n856) );
  XNOR U986 ( .A(n915), .B(n920), .Z(n869) );
  NOR U987 ( .A(n921), .B(n922), .Z(n920) );
  ANDN U988 ( .A(n923), .B(n924), .Z(n915) );
  XNOR U989 ( .A(n925), .B(n855), .Z(n911) );
  OR U990 ( .A(n895), .B(n926), .Z(n855) );
  XOR U991 ( .A(n919), .B(n881), .Z(n895) );
  XOR U992 ( .A(n927), .B(n928), .Z(n919) );
  ANDN U993 ( .A(n929), .B(n922), .Z(n928) );
  OR U994 ( .A(n881), .B(n930), .Z(n925) );
  XOR U995 ( .A(n931), .B(n927), .Z(n881) );
  XOR U996 ( .A(n922), .B(n918), .Z(n923) );
  XNOR U997 ( .A(n933), .B(n934), .Z(n922) );
  XNOR U998 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U999 ( .B(n937), .A(n917), .Z(n935) );
  OR U1000 ( .A(n918), .B(n937), .Z(n931) );
  XOR U1001 ( .A(n938), .B(n939), .Z(n918) );
  XOR U1002 ( .A(n940), .B(n941), .Z(n939) );
  XNOR U1003 ( .A(n936), .B(n942), .Z(n941) );
  ANDN U1004 ( .A(n929), .B(n921), .Z(n942) );
  OR U1005 ( .A(n924), .B(n932), .Z(n936) );
  XNOR U1006 ( .A(n943), .B(n929), .Z(n932) );
  XOR U1007 ( .A(n917), .B(n921), .Z(n924) );
  IV U1008 ( .A(n940), .Z(n921) );
  XNOR U1009 ( .A(n944), .B(n945), .Z(n940) );
  XNOR U1010 ( .A(n930), .B(n946), .Z(n945) );
  XNOR U1011 ( .A(n947), .B(n948), .Z(n946) );
  ANDN U1012 ( .A(n857), .B(n949), .Z(n947) );
  XNOR U1013 ( .A(n950), .B(n951), .Z(n944) );
  XOR U1014 ( .A(n952), .B(n880), .Z(n950) );
  XOR U1015 ( .A(n934), .B(n929), .Z(n938) );
  XNOR U1016 ( .A(n953), .B(n954), .Z(n929) );
  XNOR U1017 ( .A(n955), .B(n956), .Z(n954) );
  ANDN U1018 ( .A(n870), .B(n909), .Z(n955) );
  XNOR U1019 ( .A(n957), .B(n952), .Z(n953) );
  XOR U1020 ( .A(n958), .B(n959), .Z(n952) );
  XNOR U1021 ( .A(n960), .B(n961), .Z(n958) );
  NANDN U1022 ( .B(n907), .A(n892), .Z(n960) );
  XNOR U1023 ( .A(n943), .B(n917), .Z(n934) );
  XNOR U1024 ( .A(n962), .B(n963), .Z(n917) );
  XOR U1025 ( .A(n857), .B(n964), .Z(n963) );
  XNOR U1026 ( .A(n965), .B(n948), .Z(n964) );
  OR U1027 ( .A(n896), .B(n926), .Z(n948) );
  XNOR U1028 ( .A(n894), .B(n880), .Z(n896) );
  IV U1029 ( .A(n949), .Z(n894) );
  ANDN U1030 ( .A(n880), .B(n930), .Z(n965) );
  XNOR U1031 ( .A(n966), .B(n957), .Z(n962) );
  XOR U1032 ( .A(n959), .B(n949), .Z(n966) );
  IV U1033 ( .A(n937), .Z(n943) );
  XOR U1034 ( .A(n967), .B(n968), .Z(n937) );
  XOR U1035 ( .A(n959), .B(n969), .Z(n968) );
  XNOR U1036 ( .A(n970), .B(n956), .Z(n969) );
  OR U1037 ( .A(n867), .B(n910), .Z(n956) );
  XNOR U1038 ( .A(n909), .B(n901), .Z(n910) );
  XNOR U1039 ( .A(n971), .B(n870), .Z(n867) );
  ANDN U1040 ( .A(n972), .B(n847), .Z(n970) );
  XNOR U1041 ( .A(n961), .B(n973), .Z(n959) );
  ANDN U1042 ( .A(n974), .B(n886), .Z(n973) );
  OR U1043 ( .A(n914), .B(n890), .Z(n961) );
  XOR U1044 ( .A(n886), .B(n892), .Z(n890) );
  XNOR U1045 ( .A(n847), .B(n880), .Z(n892) );
  XNOR U1046 ( .A(n975), .B(n870), .Z(n880) );
  XNOR U1047 ( .A(n976), .B(n977), .Z(n975) );
  XOR U1048 ( .A(n949), .B(n870), .Z(n886) );
  XOR U1049 ( .A(n978), .B(n979), .Z(n949) );
  XNOR U1050 ( .A(n980), .B(n981), .Z(n978) );
  XOR U1051 ( .A(n974), .B(n907), .Z(n914) );
  XOR U1052 ( .A(n972), .B(n930), .Z(n907) );
  XOR U1053 ( .A(n982), .B(n983), .Z(n930) );
  XNOR U1054 ( .A(n984), .B(n857), .Z(n983) );
  XNOR U1055 ( .A(n985), .B(n980), .Z(n982) );
  XOR U1056 ( .A(g_input[20]), .B(state[20]), .Z(n980) );
  IV U1057 ( .A(n913), .Z(n974) );
  XOR U1058 ( .A(n909), .B(n857), .Z(n913) );
  XNOR U1059 ( .A(n957), .B(n951), .Z(n967) );
  XNOR U1060 ( .A(n971), .B(n972), .Z(n951) );
  IV U1061 ( .A(n901), .Z(n972) );
  IV U1062 ( .A(n847), .Z(n971) );
  XOR U1063 ( .A(n986), .B(n979), .Z(n847) );
  XNOR U1064 ( .A(n977), .B(n981), .Z(n986) );
  XOR U1065 ( .A(n870), .B(n909), .Z(n957) );
  XNOR U1066 ( .A(n976), .B(n987), .Z(n909) );
  XNOR U1067 ( .A(n984), .B(n981), .Z(n987) );
  XOR U1068 ( .A(n988), .B(n977), .Z(n984) );
  XOR U1069 ( .A(g_input[17]), .B(state[17]), .Z(n977) );
  XNOR U1070 ( .A(g_input[19]), .B(state[19]), .Z(n988) );
  XOR U1071 ( .A(g_input[18]), .B(state[18]), .Z(n976) );
  XNOR U1072 ( .A(n989), .B(n979), .Z(n870) );
  XOR U1073 ( .A(g_input[21]), .B(state[21]), .Z(n979) );
  XNOR U1074 ( .A(n985), .B(n981), .Z(n989) );
  XNOR U1075 ( .A(n990), .B(n857), .Z(n981) );
  XOR U1076 ( .A(g_input[16]), .B(state[16]), .Z(n857) );
  XNOR U1077 ( .A(g_input[22]), .B(state[22]), .Z(n990) );
  XOR U1078 ( .A(g_input[23]), .B(state[23]), .Z(n985) );
  XOR U1079 ( .A(n991), .B(n992), .Z(o[47]) );
  XOR U1080 ( .A(n993), .B(n994), .Z(n992) );
  XOR U1081 ( .A(g_input[47]), .B(n995), .Z(n994) );
  XOR U1082 ( .A(n996), .B(n997), .Z(n991) );
  XNOR U1083 ( .A(n998), .B(n999), .Z(o[46]) );
  XNOR U1084 ( .A(n995), .B(g_input[46]), .Z(n998) );
  XOR U1085 ( .A(n1000), .B(n1001), .Z(o[45]) );
  XOR U1086 ( .A(n1002), .B(n1003), .Z(n1001) );
  XNOR U1087 ( .A(g_input[45]), .B(n1004), .Z(n1003) );
  NOR U1088 ( .A(n1005), .B(n1006), .Z(n1002) );
  XNOR U1089 ( .A(n1007), .B(n1008), .Z(n1000) );
  XOR U1090 ( .A(n996), .B(n1009), .Z(n1007) );
  XNOR U1091 ( .A(n1010), .B(n1011), .Z(n996) );
  XNOR U1092 ( .A(n1012), .B(n1013), .Z(n1010) );
  NANDN U1093 ( .B(n1014), .A(n1015), .Z(n1012) );
  XNOR U1094 ( .A(n1016), .B(n1017), .Z(o[44]) );
  XOR U1095 ( .A(n1008), .B(g_input[44]), .Z(n1016) );
  XOR U1096 ( .A(n1018), .B(n1019), .Z(o[43]) );
  XOR U1097 ( .A(n993), .B(n1020), .Z(n1019) );
  XNOR U1098 ( .A(g_input[43]), .B(n1021), .Z(n1020) );
  XNOR U1099 ( .A(n999), .B(n997), .Z(n1018) );
  XNOR U1100 ( .A(n1022), .B(n1023), .Z(n999) );
  XNOR U1101 ( .A(n1024), .B(n1004), .Z(n1022) );
  NANDN U1102 ( .B(n1025), .A(n1026), .Z(n1004) );
  NANDN U1103 ( .B(n1027), .A(n1028), .Z(n1024) );
  XOR U1104 ( .A(n1017), .B(g_input[42]), .Z(o[42]) );
  XOR U1105 ( .A(n1029), .B(n1030), .Z(n1017) );
  XOR U1106 ( .A(n1031), .B(n1032), .Z(o[41]) );
  XOR U1107 ( .A(g_input[41]), .B(n995), .Z(n1032) );
  XOR U1108 ( .A(n1021), .B(n1030), .Z(n995) );
  XNOR U1109 ( .A(n1033), .B(n1009), .Z(n1021) );
  XOR U1110 ( .A(n1034), .B(n1035), .Z(n1033) );
  ANDN U1111 ( .A(n1036), .B(n1037), .Z(n1035) );
  XNOR U1112 ( .A(n1029), .B(n993), .Z(n1031) );
  XOR U1113 ( .A(n1038), .B(n1023), .Z(n993) );
  XNOR U1114 ( .A(n1039), .B(n1009), .Z(n1023) );
  XNOR U1115 ( .A(n1040), .B(n1041), .Z(n1009) );
  NOR U1116 ( .A(n1042), .B(n1043), .Z(n1041) );
  XOR U1117 ( .A(n1044), .B(n1040), .Z(n1039) );
  NOR U1118 ( .A(n1045), .B(n1046), .Z(n1040) );
  NANDN U1119 ( .B(n1047), .A(n1048), .Z(n1044) );
  XOR U1120 ( .A(n1034), .B(n1049), .Z(n1038) );
  ANDN U1121 ( .A(n1050), .B(n1014), .Z(n1049) );
  OR U1122 ( .A(n1051), .B(n1052), .Z(n1034) );
  IV U1123 ( .A(n997), .Z(n1029) );
  XNOR U1124 ( .A(n1053), .B(n1054), .Z(n997) );
  XNOR U1125 ( .A(n1055), .B(n1056), .Z(n1053) );
  NOR U1126 ( .A(n1057), .B(n1006), .Z(n1056) );
  XNOR U1127 ( .A(n1058), .B(n1008), .Z(o[40]) );
  XOR U1128 ( .A(n1059), .B(n1011), .Z(n1008) );
  XOR U1129 ( .A(n1060), .B(n1054), .Z(n1011) );
  XNOR U1130 ( .A(n1061), .B(n1062), .Z(n1060) );
  NOR U1131 ( .A(n1047), .B(n1063), .Z(n1062) );
  XNOR U1132 ( .A(n1055), .B(n1064), .Z(n1059) );
  NOR U1133 ( .A(n1027), .B(n1065), .Z(n1064) );
  ANDN U1134 ( .A(n1026), .B(n1066), .Z(n1055) );
  XOR U1135 ( .A(n1027), .B(n1006), .Z(n1026) );
  XOR U1136 ( .A(n1030), .B(g_input[40]), .Z(n1058) );
  XNOR U1137 ( .A(n1067), .B(n1054), .Z(n1030) );
  XNOR U1138 ( .A(n1061), .B(n1068), .Z(n1054) );
  NOR U1139 ( .A(n1069), .B(n1043), .Z(n1068) );
  NOR U1140 ( .A(n1045), .B(n1070), .Z(n1061) );
  XNOR U1141 ( .A(n1037), .B(n1006), .Z(n1047) );
  XNOR U1142 ( .A(n1071), .B(n1072), .Z(n1006) );
  ANDN U1143 ( .A(n1073), .B(n1074), .Z(n1072) );
  IV U1144 ( .A(n1075), .Z(n1014) );
  XNOR U1145 ( .A(n1071), .B(n1076), .Z(n1027) );
  NOR U1146 ( .A(n1077), .B(n1078), .Z(n1076) );
  ANDN U1147 ( .A(n1079), .B(n1080), .Z(n1071) );
  XNOR U1148 ( .A(n1081), .B(n1013), .Z(n1067) );
  OR U1149 ( .A(n1051), .B(n1082), .Z(n1013) );
  XOR U1150 ( .A(n1075), .B(n1037), .Z(n1051) );
  XOR U1151 ( .A(n1083), .B(n1084), .Z(n1075) );
  ANDN U1152 ( .A(n1085), .B(n1078), .Z(n1084) );
  OR U1153 ( .A(n1037), .B(n1086), .Z(n1081) );
  XOR U1154 ( .A(n1087), .B(n1083), .Z(n1037) );
  XOR U1155 ( .A(n1078), .B(n1074), .Z(n1079) );
  XNOR U1156 ( .A(n1089), .B(n1090), .Z(n1078) );
  XNOR U1157 ( .A(n1091), .B(n1092), .Z(n1089) );
  NANDN U1158 ( .B(n1093), .A(n1073), .Z(n1091) );
  OR U1159 ( .A(n1074), .B(n1093), .Z(n1087) );
  XOR U1160 ( .A(n1094), .B(n1095), .Z(n1074) );
  XOR U1161 ( .A(n1096), .B(n1097), .Z(n1095) );
  XNOR U1162 ( .A(n1092), .B(n1098), .Z(n1097) );
  ANDN U1163 ( .A(n1085), .B(n1077), .Z(n1098) );
  OR U1164 ( .A(n1080), .B(n1088), .Z(n1092) );
  XNOR U1165 ( .A(n1099), .B(n1085), .Z(n1088) );
  XOR U1166 ( .A(n1073), .B(n1077), .Z(n1080) );
  IV U1167 ( .A(n1096), .Z(n1077) );
  XNOR U1168 ( .A(n1100), .B(n1101), .Z(n1096) );
  XNOR U1169 ( .A(n1086), .B(n1102), .Z(n1101) );
  XNOR U1170 ( .A(n1103), .B(n1104), .Z(n1102) );
  ANDN U1171 ( .A(n1015), .B(n1105), .Z(n1103) );
  XNOR U1172 ( .A(n1106), .B(n1107), .Z(n1100) );
  XOR U1173 ( .A(n1108), .B(n1036), .Z(n1106) );
  XOR U1174 ( .A(n1090), .B(n1085), .Z(n1094) );
  XNOR U1175 ( .A(n1109), .B(n1110), .Z(n1085) );
  XNOR U1176 ( .A(n1111), .B(n1112), .Z(n1110) );
  ANDN U1177 ( .A(n1028), .B(n1065), .Z(n1111) );
  XNOR U1178 ( .A(n1113), .B(n1108), .Z(n1109) );
  XOR U1179 ( .A(n1114), .B(n1115), .Z(n1108) );
  XNOR U1180 ( .A(n1116), .B(n1117), .Z(n1114) );
  NANDN U1181 ( .B(n1063), .A(n1048), .Z(n1116) );
  XNOR U1182 ( .A(n1099), .B(n1073), .Z(n1090) );
  XNOR U1183 ( .A(n1118), .B(n1119), .Z(n1073) );
  XOR U1184 ( .A(n1015), .B(n1120), .Z(n1119) );
  XNOR U1185 ( .A(n1121), .B(n1104), .Z(n1120) );
  OR U1186 ( .A(n1052), .B(n1082), .Z(n1104) );
  XNOR U1187 ( .A(n1050), .B(n1036), .Z(n1052) );
  IV U1188 ( .A(n1105), .Z(n1050) );
  ANDN U1189 ( .A(n1036), .B(n1086), .Z(n1121) );
  XNOR U1190 ( .A(n1122), .B(n1113), .Z(n1118) );
  XOR U1191 ( .A(n1115), .B(n1105), .Z(n1122) );
  IV U1192 ( .A(n1093), .Z(n1099) );
  XOR U1193 ( .A(n1123), .B(n1124), .Z(n1093) );
  XOR U1194 ( .A(n1115), .B(n1125), .Z(n1124) );
  XNOR U1195 ( .A(n1126), .B(n1112), .Z(n1125) );
  OR U1196 ( .A(n1025), .B(n1066), .Z(n1112) );
  XNOR U1197 ( .A(n1065), .B(n1057), .Z(n1066) );
  XNOR U1198 ( .A(n1127), .B(n1028), .Z(n1025) );
  ANDN U1199 ( .A(n1128), .B(n1005), .Z(n1126) );
  XNOR U1200 ( .A(n1117), .B(n1129), .Z(n1115) );
  ANDN U1201 ( .A(n1130), .B(n1042), .Z(n1129) );
  OR U1202 ( .A(n1070), .B(n1046), .Z(n1117) );
  XOR U1203 ( .A(n1042), .B(n1048), .Z(n1046) );
  XNOR U1204 ( .A(n1005), .B(n1036), .Z(n1048) );
  XNOR U1205 ( .A(n1131), .B(n1028), .Z(n1036) );
  XNOR U1206 ( .A(n1132), .B(n1133), .Z(n1131) );
  XOR U1207 ( .A(n1105), .B(n1028), .Z(n1042) );
  XOR U1208 ( .A(n1134), .B(n1135), .Z(n1105) );
  XNOR U1209 ( .A(n1136), .B(n1137), .Z(n1134) );
  XOR U1210 ( .A(n1130), .B(n1063), .Z(n1070) );
  XOR U1211 ( .A(n1128), .B(n1086), .Z(n1063) );
  XOR U1212 ( .A(n1138), .B(n1139), .Z(n1086) );
  XNOR U1213 ( .A(n1140), .B(n1015), .Z(n1139) );
  XNOR U1214 ( .A(n1141), .B(n1136), .Z(n1138) );
  XOR U1215 ( .A(g_input[108]), .B(state[108]), .Z(n1136) );
  IV U1216 ( .A(n1069), .Z(n1130) );
  XOR U1217 ( .A(n1065), .B(n1015), .Z(n1069) );
  XNOR U1218 ( .A(n1113), .B(n1107), .Z(n1123) );
  XNOR U1219 ( .A(n1127), .B(n1128), .Z(n1107) );
  IV U1220 ( .A(n1057), .Z(n1128) );
  IV U1221 ( .A(n1005), .Z(n1127) );
  XOR U1222 ( .A(n1142), .B(n1135), .Z(n1005) );
  XNOR U1223 ( .A(n1133), .B(n1137), .Z(n1142) );
  XOR U1224 ( .A(n1028), .B(n1065), .Z(n1113) );
  XNOR U1225 ( .A(n1132), .B(n1143), .Z(n1065) );
  XNOR U1226 ( .A(n1140), .B(n1137), .Z(n1143) );
  XOR U1227 ( .A(n1144), .B(n1133), .Z(n1140) );
  XOR U1228 ( .A(g_input[105]), .B(state[105]), .Z(n1133) );
  XNOR U1229 ( .A(g_input[107]), .B(state[107]), .Z(n1144) );
  XOR U1230 ( .A(g_input[106]), .B(state[106]), .Z(n1132) );
  XNOR U1231 ( .A(n1145), .B(n1135), .Z(n1028) );
  XOR U1232 ( .A(g_input[109]), .B(state[109]), .Z(n1135) );
  XNOR U1233 ( .A(n1141), .B(n1137), .Z(n1145) );
  XNOR U1234 ( .A(n1146), .B(n1015), .Z(n1137) );
  XOR U1235 ( .A(g_input[104]), .B(state[104]), .Z(n1015) );
  XNOR U1236 ( .A(g_input[110]), .B(state[110]), .Z(n1146) );
  XOR U1237 ( .A(g_input[111]), .B(state[111]), .Z(n1141) );
  XOR U1238 ( .A(n1147), .B(n1148), .Z(o[3]) );
  XOR U1239 ( .A(n337), .B(n1149), .Z(n1148) );
  XNOR U1240 ( .A(g_input[3]), .B(n1150), .Z(n1149) );
  XNOR U1241 ( .A(n514), .B(n341), .Z(n1147) );
  XNOR U1242 ( .A(n1151), .B(n1152), .Z(n514) );
  XNOR U1243 ( .A(n1153), .B(n692), .Z(n1151) );
  NANDN U1244 ( .B(n1154), .A(n1155), .Z(n692) );
  NANDN U1245 ( .B(n1156), .A(n1157), .Z(n1153) );
  XOR U1246 ( .A(n1158), .B(n1159), .Z(o[39]) );
  XOR U1247 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U1248 ( .A(n1163), .B(n1164), .Z(n1158) );
  XNOR U1249 ( .A(n1165), .B(n1166), .Z(o[38]) );
  XNOR U1250 ( .A(n1162), .B(g_input[38]), .Z(n1165) );
  XOR U1251 ( .A(n1167), .B(n1168), .Z(o[37]) );
  XOR U1252 ( .A(n1169), .B(n1170), .Z(n1168) );
  XNOR U1253 ( .A(g_input[37]), .B(n1171), .Z(n1170) );
  NOR U1254 ( .A(n1172), .B(n1173), .Z(n1169) );
  XNOR U1255 ( .A(n1174), .B(n1175), .Z(n1167) );
  XOR U1256 ( .A(n1163), .B(n1176), .Z(n1174) );
  XNOR U1257 ( .A(n1177), .B(n1178), .Z(n1163) );
  XNOR U1258 ( .A(n1179), .B(n1180), .Z(n1177) );
  NANDN U1259 ( .B(n1181), .A(n1182), .Z(n1179) );
  XNOR U1260 ( .A(n1183), .B(n1184), .Z(o[36]) );
  XOR U1261 ( .A(n1175), .B(g_input[36]), .Z(n1183) );
  XOR U1262 ( .A(n1185), .B(n1186), .Z(o[35]) );
  XOR U1263 ( .A(n1160), .B(n1187), .Z(n1186) );
  XNOR U1264 ( .A(g_input[35]), .B(n1188), .Z(n1187) );
  XNOR U1265 ( .A(n1166), .B(n1164), .Z(n1185) );
  XNOR U1266 ( .A(n1189), .B(n1190), .Z(n1166) );
  XNOR U1267 ( .A(n1191), .B(n1171), .Z(n1189) );
  NANDN U1268 ( .B(n1192), .A(n1193), .Z(n1171) );
  NANDN U1269 ( .B(n1194), .A(n1195), .Z(n1191) );
  XOR U1270 ( .A(n1184), .B(g_input[34]), .Z(o[34]) );
  XOR U1271 ( .A(n1196), .B(n1197), .Z(n1184) );
  XOR U1272 ( .A(n1198), .B(n1199), .Z(o[33]) );
  XOR U1273 ( .A(g_input[33]), .B(n1162), .Z(n1199) );
  XOR U1274 ( .A(n1188), .B(n1197), .Z(n1162) );
  XNOR U1275 ( .A(n1200), .B(n1176), .Z(n1188) );
  XOR U1276 ( .A(n1201), .B(n1202), .Z(n1200) );
  ANDN U1277 ( .A(n1203), .B(n1204), .Z(n1202) );
  XNOR U1278 ( .A(n1196), .B(n1160), .Z(n1198) );
  XOR U1279 ( .A(n1205), .B(n1190), .Z(n1160) );
  XNOR U1280 ( .A(n1206), .B(n1176), .Z(n1190) );
  XNOR U1281 ( .A(n1207), .B(n1208), .Z(n1176) );
  NOR U1282 ( .A(n1209), .B(n1210), .Z(n1208) );
  XOR U1283 ( .A(n1211), .B(n1207), .Z(n1206) );
  NOR U1284 ( .A(n1212), .B(n1213), .Z(n1207) );
  NANDN U1285 ( .B(n1214), .A(n1215), .Z(n1211) );
  XOR U1286 ( .A(n1201), .B(n1216), .Z(n1205) );
  ANDN U1287 ( .A(n1217), .B(n1181), .Z(n1216) );
  OR U1288 ( .A(n1218), .B(n1219), .Z(n1201) );
  IV U1289 ( .A(n1164), .Z(n1196) );
  XNOR U1290 ( .A(n1220), .B(n1221), .Z(n1164) );
  XNOR U1291 ( .A(n1222), .B(n1223), .Z(n1220) );
  NOR U1292 ( .A(n1224), .B(n1173), .Z(n1223) );
  XNOR U1293 ( .A(n1225), .B(n1175), .Z(o[32]) );
  XOR U1294 ( .A(n1226), .B(n1178), .Z(n1175) );
  XOR U1295 ( .A(n1227), .B(n1221), .Z(n1178) );
  XNOR U1296 ( .A(n1228), .B(n1229), .Z(n1227) );
  NOR U1297 ( .A(n1214), .B(n1230), .Z(n1229) );
  XNOR U1298 ( .A(n1222), .B(n1231), .Z(n1226) );
  NOR U1299 ( .A(n1194), .B(n1232), .Z(n1231) );
  ANDN U1300 ( .A(n1193), .B(n1233), .Z(n1222) );
  XOR U1301 ( .A(n1194), .B(n1173), .Z(n1193) );
  XOR U1302 ( .A(n1197), .B(g_input[32]), .Z(n1225) );
  XNOR U1303 ( .A(n1234), .B(n1221), .Z(n1197) );
  XNOR U1304 ( .A(n1228), .B(n1235), .Z(n1221) );
  NOR U1305 ( .A(n1236), .B(n1210), .Z(n1235) );
  NOR U1306 ( .A(n1212), .B(n1237), .Z(n1228) );
  XNOR U1307 ( .A(n1204), .B(n1173), .Z(n1214) );
  XNOR U1308 ( .A(n1238), .B(n1239), .Z(n1173) );
  ANDN U1309 ( .A(n1240), .B(n1241), .Z(n1239) );
  IV U1310 ( .A(n1242), .Z(n1181) );
  XNOR U1311 ( .A(n1238), .B(n1243), .Z(n1194) );
  NOR U1312 ( .A(n1244), .B(n1245), .Z(n1243) );
  ANDN U1313 ( .A(n1246), .B(n1247), .Z(n1238) );
  XNOR U1314 ( .A(n1248), .B(n1180), .Z(n1234) );
  OR U1315 ( .A(n1218), .B(n1249), .Z(n1180) );
  XOR U1316 ( .A(n1242), .B(n1204), .Z(n1218) );
  XOR U1317 ( .A(n1250), .B(n1251), .Z(n1242) );
  ANDN U1318 ( .A(n1252), .B(n1245), .Z(n1251) );
  OR U1319 ( .A(n1204), .B(n1253), .Z(n1248) );
  XOR U1320 ( .A(n1254), .B(n1250), .Z(n1204) );
  XOR U1321 ( .A(n1245), .B(n1241), .Z(n1246) );
  XNOR U1322 ( .A(n1256), .B(n1257), .Z(n1245) );
  XNOR U1323 ( .A(n1258), .B(n1259), .Z(n1256) );
  NANDN U1324 ( .B(n1260), .A(n1240), .Z(n1258) );
  OR U1325 ( .A(n1241), .B(n1260), .Z(n1254) );
  XOR U1326 ( .A(n1261), .B(n1262), .Z(n1241) );
  XOR U1327 ( .A(n1263), .B(n1264), .Z(n1262) );
  XNOR U1328 ( .A(n1259), .B(n1265), .Z(n1264) );
  ANDN U1329 ( .A(n1252), .B(n1244), .Z(n1265) );
  OR U1330 ( .A(n1247), .B(n1255), .Z(n1259) );
  XNOR U1331 ( .A(n1266), .B(n1252), .Z(n1255) );
  XOR U1332 ( .A(n1240), .B(n1244), .Z(n1247) );
  IV U1333 ( .A(n1263), .Z(n1244) );
  XNOR U1334 ( .A(n1267), .B(n1268), .Z(n1263) );
  XNOR U1335 ( .A(n1253), .B(n1269), .Z(n1268) );
  XNOR U1336 ( .A(n1270), .B(n1271), .Z(n1269) );
  ANDN U1337 ( .A(n1182), .B(n1272), .Z(n1270) );
  XNOR U1338 ( .A(n1273), .B(n1274), .Z(n1267) );
  XOR U1339 ( .A(n1275), .B(n1203), .Z(n1273) );
  XOR U1340 ( .A(n1257), .B(n1252), .Z(n1261) );
  XNOR U1341 ( .A(n1276), .B(n1277), .Z(n1252) );
  XNOR U1342 ( .A(n1278), .B(n1279), .Z(n1277) );
  ANDN U1343 ( .A(n1195), .B(n1232), .Z(n1278) );
  XNOR U1344 ( .A(n1280), .B(n1275), .Z(n1276) );
  XOR U1345 ( .A(n1281), .B(n1282), .Z(n1275) );
  XNOR U1346 ( .A(n1283), .B(n1284), .Z(n1281) );
  NANDN U1347 ( .B(n1230), .A(n1215), .Z(n1283) );
  XNOR U1348 ( .A(n1266), .B(n1240), .Z(n1257) );
  XNOR U1349 ( .A(n1285), .B(n1286), .Z(n1240) );
  XOR U1350 ( .A(n1182), .B(n1287), .Z(n1286) );
  XNOR U1351 ( .A(n1288), .B(n1271), .Z(n1287) );
  OR U1352 ( .A(n1219), .B(n1249), .Z(n1271) );
  XNOR U1353 ( .A(n1217), .B(n1203), .Z(n1219) );
  IV U1354 ( .A(n1272), .Z(n1217) );
  ANDN U1355 ( .A(n1203), .B(n1253), .Z(n1288) );
  XNOR U1356 ( .A(n1289), .B(n1280), .Z(n1285) );
  XOR U1357 ( .A(n1282), .B(n1272), .Z(n1289) );
  IV U1358 ( .A(n1260), .Z(n1266) );
  XOR U1359 ( .A(n1290), .B(n1291), .Z(n1260) );
  XOR U1360 ( .A(n1282), .B(n1292), .Z(n1291) );
  XNOR U1361 ( .A(n1293), .B(n1279), .Z(n1292) );
  OR U1362 ( .A(n1192), .B(n1233), .Z(n1279) );
  XNOR U1363 ( .A(n1232), .B(n1224), .Z(n1233) );
  XNOR U1364 ( .A(n1294), .B(n1195), .Z(n1192) );
  ANDN U1365 ( .A(n1295), .B(n1172), .Z(n1293) );
  XNOR U1366 ( .A(n1284), .B(n1296), .Z(n1282) );
  ANDN U1367 ( .A(n1297), .B(n1209), .Z(n1296) );
  OR U1368 ( .A(n1237), .B(n1213), .Z(n1284) );
  XOR U1369 ( .A(n1209), .B(n1215), .Z(n1213) );
  XNOR U1370 ( .A(n1172), .B(n1203), .Z(n1215) );
  XNOR U1371 ( .A(n1298), .B(n1195), .Z(n1203) );
  XOR U1372 ( .A(n1299), .B(n1300), .Z(n1298) );
  IV U1373 ( .A(n1294), .Z(n1172) );
  XOR U1374 ( .A(n1272), .B(n1195), .Z(n1209) );
  XOR U1375 ( .A(n1301), .B(n1302), .Z(n1272) );
  XOR U1376 ( .A(n1303), .B(n1304), .Z(n1301) );
  XOR U1377 ( .A(n1297), .B(n1230), .Z(n1237) );
  XOR U1378 ( .A(n1295), .B(n1253), .Z(n1230) );
  XOR U1379 ( .A(n1305), .B(n1306), .Z(n1253) );
  XNOR U1380 ( .A(n1307), .B(n1182), .Z(n1306) );
  XNOR U1381 ( .A(n1308), .B(n1303), .Z(n1305) );
  XNOR U1382 ( .A(g_input[68]), .B(state[68]), .Z(n1303) );
  IV U1383 ( .A(n1236), .Z(n1297) );
  XOR U1384 ( .A(n1232), .B(n1182), .Z(n1236) );
  XNOR U1385 ( .A(n1280), .B(n1274), .Z(n1290) );
  XNOR U1386 ( .A(n1294), .B(n1295), .Z(n1274) );
  IV U1387 ( .A(n1224), .Z(n1295) );
  XOR U1388 ( .A(n1309), .B(n1304), .Z(n1224) );
  XOR U1389 ( .A(n1310), .B(n1309), .Z(n1294) );
  IV U1390 ( .A(n1302), .Z(n1309) );
  XNOR U1391 ( .A(n1300), .B(n1304), .Z(n1310) );
  XOR U1392 ( .A(n1195), .B(n1232), .Z(n1280) );
  XOR U1393 ( .A(n1299), .B(n1311), .Z(n1232) );
  XNOR U1394 ( .A(n1307), .B(n1304), .Z(n1311) );
  XOR U1395 ( .A(n1312), .B(n1300), .Z(n1307) );
  XOR U1396 ( .A(g_input[65]), .B(state[65]), .Z(n1300) );
  XNOR U1397 ( .A(g_input[67]), .B(state[67]), .Z(n1312) );
  XNOR U1398 ( .A(g_input[66]), .B(state[66]), .Z(n1299) );
  XNOR U1399 ( .A(n1313), .B(n1302), .Z(n1195) );
  XOR U1400 ( .A(g_input[69]), .B(state[69]), .Z(n1302) );
  XOR U1401 ( .A(n1308), .B(n1304), .Z(n1313) );
  XNOR U1402 ( .A(n1314), .B(n1182), .Z(n1304) );
  XOR U1403 ( .A(g_input[64]), .B(state[64]), .Z(n1182) );
  XNOR U1404 ( .A(g_input[70]), .B(state[70]), .Z(n1314) );
  XNOR U1405 ( .A(g_input[71]), .B(state[71]), .Z(n1308) );
  XOR U1406 ( .A(n1315), .B(n1316), .Z(o[31]) );
  XOR U1407 ( .A(n1317), .B(n1318), .Z(n1316) );
  XOR U1408 ( .A(n1320), .B(n1321), .Z(n1315) );
  XNOR U1409 ( .A(n1322), .B(n1323), .Z(o[30]) );
  XNOR U1410 ( .A(n1319), .B(g_input[30]), .Z(n1322) );
  XOR U1411 ( .A(n874), .B(g_input[2]), .Z(o[2]) );
  XOR U1412 ( .A(n1324), .B(n1325), .Z(n874) );
  XOR U1413 ( .A(n1326), .B(n1327), .Z(o[29]) );
  XOR U1414 ( .A(n1328), .B(n1329), .Z(n1327) );
  XNOR U1415 ( .A(g_input[29]), .B(n1330), .Z(n1329) );
  NOR U1416 ( .A(n1331), .B(n1332), .Z(n1328) );
  XNOR U1417 ( .A(n1333), .B(n1334), .Z(n1326) );
  XOR U1418 ( .A(n1320), .B(n1335), .Z(n1333) );
  XNOR U1419 ( .A(n1336), .B(n1337), .Z(n1320) );
  XNOR U1420 ( .A(n1338), .B(n1339), .Z(n1336) );
  NANDN U1421 ( .B(n1340), .A(n1341), .Z(n1338) );
  XNOR U1422 ( .A(n1342), .B(n1343), .Z(o[28]) );
  XOR U1423 ( .A(n1334), .B(g_input[28]), .Z(n1342) );
  XOR U1424 ( .A(n1344), .B(n1345), .Z(o[27]) );
  XOR U1425 ( .A(n1317), .B(n1346), .Z(n1345) );
  XNOR U1426 ( .A(g_input[27]), .B(n1347), .Z(n1346) );
  XNOR U1427 ( .A(n1323), .B(n1321), .Z(n1344) );
  XNOR U1428 ( .A(n1348), .B(n1349), .Z(n1323) );
  XNOR U1429 ( .A(n1350), .B(n1330), .Z(n1348) );
  NANDN U1430 ( .B(n1351), .A(n1352), .Z(n1330) );
  NANDN U1431 ( .B(n1353), .A(n1354), .Z(n1350) );
  XOR U1432 ( .A(n1343), .B(g_input[26]), .Z(o[26]) );
  XOR U1433 ( .A(n1355), .B(n1356), .Z(n1343) );
  XOR U1434 ( .A(n1357), .B(n1358), .Z(o[25]) );
  XOR U1435 ( .A(g_input[25]), .B(n1319), .Z(n1358) );
  XOR U1436 ( .A(n1347), .B(n1356), .Z(n1319) );
  XNOR U1437 ( .A(n1359), .B(n1335), .Z(n1347) );
  XOR U1438 ( .A(n1360), .B(n1361), .Z(n1359) );
  ANDN U1439 ( .A(n1362), .B(n1363), .Z(n1361) );
  XNOR U1440 ( .A(n1355), .B(n1317), .Z(n1357) );
  XOR U1441 ( .A(n1364), .B(n1349), .Z(n1317) );
  XNOR U1442 ( .A(n1365), .B(n1335), .Z(n1349) );
  XNOR U1443 ( .A(n1366), .B(n1367), .Z(n1335) );
  NOR U1444 ( .A(n1368), .B(n1369), .Z(n1367) );
  XOR U1445 ( .A(n1370), .B(n1366), .Z(n1365) );
  NOR U1446 ( .A(n1371), .B(n1372), .Z(n1366) );
  NANDN U1447 ( .B(n1373), .A(n1374), .Z(n1370) );
  XOR U1448 ( .A(n1360), .B(n1375), .Z(n1364) );
  ANDN U1449 ( .A(n1376), .B(n1340), .Z(n1375) );
  OR U1450 ( .A(n1377), .B(n1378), .Z(n1360) );
  IV U1451 ( .A(n1321), .Z(n1355) );
  XNOR U1452 ( .A(n1379), .B(n1380), .Z(n1321) );
  XNOR U1453 ( .A(n1381), .B(n1382), .Z(n1379) );
  NOR U1454 ( .A(n1383), .B(n1332), .Z(n1382) );
  XNOR U1455 ( .A(n1384), .B(n1334), .Z(o[24]) );
  XOR U1456 ( .A(n1385), .B(n1337), .Z(n1334) );
  XOR U1457 ( .A(n1386), .B(n1380), .Z(n1337) );
  XNOR U1458 ( .A(n1387), .B(n1388), .Z(n1386) );
  NOR U1459 ( .A(n1373), .B(n1389), .Z(n1388) );
  XNOR U1460 ( .A(n1381), .B(n1390), .Z(n1385) );
  NOR U1461 ( .A(n1353), .B(n1391), .Z(n1390) );
  ANDN U1462 ( .A(n1352), .B(n1392), .Z(n1381) );
  XOR U1463 ( .A(n1353), .B(n1332), .Z(n1352) );
  XOR U1464 ( .A(n1356), .B(g_input[24]), .Z(n1384) );
  XNOR U1465 ( .A(n1393), .B(n1380), .Z(n1356) );
  XNOR U1466 ( .A(n1387), .B(n1394), .Z(n1380) );
  NOR U1467 ( .A(n1395), .B(n1369), .Z(n1394) );
  NOR U1468 ( .A(n1371), .B(n1396), .Z(n1387) );
  XNOR U1469 ( .A(n1363), .B(n1332), .Z(n1373) );
  XNOR U1470 ( .A(n1397), .B(n1398), .Z(n1332) );
  ANDN U1471 ( .A(n1399), .B(n1400), .Z(n1398) );
  IV U1472 ( .A(n1401), .Z(n1340) );
  XNOR U1473 ( .A(n1397), .B(n1402), .Z(n1353) );
  NOR U1474 ( .A(n1403), .B(n1404), .Z(n1402) );
  ANDN U1475 ( .A(n1405), .B(n1406), .Z(n1397) );
  XNOR U1476 ( .A(n1407), .B(n1339), .Z(n1393) );
  OR U1477 ( .A(n1377), .B(n1408), .Z(n1339) );
  XOR U1478 ( .A(n1401), .B(n1363), .Z(n1377) );
  XOR U1479 ( .A(n1409), .B(n1410), .Z(n1401) );
  ANDN U1480 ( .A(n1411), .B(n1404), .Z(n1410) );
  OR U1481 ( .A(n1363), .B(n1412), .Z(n1407) );
  XOR U1482 ( .A(n1413), .B(n1409), .Z(n1363) );
  XOR U1483 ( .A(n1404), .B(n1400), .Z(n1405) );
  XNOR U1484 ( .A(n1415), .B(n1416), .Z(n1404) );
  XNOR U1485 ( .A(n1417), .B(n1418), .Z(n1415) );
  NANDN U1486 ( .B(n1419), .A(n1399), .Z(n1417) );
  OR U1487 ( .A(n1400), .B(n1419), .Z(n1413) );
  XOR U1488 ( .A(n1420), .B(n1421), .Z(n1400) );
  XOR U1489 ( .A(n1422), .B(n1423), .Z(n1421) );
  XNOR U1490 ( .A(n1418), .B(n1424), .Z(n1423) );
  ANDN U1491 ( .A(n1411), .B(n1403), .Z(n1424) );
  OR U1492 ( .A(n1406), .B(n1414), .Z(n1418) );
  XNOR U1493 ( .A(n1425), .B(n1411), .Z(n1414) );
  XOR U1494 ( .A(n1399), .B(n1403), .Z(n1406) );
  IV U1495 ( .A(n1422), .Z(n1403) );
  XNOR U1496 ( .A(n1426), .B(n1427), .Z(n1422) );
  XNOR U1497 ( .A(n1412), .B(n1428), .Z(n1427) );
  XNOR U1498 ( .A(n1429), .B(n1430), .Z(n1428) );
  ANDN U1499 ( .A(n1341), .B(n1431), .Z(n1429) );
  XNOR U1500 ( .A(n1432), .B(n1433), .Z(n1426) );
  XOR U1501 ( .A(n1434), .B(n1362), .Z(n1432) );
  XOR U1502 ( .A(n1416), .B(n1411), .Z(n1420) );
  XNOR U1503 ( .A(n1435), .B(n1436), .Z(n1411) );
  XNOR U1504 ( .A(n1437), .B(n1438), .Z(n1436) );
  ANDN U1505 ( .A(n1354), .B(n1391), .Z(n1437) );
  XNOR U1506 ( .A(n1439), .B(n1434), .Z(n1435) );
  XOR U1507 ( .A(n1440), .B(n1441), .Z(n1434) );
  XNOR U1508 ( .A(n1442), .B(n1443), .Z(n1440) );
  NANDN U1509 ( .B(n1389), .A(n1374), .Z(n1442) );
  XNOR U1510 ( .A(n1425), .B(n1399), .Z(n1416) );
  XNOR U1511 ( .A(n1444), .B(n1445), .Z(n1399) );
  XOR U1512 ( .A(n1341), .B(n1446), .Z(n1445) );
  XNOR U1513 ( .A(n1447), .B(n1430), .Z(n1446) );
  OR U1514 ( .A(n1378), .B(n1408), .Z(n1430) );
  XNOR U1515 ( .A(n1376), .B(n1362), .Z(n1378) );
  IV U1516 ( .A(n1431), .Z(n1376) );
  ANDN U1517 ( .A(n1362), .B(n1412), .Z(n1447) );
  XNOR U1518 ( .A(n1448), .B(n1439), .Z(n1444) );
  XOR U1519 ( .A(n1441), .B(n1431), .Z(n1448) );
  IV U1520 ( .A(n1419), .Z(n1425) );
  XOR U1521 ( .A(n1449), .B(n1450), .Z(n1419) );
  XOR U1522 ( .A(n1441), .B(n1451), .Z(n1450) );
  XNOR U1523 ( .A(n1452), .B(n1438), .Z(n1451) );
  OR U1524 ( .A(n1351), .B(n1392), .Z(n1438) );
  XNOR U1525 ( .A(n1391), .B(n1383), .Z(n1392) );
  XNOR U1526 ( .A(n1453), .B(n1354), .Z(n1351) );
  ANDN U1527 ( .A(n1454), .B(n1331), .Z(n1452) );
  XNOR U1528 ( .A(n1443), .B(n1455), .Z(n1441) );
  ANDN U1529 ( .A(n1456), .B(n1368), .Z(n1455) );
  OR U1530 ( .A(n1396), .B(n1372), .Z(n1443) );
  XOR U1531 ( .A(n1368), .B(n1374), .Z(n1372) );
  XNOR U1532 ( .A(n1331), .B(n1362), .Z(n1374) );
  XNOR U1533 ( .A(n1457), .B(n1354), .Z(n1362) );
  XNOR U1534 ( .A(n1458), .B(n1459), .Z(n1457) );
  XOR U1535 ( .A(n1431), .B(n1354), .Z(n1368) );
  XOR U1536 ( .A(n1460), .B(n1461), .Z(n1431) );
  XNOR U1537 ( .A(n1462), .B(n1463), .Z(n1460) );
  XOR U1538 ( .A(n1456), .B(n1389), .Z(n1396) );
  XOR U1539 ( .A(n1454), .B(n1412), .Z(n1389) );
  XOR U1540 ( .A(n1464), .B(n1465), .Z(n1412) );
  XNOR U1541 ( .A(n1466), .B(n1341), .Z(n1465) );
  XNOR U1542 ( .A(n1467), .B(n1462), .Z(n1464) );
  XOR U1543 ( .A(g_input[28]), .B(state[28]), .Z(n1462) );
  IV U1544 ( .A(n1395), .Z(n1456) );
  XOR U1545 ( .A(n1391), .B(n1341), .Z(n1395) );
  XNOR U1546 ( .A(n1439), .B(n1433), .Z(n1449) );
  XNOR U1547 ( .A(n1453), .B(n1454), .Z(n1433) );
  IV U1548 ( .A(n1383), .Z(n1454) );
  IV U1549 ( .A(n1331), .Z(n1453) );
  XOR U1550 ( .A(n1468), .B(n1461), .Z(n1331) );
  XNOR U1551 ( .A(n1459), .B(n1463), .Z(n1468) );
  XOR U1552 ( .A(n1354), .B(n1391), .Z(n1439) );
  XNOR U1553 ( .A(n1458), .B(n1469), .Z(n1391) );
  XNOR U1554 ( .A(n1466), .B(n1463), .Z(n1469) );
  XOR U1555 ( .A(n1470), .B(n1459), .Z(n1466) );
  XOR U1556 ( .A(g_input[25]), .B(state[25]), .Z(n1459) );
  XNOR U1557 ( .A(g_input[27]), .B(state[27]), .Z(n1470) );
  XOR U1558 ( .A(g_input[26]), .B(state[26]), .Z(n1458) );
  XNOR U1559 ( .A(n1471), .B(n1461), .Z(n1354) );
  XOR U1560 ( .A(g_input[29]), .B(state[29]), .Z(n1461) );
  XNOR U1561 ( .A(n1467), .B(n1463), .Z(n1471) );
  XNOR U1562 ( .A(n1472), .B(n1341), .Z(n1463) );
  XOR U1563 ( .A(g_input[24]), .B(state[24]), .Z(n1341) );
  XNOR U1564 ( .A(g_input[30]), .B(state[30]), .Z(n1472) );
  XOR U1565 ( .A(g_input[31]), .B(state[31]), .Z(n1467) );
  XOR U1566 ( .A(n1473), .B(n1474), .Z(o[23]) );
  XOR U1567 ( .A(n1475), .B(n1476), .Z(n1474) );
  XOR U1568 ( .A(n1478), .B(n1479), .Z(n1473) );
  XNOR U1569 ( .A(n1480), .B(n1481), .Z(o[22]) );
  XNOR U1570 ( .A(n1477), .B(g_input[22]), .Z(n1480) );
  XOR U1571 ( .A(n1482), .B(n1483), .Z(o[21]) );
  XOR U1572 ( .A(n1484), .B(n1485), .Z(n1483) );
  XNOR U1573 ( .A(g_input[21]), .B(n1486), .Z(n1485) );
  NOR U1574 ( .A(n1487), .B(n1488), .Z(n1484) );
  XNOR U1575 ( .A(n1489), .B(n1490), .Z(n1482) );
  XOR U1576 ( .A(n1478), .B(n1491), .Z(n1489) );
  XNOR U1577 ( .A(n1492), .B(n1493), .Z(n1478) );
  XNOR U1578 ( .A(n1494), .B(n1495), .Z(n1492) );
  NANDN U1579 ( .B(n1496), .A(n1497), .Z(n1494) );
  XNOR U1580 ( .A(n1498), .B(n1499), .Z(o[20]) );
  XOR U1581 ( .A(n1490), .B(g_input[20]), .Z(n1498) );
  XOR U1582 ( .A(n1500), .B(n1501), .Z(o[1]) );
  XOR U1583 ( .A(g_input[1]), .B(n339), .Z(n1501) );
  XOR U1584 ( .A(n1150), .B(n1325), .Z(n339) );
  XNOR U1585 ( .A(n1502), .B(n697), .Z(n1150) );
  XOR U1586 ( .A(n1503), .B(n1504), .Z(n1502) );
  ANDN U1587 ( .A(n1505), .B(n1506), .Z(n1504) );
  XNOR U1588 ( .A(n1324), .B(n337), .Z(n1500) );
  XOR U1589 ( .A(n1507), .B(n1152), .Z(n337) );
  XNOR U1590 ( .A(n1508), .B(n697), .Z(n1152) );
  XNOR U1591 ( .A(n1509), .B(n1510), .Z(n697) );
  NOR U1592 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U1593 ( .A(n1513), .B(n1509), .Z(n1508) );
  NOR U1594 ( .A(n1514), .B(n1515), .Z(n1509) );
  NANDN U1595 ( .B(n1516), .A(n1517), .Z(n1513) );
  XOR U1596 ( .A(n1503), .B(n1518), .Z(n1507) );
  ANDN U1597 ( .A(n1519), .B(n702), .Z(n1518) );
  OR U1598 ( .A(n1520), .B(n1521), .Z(n1503) );
  IV U1599 ( .A(n341), .Z(n1324) );
  XNOR U1600 ( .A(n1522), .B(n1523), .Z(n341) );
  XNOR U1601 ( .A(n1524), .B(n1525), .Z(n1522) );
  NOR U1602 ( .A(n1526), .B(n694), .Z(n1525) );
  XOR U1603 ( .A(n1527), .B(n1528), .Z(o[19]) );
  XOR U1604 ( .A(n1475), .B(n1529), .Z(n1528) );
  XNOR U1605 ( .A(g_input[19]), .B(n1530), .Z(n1529) );
  XNOR U1606 ( .A(n1481), .B(n1479), .Z(n1527) );
  XNOR U1607 ( .A(n1531), .B(n1532), .Z(n1481) );
  XNOR U1608 ( .A(n1533), .B(n1486), .Z(n1531) );
  NANDN U1609 ( .B(n1534), .A(n1535), .Z(n1486) );
  NANDN U1610 ( .B(n1536), .A(n1537), .Z(n1533) );
  XOR U1611 ( .A(n1499), .B(g_input[18]), .Z(o[18]) );
  XOR U1612 ( .A(n1538), .B(n1539), .Z(n1499) );
  XOR U1613 ( .A(n1540), .B(n1541), .Z(o[17]) );
  XOR U1614 ( .A(g_input[17]), .B(n1477), .Z(n1541) );
  XOR U1615 ( .A(n1530), .B(n1539), .Z(n1477) );
  XNOR U1616 ( .A(n1542), .B(n1491), .Z(n1530) );
  XOR U1617 ( .A(n1543), .B(n1544), .Z(n1542) );
  ANDN U1618 ( .A(n1545), .B(n1546), .Z(n1544) );
  XNOR U1619 ( .A(n1538), .B(n1475), .Z(n1540) );
  XOR U1620 ( .A(n1547), .B(n1532), .Z(n1475) );
  XNOR U1621 ( .A(n1548), .B(n1491), .Z(n1532) );
  XNOR U1622 ( .A(n1549), .B(n1550), .Z(n1491) );
  NOR U1623 ( .A(n1551), .B(n1552), .Z(n1550) );
  XOR U1624 ( .A(n1553), .B(n1549), .Z(n1548) );
  NOR U1625 ( .A(n1554), .B(n1555), .Z(n1549) );
  NANDN U1626 ( .B(n1556), .A(n1557), .Z(n1553) );
  XOR U1627 ( .A(n1543), .B(n1558), .Z(n1547) );
  ANDN U1628 ( .A(n1559), .B(n1496), .Z(n1558) );
  OR U1629 ( .A(n1560), .B(n1561), .Z(n1543) );
  IV U1630 ( .A(n1479), .Z(n1538) );
  XNOR U1631 ( .A(n1562), .B(n1563), .Z(n1479) );
  XNOR U1632 ( .A(n1564), .B(n1565), .Z(n1562) );
  NOR U1633 ( .A(n1566), .B(n1488), .Z(n1565) );
  XNOR U1634 ( .A(n1567), .B(n1490), .Z(o[16]) );
  XOR U1635 ( .A(n1568), .B(n1493), .Z(n1490) );
  XOR U1636 ( .A(n1569), .B(n1563), .Z(n1493) );
  XNOR U1637 ( .A(n1570), .B(n1571), .Z(n1569) );
  NOR U1638 ( .A(n1556), .B(n1572), .Z(n1571) );
  XNOR U1639 ( .A(n1564), .B(n1573), .Z(n1568) );
  NOR U1640 ( .A(n1536), .B(n1574), .Z(n1573) );
  ANDN U1641 ( .A(n1535), .B(n1575), .Z(n1564) );
  XOR U1642 ( .A(n1536), .B(n1488), .Z(n1535) );
  XOR U1643 ( .A(n1539), .B(g_input[16]), .Z(n1567) );
  XNOR U1644 ( .A(n1576), .B(n1563), .Z(n1539) );
  XNOR U1645 ( .A(n1570), .B(n1577), .Z(n1563) );
  NOR U1646 ( .A(n1578), .B(n1552), .Z(n1577) );
  NOR U1647 ( .A(n1554), .B(n1579), .Z(n1570) );
  XNOR U1648 ( .A(n1546), .B(n1488), .Z(n1556) );
  XNOR U1649 ( .A(n1580), .B(n1581), .Z(n1488) );
  ANDN U1650 ( .A(n1582), .B(n1583), .Z(n1581) );
  IV U1651 ( .A(n1584), .Z(n1496) );
  XNOR U1652 ( .A(n1580), .B(n1585), .Z(n1536) );
  NOR U1653 ( .A(n1586), .B(n1587), .Z(n1585) );
  ANDN U1654 ( .A(n1588), .B(n1589), .Z(n1580) );
  XNOR U1655 ( .A(n1590), .B(n1495), .Z(n1576) );
  OR U1656 ( .A(n1560), .B(n1591), .Z(n1495) );
  XOR U1657 ( .A(n1584), .B(n1546), .Z(n1560) );
  XOR U1658 ( .A(n1592), .B(n1593), .Z(n1584) );
  ANDN U1659 ( .A(n1594), .B(n1587), .Z(n1593) );
  OR U1660 ( .A(n1546), .B(n1595), .Z(n1590) );
  XOR U1661 ( .A(n1596), .B(n1592), .Z(n1546) );
  XOR U1662 ( .A(n1587), .B(n1583), .Z(n1588) );
  XNOR U1663 ( .A(n1598), .B(n1599), .Z(n1587) );
  XNOR U1664 ( .A(n1600), .B(n1601), .Z(n1598) );
  NANDN U1665 ( .B(n1602), .A(n1582), .Z(n1600) );
  OR U1666 ( .A(n1583), .B(n1602), .Z(n1596) );
  XOR U1667 ( .A(n1603), .B(n1604), .Z(n1583) );
  XOR U1668 ( .A(n1605), .B(n1606), .Z(n1604) );
  XNOR U1669 ( .A(n1601), .B(n1607), .Z(n1606) );
  ANDN U1670 ( .A(n1594), .B(n1586), .Z(n1607) );
  OR U1671 ( .A(n1589), .B(n1597), .Z(n1601) );
  XNOR U1672 ( .A(n1608), .B(n1594), .Z(n1597) );
  XOR U1673 ( .A(n1582), .B(n1586), .Z(n1589) );
  IV U1674 ( .A(n1605), .Z(n1586) );
  XNOR U1675 ( .A(n1609), .B(n1610), .Z(n1605) );
  XNOR U1676 ( .A(n1595), .B(n1611), .Z(n1610) );
  XNOR U1677 ( .A(n1612), .B(n1613), .Z(n1611) );
  ANDN U1678 ( .A(n1497), .B(n1614), .Z(n1612) );
  XNOR U1679 ( .A(n1615), .B(n1616), .Z(n1609) );
  XOR U1680 ( .A(n1617), .B(n1545), .Z(n1615) );
  XOR U1681 ( .A(n1599), .B(n1594), .Z(n1603) );
  XNOR U1682 ( .A(n1618), .B(n1619), .Z(n1594) );
  XNOR U1683 ( .A(n1620), .B(n1621), .Z(n1619) );
  ANDN U1684 ( .A(n1537), .B(n1574), .Z(n1620) );
  XNOR U1685 ( .A(n1622), .B(n1617), .Z(n1618) );
  XOR U1686 ( .A(n1623), .B(n1624), .Z(n1617) );
  XNOR U1687 ( .A(n1625), .B(n1626), .Z(n1623) );
  NANDN U1688 ( .B(n1572), .A(n1557), .Z(n1625) );
  XNOR U1689 ( .A(n1608), .B(n1582), .Z(n1599) );
  XNOR U1690 ( .A(n1627), .B(n1628), .Z(n1582) );
  XOR U1691 ( .A(n1497), .B(n1629), .Z(n1628) );
  XNOR U1692 ( .A(n1630), .B(n1613), .Z(n1629) );
  OR U1693 ( .A(n1561), .B(n1591), .Z(n1613) );
  XNOR U1694 ( .A(n1559), .B(n1545), .Z(n1561) );
  IV U1695 ( .A(n1614), .Z(n1559) );
  ANDN U1696 ( .A(n1545), .B(n1595), .Z(n1630) );
  XNOR U1697 ( .A(n1631), .B(n1622), .Z(n1627) );
  XOR U1698 ( .A(n1624), .B(n1614), .Z(n1631) );
  IV U1699 ( .A(n1602), .Z(n1608) );
  XOR U1700 ( .A(n1632), .B(n1633), .Z(n1602) );
  XOR U1701 ( .A(n1624), .B(n1634), .Z(n1633) );
  XNOR U1702 ( .A(n1635), .B(n1621), .Z(n1634) );
  OR U1703 ( .A(n1534), .B(n1575), .Z(n1621) );
  XNOR U1704 ( .A(n1574), .B(n1566), .Z(n1575) );
  XNOR U1705 ( .A(n1636), .B(n1537), .Z(n1534) );
  ANDN U1706 ( .A(n1637), .B(n1487), .Z(n1635) );
  XNOR U1707 ( .A(n1626), .B(n1638), .Z(n1624) );
  ANDN U1708 ( .A(n1639), .B(n1551), .Z(n1638) );
  OR U1709 ( .A(n1579), .B(n1555), .Z(n1626) );
  XOR U1710 ( .A(n1551), .B(n1557), .Z(n1555) );
  XNOR U1711 ( .A(n1487), .B(n1545), .Z(n1557) );
  XNOR U1712 ( .A(n1640), .B(n1537), .Z(n1545) );
  XNOR U1713 ( .A(n1641), .B(n1642), .Z(n1640) );
  XOR U1714 ( .A(n1614), .B(n1537), .Z(n1551) );
  XOR U1715 ( .A(n1643), .B(n1644), .Z(n1614) );
  XNOR U1716 ( .A(n1645), .B(n1646), .Z(n1643) );
  XOR U1717 ( .A(n1639), .B(n1572), .Z(n1579) );
  XOR U1718 ( .A(n1637), .B(n1595), .Z(n1572) );
  XOR U1719 ( .A(n1647), .B(n1648), .Z(n1595) );
  XNOR U1720 ( .A(n1649), .B(n1497), .Z(n1648) );
  XNOR U1721 ( .A(n1650), .B(n1645), .Z(n1647) );
  XOR U1722 ( .A(g_input[116]), .B(state[116]), .Z(n1645) );
  IV U1723 ( .A(n1578), .Z(n1639) );
  XOR U1724 ( .A(n1574), .B(n1497), .Z(n1578) );
  XNOR U1725 ( .A(n1622), .B(n1616), .Z(n1632) );
  XNOR U1726 ( .A(n1636), .B(n1637), .Z(n1616) );
  IV U1727 ( .A(n1566), .Z(n1637) );
  IV U1728 ( .A(n1487), .Z(n1636) );
  XOR U1729 ( .A(n1651), .B(n1644), .Z(n1487) );
  XNOR U1730 ( .A(n1642), .B(n1646), .Z(n1651) );
  XOR U1731 ( .A(n1537), .B(n1574), .Z(n1622) );
  XNOR U1732 ( .A(n1641), .B(n1652), .Z(n1574) );
  XNOR U1733 ( .A(n1649), .B(n1646), .Z(n1652) );
  XOR U1734 ( .A(n1653), .B(n1642), .Z(n1649) );
  XOR U1735 ( .A(g_input[113]), .B(state[113]), .Z(n1642) );
  XNOR U1736 ( .A(g_input[115]), .B(state[115]), .Z(n1653) );
  XOR U1737 ( .A(g_input[114]), .B(state[114]), .Z(n1641) );
  XNOR U1738 ( .A(n1654), .B(n1644), .Z(n1537) );
  XOR U1739 ( .A(g_input[117]), .B(state[117]), .Z(n1644) );
  XNOR U1740 ( .A(n1650), .B(n1646), .Z(n1654) );
  XNOR U1741 ( .A(n1655), .B(n1497), .Z(n1646) );
  XOR U1742 ( .A(g_input[112]), .B(state[112]), .Z(n1497) );
  XNOR U1743 ( .A(g_input[118]), .B(state[118]), .Z(n1655) );
  XOR U1744 ( .A(g_input[119]), .B(state[119]), .Z(n1650) );
  XOR U1745 ( .A(n1656), .B(n1657), .Z(o[15]) );
  XNOR U1746 ( .A(n5), .B(n1658), .Z(n1657) );
  XOR U1747 ( .A(g_input[15]), .B(n3), .Z(n1658) );
  IV U1748 ( .A(n1659), .Z(n5) );
  XOR U1749 ( .A(n1660), .B(n4), .Z(n1656) );
  XNOR U1750 ( .A(n1661), .B(n1662), .Z(o[14]) );
  XNOR U1751 ( .A(n1659), .B(g_input[14]), .Z(n1661) );
  XOR U1752 ( .A(n1663), .B(n62), .Z(n1659) );
  XOR U1753 ( .A(n1664), .B(n1665), .Z(o[13]) );
  XOR U1754 ( .A(n1666), .B(n1667), .Z(n1665) );
  XNOR U1755 ( .A(g_input[13]), .B(n1668), .Z(n1667) );
  ANDN U1756 ( .A(n1669), .B(n1670), .Z(n1666) );
  XNOR U1757 ( .A(n1671), .B(n1660), .Z(n1664) );
  XNOR U1758 ( .A(n1672), .B(n1673), .Z(n1660) );
  XNOR U1759 ( .A(n1674), .B(n1675), .Z(n1672) );
  NANDN U1760 ( .B(n1676), .A(n1677), .Z(n1674) );
  XNOR U1761 ( .A(n61), .B(n1678), .Z(n1671) );
  XNOR U1762 ( .A(n1679), .B(n1680), .Z(o[12]) );
  XOR U1763 ( .A(n61), .B(g_input[12]), .Z(n1679) );
  XNOR U1764 ( .A(n1681), .B(n1673), .Z(n61) );
  XNOR U1765 ( .A(n1682), .B(n1683), .Z(n1673) );
  XNOR U1766 ( .A(n1684), .B(n1685), .Z(n1682) );
  NANDN U1767 ( .B(n1686), .A(n1687), .Z(n1684) );
  XOR U1768 ( .A(n1688), .B(n1689), .Z(n1681) );
  ANDN U1769 ( .A(n1690), .B(n1691), .Z(n1689) );
  XOR U1770 ( .A(n1692), .B(n1693), .Z(o[127]) );
  XOR U1771 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U1772 ( .A(n1697), .B(n1698), .Z(n1692) );
  XNOR U1773 ( .A(n1699), .B(n1700), .Z(o[126]) );
  XNOR U1774 ( .A(n1696), .B(g_input[126]), .Z(n1699) );
  XOR U1775 ( .A(n1701), .B(n1702), .Z(o[125]) );
  XOR U1776 ( .A(n1703), .B(n1704), .Z(n1702) );
  XNOR U1777 ( .A(g_input[125]), .B(n1705), .Z(n1704) );
  NOR U1778 ( .A(n1706), .B(n1707), .Z(n1703) );
  XNOR U1779 ( .A(n1708), .B(n1709), .Z(n1701) );
  XOR U1780 ( .A(n1697), .B(n1710), .Z(n1708) );
  XNOR U1781 ( .A(n1711), .B(n1712), .Z(n1697) );
  XNOR U1782 ( .A(n1713), .B(n1714), .Z(n1711) );
  NANDN U1783 ( .B(n1715), .A(n1716), .Z(n1713) );
  XNOR U1784 ( .A(n1717), .B(n1718), .Z(o[124]) );
  XOR U1785 ( .A(n1709), .B(g_input[124]), .Z(n1717) );
  XOR U1786 ( .A(n1719), .B(n1720), .Z(o[123]) );
  XOR U1787 ( .A(n1694), .B(n1721), .Z(n1720) );
  XNOR U1788 ( .A(g_input[123]), .B(n1722), .Z(n1721) );
  XNOR U1789 ( .A(n1700), .B(n1698), .Z(n1719) );
  XNOR U1790 ( .A(n1723), .B(n1724), .Z(n1700) );
  XNOR U1791 ( .A(n1725), .B(n1705), .Z(n1723) );
  NANDN U1792 ( .B(n1726), .A(n1727), .Z(n1705) );
  NANDN U1793 ( .B(n1728), .A(n1729), .Z(n1725) );
  XOR U1794 ( .A(n1718), .B(g_input[122]), .Z(o[122]) );
  XOR U1795 ( .A(n1730), .B(n1731), .Z(n1718) );
  XOR U1796 ( .A(n1732), .B(n1733), .Z(o[121]) );
  XOR U1797 ( .A(g_input[121]), .B(n1696), .Z(n1733) );
  XOR U1798 ( .A(n1722), .B(n1731), .Z(n1696) );
  XNOR U1799 ( .A(n1734), .B(n1710), .Z(n1722) );
  XOR U1800 ( .A(n1735), .B(n1736), .Z(n1734) );
  ANDN U1801 ( .A(n1737), .B(n1738), .Z(n1736) );
  XNOR U1802 ( .A(n1730), .B(n1694), .Z(n1732) );
  XOR U1803 ( .A(n1739), .B(n1724), .Z(n1694) );
  XNOR U1804 ( .A(n1740), .B(n1710), .Z(n1724) );
  XNOR U1805 ( .A(n1741), .B(n1742), .Z(n1710) );
  NOR U1806 ( .A(n1743), .B(n1744), .Z(n1742) );
  XOR U1807 ( .A(n1745), .B(n1741), .Z(n1740) );
  NOR U1808 ( .A(n1746), .B(n1747), .Z(n1741) );
  NANDN U1809 ( .B(n1748), .A(n1749), .Z(n1745) );
  XOR U1810 ( .A(n1735), .B(n1750), .Z(n1739) );
  ANDN U1811 ( .A(n1751), .B(n1715), .Z(n1750) );
  OR U1812 ( .A(n1752), .B(n1753), .Z(n1735) );
  IV U1813 ( .A(n1698), .Z(n1730) );
  XNOR U1814 ( .A(n1754), .B(n1755), .Z(n1698) );
  XNOR U1815 ( .A(n1756), .B(n1757), .Z(n1754) );
  NOR U1816 ( .A(n1758), .B(n1707), .Z(n1757) );
  XNOR U1817 ( .A(n1759), .B(n1709), .Z(o[120]) );
  XOR U1818 ( .A(n1760), .B(n1712), .Z(n1709) );
  XOR U1819 ( .A(n1761), .B(n1755), .Z(n1712) );
  XNOR U1820 ( .A(n1762), .B(n1763), .Z(n1761) );
  NOR U1821 ( .A(n1748), .B(n1764), .Z(n1763) );
  XNOR U1822 ( .A(n1756), .B(n1765), .Z(n1760) );
  NOR U1823 ( .A(n1728), .B(n1766), .Z(n1765) );
  ANDN U1824 ( .A(n1727), .B(n1767), .Z(n1756) );
  XOR U1825 ( .A(n1728), .B(n1707), .Z(n1727) );
  XOR U1826 ( .A(n1731), .B(g_input[120]), .Z(n1759) );
  XNOR U1827 ( .A(n1768), .B(n1755), .Z(n1731) );
  XNOR U1828 ( .A(n1762), .B(n1769), .Z(n1755) );
  NOR U1829 ( .A(n1770), .B(n1744), .Z(n1769) );
  NOR U1830 ( .A(n1746), .B(n1771), .Z(n1762) );
  XNOR U1831 ( .A(n1738), .B(n1707), .Z(n1748) );
  XNOR U1832 ( .A(n1772), .B(n1773), .Z(n1707) );
  ANDN U1833 ( .A(n1774), .B(n1775), .Z(n1773) );
  IV U1834 ( .A(n1776), .Z(n1715) );
  XNOR U1835 ( .A(n1772), .B(n1777), .Z(n1728) );
  NOR U1836 ( .A(n1778), .B(n1779), .Z(n1777) );
  ANDN U1837 ( .A(n1780), .B(n1781), .Z(n1772) );
  XNOR U1838 ( .A(n1782), .B(n1714), .Z(n1768) );
  OR U1839 ( .A(n1752), .B(n1783), .Z(n1714) );
  XOR U1840 ( .A(n1776), .B(n1738), .Z(n1752) );
  XOR U1841 ( .A(n1784), .B(n1785), .Z(n1776) );
  ANDN U1842 ( .A(n1786), .B(n1779), .Z(n1785) );
  OR U1843 ( .A(n1738), .B(n1787), .Z(n1782) );
  XOR U1844 ( .A(n1788), .B(n1784), .Z(n1738) );
  XOR U1845 ( .A(n1779), .B(n1775), .Z(n1780) );
  XNOR U1846 ( .A(n1790), .B(n1791), .Z(n1779) );
  XNOR U1847 ( .A(n1792), .B(n1793), .Z(n1790) );
  NANDN U1848 ( .B(n1794), .A(n1774), .Z(n1792) );
  OR U1849 ( .A(n1775), .B(n1794), .Z(n1788) );
  XOR U1850 ( .A(n1795), .B(n1796), .Z(n1775) );
  XOR U1851 ( .A(n1797), .B(n1798), .Z(n1796) );
  XNOR U1852 ( .A(n1793), .B(n1799), .Z(n1798) );
  ANDN U1853 ( .A(n1786), .B(n1778), .Z(n1799) );
  OR U1854 ( .A(n1781), .B(n1789), .Z(n1793) );
  XNOR U1855 ( .A(n1800), .B(n1786), .Z(n1789) );
  XOR U1856 ( .A(n1774), .B(n1778), .Z(n1781) );
  IV U1857 ( .A(n1797), .Z(n1778) );
  XNOR U1858 ( .A(n1801), .B(n1802), .Z(n1797) );
  XNOR U1859 ( .A(n1787), .B(n1803), .Z(n1802) );
  XNOR U1860 ( .A(n1804), .B(n1805), .Z(n1803) );
  ANDN U1861 ( .A(n1716), .B(n1806), .Z(n1804) );
  XNOR U1862 ( .A(n1807), .B(n1808), .Z(n1801) );
  XOR U1863 ( .A(n1809), .B(n1737), .Z(n1807) );
  XOR U1864 ( .A(n1791), .B(n1786), .Z(n1795) );
  XNOR U1865 ( .A(n1810), .B(n1811), .Z(n1786) );
  XNOR U1866 ( .A(n1812), .B(n1813), .Z(n1811) );
  ANDN U1867 ( .A(n1729), .B(n1766), .Z(n1812) );
  XNOR U1868 ( .A(n1814), .B(n1809), .Z(n1810) );
  XOR U1869 ( .A(n1815), .B(n1816), .Z(n1809) );
  XNOR U1870 ( .A(n1817), .B(n1818), .Z(n1815) );
  NANDN U1871 ( .B(n1764), .A(n1749), .Z(n1817) );
  XNOR U1872 ( .A(n1800), .B(n1774), .Z(n1791) );
  XNOR U1873 ( .A(n1819), .B(n1820), .Z(n1774) );
  XOR U1874 ( .A(n1716), .B(n1821), .Z(n1820) );
  XNOR U1875 ( .A(n1822), .B(n1805), .Z(n1821) );
  OR U1876 ( .A(n1753), .B(n1783), .Z(n1805) );
  XNOR U1877 ( .A(n1751), .B(n1737), .Z(n1753) );
  IV U1878 ( .A(n1806), .Z(n1751) );
  ANDN U1879 ( .A(n1737), .B(n1787), .Z(n1822) );
  XNOR U1880 ( .A(n1823), .B(n1814), .Z(n1819) );
  XOR U1881 ( .A(n1816), .B(n1806), .Z(n1823) );
  IV U1882 ( .A(n1794), .Z(n1800) );
  XOR U1883 ( .A(n1824), .B(n1825), .Z(n1794) );
  XOR U1884 ( .A(n1816), .B(n1826), .Z(n1825) );
  XNOR U1885 ( .A(n1827), .B(n1813), .Z(n1826) );
  OR U1886 ( .A(n1726), .B(n1767), .Z(n1813) );
  XNOR U1887 ( .A(n1766), .B(n1758), .Z(n1767) );
  XNOR U1888 ( .A(n1828), .B(n1729), .Z(n1726) );
  ANDN U1889 ( .A(n1829), .B(n1706), .Z(n1827) );
  XNOR U1890 ( .A(n1818), .B(n1830), .Z(n1816) );
  ANDN U1891 ( .A(n1831), .B(n1743), .Z(n1830) );
  OR U1892 ( .A(n1771), .B(n1747), .Z(n1818) );
  XOR U1893 ( .A(n1743), .B(n1749), .Z(n1747) );
  XNOR U1894 ( .A(n1706), .B(n1737), .Z(n1749) );
  XNOR U1895 ( .A(n1832), .B(n1729), .Z(n1737) );
  XNOR U1896 ( .A(n1833), .B(n1834), .Z(n1832) );
  XOR U1897 ( .A(n1806), .B(n1729), .Z(n1743) );
  XOR U1898 ( .A(n1835), .B(n1836), .Z(n1806) );
  XNOR U1899 ( .A(n1837), .B(n1838), .Z(n1835) );
  XOR U1900 ( .A(n1831), .B(n1764), .Z(n1771) );
  XOR U1901 ( .A(n1829), .B(n1787), .Z(n1764) );
  XOR U1902 ( .A(n1839), .B(n1840), .Z(n1787) );
  XNOR U1903 ( .A(n1841), .B(n1716), .Z(n1840) );
  XNOR U1904 ( .A(n1842), .B(n1837), .Z(n1839) );
  XOR U1905 ( .A(g_input[124]), .B(state[124]), .Z(n1837) );
  IV U1906 ( .A(n1770), .Z(n1831) );
  XOR U1907 ( .A(n1766), .B(n1716), .Z(n1770) );
  XNOR U1908 ( .A(n1814), .B(n1808), .Z(n1824) );
  XNOR U1909 ( .A(n1828), .B(n1829), .Z(n1808) );
  IV U1910 ( .A(n1758), .Z(n1829) );
  IV U1911 ( .A(n1706), .Z(n1828) );
  XOR U1912 ( .A(n1843), .B(n1836), .Z(n1706) );
  XNOR U1913 ( .A(n1834), .B(n1838), .Z(n1843) );
  XOR U1914 ( .A(n1729), .B(n1766), .Z(n1814) );
  XNOR U1915 ( .A(n1833), .B(n1844), .Z(n1766) );
  XNOR U1916 ( .A(n1841), .B(n1838), .Z(n1844) );
  XOR U1917 ( .A(n1845), .B(n1834), .Z(n1841) );
  XOR U1918 ( .A(g_input[121]), .B(state[121]), .Z(n1834) );
  XNOR U1919 ( .A(g_input[123]), .B(state[123]), .Z(n1845) );
  XOR U1920 ( .A(g_input[122]), .B(state[122]), .Z(n1833) );
  XNOR U1921 ( .A(n1846), .B(n1836), .Z(n1729) );
  XOR U1922 ( .A(g_input[125]), .B(state[125]), .Z(n1836) );
  XNOR U1923 ( .A(n1842), .B(n1838), .Z(n1846) );
  XNOR U1924 ( .A(n1847), .B(n1716), .Z(n1838) );
  XOR U1925 ( .A(g_input[120]), .B(state[120]), .Z(n1716) );
  XNOR U1926 ( .A(g_input[126]), .B(state[126]), .Z(n1847) );
  XOR U1927 ( .A(g_input[127]), .B(state[127]), .Z(n1842) );
  XOR U1928 ( .A(n1848), .B(n1849), .Z(o[11]) );
  XNOR U1929 ( .A(n1663), .B(n1850), .Z(n1849) );
  XOR U1930 ( .A(g_input[11]), .B(n3), .Z(n1850) );
  XNOR U1931 ( .A(n1851), .B(n1678), .Z(n1663) );
  XNOR U1932 ( .A(n1852), .B(n1853), .Z(n1851) );
  NANDN U1933 ( .B(n1854), .A(n1855), .Z(n1852) );
  XOR U1934 ( .A(n1662), .B(n4), .Z(n1848) );
  XOR U1935 ( .A(n1856), .B(n1857), .Z(n4) );
  XOR U1936 ( .A(n1853), .B(n1858), .Z(n1856) );
  ANDN U1937 ( .A(n1677), .B(n1859), .Z(n1858) );
  OR U1938 ( .A(n1860), .B(n1861), .Z(n1853) );
  XNOR U1939 ( .A(n1862), .B(n1857), .Z(n1662) );
  XNOR U1940 ( .A(n1863), .B(n1678), .Z(n1857) );
  XNOR U1941 ( .A(n1864), .B(n1865), .Z(n1678) );
  NOR U1942 ( .A(n1866), .B(n1867), .Z(n1865) );
  XNOR U1943 ( .A(n1864), .B(n1868), .Z(n1863) );
  ANDN U1944 ( .A(n1869), .B(n1686), .Z(n1868) );
  NOR U1945 ( .A(n1870), .B(n1871), .Z(n1864) );
  XNOR U1946 ( .A(n1872), .B(n1668), .Z(n1862) );
  OR U1947 ( .A(n1873), .B(n1874), .Z(n1668) );
  NANDN U1948 ( .B(n1875), .A(n1690), .Z(n1872) );
  XOR U1949 ( .A(n1876), .B(n1877), .Z(o[119]) );
  XOR U1950 ( .A(n1878), .B(n1879), .Z(n1877) );
  XOR U1951 ( .A(n1881), .B(n1882), .Z(n1876) );
  XNOR U1952 ( .A(n1883), .B(n1884), .Z(o[118]) );
  XNOR U1953 ( .A(n1880), .B(g_input[118]), .Z(n1883) );
  XOR U1954 ( .A(n1885), .B(n1886), .Z(o[117]) );
  XOR U1955 ( .A(n1887), .B(n1888), .Z(n1886) );
  XNOR U1956 ( .A(g_input[117]), .B(n1889), .Z(n1888) );
  NOR U1957 ( .A(n1890), .B(n1891), .Z(n1887) );
  XNOR U1958 ( .A(n1892), .B(n1893), .Z(n1885) );
  XOR U1959 ( .A(n1881), .B(n1894), .Z(n1892) );
  XNOR U1960 ( .A(n1895), .B(n1896), .Z(n1881) );
  XNOR U1961 ( .A(n1897), .B(n1898), .Z(n1895) );
  NANDN U1962 ( .B(n1899), .A(n1900), .Z(n1897) );
  XNOR U1963 ( .A(n1901), .B(n1902), .Z(o[116]) );
  XOR U1964 ( .A(n1893), .B(g_input[116]), .Z(n1901) );
  XOR U1965 ( .A(n1903), .B(n1904), .Z(o[115]) );
  XOR U1966 ( .A(n1878), .B(n1905), .Z(n1904) );
  XNOR U1967 ( .A(g_input[115]), .B(n1906), .Z(n1905) );
  XNOR U1968 ( .A(n1884), .B(n1882), .Z(n1903) );
  XNOR U1969 ( .A(n1907), .B(n1908), .Z(n1884) );
  XNOR U1970 ( .A(n1909), .B(n1889), .Z(n1907) );
  NANDN U1971 ( .B(n1910), .A(n1911), .Z(n1889) );
  NANDN U1972 ( .B(n1912), .A(n1913), .Z(n1909) );
  XOR U1973 ( .A(n1902), .B(g_input[114]), .Z(o[114]) );
  XOR U1974 ( .A(n1914), .B(n1915), .Z(n1902) );
  XOR U1975 ( .A(n1916), .B(n1917), .Z(o[113]) );
  XOR U1976 ( .A(g_input[113]), .B(n1880), .Z(n1917) );
  XOR U1977 ( .A(n1906), .B(n1915), .Z(n1880) );
  XNOR U1978 ( .A(n1918), .B(n1894), .Z(n1906) );
  XOR U1979 ( .A(n1919), .B(n1920), .Z(n1918) );
  ANDN U1980 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1981 ( .A(n1914), .B(n1878), .Z(n1916) );
  XOR U1982 ( .A(n1923), .B(n1908), .Z(n1878) );
  XNOR U1983 ( .A(n1924), .B(n1894), .Z(n1908) );
  XNOR U1984 ( .A(n1925), .B(n1926), .Z(n1894) );
  NOR U1985 ( .A(n1927), .B(n1928), .Z(n1926) );
  XOR U1986 ( .A(n1929), .B(n1925), .Z(n1924) );
  NOR U1987 ( .A(n1930), .B(n1931), .Z(n1925) );
  NANDN U1988 ( .B(n1932), .A(n1933), .Z(n1929) );
  XOR U1989 ( .A(n1919), .B(n1934), .Z(n1923) );
  ANDN U1990 ( .A(n1935), .B(n1899), .Z(n1934) );
  OR U1991 ( .A(n1936), .B(n1937), .Z(n1919) );
  IV U1992 ( .A(n1882), .Z(n1914) );
  XNOR U1993 ( .A(n1938), .B(n1939), .Z(n1882) );
  XNOR U1994 ( .A(n1940), .B(n1941), .Z(n1938) );
  NOR U1995 ( .A(n1942), .B(n1891), .Z(n1941) );
  XNOR U1996 ( .A(n1943), .B(n1893), .Z(o[112]) );
  XOR U1997 ( .A(n1944), .B(n1896), .Z(n1893) );
  XOR U1998 ( .A(n1945), .B(n1939), .Z(n1896) );
  XNOR U1999 ( .A(n1946), .B(n1947), .Z(n1945) );
  NOR U2000 ( .A(n1932), .B(n1948), .Z(n1947) );
  XNOR U2001 ( .A(n1940), .B(n1949), .Z(n1944) );
  NOR U2002 ( .A(n1912), .B(n1950), .Z(n1949) );
  ANDN U2003 ( .A(n1911), .B(n1951), .Z(n1940) );
  XOR U2004 ( .A(n1912), .B(n1891), .Z(n1911) );
  XOR U2005 ( .A(n1915), .B(g_input[112]), .Z(n1943) );
  XNOR U2006 ( .A(n1952), .B(n1939), .Z(n1915) );
  XNOR U2007 ( .A(n1946), .B(n1953), .Z(n1939) );
  NOR U2008 ( .A(n1954), .B(n1928), .Z(n1953) );
  NOR U2009 ( .A(n1930), .B(n1955), .Z(n1946) );
  XNOR U2010 ( .A(n1922), .B(n1891), .Z(n1932) );
  XNOR U2011 ( .A(n1956), .B(n1957), .Z(n1891) );
  ANDN U2012 ( .A(n1958), .B(n1959), .Z(n1957) );
  IV U2013 ( .A(n1960), .Z(n1899) );
  XNOR U2014 ( .A(n1956), .B(n1961), .Z(n1912) );
  NOR U2015 ( .A(n1962), .B(n1963), .Z(n1961) );
  ANDN U2016 ( .A(n1964), .B(n1965), .Z(n1956) );
  XNOR U2017 ( .A(n1966), .B(n1898), .Z(n1952) );
  OR U2018 ( .A(n1936), .B(n1967), .Z(n1898) );
  XOR U2019 ( .A(n1960), .B(n1922), .Z(n1936) );
  XOR U2020 ( .A(n1968), .B(n1969), .Z(n1960) );
  ANDN U2021 ( .A(n1970), .B(n1963), .Z(n1969) );
  OR U2022 ( .A(n1922), .B(n1971), .Z(n1966) );
  XOR U2023 ( .A(n1972), .B(n1968), .Z(n1922) );
  XOR U2024 ( .A(n1963), .B(n1959), .Z(n1964) );
  XNOR U2025 ( .A(n1974), .B(n1975), .Z(n1963) );
  XNOR U2026 ( .A(n1976), .B(n1977), .Z(n1974) );
  NANDN U2027 ( .B(n1978), .A(n1958), .Z(n1976) );
  OR U2028 ( .A(n1959), .B(n1978), .Z(n1972) );
  XOR U2029 ( .A(n1979), .B(n1980), .Z(n1959) );
  XOR U2030 ( .A(n1981), .B(n1982), .Z(n1980) );
  XNOR U2031 ( .A(n1977), .B(n1983), .Z(n1982) );
  ANDN U2032 ( .A(n1970), .B(n1962), .Z(n1983) );
  OR U2033 ( .A(n1965), .B(n1973), .Z(n1977) );
  XNOR U2034 ( .A(n1984), .B(n1970), .Z(n1973) );
  XOR U2035 ( .A(n1958), .B(n1962), .Z(n1965) );
  IV U2036 ( .A(n1981), .Z(n1962) );
  XNOR U2037 ( .A(n1985), .B(n1986), .Z(n1981) );
  XNOR U2038 ( .A(n1971), .B(n1987), .Z(n1986) );
  XNOR U2039 ( .A(n1988), .B(n1989), .Z(n1987) );
  ANDN U2040 ( .A(n1900), .B(n1990), .Z(n1988) );
  XNOR U2041 ( .A(n1991), .B(n1992), .Z(n1985) );
  XOR U2042 ( .A(n1993), .B(n1921), .Z(n1991) );
  XOR U2043 ( .A(n1975), .B(n1970), .Z(n1979) );
  XNOR U2044 ( .A(n1994), .B(n1995), .Z(n1970) );
  XNOR U2045 ( .A(n1996), .B(n1997), .Z(n1995) );
  ANDN U2046 ( .A(n1913), .B(n1950), .Z(n1996) );
  XNOR U2047 ( .A(n1998), .B(n1993), .Z(n1994) );
  XOR U2048 ( .A(n1999), .B(n2000), .Z(n1993) );
  XNOR U2049 ( .A(n2001), .B(n2002), .Z(n1999) );
  NANDN U2050 ( .B(n1948), .A(n1933), .Z(n2001) );
  XNOR U2051 ( .A(n1984), .B(n1958), .Z(n1975) );
  XNOR U2052 ( .A(n2003), .B(n2004), .Z(n1958) );
  XOR U2053 ( .A(n1900), .B(n2005), .Z(n2004) );
  XNOR U2054 ( .A(n2006), .B(n1989), .Z(n2005) );
  OR U2055 ( .A(n1937), .B(n1967), .Z(n1989) );
  XNOR U2056 ( .A(n1935), .B(n1921), .Z(n1937) );
  IV U2057 ( .A(n1990), .Z(n1935) );
  ANDN U2058 ( .A(n1921), .B(n1971), .Z(n2006) );
  XNOR U2059 ( .A(n2007), .B(n1998), .Z(n2003) );
  XOR U2060 ( .A(n2000), .B(n1990), .Z(n2007) );
  IV U2061 ( .A(n1978), .Z(n1984) );
  XOR U2062 ( .A(n2008), .B(n2009), .Z(n1978) );
  XOR U2063 ( .A(n2000), .B(n2010), .Z(n2009) );
  XNOR U2064 ( .A(n2011), .B(n1997), .Z(n2010) );
  OR U2065 ( .A(n1910), .B(n1951), .Z(n1997) );
  XNOR U2066 ( .A(n1950), .B(n1942), .Z(n1951) );
  XNOR U2067 ( .A(n2012), .B(n1913), .Z(n1910) );
  ANDN U2068 ( .A(n2013), .B(n1890), .Z(n2011) );
  XNOR U2069 ( .A(n2002), .B(n2014), .Z(n2000) );
  ANDN U2070 ( .A(n2015), .B(n1927), .Z(n2014) );
  OR U2071 ( .A(n1955), .B(n1931), .Z(n2002) );
  XOR U2072 ( .A(n1927), .B(n1933), .Z(n1931) );
  XNOR U2073 ( .A(n1890), .B(n1921), .Z(n1933) );
  XNOR U2074 ( .A(n2016), .B(n1913), .Z(n1921) );
  XOR U2075 ( .A(n2017), .B(n2018), .Z(n2016) );
  IV U2076 ( .A(n2012), .Z(n1890) );
  XOR U2077 ( .A(n1990), .B(n1913), .Z(n1927) );
  XOR U2078 ( .A(n2019), .B(n2020), .Z(n1990) );
  XOR U2079 ( .A(n2021), .B(n2022), .Z(n2019) );
  XOR U2080 ( .A(n2015), .B(n1948), .Z(n1955) );
  XOR U2081 ( .A(n2013), .B(n1971), .Z(n1948) );
  XOR U2082 ( .A(n2023), .B(n2024), .Z(n1971) );
  XNOR U2083 ( .A(n2025), .B(n1900), .Z(n2024) );
  XNOR U2084 ( .A(n2026), .B(n2021), .Z(n2023) );
  XNOR U2085 ( .A(g_input[84]), .B(state[84]), .Z(n2021) );
  IV U2086 ( .A(n1954), .Z(n2015) );
  XOR U2087 ( .A(n1950), .B(n1900), .Z(n1954) );
  XNOR U2088 ( .A(n1998), .B(n1992), .Z(n2008) );
  XNOR U2089 ( .A(n2012), .B(n2013), .Z(n1992) );
  IV U2090 ( .A(n1942), .Z(n2013) );
  XOR U2091 ( .A(n2027), .B(n2022), .Z(n1942) );
  XOR U2092 ( .A(n2028), .B(n2027), .Z(n2012) );
  IV U2093 ( .A(n2020), .Z(n2027) );
  XNOR U2094 ( .A(n2018), .B(n2022), .Z(n2028) );
  XOR U2095 ( .A(n1913), .B(n1950), .Z(n1998) );
  XOR U2096 ( .A(n2017), .B(n2029), .Z(n1950) );
  XNOR U2097 ( .A(n2025), .B(n2022), .Z(n2029) );
  XOR U2098 ( .A(n2030), .B(n2018), .Z(n2025) );
  XOR U2099 ( .A(g_input[81]), .B(state[81]), .Z(n2018) );
  XNOR U2100 ( .A(g_input[83]), .B(state[83]), .Z(n2030) );
  XNOR U2101 ( .A(g_input[82]), .B(state[82]), .Z(n2017) );
  XNOR U2102 ( .A(n2031), .B(n2020), .Z(n1913) );
  XOR U2103 ( .A(g_input[85]), .B(state[85]), .Z(n2020) );
  XOR U2104 ( .A(n2026), .B(n2022), .Z(n2031) );
  XNOR U2105 ( .A(n2032), .B(n1900), .Z(n2022) );
  XOR U2106 ( .A(g_input[80]), .B(state[80]), .Z(n1900) );
  XNOR U2107 ( .A(g_input[86]), .B(state[86]), .Z(n2032) );
  XNOR U2108 ( .A(g_input[87]), .B(state[87]), .Z(n2026) );
  XOR U2109 ( .A(n2033), .B(n2034), .Z(o[111]) );
  XOR U2110 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U2111 ( .A(n2038), .B(n2039), .Z(n2033) );
  XNOR U2112 ( .A(n2040), .B(n2041), .Z(o[110]) );
  XNOR U2113 ( .A(n2037), .B(g_input[110]), .Z(n2040) );
  XOR U2114 ( .A(n1680), .B(g_input[10]), .Z(o[10]) );
  XOR U2115 ( .A(n62), .B(n3), .Z(n1680) );
  XOR U2116 ( .A(n2042), .B(n1683), .Z(n3) );
  XOR U2117 ( .A(n1688), .B(n2043), .Z(n2042) );
  ANDN U2118 ( .A(n2044), .B(n1670), .Z(n2043) );
  OR U2119 ( .A(n2045), .B(n1873), .Z(n1688) );
  XNOR U2120 ( .A(n2046), .B(n1683), .Z(n62) );
  XOR U2121 ( .A(n1685), .B(n2047), .Z(n1683) );
  NOR U2122 ( .A(n1866), .B(n2048), .Z(n2047) );
  OR U2123 ( .A(n1871), .B(n2049), .Z(n1685) );
  XNOR U2124 ( .A(n1686), .B(n1866), .Z(n1871) );
  XNOR U2125 ( .A(n1690), .B(n1677), .Z(n1866) );
  XOR U2126 ( .A(n2050), .B(n2051), .Z(n1690) );
  NOR U2127 ( .A(n2052), .B(n2053), .Z(n2051) );
  XOR U2128 ( .A(n1855), .B(n1670), .Z(n1686) );
  XNOR U2129 ( .A(n2050), .B(n2054), .Z(n1670) );
  ANDN U2130 ( .A(n2055), .B(n2056), .Z(n2054) );
  AND U2131 ( .A(n2057), .B(n2058), .Z(n2050) );
  XNOR U2132 ( .A(n2059), .B(n1675), .Z(n2046) );
  OR U2133 ( .A(n1861), .B(n2060), .Z(n1675) );
  XNOR U2134 ( .A(n1855), .B(n1677), .Z(n1861) );
  XNOR U2135 ( .A(n2061), .B(n2062), .Z(n1677) );
  NOR U2136 ( .A(n2063), .B(n2053), .Z(n2062) );
  NANDN U2137 ( .B(n2064), .A(n1855), .Z(n2059) );
  XOR U2138 ( .A(n2065), .B(n2061), .Z(n1855) );
  NANDN U2139 ( .B(n2066), .A(n2057), .Z(n2061) );
  XNOR U2140 ( .A(n2053), .B(n2055), .Z(n2057) );
  XNOR U2141 ( .A(n2067), .B(n2068), .Z(n2053) );
  XNOR U2142 ( .A(n2069), .B(n2070), .Z(n2067) );
  NANDN U2143 ( .B(n2071), .A(n2072), .Z(n2069) );
  NANDN U2144 ( .B(n2071), .A(n2055), .Z(n2065) );
  XNOR U2145 ( .A(n2073), .B(n2074), .Z(n2055) );
  XOR U2146 ( .A(n2075), .B(n2076), .Z(n2074) );
  XNOR U2147 ( .A(n2070), .B(n2077), .Z(n2076) );
  ANDN U2148 ( .A(n2078), .B(n2063), .Z(n2077) );
  IV U2149 ( .A(n2075), .Z(n2063) );
  NANDN U2150 ( .B(n2066), .A(n2058), .Z(n2070) );
  XOR U2151 ( .A(n2056), .B(n2052), .Z(n2058) );
  XNOR U2152 ( .A(n2079), .B(n2080), .Z(n2075) );
  XNOR U2153 ( .A(n2081), .B(n2082), .Z(n2080) );
  NOR U2154 ( .A(n1875), .B(n1691), .Z(n2081) );
  XOR U2155 ( .A(n2083), .B(n2084), .Z(n2079) );
  XNOR U2156 ( .A(n2068), .B(n2052), .Z(n2073) );
  IV U2157 ( .A(n2078), .Z(n2052) );
  XNOR U2158 ( .A(n2085), .B(n2086), .Z(n2078) );
  XNOR U2159 ( .A(n2064), .B(n2087), .Z(n2086) );
  XNOR U2160 ( .A(n2088), .B(n2089), .Z(n2087) );
  ANDN U2161 ( .A(n2090), .B(n1859), .Z(n2088) );
  XOR U2162 ( .A(n2091), .B(n2092), .Z(n2085) );
  XNOR U2163 ( .A(n2084), .B(n1854), .Z(n2091) );
  XOR U2164 ( .A(n2093), .B(n2094), .Z(n2084) );
  XNOR U2165 ( .A(n2095), .B(n2096), .Z(n2093) );
  NAND U2166 ( .A(n1687), .B(n1869), .Z(n2095) );
  XOR U2167 ( .A(n2072), .B(n2071), .Z(n2068) );
  IV U2168 ( .A(n2056), .Z(n2072) );
  XOR U2169 ( .A(n2097), .B(n2098), .Z(n2056) );
  XNOR U2170 ( .A(n1676), .B(n2099), .Z(n2098) );
  XNOR U2171 ( .A(n2100), .B(n2089), .Z(n2099) );
  OR U2172 ( .A(n1860), .B(n2060), .Z(n2089) );
  XNOR U2173 ( .A(n2101), .B(n2090), .Z(n2060) );
  ANDN U2174 ( .A(n2101), .B(n1854), .Z(n2100) );
  XOR U2175 ( .A(n2094), .B(n1859), .Z(n2102) );
  XOR U2176 ( .A(n2103), .B(n2104), .Z(n2071) );
  XOR U2177 ( .A(n2094), .B(n2105), .Z(n2104) );
  XNOR U2178 ( .A(n2106), .B(n2082), .Z(n2105) );
  OR U2179 ( .A(n1874), .B(n2045), .Z(n2082) );
  XOR U2180 ( .A(n2044), .B(n1691), .Z(n2045) );
  XNOR U2181 ( .A(n1669), .B(n2107), .Z(n1874) );
  ANDN U2182 ( .A(n1669), .B(n2108), .Z(n2106) );
  XNOR U2183 ( .A(n2096), .B(n2109), .Z(n2094) );
  NOR U2184 ( .A(n2048), .B(n1867), .Z(n2109) );
  OR U2185 ( .A(n2049), .B(n1870), .Z(n2096) );
  XOR U2186 ( .A(n1869), .B(n1867), .Z(n1870) );
  XOR U2187 ( .A(n2110), .B(n2111), .Z(n1859) );
  XOR U2188 ( .A(n2112), .B(n2113), .Z(n2110) );
  XNOR U2189 ( .A(n1854), .B(n1669), .Z(n1869) );
  XOR U2190 ( .A(n2114), .B(n2107), .Z(n1854) );
  IV U2191 ( .A(n1875), .Z(n2107) );
  XNOR U2192 ( .A(n2115), .B(n2116), .Z(n2114) );
  XOR U2193 ( .A(n1687), .B(n2048), .Z(n2049) );
  XOR U2194 ( .A(n1691), .B(n2090), .Z(n2048) );
  XNOR U2195 ( .A(n2108), .B(n2101), .Z(n1687) );
  IV U2196 ( .A(n2064), .Z(n2101) );
  IV U2197 ( .A(n2044), .Z(n2108) );
  XNOR U2198 ( .A(n2092), .B(n2083), .Z(n2103) );
  XOR U2199 ( .A(n1875), .B(n1691), .Z(n2083) );
  XNOR U2200 ( .A(n2117), .B(n2113), .Z(n1691) );
  XNOR U2201 ( .A(n2116), .B(n2118), .Z(n2117) );
  XOR U2202 ( .A(g_input[74]), .B(state[74]), .Z(n2116) );
  XOR U2203 ( .A(n2119), .B(n2111), .Z(n1875) );
  XOR U2204 ( .A(n2120), .B(n2113), .Z(n2119) );
  XOR U2205 ( .A(n1669), .B(n2044), .Z(n2092) );
  XNOR U2206 ( .A(n2121), .B(n2111), .Z(n1669) );
  XOR U2207 ( .A(g_input[77]), .B(state[77]), .Z(n2111) );
  XOR U2208 ( .A(n2115), .B(n2113), .Z(n2121) );
  XOR U2209 ( .A(n2122), .B(n2090), .Z(n2113) );
  XNOR U2210 ( .A(g_input[78]), .B(state[78]), .Z(n2122) );
  XOR U2211 ( .A(n2123), .B(n2124), .Z(n2064) );
  XNOR U2212 ( .A(n1676), .B(n2118), .Z(n2124) );
  XNOR U2213 ( .A(n2125), .B(n2115), .Z(n2118) );
  XOR U2214 ( .A(g_input[73]), .B(state[73]), .Z(n2115) );
  XNOR U2215 ( .A(g_input[75]), .B(state[75]), .Z(n2125) );
  IV U2216 ( .A(n2090), .Z(n1676) );
  XOR U2217 ( .A(g_input[72]), .B(state[72]), .Z(n2090) );
  XNOR U2218 ( .A(n2120), .B(n2112), .Z(n2123) );
  XOR U2219 ( .A(g_input[76]), .B(state[76]), .Z(n2112) );
  XOR U2220 ( .A(g_input[79]), .B(state[79]), .Z(n2120) );
  XOR U2221 ( .A(n2126), .B(n2127), .Z(o[109]) );
  XOR U2222 ( .A(n2128), .B(n2129), .Z(n2127) );
  XNOR U2223 ( .A(g_input[109]), .B(n2130), .Z(n2129) );
  NOR U2224 ( .A(n2131), .B(n2132), .Z(n2128) );
  XNOR U2225 ( .A(n2133), .B(n2134), .Z(n2126) );
  XOR U2226 ( .A(n2038), .B(n2135), .Z(n2133) );
  XNOR U2227 ( .A(n2136), .B(n2137), .Z(n2038) );
  XNOR U2228 ( .A(n2138), .B(n2139), .Z(n2136) );
  NANDN U2229 ( .B(n2140), .A(n2141), .Z(n2138) );
  XNOR U2230 ( .A(n2142), .B(n2143), .Z(o[108]) );
  XOR U2231 ( .A(n2134), .B(g_input[108]), .Z(n2142) );
  XOR U2232 ( .A(n2144), .B(n2145), .Z(o[107]) );
  XOR U2233 ( .A(n2035), .B(n2146), .Z(n2145) );
  XNOR U2234 ( .A(g_input[107]), .B(n2147), .Z(n2146) );
  XNOR U2235 ( .A(n2041), .B(n2039), .Z(n2144) );
  XNOR U2236 ( .A(n2148), .B(n2149), .Z(n2041) );
  XNOR U2237 ( .A(n2150), .B(n2130), .Z(n2148) );
  NANDN U2238 ( .B(n2151), .A(n2152), .Z(n2130) );
  NANDN U2239 ( .B(n2153), .A(n2154), .Z(n2150) );
  XOR U2240 ( .A(n2143), .B(g_input[106]), .Z(o[106]) );
  XOR U2241 ( .A(n2155), .B(n2156), .Z(n2143) );
  XOR U2242 ( .A(n2157), .B(n2158), .Z(o[105]) );
  XOR U2243 ( .A(g_input[105]), .B(n2037), .Z(n2158) );
  XOR U2244 ( .A(n2147), .B(n2156), .Z(n2037) );
  XNOR U2245 ( .A(n2159), .B(n2135), .Z(n2147) );
  XOR U2246 ( .A(n2160), .B(n2161), .Z(n2159) );
  ANDN U2247 ( .A(n2162), .B(n2163), .Z(n2161) );
  XNOR U2248 ( .A(n2155), .B(n2035), .Z(n2157) );
  XOR U2249 ( .A(n2164), .B(n2149), .Z(n2035) );
  XNOR U2250 ( .A(n2165), .B(n2135), .Z(n2149) );
  XNOR U2251 ( .A(n2166), .B(n2167), .Z(n2135) );
  NOR U2252 ( .A(n2168), .B(n2169), .Z(n2167) );
  XOR U2253 ( .A(n2170), .B(n2166), .Z(n2165) );
  NOR U2254 ( .A(n2171), .B(n2172), .Z(n2166) );
  NANDN U2255 ( .B(n2173), .A(n2174), .Z(n2170) );
  XOR U2256 ( .A(n2160), .B(n2175), .Z(n2164) );
  ANDN U2257 ( .A(n2176), .B(n2140), .Z(n2175) );
  OR U2258 ( .A(n2177), .B(n2178), .Z(n2160) );
  IV U2259 ( .A(n2039), .Z(n2155) );
  XNOR U2260 ( .A(n2179), .B(n2180), .Z(n2039) );
  XNOR U2261 ( .A(n2181), .B(n2182), .Z(n2179) );
  NOR U2262 ( .A(n2183), .B(n2132), .Z(n2182) );
  XNOR U2263 ( .A(n2184), .B(n2134), .Z(o[104]) );
  XOR U2264 ( .A(n2185), .B(n2137), .Z(n2134) );
  XOR U2265 ( .A(n2186), .B(n2180), .Z(n2137) );
  XNOR U2266 ( .A(n2187), .B(n2188), .Z(n2186) );
  NOR U2267 ( .A(n2173), .B(n2189), .Z(n2188) );
  XNOR U2268 ( .A(n2181), .B(n2190), .Z(n2185) );
  NOR U2269 ( .A(n2153), .B(n2191), .Z(n2190) );
  ANDN U2270 ( .A(n2152), .B(n2192), .Z(n2181) );
  XOR U2271 ( .A(n2153), .B(n2132), .Z(n2152) );
  XOR U2272 ( .A(n2156), .B(g_input[104]), .Z(n2184) );
  XNOR U2273 ( .A(n2193), .B(n2180), .Z(n2156) );
  XNOR U2274 ( .A(n2187), .B(n2194), .Z(n2180) );
  NOR U2275 ( .A(n2195), .B(n2169), .Z(n2194) );
  NOR U2276 ( .A(n2171), .B(n2196), .Z(n2187) );
  XNOR U2277 ( .A(n2163), .B(n2132), .Z(n2173) );
  XNOR U2278 ( .A(n2197), .B(n2198), .Z(n2132) );
  ANDN U2279 ( .A(n2199), .B(n2200), .Z(n2198) );
  IV U2280 ( .A(n2201), .Z(n2140) );
  XNOR U2281 ( .A(n2197), .B(n2202), .Z(n2153) );
  NOR U2282 ( .A(n2203), .B(n2204), .Z(n2202) );
  ANDN U2283 ( .A(n2205), .B(n2206), .Z(n2197) );
  XNOR U2284 ( .A(n2207), .B(n2139), .Z(n2193) );
  OR U2285 ( .A(n2177), .B(n2208), .Z(n2139) );
  XOR U2286 ( .A(n2201), .B(n2163), .Z(n2177) );
  XOR U2287 ( .A(n2209), .B(n2210), .Z(n2201) );
  ANDN U2288 ( .A(n2211), .B(n2204), .Z(n2210) );
  OR U2289 ( .A(n2163), .B(n2212), .Z(n2207) );
  XOR U2290 ( .A(n2213), .B(n2209), .Z(n2163) );
  XOR U2291 ( .A(n2204), .B(n2200), .Z(n2205) );
  XNOR U2292 ( .A(n2215), .B(n2216), .Z(n2204) );
  XNOR U2293 ( .A(n2217), .B(n2218), .Z(n2215) );
  NANDN U2294 ( .B(n2219), .A(n2199), .Z(n2217) );
  OR U2295 ( .A(n2200), .B(n2219), .Z(n2213) );
  XOR U2296 ( .A(n2220), .B(n2221), .Z(n2200) );
  XOR U2297 ( .A(n2222), .B(n2223), .Z(n2221) );
  XNOR U2298 ( .A(n2218), .B(n2224), .Z(n2223) );
  ANDN U2299 ( .A(n2211), .B(n2203), .Z(n2224) );
  OR U2300 ( .A(n2206), .B(n2214), .Z(n2218) );
  XNOR U2301 ( .A(n2225), .B(n2211), .Z(n2214) );
  XOR U2302 ( .A(n2199), .B(n2203), .Z(n2206) );
  IV U2303 ( .A(n2222), .Z(n2203) );
  XNOR U2304 ( .A(n2226), .B(n2227), .Z(n2222) );
  XNOR U2305 ( .A(n2212), .B(n2228), .Z(n2227) );
  XNOR U2306 ( .A(n2229), .B(n2230), .Z(n2228) );
  ANDN U2307 ( .A(n2141), .B(n2231), .Z(n2229) );
  XNOR U2308 ( .A(n2232), .B(n2233), .Z(n2226) );
  XOR U2309 ( .A(n2234), .B(n2162), .Z(n2232) );
  XOR U2310 ( .A(n2216), .B(n2211), .Z(n2220) );
  XNOR U2311 ( .A(n2235), .B(n2236), .Z(n2211) );
  XNOR U2312 ( .A(n2237), .B(n2238), .Z(n2236) );
  ANDN U2313 ( .A(n2154), .B(n2191), .Z(n2237) );
  XNOR U2314 ( .A(n2239), .B(n2234), .Z(n2235) );
  XOR U2315 ( .A(n2240), .B(n2241), .Z(n2234) );
  XNOR U2316 ( .A(n2242), .B(n2243), .Z(n2240) );
  NANDN U2317 ( .B(n2189), .A(n2174), .Z(n2242) );
  XNOR U2318 ( .A(n2225), .B(n2199), .Z(n2216) );
  XNOR U2319 ( .A(n2244), .B(n2245), .Z(n2199) );
  XOR U2320 ( .A(n2141), .B(n2246), .Z(n2245) );
  XNOR U2321 ( .A(n2247), .B(n2230), .Z(n2246) );
  OR U2322 ( .A(n2178), .B(n2208), .Z(n2230) );
  XNOR U2323 ( .A(n2176), .B(n2162), .Z(n2178) );
  IV U2324 ( .A(n2231), .Z(n2176) );
  ANDN U2325 ( .A(n2162), .B(n2212), .Z(n2247) );
  XNOR U2326 ( .A(n2248), .B(n2239), .Z(n2244) );
  XOR U2327 ( .A(n2241), .B(n2231), .Z(n2248) );
  IV U2328 ( .A(n2219), .Z(n2225) );
  XOR U2329 ( .A(n2249), .B(n2250), .Z(n2219) );
  XOR U2330 ( .A(n2241), .B(n2251), .Z(n2250) );
  XNOR U2331 ( .A(n2252), .B(n2238), .Z(n2251) );
  OR U2332 ( .A(n2151), .B(n2192), .Z(n2238) );
  XNOR U2333 ( .A(n2191), .B(n2183), .Z(n2192) );
  XNOR U2334 ( .A(n2253), .B(n2154), .Z(n2151) );
  ANDN U2335 ( .A(n2254), .B(n2131), .Z(n2252) );
  XNOR U2336 ( .A(n2243), .B(n2255), .Z(n2241) );
  ANDN U2337 ( .A(n2256), .B(n2168), .Z(n2255) );
  OR U2338 ( .A(n2196), .B(n2172), .Z(n2243) );
  XOR U2339 ( .A(n2168), .B(n2174), .Z(n2172) );
  XNOR U2340 ( .A(n2131), .B(n2162), .Z(n2174) );
  XNOR U2341 ( .A(n2257), .B(n2154), .Z(n2162) );
  XOR U2342 ( .A(n2258), .B(n2259), .Z(n2257) );
  IV U2343 ( .A(n2253), .Z(n2131) );
  XOR U2344 ( .A(n2231), .B(n2154), .Z(n2168) );
  XOR U2345 ( .A(n2260), .B(n2261), .Z(n2231) );
  XOR U2346 ( .A(n2262), .B(n2263), .Z(n2260) );
  XOR U2347 ( .A(n2256), .B(n2189), .Z(n2196) );
  XOR U2348 ( .A(n2254), .B(n2212), .Z(n2189) );
  XOR U2349 ( .A(n2264), .B(n2265), .Z(n2212) );
  XNOR U2350 ( .A(n2266), .B(n2141), .Z(n2265) );
  XNOR U2351 ( .A(n2267), .B(n2262), .Z(n2264) );
  XNOR U2352 ( .A(g_input[44]), .B(state[44]), .Z(n2262) );
  IV U2353 ( .A(n2195), .Z(n2256) );
  XOR U2354 ( .A(n2191), .B(n2141), .Z(n2195) );
  XNOR U2355 ( .A(n2239), .B(n2233), .Z(n2249) );
  XNOR U2356 ( .A(n2253), .B(n2254), .Z(n2233) );
  IV U2357 ( .A(n2183), .Z(n2254) );
  XOR U2358 ( .A(n2268), .B(n2263), .Z(n2183) );
  XOR U2359 ( .A(n2269), .B(n2268), .Z(n2253) );
  IV U2360 ( .A(n2261), .Z(n2268) );
  XNOR U2361 ( .A(n2259), .B(n2263), .Z(n2269) );
  XOR U2362 ( .A(n2154), .B(n2191), .Z(n2239) );
  XOR U2363 ( .A(n2258), .B(n2270), .Z(n2191) );
  XNOR U2364 ( .A(n2266), .B(n2263), .Z(n2270) );
  XOR U2365 ( .A(n2271), .B(n2259), .Z(n2266) );
  XOR U2366 ( .A(g_input[41]), .B(state[41]), .Z(n2259) );
  XNOR U2367 ( .A(g_input[43]), .B(state[43]), .Z(n2271) );
  XNOR U2368 ( .A(g_input[42]), .B(state[42]), .Z(n2258) );
  XNOR U2369 ( .A(n2272), .B(n2261), .Z(n2154) );
  XOR U2370 ( .A(g_input[45]), .B(state[45]), .Z(n2261) );
  XOR U2371 ( .A(n2267), .B(n2263), .Z(n2272) );
  XNOR U2372 ( .A(n2273), .B(n2141), .Z(n2263) );
  XOR U2373 ( .A(g_input[40]), .B(state[40]), .Z(n2141) );
  XNOR U2374 ( .A(g_input[46]), .B(state[46]), .Z(n2273) );
  XNOR U2375 ( .A(g_input[47]), .B(state[47]), .Z(n2267) );
  XOR U2376 ( .A(n2274), .B(n2275), .Z(o[103]) );
  XOR U2377 ( .A(n12), .B(n2276), .Z(n2275) );
  XNOR U2378 ( .A(g_input[103]), .B(n8), .Z(n2276) );
  XOR U2379 ( .A(n2277), .B(n2278), .Z(n8) );
  XNOR U2380 ( .A(n2279), .B(n2280), .Z(n2277) );
  ANDN U2381 ( .A(n2281), .B(n2282), .Z(n2280) );
  XNOR U2382 ( .A(n2283), .B(n16), .Z(n2274) );
  IV U2383 ( .A(n2284), .Z(n16) );
  XOR U2384 ( .A(n2285), .B(n2284), .Z(o[102]) );
  XNOR U2385 ( .A(n19), .B(n10), .Z(n2284) );
  XNOR U2386 ( .A(n2286), .B(n2287), .Z(n10) );
  XNOR U2387 ( .A(n2279), .B(n2288), .Z(n2286) );
  ANDN U2388 ( .A(n2289), .B(n2290), .Z(n2288) );
  ANDN U2389 ( .A(n2291), .B(n2292), .Z(n2279) );
  XNOR U2390 ( .A(n11), .B(g_input[102]), .Z(n2285) );
  XNOR U2391 ( .A(n2293), .B(n2278), .Z(n11) );
  XOR U2392 ( .A(n2294), .B(n2287), .Z(n2278) );
  XNOR U2393 ( .A(n2295), .B(n2296), .Z(n2294) );
  ANDN U2394 ( .A(n2297), .B(n2298), .Z(n2296) );
  XNOR U2395 ( .A(n2299), .B(n2300), .Z(n2293) );
  NANDN U2396 ( .B(n2301), .A(n2302), .Z(n2299) );
  XOR U2397 ( .A(n2303), .B(n2304), .Z(o[101]) );
  XOR U2398 ( .A(n2305), .B(n2306), .Z(n2304) );
  XNOR U2399 ( .A(g_input[101]), .B(n2300), .Z(n2306) );
  OR U2400 ( .A(n2307), .B(n2308), .Z(n2300) );
  NOR U2401 ( .A(n2309), .B(n2310), .Z(n2305) );
  XNOR U2402 ( .A(n2311), .B(n2283), .Z(n2303) );
  XNOR U2403 ( .A(n2312), .B(n2313), .Z(n2283) );
  XNOR U2404 ( .A(n2314), .B(n2315), .Z(n2312) );
  OR U2405 ( .A(n2282), .B(n2316), .Z(n2314) );
  XOR U2406 ( .A(n18), .B(n2287), .Z(n2311) );
  XNOR U2407 ( .A(n2295), .B(n2317), .Z(n2287) );
  ANDN U2408 ( .A(n2318), .B(n2319), .Z(n2317) );
  NOR U2409 ( .A(n2320), .B(n2321), .Z(n2295) );
  XOR U2410 ( .A(n2322), .B(n18), .Z(o[100]) );
  XOR U2411 ( .A(n2323), .B(n2313), .Z(n18) );
  XNOR U2412 ( .A(n2324), .B(n2325), .Z(n2313) );
  XNOR U2413 ( .A(n2326), .B(n2327), .Z(n2324) );
  NANDN U2414 ( .B(n2298), .A(n2328), .Z(n2326) );
  XNOR U2415 ( .A(n2329), .B(n2330), .Z(n2323) );
  ANDN U2416 ( .A(n2302), .B(n2331), .Z(n2330) );
  XNOR U2417 ( .A(n13), .B(g_input[100]), .Z(n2322) );
  XOR U2418 ( .A(n19), .B(n12), .Z(n13) );
  XOR U2419 ( .A(n2332), .B(n2325), .Z(n12) );
  XNOR U2420 ( .A(n2329), .B(n2333), .Z(n2332) );
  NOR U2421 ( .A(n2397), .B(n2310), .Z(n2333) );
  NOR U2422 ( .A(n2308), .B(n2334), .Z(n2329) );
  XOR U2423 ( .A(n2310), .B(n2302), .Z(n2308) );
  XOR U2424 ( .A(n2335), .B(n2325), .Z(n19) );
  XOR U2425 ( .A(n2327), .B(n2336), .Z(n2325) );
  NOR U2426 ( .A(n2319), .B(n2337), .Z(n2336) );
  OR U2427 ( .A(n2321), .B(n2338), .Z(n2327) );
  XOR U2428 ( .A(n2302), .B(n2282), .Z(n2319) );
  XOR U2429 ( .A(n2339), .B(n2340), .Z(n2302) );
  ANDN U2430 ( .A(n2341), .B(n2342), .Z(n2340) );
  XOR U2431 ( .A(n2343), .B(n2339), .Z(n2310) );
  OR U2432 ( .A(n2346), .B(n2347), .Z(n2343) );
  XNOR U2433 ( .A(n2348), .B(n2315), .Z(n2335) );
  NANDN U2434 ( .B(n2349), .A(n2291), .Z(n2315) );
  XOR U2435 ( .A(n2290), .B(n2282), .Z(n2291) );
  XNOR U2436 ( .A(n2350), .B(n2351), .Z(n2282) );
  NOR U2437 ( .A(n2352), .B(n2342), .Z(n2351) );
  NANDN U2438 ( .B(n2290), .A(n2353), .Z(n2348) );
  XNOR U2439 ( .A(n2350), .B(n2354), .Z(n2290) );
  ANDN U2440 ( .A(n2355), .B(n2346), .Z(n2354) );
  ANDN U2441 ( .A(n2345), .B(n2356), .Z(n2350) );
  XOR U2442 ( .A(n2342), .B(n2346), .Z(n2345) );
  XOR U2443 ( .A(n2357), .B(n2358), .Z(n2346) );
  XOR U2444 ( .A(n2359), .B(n2360), .Z(n2358) );
  XNOR U2445 ( .A(n2361), .B(n2362), .Z(n2360) );
  ANDN U2446 ( .A(n2341), .B(n2352), .Z(n2362) );
  XOR U2447 ( .A(n2363), .B(n2341), .Z(n2357) );
  XNOR U2448 ( .A(n2364), .B(n2363), .Z(n2342) );
  XNOR U2449 ( .A(n2365), .B(n2355), .Z(n2363) );
  XNOR U2450 ( .A(n2366), .B(n2361), .Z(n2364) );
  OR U2451 ( .A(n2356), .B(n2344), .Z(n2361) );
  XNOR U2452 ( .A(n2365), .B(n2341), .Z(n2344) );
  XNOR U2453 ( .A(n2367), .B(n2368), .Z(n2341) );
  XNOR U2454 ( .A(n2369), .B(n2370), .Z(n2368) );
  XNOR U2455 ( .A(n2371), .B(n2372), .Z(n2370) );
  ANDN U2456 ( .A(n2281), .B(n2316), .Z(n2371) );
  XOR U2457 ( .A(n2373), .B(n2374), .Z(n2367) );
  XNOR U2458 ( .A(n2375), .B(n2353), .Z(n2373) );
  IV U2459 ( .A(n2347), .Z(n2365) );
  XOR U2460 ( .A(n2355), .B(n2352), .Z(n2356) );
  IV U2461 ( .A(n2359), .Z(n2352) );
  XNOR U2462 ( .A(n2376), .B(n2377), .Z(n2359) );
  XNOR U2463 ( .A(n2378), .B(n2379), .Z(n2377) );
  XOR U2464 ( .A(n2380), .B(n2375), .Z(n2376) );
  XNOR U2465 ( .A(n2381), .B(n2382), .Z(n2375) );
  XNOR U2466 ( .A(n2383), .B(n2384), .Z(n2381) );
  AND U2467 ( .A(n2328), .B(n2297), .Z(n2384) );
  NANDN U2468 ( .B(n2347), .A(n2355), .Z(n2366) );
  XNOR U2469 ( .A(n2385), .B(n2386), .Z(n2355) );
  XOR U2470 ( .A(n2382), .B(n2387), .Z(n2386) );
  XNOR U2471 ( .A(n2388), .B(n2379), .Z(n2387) );
  OR U2472 ( .A(n2307), .B(n2334), .Z(n2379) );
  XNOR U2473 ( .A(n2389), .B(n2390), .Z(n2334) );
  ANDN U2474 ( .A(n2389), .B(n2309), .Z(n2388) );
  XOR U2475 ( .A(n2374), .B(n2380), .Z(n2385) );
  XOR U2476 ( .A(n2397), .B(n2309), .Z(n2374) );
  XOR U2477 ( .A(n2391), .B(n2392), .Z(n2347) );
  XNOR U2478 ( .A(n2316), .B(n2393), .Z(n2392) );
  XNOR U2479 ( .A(n2394), .B(n2372), .Z(n2393) );
  OR U2480 ( .A(n2292), .B(n2349), .Z(n2372) );
  XOR U2481 ( .A(n2353), .B(n2316), .Z(n2349) );
  XNOR U2482 ( .A(n2289), .B(n2281), .Z(n2292) );
  ANDN U2483 ( .A(n2353), .B(n2369), .Z(n2394) );
  IV U2484 ( .A(n2289), .Z(n2369) );
  XNOR U2485 ( .A(n2395), .B(n2380), .Z(n2391) );
  XOR U2486 ( .A(n2390), .B(n2301), .Z(n2380) );
  XNOR U2487 ( .A(n2382), .B(n2281), .Z(n2395) );
  XOR U2488 ( .A(n2383), .B(n2396), .Z(n2382) );
  ANDN U2489 ( .A(n2318), .B(n2337), .Z(n2396) );
  NOR U2490 ( .A(n2338), .B(n2320), .Z(n2383) );
  XNOR U2491 ( .A(n2297), .B(n2318), .Z(n2320) );
  XNOR U2492 ( .A(n2301), .B(n2281), .Z(n2318) );
  XNOR U2493 ( .A(n2397), .B(n2398), .Z(n2281) );
  XNOR U2494 ( .A(n2399), .B(n2400), .Z(n2397) );
  XNOR U2495 ( .A(n2309), .B(n2289), .Z(n2297) );
  XNOR U2496 ( .A(n2401), .B(n2402), .Z(n2289) );
  XOR U2497 ( .A(n2403), .B(n2301), .Z(n2401) );
  XNOR U2498 ( .A(n2404), .B(n2405), .Z(n2301) );
  XOR U2499 ( .A(n2404), .B(n2402), .Z(n2309) );
  XOR U2500 ( .A(n2399), .B(n2406), .Z(n2404) );
  XOR U2501 ( .A(n2328), .B(n2337), .Z(n2338) );
  XOR U2502 ( .A(n2390), .B(n2316), .Z(n2337) );
  IV U2503 ( .A(n2331), .Z(n2390) );
  XOR U2504 ( .A(n2407), .B(n2408), .Z(n2331) );
  XOR U2505 ( .A(n2403), .B(n2406), .Z(n2407) );
  XOR U2506 ( .A(g_input[2]), .B(state[2]), .Z(n2403) );
  XOR U2507 ( .A(n2353), .B(n2389), .Z(n2328) );
  XOR U2508 ( .A(n2399), .B(n2400), .Z(n2389) );
  IV U2509 ( .A(n2406), .Z(n2400) );
  XNOR U2510 ( .A(n2409), .B(n2316), .Z(n2406) );
  XNOR U2511 ( .A(g_input[6]), .B(state[6]), .Z(n2409) );
  XOR U2512 ( .A(g_input[5]), .B(state[5]), .Z(n2399) );
  XNOR U2513 ( .A(n2410), .B(n2411), .Z(n2353) );
  XNOR U2514 ( .A(n2316), .B(n2398), .Z(n2411) );
  XOR U2515 ( .A(g_input[4]), .B(state[4]), .Z(n2398) );
  XNOR U2516 ( .A(g_input[0]), .B(state[0]), .Z(n2316) );
  XOR U2517 ( .A(n2405), .B(n2408), .Z(n2410) );
  XNOR U2518 ( .A(n2412), .B(n2402), .Z(n2408) );
  XOR U2519 ( .A(g_input[1]), .B(state[1]), .Z(n2402) );
  XNOR U2520 ( .A(g_input[3]), .B(state[3]), .Z(n2412) );
  XNOR U2521 ( .A(g_input[7]), .B(state[7]), .Z(n2405) );
  XNOR U2522 ( .A(n2413), .B(n696), .Z(o[0]) );
  XOR U2523 ( .A(n2414), .B(n699), .Z(n696) );
  XOR U2524 ( .A(n2415), .B(n1523), .Z(n699) );
  XNOR U2525 ( .A(n2416), .B(n2417), .Z(n2415) );
  NOR U2526 ( .A(n1516), .B(n2418), .Z(n2417) );
  XNOR U2527 ( .A(n1524), .B(n2419), .Z(n2414) );
  NOR U2528 ( .A(n1156), .B(n2420), .Z(n2419) );
  ANDN U2529 ( .A(n1155), .B(n2421), .Z(n1524) );
  XOR U2530 ( .A(n1156), .B(n694), .Z(n1155) );
  XOR U2531 ( .A(n1325), .B(g_input[0]), .Z(n2413) );
  XNOR U2532 ( .A(n2422), .B(n1523), .Z(n1325) );
  XNOR U2533 ( .A(n2416), .B(n2423), .Z(n1523) );
  NOR U2534 ( .A(n2424), .B(n1512), .Z(n2423) );
  NOR U2535 ( .A(n1514), .B(n2425), .Z(n2416) );
  XNOR U2536 ( .A(n1506), .B(n694), .Z(n1516) );
  XNOR U2537 ( .A(n2426), .B(n2427), .Z(n694) );
  ANDN U2538 ( .A(n2428), .B(n2429), .Z(n2427) );
  IV U2539 ( .A(n2430), .Z(n702) );
  XNOR U2540 ( .A(n2426), .B(n2431), .Z(n1156) );
  NOR U2541 ( .A(n2432), .B(n2433), .Z(n2431) );
  ANDN U2542 ( .A(n2434), .B(n2435), .Z(n2426) );
  XNOR U2543 ( .A(n2436), .B(n701), .Z(n2422) );
  OR U2544 ( .A(n1520), .B(n2437), .Z(n701) );
  XOR U2545 ( .A(n2430), .B(n1506), .Z(n1520) );
  XOR U2546 ( .A(n2438), .B(n2439), .Z(n2430) );
  ANDN U2547 ( .A(n2440), .B(n2433), .Z(n2439) );
  OR U2548 ( .A(n1506), .B(n2441), .Z(n2436) );
  XOR U2549 ( .A(n2442), .B(n2438), .Z(n1506) );
  XOR U2550 ( .A(n2433), .B(n2429), .Z(n2434) );
  XNOR U2551 ( .A(n2444), .B(n2445), .Z(n2433) );
  XNOR U2552 ( .A(n2446), .B(n2447), .Z(n2444) );
  NANDN U2553 ( .B(n2448), .A(n2428), .Z(n2446) );
  OR U2554 ( .A(n2429), .B(n2448), .Z(n2442) );
  XOR U2555 ( .A(n2449), .B(n2450), .Z(n2429) );
  XOR U2556 ( .A(n2451), .B(n2452), .Z(n2450) );
  XNOR U2557 ( .A(n2447), .B(n2453), .Z(n2452) );
  ANDN U2558 ( .A(n2440), .B(n2432), .Z(n2453) );
  OR U2559 ( .A(n2435), .B(n2443), .Z(n2447) );
  XNOR U2560 ( .A(n2454), .B(n2440), .Z(n2443) );
  XOR U2561 ( .A(n2428), .B(n2432), .Z(n2435) );
  IV U2562 ( .A(n2451), .Z(n2432) );
  XNOR U2563 ( .A(n2455), .B(n2456), .Z(n2451) );
  XNOR U2564 ( .A(n2441), .B(n2457), .Z(n2456) );
  XNOR U2565 ( .A(n2458), .B(n2459), .Z(n2457) );
  ANDN U2566 ( .A(n703), .B(n2460), .Z(n2458) );
  XNOR U2567 ( .A(n2461), .B(n2462), .Z(n2455) );
  XOR U2568 ( .A(n2463), .B(n1505), .Z(n2461) );
  XOR U2569 ( .A(n2445), .B(n2440), .Z(n2449) );
  XNOR U2570 ( .A(n2464), .B(n2465), .Z(n2440) );
  XNOR U2571 ( .A(n2466), .B(n2467), .Z(n2465) );
  ANDN U2572 ( .A(n1157), .B(n2420), .Z(n2466) );
  XNOR U2573 ( .A(n2468), .B(n2463), .Z(n2464) );
  XOR U2574 ( .A(n2469), .B(n2470), .Z(n2463) );
  XNOR U2575 ( .A(n2471), .B(n2472), .Z(n2469) );
  NANDN U2576 ( .B(n2418), .A(n1517), .Z(n2471) );
  XNOR U2577 ( .A(n2454), .B(n2428), .Z(n2445) );
  XNOR U2578 ( .A(n2473), .B(n2474), .Z(n2428) );
  XOR U2579 ( .A(n703), .B(n2475), .Z(n2474) );
  XNOR U2580 ( .A(n2476), .B(n2459), .Z(n2475) );
  OR U2581 ( .A(n1521), .B(n2437), .Z(n2459) );
  XNOR U2582 ( .A(n1519), .B(n1505), .Z(n1521) );
  IV U2583 ( .A(n2460), .Z(n1519) );
  ANDN U2584 ( .A(n1505), .B(n2441), .Z(n2476) );
  XNOR U2585 ( .A(n2477), .B(n2468), .Z(n2473) );
  XOR U2586 ( .A(n2470), .B(n2460), .Z(n2477) );
  IV U2587 ( .A(n2448), .Z(n2454) );
  XOR U2588 ( .A(n2478), .B(n2479), .Z(n2448) );
  XOR U2589 ( .A(n2470), .B(n2480), .Z(n2479) );
  XNOR U2590 ( .A(n2481), .B(n2467), .Z(n2480) );
  OR U2591 ( .A(n1154), .B(n2421), .Z(n2467) );
  XNOR U2592 ( .A(n2420), .B(n1526), .Z(n2421) );
  XNOR U2593 ( .A(n2482), .B(n1157), .Z(n1154) );
  ANDN U2594 ( .A(n2483), .B(n693), .Z(n2481) );
  XNOR U2595 ( .A(n2472), .B(n2484), .Z(n2470) );
  ANDN U2596 ( .A(n2485), .B(n1511), .Z(n2484) );
  OR U2597 ( .A(n2425), .B(n1515), .Z(n2472) );
  XOR U2598 ( .A(n1511), .B(n1517), .Z(n1515) );
  XNOR U2599 ( .A(n693), .B(n1505), .Z(n1517) );
  XNOR U2600 ( .A(n2486), .B(n1157), .Z(n1505) );
  XNOR U2601 ( .A(n2487), .B(n2488), .Z(n2486) );
  XOR U2602 ( .A(n2460), .B(n1157), .Z(n1511) );
  XOR U2603 ( .A(n2489), .B(n2490), .Z(n2460) );
  XNOR U2604 ( .A(n2491), .B(n2492), .Z(n2489) );
  XOR U2605 ( .A(n2485), .B(n2418), .Z(n2425) );
  XOR U2606 ( .A(n2483), .B(n2441), .Z(n2418) );
  XOR U2607 ( .A(n2493), .B(n2494), .Z(n2441) );
  XNOR U2608 ( .A(n2495), .B(n703), .Z(n2494) );
  XNOR U2609 ( .A(n2496), .B(n2491), .Z(n2493) );
  XOR U2610 ( .A(g_input[36]), .B(state[36]), .Z(n2491) );
  IV U2611 ( .A(n2424), .Z(n2485) );
  XOR U2612 ( .A(n2420), .B(n703), .Z(n2424) );
  XNOR U2613 ( .A(n2468), .B(n2462), .Z(n2478) );
  XNOR U2614 ( .A(n2482), .B(n2483), .Z(n2462) );
  IV U2615 ( .A(n1526), .Z(n2483) );
  IV U2616 ( .A(n693), .Z(n2482) );
  XOR U2617 ( .A(n2497), .B(n2490), .Z(n693) );
  XNOR U2618 ( .A(n2488), .B(n2492), .Z(n2497) );
  XOR U2619 ( .A(n1157), .B(n2420), .Z(n2468) );
  XNOR U2620 ( .A(n2487), .B(n2498), .Z(n2420) );
  XNOR U2621 ( .A(n2495), .B(n2492), .Z(n2498) );
  XOR U2622 ( .A(n2499), .B(n2488), .Z(n2495) );
  XOR U2623 ( .A(g_input[33]), .B(state[33]), .Z(n2488) );
  XNOR U2624 ( .A(g_input[35]), .B(state[35]), .Z(n2499) );
  XOR U2625 ( .A(g_input[34]), .B(state[34]), .Z(n2487) );
  XNOR U2626 ( .A(n2500), .B(n2490), .Z(n1157) );
  XOR U2627 ( .A(g_input[37]), .B(state[37]), .Z(n2490) );
  XNOR U2628 ( .A(n2496), .B(n2492), .Z(n2500) );
  XNOR U2629 ( .A(n2501), .B(n703), .Z(n2492) );
  XOR U2630 ( .A(g_input[32]), .B(state[32]), .Z(n703) );
  XNOR U2631 ( .A(g_input[38]), .B(state[38]), .Z(n2501) );
  XOR U2632 ( .A(g_input[39]), .B(state[39]), .Z(n2496) );
endmodule

