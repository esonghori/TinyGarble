
module mult_N128_CC32 ( clk, rst, a, b, c );
  input [127:0] a;
  input [3:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179;
  wire   [255:0] sreg;

  DFF \sreg_reg[251]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U7 ( .A(sreg[128]), .B(n440), .Z(n1) );
  XOR U8 ( .A(sreg[128]), .B(n440), .Z(n2) );
  NANDN U9 ( .A(n439), .B(n2), .Z(n3) );
  NAND U10 ( .A(n1), .B(n3), .Z(n461) );
  XOR U11 ( .A(sreg[132]), .B(n527), .Z(n4) );
  NANDN U12 ( .A(n528), .B(n4), .Z(n5) );
  NAND U13 ( .A(sreg[132]), .B(n527), .Z(n6) );
  AND U14 ( .A(n5), .B(n6), .Z(n549) );
  NAND U15 ( .A(n615), .B(n616), .Z(n7) );
  XOR U16 ( .A(n615), .B(n616), .Z(n8) );
  NAND U17 ( .A(n8), .B(sreg[136]), .Z(n9) );
  NAND U18 ( .A(n7), .B(n9), .Z(n637) );
  NAND U19 ( .A(n703), .B(n704), .Z(n10) );
  XOR U20 ( .A(n703), .B(n704), .Z(n11) );
  NAND U21 ( .A(n11), .B(sreg[140]), .Z(n12) );
  NAND U22 ( .A(n10), .B(n12), .Z(n725) );
  NAND U23 ( .A(n791), .B(n792), .Z(n13) );
  XOR U24 ( .A(n791), .B(n792), .Z(n14) );
  NAND U25 ( .A(n14), .B(sreg[144]), .Z(n15) );
  NAND U26 ( .A(n13), .B(n15), .Z(n813) );
  NAND U27 ( .A(sreg[148]), .B(n880), .Z(n16) );
  XOR U28 ( .A(sreg[148]), .B(n880), .Z(n17) );
  NANDN U29 ( .A(n879), .B(n17), .Z(n18) );
  NAND U30 ( .A(n16), .B(n18), .Z(n901) );
  XOR U31 ( .A(sreg[152]), .B(n967), .Z(n19) );
  NANDN U32 ( .A(n968), .B(n19), .Z(n20) );
  NAND U33 ( .A(sreg[152]), .B(n967), .Z(n21) );
  AND U34 ( .A(n20), .B(n21), .Z(n989) );
  XOR U35 ( .A(sreg[156]), .B(n1055), .Z(n22) );
  NANDN U36 ( .A(n1056), .B(n22), .Z(n23) );
  NAND U37 ( .A(sreg[156]), .B(n1055), .Z(n24) );
  AND U38 ( .A(n23), .B(n24), .Z(n1077) );
  NAND U39 ( .A(n1143), .B(n1144), .Z(n25) );
  XOR U40 ( .A(n1143), .B(n1144), .Z(n26) );
  NAND U41 ( .A(n26), .B(sreg[160]), .Z(n27) );
  NAND U42 ( .A(n25), .B(n27), .Z(n1165) );
  NAND U43 ( .A(sreg[164]), .B(n1232), .Z(n28) );
  XOR U44 ( .A(sreg[164]), .B(n1232), .Z(n29) );
  NANDN U45 ( .A(n1231), .B(n29), .Z(n30) );
  NAND U46 ( .A(n28), .B(n30), .Z(n1253) );
  NAND U47 ( .A(n1319), .B(n1320), .Z(n31) );
  XOR U48 ( .A(n1319), .B(n1320), .Z(n32) );
  NAND U49 ( .A(n32), .B(sreg[168]), .Z(n33) );
  NAND U50 ( .A(n31), .B(n33), .Z(n1341) );
  NAND U51 ( .A(n1407), .B(n1408), .Z(n34) );
  XOR U52 ( .A(n1407), .B(n1408), .Z(n35) );
  NAND U53 ( .A(n35), .B(sreg[172]), .Z(n36) );
  NAND U54 ( .A(n34), .B(n36), .Z(n1429) );
  NAND U55 ( .A(n1495), .B(n1496), .Z(n37) );
  XOR U56 ( .A(n1495), .B(n1496), .Z(n38) );
  NAND U57 ( .A(n38), .B(sreg[176]), .Z(n39) );
  NAND U58 ( .A(n37), .B(n39), .Z(n1517) );
  NAND U59 ( .A(sreg[180]), .B(n1584), .Z(n40) );
  XOR U60 ( .A(sreg[180]), .B(n1584), .Z(n41) );
  NANDN U61 ( .A(n1583), .B(n41), .Z(n42) );
  NAND U62 ( .A(n40), .B(n42), .Z(n1605) );
  NAND U63 ( .A(n1671), .B(n1672), .Z(n43) );
  XOR U64 ( .A(n1671), .B(n1672), .Z(n44) );
  NAND U65 ( .A(n44), .B(sreg[184]), .Z(n45) );
  NAND U66 ( .A(n43), .B(n45), .Z(n1693) );
  NAND U67 ( .A(n1759), .B(n1760), .Z(n46) );
  XOR U68 ( .A(n1759), .B(n1760), .Z(n47) );
  NAND U69 ( .A(n47), .B(sreg[188]), .Z(n48) );
  NAND U70 ( .A(n46), .B(n48), .Z(n1781) );
  NAND U71 ( .A(sreg[192]), .B(n1848), .Z(n49) );
  XOR U72 ( .A(sreg[192]), .B(n1848), .Z(n50) );
  NANDN U73 ( .A(n1847), .B(n50), .Z(n51) );
  NAND U74 ( .A(n49), .B(n51), .Z(n1869) );
  NAND U75 ( .A(sreg[196]), .B(n1936), .Z(n52) );
  XOR U76 ( .A(sreg[196]), .B(n1936), .Z(n53) );
  NANDN U77 ( .A(n1935), .B(n53), .Z(n54) );
  NAND U78 ( .A(n52), .B(n54), .Z(n1957) );
  NAND U79 ( .A(n2023), .B(n2024), .Z(n55) );
  XOR U80 ( .A(n2023), .B(n2024), .Z(n56) );
  NAND U81 ( .A(n56), .B(sreg[200]), .Z(n57) );
  NAND U82 ( .A(n55), .B(n57), .Z(n2045) );
  XOR U83 ( .A(sreg[204]), .B(n2111), .Z(n58) );
  NANDN U84 ( .A(n2112), .B(n58), .Z(n59) );
  NAND U85 ( .A(sreg[204]), .B(n2111), .Z(n60) );
  AND U86 ( .A(n59), .B(n60), .Z(n2133) );
  NAND U87 ( .A(n2199), .B(n2200), .Z(n61) );
  XOR U88 ( .A(n2199), .B(n2200), .Z(n62) );
  NAND U89 ( .A(n62), .B(sreg[208]), .Z(n63) );
  NAND U90 ( .A(n61), .B(n63), .Z(n2221) );
  NAND U91 ( .A(sreg[212]), .B(n2288), .Z(n64) );
  XOR U92 ( .A(sreg[212]), .B(n2288), .Z(n65) );
  NANDN U93 ( .A(n2287), .B(n65), .Z(n66) );
  NAND U94 ( .A(n64), .B(n66), .Z(n2309) );
  NAND U95 ( .A(n2375), .B(n2376), .Z(n67) );
  XOR U96 ( .A(n2375), .B(n2376), .Z(n68) );
  NAND U97 ( .A(n68), .B(sreg[216]), .Z(n69) );
  NAND U98 ( .A(n67), .B(n69), .Z(n2397) );
  XOR U99 ( .A(sreg[220]), .B(n2463), .Z(n70) );
  NANDN U100 ( .A(n2464), .B(n70), .Z(n71) );
  NAND U101 ( .A(sreg[220]), .B(n2463), .Z(n72) );
  AND U102 ( .A(n71), .B(n72), .Z(n2485) );
  NAND U103 ( .A(n2551), .B(n2552), .Z(n73) );
  XOR U104 ( .A(n2551), .B(n2552), .Z(n74) );
  NAND U105 ( .A(n74), .B(sreg[224]), .Z(n75) );
  NAND U106 ( .A(n73), .B(n75), .Z(n2573) );
  NAND U107 ( .A(n2639), .B(n2640), .Z(n76) );
  XOR U108 ( .A(n2639), .B(n2640), .Z(n77) );
  NAND U109 ( .A(n77), .B(sreg[228]), .Z(n78) );
  NAND U110 ( .A(n76), .B(n78), .Z(n2661) );
  NAND U111 ( .A(n2727), .B(n2728), .Z(n79) );
  XOR U112 ( .A(n2727), .B(n2728), .Z(n80) );
  NAND U113 ( .A(n80), .B(sreg[232]), .Z(n81) );
  NAND U114 ( .A(n79), .B(n81), .Z(n2749) );
  NAND U115 ( .A(n2815), .B(n2816), .Z(n82) );
  XOR U116 ( .A(n2815), .B(n2816), .Z(n83) );
  NAND U117 ( .A(n83), .B(sreg[236]), .Z(n84) );
  NAND U118 ( .A(n82), .B(n84), .Z(n2837) );
  NAND U119 ( .A(n2903), .B(n2904), .Z(n85) );
  XOR U120 ( .A(n2903), .B(n2904), .Z(n86) );
  NAND U121 ( .A(n86), .B(sreg[240]), .Z(n87) );
  NAND U122 ( .A(n85), .B(n87), .Z(n2925) );
  NAND U123 ( .A(sreg[244]), .B(n2992), .Z(n88) );
  XOR U124 ( .A(sreg[244]), .B(n2992), .Z(n89) );
  NANDN U125 ( .A(n2991), .B(n89), .Z(n90) );
  NAND U126 ( .A(n88), .B(n90), .Z(n3013) );
  NAND U127 ( .A(n3079), .B(n3080), .Z(n91) );
  XOR U128 ( .A(n3079), .B(n3080), .Z(n92) );
  NAND U129 ( .A(n92), .B(sreg[248]), .Z(n93) );
  NAND U130 ( .A(n91), .B(n93), .Z(n3101) );
  NANDN U131 ( .A(n3152), .B(n3162), .Z(n94) );
  XNOR U132 ( .A(n3160), .B(n94), .Z(n3163) );
  XOR U133 ( .A(sreg[129]), .B(n461), .Z(n95) );
  NANDN U134 ( .A(n462), .B(n95), .Z(n96) );
  NAND U135 ( .A(sreg[129]), .B(n461), .Z(n97) );
  AND U136 ( .A(n96), .B(n97), .Z(n483) );
  NAND U137 ( .A(sreg[133]), .B(n550), .Z(n98) );
  XOR U138 ( .A(sreg[133]), .B(n550), .Z(n99) );
  NANDN U139 ( .A(n549), .B(n99), .Z(n100) );
  NAND U140 ( .A(n98), .B(n100), .Z(n571) );
  NAND U141 ( .A(n637), .B(n638), .Z(n101) );
  XOR U142 ( .A(n637), .B(n638), .Z(n102) );
  NAND U143 ( .A(n102), .B(sreg[137]), .Z(n103) );
  NAND U144 ( .A(n101), .B(n103), .Z(n659) );
  NAND U145 ( .A(n725), .B(n726), .Z(n104) );
  XOR U146 ( .A(n725), .B(n726), .Z(n105) );
  NAND U147 ( .A(n105), .B(sreg[141]), .Z(n106) );
  NAND U148 ( .A(n104), .B(n106), .Z(n747) );
  NAND U149 ( .A(n813), .B(n814), .Z(n107) );
  XOR U150 ( .A(n813), .B(n814), .Z(n108) );
  NAND U151 ( .A(n108), .B(sreg[145]), .Z(n109) );
  NAND U152 ( .A(n107), .B(n109), .Z(n835) );
  XOR U153 ( .A(sreg[149]), .B(n901), .Z(n110) );
  NANDN U154 ( .A(n902), .B(n110), .Z(n111) );
  NAND U155 ( .A(sreg[149]), .B(n901), .Z(n112) );
  AND U156 ( .A(n111), .B(n112), .Z(n923) );
  NAND U157 ( .A(n989), .B(n990), .Z(n113) );
  XOR U158 ( .A(n989), .B(n990), .Z(n114) );
  NANDN U159 ( .A(sreg[153]), .B(n114), .Z(n115) );
  NAND U160 ( .A(n113), .B(n115), .Z(n1011) );
  NAND U161 ( .A(sreg[157]), .B(n1078), .Z(n116) );
  XOR U162 ( .A(sreg[157]), .B(n1078), .Z(n117) );
  NANDN U163 ( .A(n1077), .B(n117), .Z(n118) );
  NAND U164 ( .A(n116), .B(n118), .Z(n1099) );
  NAND U165 ( .A(n1165), .B(n1166), .Z(n119) );
  XOR U166 ( .A(n1165), .B(n1166), .Z(n120) );
  NAND U167 ( .A(n120), .B(sreg[161]), .Z(n121) );
  NAND U168 ( .A(n119), .B(n121), .Z(n1187) );
  XOR U169 ( .A(sreg[165]), .B(n1253), .Z(n122) );
  NANDN U170 ( .A(n1254), .B(n122), .Z(n123) );
  NAND U171 ( .A(sreg[165]), .B(n1253), .Z(n124) );
  AND U172 ( .A(n123), .B(n124), .Z(n1275) );
  NAND U173 ( .A(n1341), .B(n1342), .Z(n125) );
  XOR U174 ( .A(n1341), .B(n1342), .Z(n126) );
  NAND U175 ( .A(n126), .B(sreg[169]), .Z(n127) );
  NAND U176 ( .A(n125), .B(n127), .Z(n1363) );
  NAND U177 ( .A(n1429), .B(n1430), .Z(n128) );
  XOR U178 ( .A(n1429), .B(n1430), .Z(n129) );
  NAND U179 ( .A(n129), .B(sreg[173]), .Z(n130) );
  NAND U180 ( .A(n128), .B(n130), .Z(n1451) );
  NAND U181 ( .A(n1517), .B(n1518), .Z(n131) );
  XOR U182 ( .A(n1517), .B(n1518), .Z(n132) );
  NAND U183 ( .A(n132), .B(sreg[177]), .Z(n133) );
  NAND U184 ( .A(n131), .B(n133), .Z(n1539) );
  NAND U185 ( .A(n1605), .B(n1606), .Z(n134) );
  XOR U186 ( .A(n1605), .B(n1606), .Z(n135) );
  NAND U187 ( .A(n135), .B(sreg[181]), .Z(n136) );
  NAND U188 ( .A(n134), .B(n136), .Z(n1627) );
  NAND U189 ( .A(n1693), .B(n1694), .Z(n137) );
  XOR U190 ( .A(n1693), .B(n1694), .Z(n138) );
  NAND U191 ( .A(n138), .B(sreg[185]), .Z(n139) );
  NAND U192 ( .A(n137), .B(n139), .Z(n1715) );
  NAND U193 ( .A(n1781), .B(n1782), .Z(n140) );
  XOR U194 ( .A(n1781), .B(n1782), .Z(n141) );
  NAND U195 ( .A(n141), .B(sreg[189]), .Z(n142) );
  NAND U196 ( .A(n140), .B(n142), .Z(n1803) );
  NAND U197 ( .A(n1869), .B(n1870), .Z(n143) );
  XOR U198 ( .A(n1869), .B(n1870), .Z(n144) );
  NAND U199 ( .A(n144), .B(sreg[193]), .Z(n145) );
  NAND U200 ( .A(n143), .B(n145), .Z(n1891) );
  XOR U201 ( .A(sreg[197]), .B(n1957), .Z(n146) );
  NANDN U202 ( .A(n1958), .B(n146), .Z(n147) );
  NAND U203 ( .A(sreg[197]), .B(n1957), .Z(n148) );
  AND U204 ( .A(n147), .B(n148), .Z(n1979) );
  NAND U205 ( .A(n2045), .B(n2046), .Z(n149) );
  XOR U206 ( .A(n2045), .B(n2046), .Z(n150) );
  NAND U207 ( .A(n150), .B(sreg[201]), .Z(n151) );
  NAND U208 ( .A(n149), .B(n151), .Z(n2067) );
  NAND U209 ( .A(sreg[205]), .B(n2134), .Z(n152) );
  XOR U210 ( .A(sreg[205]), .B(n2134), .Z(n153) );
  NANDN U211 ( .A(n2133), .B(n153), .Z(n154) );
  NAND U212 ( .A(n152), .B(n154), .Z(n2155) );
  NAND U213 ( .A(n2221), .B(n2222), .Z(n155) );
  XOR U214 ( .A(n2221), .B(n2222), .Z(n156) );
  NAND U215 ( .A(n156), .B(sreg[209]), .Z(n157) );
  NAND U216 ( .A(n155), .B(n157), .Z(n2243) );
  XOR U217 ( .A(sreg[213]), .B(n2309), .Z(n158) );
  NANDN U218 ( .A(n2310), .B(n158), .Z(n159) );
  NAND U219 ( .A(sreg[213]), .B(n2309), .Z(n160) );
  AND U220 ( .A(n159), .B(n160), .Z(n2331) );
  NAND U221 ( .A(n2397), .B(n2398), .Z(n161) );
  XOR U222 ( .A(n2397), .B(n2398), .Z(n162) );
  NAND U223 ( .A(n162), .B(sreg[217]), .Z(n163) );
  NAND U224 ( .A(n161), .B(n163), .Z(n2419) );
  NAND U225 ( .A(sreg[221]), .B(n2486), .Z(n164) );
  XOR U226 ( .A(sreg[221]), .B(n2486), .Z(n165) );
  NANDN U227 ( .A(n2485), .B(n165), .Z(n166) );
  NAND U228 ( .A(n164), .B(n166), .Z(n2507) );
  NAND U229 ( .A(n2573), .B(n2574), .Z(n167) );
  XOR U230 ( .A(n2573), .B(n2574), .Z(n168) );
  NAND U231 ( .A(n168), .B(sreg[225]), .Z(n169) );
  NAND U232 ( .A(n167), .B(n169), .Z(n2595) );
  NAND U233 ( .A(n2661), .B(n2662), .Z(n170) );
  XOR U234 ( .A(n2661), .B(n2662), .Z(n171) );
  NAND U235 ( .A(n171), .B(sreg[229]), .Z(n172) );
  NAND U236 ( .A(n170), .B(n172), .Z(n2683) );
  NAND U237 ( .A(n2749), .B(n2750), .Z(n173) );
  XOR U238 ( .A(n2749), .B(n2750), .Z(n174) );
  NAND U239 ( .A(n174), .B(sreg[233]), .Z(n175) );
  NAND U240 ( .A(n173), .B(n175), .Z(n2771) );
  NAND U241 ( .A(n2837), .B(n2838), .Z(n176) );
  XOR U242 ( .A(n2837), .B(n2838), .Z(n177) );
  NAND U243 ( .A(n177), .B(sreg[237]), .Z(n178) );
  NAND U244 ( .A(n176), .B(n178), .Z(n2859) );
  NAND U245 ( .A(n2925), .B(n2926), .Z(n179) );
  XOR U246 ( .A(n2925), .B(n2926), .Z(n180) );
  NAND U247 ( .A(n180), .B(sreg[241]), .Z(n181) );
  NAND U248 ( .A(n179), .B(n181), .Z(n2947) );
  XOR U249 ( .A(sreg[245]), .B(n3013), .Z(n182) );
  NANDN U250 ( .A(n3014), .B(n182), .Z(n183) );
  NAND U251 ( .A(sreg[245]), .B(n3013), .Z(n184) );
  AND U252 ( .A(n183), .B(n184), .Z(n3035) );
  NAND U253 ( .A(n3101), .B(n3102), .Z(n185) );
  XOR U254 ( .A(n3101), .B(n3102), .Z(n186) );
  NAND U255 ( .A(n186), .B(sreg[249]), .Z(n187) );
  NAND U256 ( .A(n185), .B(n187), .Z(n3123) );
  XNOR U257 ( .A(n418), .B(n417), .Z(n392) );
  NAND U258 ( .A(n3148), .B(n3149), .Z(n188) );
  NANDN U259 ( .A(n3151), .B(n3150), .Z(n189) );
  AND U260 ( .A(n188), .B(n189), .Z(n3166) );
  NAND U261 ( .A(sreg[131]), .B(n506), .Z(n190) );
  XOR U262 ( .A(sreg[131]), .B(n506), .Z(n191) );
  NANDN U263 ( .A(n505), .B(n191), .Z(n192) );
  NAND U264 ( .A(n190), .B(n192), .Z(n527) );
  NAND U265 ( .A(n593), .B(n594), .Z(n193) );
  XOR U266 ( .A(n593), .B(n594), .Z(n194) );
  NAND U267 ( .A(n194), .B(sreg[135]), .Z(n195) );
  NAND U268 ( .A(n193), .B(n195), .Z(n615) );
  NAND U269 ( .A(n681), .B(n682), .Z(n196) );
  XOR U270 ( .A(n681), .B(n682), .Z(n197) );
  NAND U271 ( .A(n197), .B(sreg[139]), .Z(n198) );
  NAND U272 ( .A(n196), .B(n198), .Z(n703) );
  NAND U273 ( .A(sreg[143]), .B(n770), .Z(n199) );
  XOR U274 ( .A(sreg[143]), .B(n770), .Z(n200) );
  NANDN U275 ( .A(n769), .B(n200), .Z(n201) );
  NAND U276 ( .A(n199), .B(n201), .Z(n791) );
  XOR U277 ( .A(sreg[147]), .B(n857), .Z(n202) );
  NANDN U278 ( .A(n858), .B(n202), .Z(n203) );
  NAND U279 ( .A(sreg[147]), .B(n857), .Z(n204) );
  AND U280 ( .A(n203), .B(n204), .Z(n879) );
  NAND U281 ( .A(n945), .B(n946), .Z(n205) );
  XOR U282 ( .A(n945), .B(n946), .Z(n206) );
  NAND U283 ( .A(n206), .B(sreg[151]), .Z(n207) );
  NAND U284 ( .A(n205), .B(n207), .Z(n967) );
  NAND U285 ( .A(n1033), .B(n1034), .Z(n208) );
  XOR U286 ( .A(n1033), .B(n1034), .Z(n209) );
  NAND U287 ( .A(n209), .B(sreg[155]), .Z(n210) );
  NAND U288 ( .A(n208), .B(n210), .Z(n1055) );
  NAND U289 ( .A(n1121), .B(n1122), .Z(n211) );
  XOR U290 ( .A(n1121), .B(n1122), .Z(n212) );
  NAND U291 ( .A(n212), .B(sreg[159]), .Z(n213) );
  NAND U292 ( .A(n211), .B(n213), .Z(n1143) );
  XOR U293 ( .A(sreg[163]), .B(n1209), .Z(n214) );
  NANDN U294 ( .A(n1210), .B(n214), .Z(n215) );
  NAND U295 ( .A(sreg[163]), .B(n1209), .Z(n216) );
  AND U296 ( .A(n215), .B(n216), .Z(n1231) );
  NAND U297 ( .A(n1297), .B(n1298), .Z(n217) );
  XOR U298 ( .A(n1297), .B(n1298), .Z(n218) );
  NAND U299 ( .A(n218), .B(sreg[167]), .Z(n219) );
  NAND U300 ( .A(n217), .B(n219), .Z(n1319) );
  NAND U301 ( .A(n1385), .B(n1386), .Z(n220) );
  XOR U302 ( .A(n1385), .B(n1386), .Z(n221) );
  NAND U303 ( .A(n221), .B(sreg[171]), .Z(n222) );
  NAND U304 ( .A(n220), .B(n222), .Z(n1407) );
  NAND U305 ( .A(sreg[175]), .B(n1474), .Z(n223) );
  XOR U306 ( .A(sreg[175]), .B(n1474), .Z(n224) );
  NANDN U307 ( .A(n1473), .B(n224), .Z(n225) );
  NAND U308 ( .A(n223), .B(n225), .Z(n1495) );
  XOR U309 ( .A(sreg[179]), .B(n1561), .Z(n226) );
  NANDN U310 ( .A(n1562), .B(n226), .Z(n227) );
  NAND U311 ( .A(sreg[179]), .B(n1561), .Z(n228) );
  AND U312 ( .A(n227), .B(n228), .Z(n1583) );
  NAND U313 ( .A(n1649), .B(n1650), .Z(n229) );
  XOR U314 ( .A(n1649), .B(n1650), .Z(n230) );
  NAND U315 ( .A(n230), .B(sreg[183]), .Z(n231) );
  NAND U316 ( .A(n229), .B(n231), .Z(n1671) );
  NAND U317 ( .A(n1737), .B(n1738), .Z(n232) );
  XOR U318 ( .A(n1737), .B(n1738), .Z(n233) );
  NAND U319 ( .A(n233), .B(sreg[187]), .Z(n234) );
  NAND U320 ( .A(n232), .B(n234), .Z(n1759) );
  NAND U321 ( .A(n1825), .B(n1826), .Z(n235) );
  XOR U322 ( .A(n1825), .B(n1826), .Z(n236) );
  NANDN U323 ( .A(sreg[191]), .B(n236), .Z(n237) );
  NAND U324 ( .A(n235), .B(n237), .Z(n1847) );
  XOR U325 ( .A(sreg[195]), .B(n1913), .Z(n238) );
  NANDN U326 ( .A(n1914), .B(n238), .Z(n239) );
  NAND U327 ( .A(sreg[195]), .B(n1913), .Z(n240) );
  AND U328 ( .A(n239), .B(n240), .Z(n1935) );
  NAND U329 ( .A(n2001), .B(n2002), .Z(n241) );
  XOR U330 ( .A(n2001), .B(n2002), .Z(n242) );
  NAND U331 ( .A(n242), .B(sreg[199]), .Z(n243) );
  NAND U332 ( .A(n241), .B(n243), .Z(n2023) );
  NAND U333 ( .A(n2089), .B(n2090), .Z(n244) );
  XOR U334 ( .A(n2089), .B(n2090), .Z(n245) );
  NAND U335 ( .A(n245), .B(sreg[203]), .Z(n246) );
  NAND U336 ( .A(n244), .B(n246), .Z(n2111) );
  NAND U337 ( .A(sreg[207]), .B(n2178), .Z(n247) );
  XOR U338 ( .A(sreg[207]), .B(n2178), .Z(n248) );
  NANDN U339 ( .A(n2177), .B(n248), .Z(n249) );
  NAND U340 ( .A(n247), .B(n249), .Z(n2199) );
  XOR U341 ( .A(sreg[211]), .B(n2265), .Z(n250) );
  NANDN U342 ( .A(n2266), .B(n250), .Z(n251) );
  NAND U343 ( .A(sreg[211]), .B(n2265), .Z(n252) );
  AND U344 ( .A(n251), .B(n252), .Z(n2287) );
  NAND U345 ( .A(sreg[215]), .B(n2354), .Z(n253) );
  XOR U346 ( .A(sreg[215]), .B(n2354), .Z(n254) );
  NANDN U347 ( .A(n2353), .B(n254), .Z(n255) );
  NAND U348 ( .A(n253), .B(n255), .Z(n2375) );
  NAND U349 ( .A(n2441), .B(n2442), .Z(n256) );
  XOR U350 ( .A(n2441), .B(n2442), .Z(n257) );
  NAND U351 ( .A(n257), .B(sreg[219]), .Z(n258) );
  NAND U352 ( .A(n256), .B(n258), .Z(n2463) );
  NAND U353 ( .A(n2529), .B(n2530), .Z(n259) );
  XOR U354 ( .A(n2529), .B(n2530), .Z(n260) );
  NAND U355 ( .A(n260), .B(sreg[223]), .Z(n261) );
  NAND U356 ( .A(n259), .B(n261), .Z(n2551) );
  NAND U357 ( .A(n2617), .B(n2618), .Z(n262) );
  XOR U358 ( .A(n2617), .B(n2618), .Z(n263) );
  NAND U359 ( .A(n263), .B(sreg[227]), .Z(n264) );
  NAND U360 ( .A(n262), .B(n264), .Z(n2639) );
  NAND U361 ( .A(n2705), .B(n2706), .Z(n265) );
  XOR U362 ( .A(n2705), .B(n2706), .Z(n266) );
  NAND U363 ( .A(n266), .B(sreg[231]), .Z(n267) );
  NAND U364 ( .A(n265), .B(n267), .Z(n2727) );
  NAND U365 ( .A(n2793), .B(n2794), .Z(n268) );
  XOR U366 ( .A(n2793), .B(n2794), .Z(n269) );
  NAND U367 ( .A(n269), .B(sreg[235]), .Z(n270) );
  NAND U368 ( .A(n268), .B(n270), .Z(n2815) );
  NAND U369 ( .A(sreg[239]), .B(n2882), .Z(n271) );
  XOR U370 ( .A(sreg[239]), .B(n2882), .Z(n272) );
  NANDN U371 ( .A(n2881), .B(n272), .Z(n273) );
  NAND U372 ( .A(n271), .B(n273), .Z(n2903) );
  XOR U373 ( .A(sreg[243]), .B(n2969), .Z(n274) );
  NANDN U374 ( .A(n2970), .B(n274), .Z(n275) );
  NAND U375 ( .A(sreg[243]), .B(n2969), .Z(n276) );
  AND U376 ( .A(n275), .B(n276), .Z(n2991) );
  NAND U377 ( .A(n3057), .B(n3058), .Z(n277) );
  XOR U378 ( .A(n3057), .B(n3058), .Z(n278) );
  NAND U379 ( .A(n278), .B(sreg[247]), .Z(n279) );
  NAND U380 ( .A(n277), .B(n279), .Z(n3079) );
  NAND U381 ( .A(n3126), .B(n3127), .Z(n280) );
  XOR U382 ( .A(n3126), .B(n3127), .Z(n281) );
  NAND U383 ( .A(n281), .B(sreg[251]), .Z(n282) );
  NAND U384 ( .A(n280), .B(n282), .Z(n3147) );
  NAND U385 ( .A(n428), .B(n432), .Z(n283) );
  NAND U386 ( .A(n430), .B(n429), .Z(n284) );
  AND U387 ( .A(n283), .B(n284), .Z(n457) );
  NAND U388 ( .A(n400), .B(n399), .Z(n285) );
  NAND U389 ( .A(n398), .B(sreg[126]), .Z(n286) );
  NAND U390 ( .A(n285), .B(n286), .Z(n402) );
  NAND U391 ( .A(n483), .B(n484), .Z(n287) );
  XOR U392 ( .A(n483), .B(n484), .Z(n288) );
  NANDN U393 ( .A(sreg[130]), .B(n288), .Z(n289) );
  NAND U394 ( .A(n287), .B(n289), .Z(n505) );
  NAND U395 ( .A(n571), .B(n572), .Z(n290) );
  XOR U396 ( .A(n571), .B(n572), .Z(n291) );
  NAND U397 ( .A(n291), .B(sreg[134]), .Z(n292) );
  NAND U398 ( .A(n290), .B(n292), .Z(n593) );
  NAND U399 ( .A(n659), .B(n660), .Z(n293) );
  XOR U400 ( .A(n659), .B(n660), .Z(n294) );
  NAND U401 ( .A(n294), .B(sreg[138]), .Z(n295) );
  NAND U402 ( .A(n293), .B(n295), .Z(n681) );
  XOR U403 ( .A(sreg[142]), .B(n747), .Z(n296) );
  NANDN U404 ( .A(n748), .B(n296), .Z(n297) );
  NAND U405 ( .A(sreg[142]), .B(n747), .Z(n298) );
  AND U406 ( .A(n297), .B(n298), .Z(n769) );
  NAND U407 ( .A(n835), .B(n836), .Z(n299) );
  XOR U408 ( .A(n835), .B(n836), .Z(n300) );
  NAND U409 ( .A(n300), .B(sreg[146]), .Z(n301) );
  NAND U410 ( .A(n299), .B(n301), .Z(n857) );
  NAND U411 ( .A(sreg[150]), .B(n924), .Z(n302) );
  XOR U412 ( .A(sreg[150]), .B(n924), .Z(n303) );
  NANDN U413 ( .A(n923), .B(n303), .Z(n304) );
  NAND U414 ( .A(n302), .B(n304), .Z(n945) );
  NAND U415 ( .A(sreg[154]), .B(n1012), .Z(n305) );
  XOR U416 ( .A(sreg[154]), .B(n1012), .Z(n306) );
  NANDN U417 ( .A(n1011), .B(n306), .Z(n307) );
  NAND U418 ( .A(n305), .B(n307), .Z(n1033) );
  NAND U419 ( .A(n1099), .B(n1100), .Z(n308) );
  XOR U420 ( .A(n1099), .B(n1100), .Z(n309) );
  NAND U421 ( .A(n309), .B(sreg[158]), .Z(n310) );
  NAND U422 ( .A(n308), .B(n310), .Z(n1121) );
  NAND U423 ( .A(n1187), .B(n1188), .Z(n311) );
  XOR U424 ( .A(n1187), .B(n1188), .Z(n312) );
  NAND U425 ( .A(n312), .B(sreg[162]), .Z(n313) );
  NAND U426 ( .A(n311), .B(n313), .Z(n1209) );
  NAND U427 ( .A(sreg[166]), .B(n1276), .Z(n314) );
  XOR U428 ( .A(sreg[166]), .B(n1276), .Z(n315) );
  NANDN U429 ( .A(n1275), .B(n315), .Z(n316) );
  NAND U430 ( .A(n314), .B(n316), .Z(n1297) );
  NAND U431 ( .A(n1363), .B(n1364), .Z(n317) );
  XOR U432 ( .A(n1363), .B(n1364), .Z(n318) );
  NAND U433 ( .A(n318), .B(sreg[170]), .Z(n319) );
  NAND U434 ( .A(n317), .B(n319), .Z(n1385) );
  XOR U435 ( .A(sreg[174]), .B(n1451), .Z(n320) );
  NANDN U436 ( .A(n1452), .B(n320), .Z(n321) );
  NAND U437 ( .A(sreg[174]), .B(n1451), .Z(n322) );
  AND U438 ( .A(n321), .B(n322), .Z(n1473) );
  NAND U439 ( .A(n1539), .B(n1540), .Z(n323) );
  XOR U440 ( .A(n1539), .B(n1540), .Z(n324) );
  NAND U441 ( .A(n324), .B(sreg[178]), .Z(n325) );
  NAND U442 ( .A(n323), .B(n325), .Z(n1561) );
  NAND U443 ( .A(n1627), .B(n1628), .Z(n326) );
  XOR U444 ( .A(n1627), .B(n1628), .Z(n327) );
  NAND U445 ( .A(n327), .B(sreg[182]), .Z(n328) );
  NAND U446 ( .A(n326), .B(n328), .Z(n1649) );
  NAND U447 ( .A(n1715), .B(n1716), .Z(n329) );
  XOR U448 ( .A(n1715), .B(n1716), .Z(n330) );
  NAND U449 ( .A(n330), .B(sreg[186]), .Z(n331) );
  NAND U450 ( .A(n329), .B(n331), .Z(n1737) );
  XOR U451 ( .A(sreg[190]), .B(n1803), .Z(n332) );
  NANDN U452 ( .A(n1804), .B(n332), .Z(n333) );
  NAND U453 ( .A(sreg[190]), .B(n1803), .Z(n334) );
  AND U454 ( .A(n333), .B(n334), .Z(n1825) );
  NAND U455 ( .A(n1891), .B(n1892), .Z(n335) );
  XOR U456 ( .A(n1891), .B(n1892), .Z(n336) );
  NAND U457 ( .A(n336), .B(sreg[194]), .Z(n337) );
  NAND U458 ( .A(n335), .B(n337), .Z(n1913) );
  NAND U459 ( .A(sreg[198]), .B(n1980), .Z(n338) );
  XOR U460 ( .A(sreg[198]), .B(n1980), .Z(n339) );
  NANDN U461 ( .A(n1979), .B(n339), .Z(n340) );
  NAND U462 ( .A(n338), .B(n340), .Z(n2001) );
  NAND U463 ( .A(n2067), .B(n2068), .Z(n341) );
  XOR U464 ( .A(n2067), .B(n2068), .Z(n342) );
  NAND U465 ( .A(n342), .B(sreg[202]), .Z(n343) );
  NAND U466 ( .A(n341), .B(n343), .Z(n2089) );
  XOR U467 ( .A(sreg[206]), .B(n2155), .Z(n344) );
  NANDN U468 ( .A(n2156), .B(n344), .Z(n345) );
  NAND U469 ( .A(sreg[206]), .B(n2155), .Z(n346) );
  AND U470 ( .A(n345), .B(n346), .Z(n2177) );
  NAND U471 ( .A(n2243), .B(n2244), .Z(n347) );
  XOR U472 ( .A(n2243), .B(n2244), .Z(n348) );
  NAND U473 ( .A(n348), .B(sreg[210]), .Z(n349) );
  NAND U474 ( .A(n347), .B(n349), .Z(n2265) );
  NAND U475 ( .A(n2331), .B(n2332), .Z(n350) );
  XOR U476 ( .A(n2331), .B(n2332), .Z(n351) );
  NANDN U477 ( .A(sreg[214]), .B(n351), .Z(n352) );
  NAND U478 ( .A(n350), .B(n352), .Z(n2353) );
  NAND U479 ( .A(n2419), .B(n2420), .Z(n353) );
  XOR U480 ( .A(n2419), .B(n2420), .Z(n354) );
  NAND U481 ( .A(n354), .B(sreg[218]), .Z(n355) );
  NAND U482 ( .A(n353), .B(n355), .Z(n2441) );
  NAND U483 ( .A(n2507), .B(n2508), .Z(n356) );
  XOR U484 ( .A(n2507), .B(n2508), .Z(n357) );
  NAND U485 ( .A(n357), .B(sreg[222]), .Z(n358) );
  NAND U486 ( .A(n356), .B(n358), .Z(n2529) );
  NAND U487 ( .A(n2595), .B(n2596), .Z(n359) );
  XOR U488 ( .A(n2595), .B(n2596), .Z(n360) );
  NAND U489 ( .A(n360), .B(sreg[226]), .Z(n361) );
  NAND U490 ( .A(n359), .B(n361), .Z(n2617) );
  NAND U491 ( .A(n2683), .B(n2684), .Z(n362) );
  XOR U492 ( .A(n2683), .B(n2684), .Z(n363) );
  NAND U493 ( .A(n363), .B(sreg[230]), .Z(n364) );
  NAND U494 ( .A(n362), .B(n364), .Z(n2705) );
  NAND U495 ( .A(n2771), .B(n2772), .Z(n365) );
  XOR U496 ( .A(n2771), .B(n2772), .Z(n366) );
  NAND U497 ( .A(n366), .B(sreg[234]), .Z(n367) );
  NAND U498 ( .A(n365), .B(n367), .Z(n2793) );
  XOR U499 ( .A(sreg[238]), .B(n2859), .Z(n368) );
  NANDN U500 ( .A(n2860), .B(n368), .Z(n369) );
  NAND U501 ( .A(sreg[238]), .B(n2859), .Z(n370) );
  AND U502 ( .A(n369), .B(n370), .Z(n2881) );
  NAND U503 ( .A(n2947), .B(n2948), .Z(n371) );
  XOR U504 ( .A(n2947), .B(n2948), .Z(n372) );
  NAND U505 ( .A(n372), .B(sreg[242]), .Z(n373) );
  NAND U506 ( .A(n371), .B(n373), .Z(n2969) );
  NAND U507 ( .A(sreg[246]), .B(n3036), .Z(n374) );
  XOR U508 ( .A(sreg[246]), .B(n3036), .Z(n375) );
  NANDN U509 ( .A(n3035), .B(n375), .Z(n376) );
  NAND U510 ( .A(n374), .B(n376), .Z(n3057) );
  NAND U511 ( .A(n3123), .B(n3124), .Z(n377) );
  XOR U512 ( .A(n3123), .B(n3124), .Z(n378) );
  NAND U513 ( .A(n378), .B(sreg[250]), .Z(n379) );
  NAND U514 ( .A(n377), .B(n379), .Z(n3126) );
  NAND U515 ( .A(n3163), .B(n3164), .Z(n380) );
  NANDN U516 ( .A(n3166), .B(n3165), .Z(n381) );
  NAND U517 ( .A(n380), .B(n381), .Z(n3170) );
  AND U518 ( .A(b[0]), .B(a[0]), .Z(n384) );
  XOR U519 ( .A(n384), .B(sreg[124]), .Z(c[124]) );
  AND U520 ( .A(a[1]), .B(b[0]), .Z(n383) );
  NAND U521 ( .A(a[0]), .B(b[1]), .Z(n382) );
  XOR U522 ( .A(n383), .B(n382), .Z(n385) );
  XNOR U523 ( .A(sreg[125]), .B(n385), .Z(n387) );
  AND U524 ( .A(n384), .B(sreg[124]), .Z(n386) );
  XOR U525 ( .A(n387), .B(n386), .Z(c[125]) );
  AND U526 ( .A(b[0]), .B(a[2]), .Z(n417) );
  NAND U527 ( .A(b[1]), .B(a[1]), .Z(n418) );
  NAND U528 ( .A(b[2]), .B(a[0]), .Z(n393) );
  XNOR U529 ( .A(n392), .B(n393), .Z(n394) );
  ANDN U530 ( .B(n384), .A(n418), .Z(n395) );
  XOR U531 ( .A(n394), .B(n395), .Z(n398) );
  XOR U532 ( .A(sreg[126]), .B(n398), .Z(n400) );
  NANDN U533 ( .A(n385), .B(sreg[125]), .Z(n389) );
  NAND U534 ( .A(n387), .B(n386), .Z(n388) );
  NAND U535 ( .A(n389), .B(n388), .Z(n399) );
  XOR U536 ( .A(n400), .B(n399), .Z(c[126]) );
  AND U537 ( .A(b[0]), .B(a[3]), .Z(n390) );
  AND U538 ( .A(a[1]), .B(b[2]), .Z(n428) );
  XOR U539 ( .A(n390), .B(n428), .Z(n407) );
  NAND U540 ( .A(b[0]), .B(a[1]), .Z(n414) );
  AND U541 ( .A(a[2]), .B(n414), .Z(n391) );
  AND U542 ( .A(b[1]), .B(n391), .Z(n416) );
  AND U543 ( .A(b[3]), .B(a[0]), .Z(n415) );
  XNOR U544 ( .A(n416), .B(n415), .Z(n406) );
  XNOR U545 ( .A(n407), .B(n406), .Z(n409) );
  NANDN U546 ( .A(n393), .B(n392), .Z(n397) );
  NAND U547 ( .A(n395), .B(n394), .Z(n396) );
  AND U548 ( .A(n397), .B(n396), .Z(n408) );
  XOR U549 ( .A(n409), .B(n408), .Z(n401) );
  XNOR U550 ( .A(n401), .B(sreg[127]), .Z(n403) );
  XOR U551 ( .A(n403), .B(n402), .Z(c[127]) );
  NANDN U552 ( .A(n401), .B(sreg[127]), .Z(n405) );
  NAND U553 ( .A(n403), .B(n402), .Z(n404) );
  NAND U554 ( .A(n405), .B(n404), .Z(n440) );
  NANDN U555 ( .A(n407), .B(n406), .Z(n411) );
  NAND U556 ( .A(n409), .B(n408), .Z(n410) );
  AND U557 ( .A(n411), .B(n410), .Z(n424) );
  AND U558 ( .A(a[1]), .B(b[3]), .Z(n413) );
  NAND U559 ( .A(a[2]), .B(b[2]), .Z(n412) );
  XNOR U560 ( .A(n413), .B(n412), .Z(n430) );
  AND U561 ( .A(b[2]), .B(a[3]), .Z(n470) );
  ANDN U562 ( .B(n470), .A(n414), .Z(n429) );
  XOR U563 ( .A(n430), .B(n429), .Z(n433) );
  NAND U564 ( .A(b[0]), .B(a[4]), .Z(n434) );
  XNOR U565 ( .A(n433), .B(n434), .Z(n436) );
  AND U566 ( .A(b[1]), .B(a[3]), .Z(n435) );
  XOR U567 ( .A(n436), .B(n435), .Z(n423) );
  NAND U568 ( .A(n416), .B(n415), .Z(n420) );
  NANDN U569 ( .A(n418), .B(n417), .Z(n419) );
  AND U570 ( .A(n420), .B(n419), .Z(n422) );
  XOR U571 ( .A(n423), .B(n422), .Z(n425) );
  XOR U572 ( .A(n424), .B(n425), .Z(n439) );
  XOR U573 ( .A(sreg[128]), .B(n439), .Z(n421) );
  XNOR U574 ( .A(n440), .B(n421), .Z(c[128]) );
  NANDN U575 ( .A(n423), .B(n422), .Z(n427) );
  OR U576 ( .A(n425), .B(n424), .Z(n426) );
  AND U577 ( .A(n427), .B(n426), .Z(n445) );
  AND U578 ( .A(b[3]), .B(a[2]), .Z(n432) );
  NAND U579 ( .A(a[3]), .B(b[2]), .Z(n431) );
  XNOR U580 ( .A(n432), .B(n431), .Z(n449) );
  NAND U581 ( .A(b[1]), .B(a[4]), .Z(n450) );
  XNOR U582 ( .A(n449), .B(n450), .Z(n455) );
  NAND U583 ( .A(b[0]), .B(a[5]), .Z(n456) );
  XOR U584 ( .A(n455), .B(n456), .Z(n458) );
  XOR U585 ( .A(n457), .B(n458), .Z(n443) );
  NANDN U586 ( .A(n434), .B(n433), .Z(n438) );
  NAND U587 ( .A(n436), .B(n435), .Z(n437) );
  AND U588 ( .A(n438), .B(n437), .Z(n442) );
  XNOR U589 ( .A(n443), .B(n442), .Z(n444) );
  XNOR U590 ( .A(n445), .B(n444), .Z(n462) );
  XOR U591 ( .A(n461), .B(sreg[129]), .Z(n441) );
  XNOR U592 ( .A(n462), .B(n441), .Z(c[129]) );
  NANDN U593 ( .A(n443), .B(n442), .Z(n447) );
  NANDN U594 ( .A(n445), .B(n444), .Z(n446) );
  AND U595 ( .A(n447), .B(n446), .Z(n467) );
  AND U596 ( .A(b[3]), .B(a[3]), .Z(n454) );
  AND U597 ( .A(b[2]), .B(a[2]), .Z(n448) );
  NAND U598 ( .A(n454), .B(n448), .Z(n452) );
  NANDN U599 ( .A(n450), .B(n449), .Z(n451) );
  AND U600 ( .A(n452), .B(n451), .Z(n479) );
  NAND U601 ( .A(a[4]), .B(b[2]), .Z(n453) );
  XNOR U602 ( .A(n454), .B(n453), .Z(n471) );
  NAND U603 ( .A(b[1]), .B(a[5]), .Z(n472) );
  XNOR U604 ( .A(n471), .B(n472), .Z(n477) );
  NAND U605 ( .A(b[0]), .B(a[6]), .Z(n478) );
  XOR U606 ( .A(n477), .B(n478), .Z(n480) );
  XOR U607 ( .A(n479), .B(n480), .Z(n465) );
  NANDN U608 ( .A(n456), .B(n455), .Z(n460) );
  OR U609 ( .A(n458), .B(n457), .Z(n459) );
  AND U610 ( .A(n460), .B(n459), .Z(n464) );
  XNOR U611 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U612 ( .A(n467), .B(n466), .Z(n484) );
  XNOR U613 ( .A(n483), .B(sreg[130]), .Z(n463) );
  XNOR U614 ( .A(n484), .B(n463), .Z(c[130]) );
  NANDN U615 ( .A(n465), .B(n464), .Z(n469) );
  NANDN U616 ( .A(n467), .B(n466), .Z(n468) );
  AND U617 ( .A(n469), .B(n468), .Z(n488) );
  AND U618 ( .A(b[3]), .B(a[4]), .Z(n476) );
  NAND U619 ( .A(n476), .B(n470), .Z(n474) );
  NANDN U620 ( .A(n472), .B(n471), .Z(n473) );
  AND U621 ( .A(n474), .B(n473), .Z(n501) );
  NAND U622 ( .A(a[5]), .B(b[2]), .Z(n475) );
  XNOR U623 ( .A(n476), .B(n475), .Z(n493) );
  NAND U624 ( .A(b[1]), .B(a[6]), .Z(n494) );
  XNOR U625 ( .A(n493), .B(n494), .Z(n499) );
  NAND U626 ( .A(b[0]), .B(a[7]), .Z(n500) );
  XOR U627 ( .A(n499), .B(n500), .Z(n502) );
  XOR U628 ( .A(n501), .B(n502), .Z(n487) );
  NANDN U629 ( .A(n478), .B(n477), .Z(n482) );
  OR U630 ( .A(n480), .B(n479), .Z(n481) );
  AND U631 ( .A(n482), .B(n481), .Z(n486) );
  XOR U632 ( .A(n487), .B(n486), .Z(n489) );
  XNOR U633 ( .A(n488), .B(n489), .Z(n506) );
  XOR U634 ( .A(sreg[131]), .B(n505), .Z(n485) );
  XNOR U635 ( .A(n506), .B(n485), .Z(c[131]) );
  NANDN U636 ( .A(n487), .B(n486), .Z(n491) );
  OR U637 ( .A(n489), .B(n488), .Z(n490) );
  AND U638 ( .A(n491), .B(n490), .Z(n511) );
  AND U639 ( .A(b[3]), .B(a[5]), .Z(n498) );
  AND U640 ( .A(b[2]), .B(a[4]), .Z(n492) );
  NAND U641 ( .A(n498), .B(n492), .Z(n496) );
  NANDN U642 ( .A(n494), .B(n493), .Z(n495) );
  AND U643 ( .A(n496), .B(n495), .Z(n523) );
  NAND U644 ( .A(a[6]), .B(b[2]), .Z(n497) );
  XNOR U645 ( .A(n498), .B(n497), .Z(n515) );
  NAND U646 ( .A(b[1]), .B(a[7]), .Z(n516) );
  XNOR U647 ( .A(n515), .B(n516), .Z(n521) );
  NAND U648 ( .A(b[0]), .B(a[8]), .Z(n522) );
  XOR U649 ( .A(n521), .B(n522), .Z(n524) );
  XOR U650 ( .A(n523), .B(n524), .Z(n509) );
  NANDN U651 ( .A(n500), .B(n499), .Z(n504) );
  OR U652 ( .A(n502), .B(n501), .Z(n503) );
  AND U653 ( .A(n504), .B(n503), .Z(n508) );
  XNOR U654 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U655 ( .A(n511), .B(n510), .Z(n528) );
  XOR U656 ( .A(n527), .B(sreg[132]), .Z(n507) );
  XNOR U657 ( .A(n528), .B(n507), .Z(c[132]) );
  NANDN U658 ( .A(n509), .B(n508), .Z(n513) );
  NANDN U659 ( .A(n511), .B(n510), .Z(n512) );
  AND U660 ( .A(n513), .B(n512), .Z(n532) );
  AND U661 ( .A(b[3]), .B(a[6]), .Z(n520) );
  AND U662 ( .A(b[2]), .B(a[5]), .Z(n514) );
  NAND U663 ( .A(n520), .B(n514), .Z(n518) );
  NANDN U664 ( .A(n516), .B(n515), .Z(n517) );
  AND U665 ( .A(n518), .B(n517), .Z(n545) );
  NAND U666 ( .A(a[7]), .B(b[2]), .Z(n519) );
  XNOR U667 ( .A(n520), .B(n519), .Z(n537) );
  NAND U668 ( .A(b[1]), .B(a[8]), .Z(n538) );
  XNOR U669 ( .A(n537), .B(n538), .Z(n543) );
  NAND U670 ( .A(b[0]), .B(a[9]), .Z(n544) );
  XOR U671 ( .A(n543), .B(n544), .Z(n546) );
  XOR U672 ( .A(n545), .B(n546), .Z(n531) );
  NANDN U673 ( .A(n522), .B(n521), .Z(n526) );
  OR U674 ( .A(n524), .B(n523), .Z(n525) );
  AND U675 ( .A(n526), .B(n525), .Z(n530) );
  XOR U676 ( .A(n531), .B(n530), .Z(n533) );
  XNOR U677 ( .A(n532), .B(n533), .Z(n550) );
  XOR U678 ( .A(sreg[133]), .B(n549), .Z(n529) );
  XNOR U679 ( .A(n550), .B(n529), .Z(c[133]) );
  NANDN U680 ( .A(n531), .B(n530), .Z(n535) );
  OR U681 ( .A(n533), .B(n532), .Z(n534) );
  AND U682 ( .A(n535), .B(n534), .Z(n554) );
  AND U683 ( .A(b[3]), .B(a[7]), .Z(n542) );
  AND U684 ( .A(b[2]), .B(a[6]), .Z(n536) );
  NAND U685 ( .A(n542), .B(n536), .Z(n540) );
  NANDN U686 ( .A(n538), .B(n537), .Z(n539) );
  AND U687 ( .A(n540), .B(n539), .Z(n567) );
  NAND U688 ( .A(a[8]), .B(b[2]), .Z(n541) );
  XNOR U689 ( .A(n542), .B(n541), .Z(n559) );
  NAND U690 ( .A(b[1]), .B(a[9]), .Z(n560) );
  XNOR U691 ( .A(n559), .B(n560), .Z(n565) );
  NAND U692 ( .A(b[0]), .B(a[10]), .Z(n566) );
  XOR U693 ( .A(n565), .B(n566), .Z(n568) );
  XOR U694 ( .A(n567), .B(n568), .Z(n553) );
  NANDN U695 ( .A(n544), .B(n543), .Z(n548) );
  OR U696 ( .A(n546), .B(n545), .Z(n547) );
  AND U697 ( .A(n548), .B(n547), .Z(n552) );
  XOR U698 ( .A(n553), .B(n552), .Z(n555) );
  XNOR U699 ( .A(n554), .B(n555), .Z(n572) );
  XNOR U700 ( .A(sreg[134]), .B(n571), .Z(n551) );
  XNOR U701 ( .A(n572), .B(n551), .Z(c[134]) );
  NANDN U702 ( .A(n553), .B(n552), .Z(n557) );
  OR U703 ( .A(n555), .B(n554), .Z(n556) );
  AND U704 ( .A(n557), .B(n556), .Z(n576) );
  AND U705 ( .A(b[3]), .B(a[8]), .Z(n564) );
  AND U706 ( .A(b[2]), .B(a[7]), .Z(n558) );
  NAND U707 ( .A(n564), .B(n558), .Z(n562) );
  NANDN U708 ( .A(n560), .B(n559), .Z(n561) );
  AND U709 ( .A(n562), .B(n561), .Z(n589) );
  NAND U710 ( .A(a[9]), .B(b[2]), .Z(n563) );
  XNOR U711 ( .A(n564), .B(n563), .Z(n581) );
  NAND U712 ( .A(b[1]), .B(a[10]), .Z(n582) );
  XNOR U713 ( .A(n581), .B(n582), .Z(n587) );
  NAND U714 ( .A(b[0]), .B(a[11]), .Z(n588) );
  XOR U715 ( .A(n587), .B(n588), .Z(n590) );
  XOR U716 ( .A(n589), .B(n590), .Z(n575) );
  NANDN U717 ( .A(n566), .B(n565), .Z(n570) );
  OR U718 ( .A(n568), .B(n567), .Z(n569) );
  AND U719 ( .A(n570), .B(n569), .Z(n574) );
  XOR U720 ( .A(n575), .B(n574), .Z(n577) );
  XNOR U721 ( .A(n576), .B(n577), .Z(n594) );
  XNOR U722 ( .A(sreg[135]), .B(n593), .Z(n573) );
  XNOR U723 ( .A(n594), .B(n573), .Z(c[135]) );
  NANDN U724 ( .A(n575), .B(n574), .Z(n579) );
  OR U725 ( .A(n577), .B(n576), .Z(n578) );
  AND U726 ( .A(n579), .B(n578), .Z(n598) );
  AND U727 ( .A(b[3]), .B(a[9]), .Z(n586) );
  AND U728 ( .A(b[2]), .B(a[8]), .Z(n580) );
  NAND U729 ( .A(n586), .B(n580), .Z(n584) );
  NANDN U730 ( .A(n582), .B(n581), .Z(n583) );
  AND U731 ( .A(n584), .B(n583), .Z(n611) );
  NAND U732 ( .A(a[10]), .B(b[2]), .Z(n585) );
  XNOR U733 ( .A(n586), .B(n585), .Z(n603) );
  NAND U734 ( .A(b[1]), .B(a[11]), .Z(n604) );
  XNOR U735 ( .A(n603), .B(n604), .Z(n609) );
  NAND U736 ( .A(b[0]), .B(a[12]), .Z(n610) );
  XOR U737 ( .A(n609), .B(n610), .Z(n612) );
  XOR U738 ( .A(n611), .B(n612), .Z(n597) );
  NANDN U739 ( .A(n588), .B(n587), .Z(n592) );
  OR U740 ( .A(n590), .B(n589), .Z(n591) );
  AND U741 ( .A(n592), .B(n591), .Z(n596) );
  XOR U742 ( .A(n597), .B(n596), .Z(n599) );
  XNOR U743 ( .A(n598), .B(n599), .Z(n616) );
  XNOR U744 ( .A(sreg[136]), .B(n615), .Z(n595) );
  XNOR U745 ( .A(n616), .B(n595), .Z(c[136]) );
  NANDN U746 ( .A(n597), .B(n596), .Z(n601) );
  OR U747 ( .A(n599), .B(n598), .Z(n600) );
  AND U748 ( .A(n601), .B(n600), .Z(n620) );
  AND U749 ( .A(b[3]), .B(a[10]), .Z(n608) );
  AND U750 ( .A(b[2]), .B(a[9]), .Z(n602) );
  NAND U751 ( .A(n608), .B(n602), .Z(n606) );
  NANDN U752 ( .A(n604), .B(n603), .Z(n605) );
  AND U753 ( .A(n606), .B(n605), .Z(n633) );
  NAND U754 ( .A(a[11]), .B(b[2]), .Z(n607) );
  XNOR U755 ( .A(n608), .B(n607), .Z(n625) );
  NAND U756 ( .A(b[1]), .B(a[12]), .Z(n626) );
  XNOR U757 ( .A(n625), .B(n626), .Z(n631) );
  NAND U758 ( .A(b[0]), .B(a[13]), .Z(n632) );
  XOR U759 ( .A(n631), .B(n632), .Z(n634) );
  XOR U760 ( .A(n633), .B(n634), .Z(n619) );
  NANDN U761 ( .A(n610), .B(n609), .Z(n614) );
  OR U762 ( .A(n612), .B(n611), .Z(n613) );
  AND U763 ( .A(n614), .B(n613), .Z(n618) );
  XOR U764 ( .A(n619), .B(n618), .Z(n621) );
  XNOR U765 ( .A(n620), .B(n621), .Z(n638) );
  XNOR U766 ( .A(sreg[137]), .B(n637), .Z(n617) );
  XNOR U767 ( .A(n638), .B(n617), .Z(c[137]) );
  NANDN U768 ( .A(n619), .B(n618), .Z(n623) );
  OR U769 ( .A(n621), .B(n620), .Z(n622) );
  AND U770 ( .A(n623), .B(n622), .Z(n642) );
  AND U771 ( .A(b[3]), .B(a[11]), .Z(n630) );
  AND U772 ( .A(b[2]), .B(a[10]), .Z(n624) );
  NAND U773 ( .A(n630), .B(n624), .Z(n628) );
  NANDN U774 ( .A(n626), .B(n625), .Z(n627) );
  AND U775 ( .A(n628), .B(n627), .Z(n655) );
  NAND U776 ( .A(a[12]), .B(b[2]), .Z(n629) );
  XNOR U777 ( .A(n630), .B(n629), .Z(n647) );
  NAND U778 ( .A(b[1]), .B(a[13]), .Z(n648) );
  XNOR U779 ( .A(n647), .B(n648), .Z(n653) );
  NAND U780 ( .A(b[0]), .B(a[14]), .Z(n654) );
  XOR U781 ( .A(n653), .B(n654), .Z(n656) );
  XOR U782 ( .A(n655), .B(n656), .Z(n641) );
  NANDN U783 ( .A(n632), .B(n631), .Z(n636) );
  OR U784 ( .A(n634), .B(n633), .Z(n635) );
  AND U785 ( .A(n636), .B(n635), .Z(n640) );
  XOR U786 ( .A(n641), .B(n640), .Z(n643) );
  XNOR U787 ( .A(n642), .B(n643), .Z(n660) );
  XNOR U788 ( .A(sreg[138]), .B(n659), .Z(n639) );
  XNOR U789 ( .A(n660), .B(n639), .Z(c[138]) );
  NANDN U790 ( .A(n641), .B(n640), .Z(n645) );
  OR U791 ( .A(n643), .B(n642), .Z(n644) );
  AND U792 ( .A(n645), .B(n644), .Z(n664) );
  AND U793 ( .A(b[3]), .B(a[12]), .Z(n652) );
  AND U794 ( .A(b[2]), .B(a[11]), .Z(n646) );
  NAND U795 ( .A(n652), .B(n646), .Z(n650) );
  NANDN U796 ( .A(n648), .B(n647), .Z(n649) );
  AND U797 ( .A(n650), .B(n649), .Z(n677) );
  NAND U798 ( .A(a[13]), .B(b[2]), .Z(n651) );
  XNOR U799 ( .A(n652), .B(n651), .Z(n669) );
  NAND U800 ( .A(b[1]), .B(a[14]), .Z(n670) );
  XNOR U801 ( .A(n669), .B(n670), .Z(n675) );
  NAND U802 ( .A(b[0]), .B(a[15]), .Z(n676) );
  XOR U803 ( .A(n675), .B(n676), .Z(n678) );
  XOR U804 ( .A(n677), .B(n678), .Z(n663) );
  NANDN U805 ( .A(n654), .B(n653), .Z(n658) );
  OR U806 ( .A(n656), .B(n655), .Z(n657) );
  AND U807 ( .A(n658), .B(n657), .Z(n662) );
  XOR U808 ( .A(n663), .B(n662), .Z(n665) );
  XNOR U809 ( .A(n664), .B(n665), .Z(n682) );
  XNOR U810 ( .A(sreg[139]), .B(n681), .Z(n661) );
  XNOR U811 ( .A(n682), .B(n661), .Z(c[139]) );
  NANDN U812 ( .A(n663), .B(n662), .Z(n667) );
  OR U813 ( .A(n665), .B(n664), .Z(n666) );
  AND U814 ( .A(n667), .B(n666), .Z(n686) );
  AND U815 ( .A(b[3]), .B(a[13]), .Z(n674) );
  AND U816 ( .A(b[2]), .B(a[12]), .Z(n668) );
  NAND U817 ( .A(n674), .B(n668), .Z(n672) );
  NANDN U818 ( .A(n670), .B(n669), .Z(n671) );
  AND U819 ( .A(n672), .B(n671), .Z(n699) );
  NAND U820 ( .A(a[14]), .B(b[2]), .Z(n673) );
  XNOR U821 ( .A(n674), .B(n673), .Z(n691) );
  NAND U822 ( .A(b[1]), .B(a[15]), .Z(n692) );
  XNOR U823 ( .A(n691), .B(n692), .Z(n697) );
  NAND U824 ( .A(b[0]), .B(a[16]), .Z(n698) );
  XOR U825 ( .A(n697), .B(n698), .Z(n700) );
  XOR U826 ( .A(n699), .B(n700), .Z(n685) );
  NANDN U827 ( .A(n676), .B(n675), .Z(n680) );
  OR U828 ( .A(n678), .B(n677), .Z(n679) );
  AND U829 ( .A(n680), .B(n679), .Z(n684) );
  XOR U830 ( .A(n685), .B(n684), .Z(n687) );
  XNOR U831 ( .A(n686), .B(n687), .Z(n704) );
  XNOR U832 ( .A(sreg[140]), .B(n703), .Z(n683) );
  XNOR U833 ( .A(n704), .B(n683), .Z(c[140]) );
  NANDN U834 ( .A(n685), .B(n684), .Z(n689) );
  OR U835 ( .A(n687), .B(n686), .Z(n688) );
  AND U836 ( .A(n689), .B(n688), .Z(n708) );
  AND U837 ( .A(b[3]), .B(a[14]), .Z(n696) );
  AND U838 ( .A(b[2]), .B(a[13]), .Z(n690) );
  NAND U839 ( .A(n696), .B(n690), .Z(n694) );
  NANDN U840 ( .A(n692), .B(n691), .Z(n693) );
  AND U841 ( .A(n694), .B(n693), .Z(n721) );
  NAND U842 ( .A(a[15]), .B(b[2]), .Z(n695) );
  XNOR U843 ( .A(n696), .B(n695), .Z(n713) );
  NAND U844 ( .A(b[1]), .B(a[16]), .Z(n714) );
  XNOR U845 ( .A(n713), .B(n714), .Z(n719) );
  NAND U846 ( .A(b[0]), .B(a[17]), .Z(n720) );
  XOR U847 ( .A(n719), .B(n720), .Z(n722) );
  XOR U848 ( .A(n721), .B(n722), .Z(n707) );
  NANDN U849 ( .A(n698), .B(n697), .Z(n702) );
  OR U850 ( .A(n700), .B(n699), .Z(n701) );
  AND U851 ( .A(n702), .B(n701), .Z(n706) );
  XOR U852 ( .A(n707), .B(n706), .Z(n709) );
  XNOR U853 ( .A(n708), .B(n709), .Z(n726) );
  XNOR U854 ( .A(sreg[141]), .B(n725), .Z(n705) );
  XNOR U855 ( .A(n726), .B(n705), .Z(c[141]) );
  NANDN U856 ( .A(n707), .B(n706), .Z(n711) );
  OR U857 ( .A(n709), .B(n708), .Z(n710) );
  AND U858 ( .A(n711), .B(n710), .Z(n731) );
  AND U859 ( .A(b[3]), .B(a[15]), .Z(n718) );
  AND U860 ( .A(b[2]), .B(a[14]), .Z(n712) );
  NAND U861 ( .A(n718), .B(n712), .Z(n716) );
  NANDN U862 ( .A(n714), .B(n713), .Z(n715) );
  AND U863 ( .A(n716), .B(n715), .Z(n743) );
  NAND U864 ( .A(a[16]), .B(b[2]), .Z(n717) );
  XNOR U865 ( .A(n718), .B(n717), .Z(n735) );
  NAND U866 ( .A(b[1]), .B(a[17]), .Z(n736) );
  XNOR U867 ( .A(n735), .B(n736), .Z(n741) );
  NAND U868 ( .A(b[0]), .B(a[18]), .Z(n742) );
  XOR U869 ( .A(n741), .B(n742), .Z(n744) );
  XOR U870 ( .A(n743), .B(n744), .Z(n729) );
  NANDN U871 ( .A(n720), .B(n719), .Z(n724) );
  OR U872 ( .A(n722), .B(n721), .Z(n723) );
  AND U873 ( .A(n724), .B(n723), .Z(n728) );
  XNOR U874 ( .A(n729), .B(n728), .Z(n730) );
  XNOR U875 ( .A(n731), .B(n730), .Z(n748) );
  XOR U876 ( .A(n747), .B(sreg[142]), .Z(n727) );
  XNOR U877 ( .A(n748), .B(n727), .Z(c[142]) );
  NANDN U878 ( .A(n729), .B(n728), .Z(n733) );
  NANDN U879 ( .A(n731), .B(n730), .Z(n732) );
  AND U880 ( .A(n733), .B(n732), .Z(n752) );
  AND U881 ( .A(b[3]), .B(a[16]), .Z(n740) );
  AND U882 ( .A(b[2]), .B(a[15]), .Z(n734) );
  NAND U883 ( .A(n740), .B(n734), .Z(n738) );
  NANDN U884 ( .A(n736), .B(n735), .Z(n737) );
  AND U885 ( .A(n738), .B(n737), .Z(n765) );
  NAND U886 ( .A(a[17]), .B(b[2]), .Z(n739) );
  XNOR U887 ( .A(n740), .B(n739), .Z(n757) );
  NAND U888 ( .A(b[1]), .B(a[18]), .Z(n758) );
  XNOR U889 ( .A(n757), .B(n758), .Z(n763) );
  NAND U890 ( .A(b[0]), .B(a[19]), .Z(n764) );
  XOR U891 ( .A(n763), .B(n764), .Z(n766) );
  XOR U892 ( .A(n765), .B(n766), .Z(n751) );
  NANDN U893 ( .A(n742), .B(n741), .Z(n746) );
  OR U894 ( .A(n744), .B(n743), .Z(n745) );
  AND U895 ( .A(n746), .B(n745), .Z(n750) );
  XOR U896 ( .A(n751), .B(n750), .Z(n753) );
  XNOR U897 ( .A(n752), .B(n753), .Z(n770) );
  XOR U898 ( .A(sreg[143]), .B(n769), .Z(n749) );
  XNOR U899 ( .A(n770), .B(n749), .Z(c[143]) );
  NANDN U900 ( .A(n751), .B(n750), .Z(n755) );
  OR U901 ( .A(n753), .B(n752), .Z(n754) );
  AND U902 ( .A(n755), .B(n754), .Z(n774) );
  AND U903 ( .A(b[3]), .B(a[17]), .Z(n762) );
  AND U904 ( .A(b[2]), .B(a[16]), .Z(n756) );
  NAND U905 ( .A(n762), .B(n756), .Z(n760) );
  NANDN U906 ( .A(n758), .B(n757), .Z(n759) );
  AND U907 ( .A(n760), .B(n759), .Z(n787) );
  NAND U908 ( .A(a[18]), .B(b[2]), .Z(n761) );
  XNOR U909 ( .A(n762), .B(n761), .Z(n779) );
  NAND U910 ( .A(b[1]), .B(a[19]), .Z(n780) );
  XNOR U911 ( .A(n779), .B(n780), .Z(n785) );
  NAND U912 ( .A(b[0]), .B(a[20]), .Z(n786) );
  XOR U913 ( .A(n785), .B(n786), .Z(n788) );
  XOR U914 ( .A(n787), .B(n788), .Z(n773) );
  NANDN U915 ( .A(n764), .B(n763), .Z(n768) );
  OR U916 ( .A(n766), .B(n765), .Z(n767) );
  AND U917 ( .A(n768), .B(n767), .Z(n772) );
  XOR U918 ( .A(n773), .B(n772), .Z(n775) );
  XNOR U919 ( .A(n774), .B(n775), .Z(n792) );
  XNOR U920 ( .A(sreg[144]), .B(n791), .Z(n771) );
  XNOR U921 ( .A(n792), .B(n771), .Z(c[144]) );
  NANDN U922 ( .A(n773), .B(n772), .Z(n777) );
  OR U923 ( .A(n775), .B(n774), .Z(n776) );
  AND U924 ( .A(n777), .B(n776), .Z(n796) );
  AND U925 ( .A(b[3]), .B(a[18]), .Z(n784) );
  AND U926 ( .A(b[2]), .B(a[17]), .Z(n778) );
  NAND U927 ( .A(n784), .B(n778), .Z(n782) );
  NANDN U928 ( .A(n780), .B(n779), .Z(n781) );
  AND U929 ( .A(n782), .B(n781), .Z(n809) );
  NAND U930 ( .A(a[19]), .B(b[2]), .Z(n783) );
  XNOR U931 ( .A(n784), .B(n783), .Z(n801) );
  NAND U932 ( .A(b[1]), .B(a[20]), .Z(n802) );
  XNOR U933 ( .A(n801), .B(n802), .Z(n807) );
  NAND U934 ( .A(b[0]), .B(a[21]), .Z(n808) );
  XOR U935 ( .A(n807), .B(n808), .Z(n810) );
  XOR U936 ( .A(n809), .B(n810), .Z(n795) );
  NANDN U937 ( .A(n786), .B(n785), .Z(n790) );
  OR U938 ( .A(n788), .B(n787), .Z(n789) );
  AND U939 ( .A(n790), .B(n789), .Z(n794) );
  XOR U940 ( .A(n795), .B(n794), .Z(n797) );
  XNOR U941 ( .A(n796), .B(n797), .Z(n814) );
  XNOR U942 ( .A(sreg[145]), .B(n813), .Z(n793) );
  XNOR U943 ( .A(n814), .B(n793), .Z(c[145]) );
  NANDN U944 ( .A(n795), .B(n794), .Z(n799) );
  OR U945 ( .A(n797), .B(n796), .Z(n798) );
  AND U946 ( .A(n799), .B(n798), .Z(n818) );
  AND U947 ( .A(b[3]), .B(a[19]), .Z(n806) );
  AND U948 ( .A(b[2]), .B(a[18]), .Z(n800) );
  NAND U949 ( .A(n806), .B(n800), .Z(n804) );
  NANDN U950 ( .A(n802), .B(n801), .Z(n803) );
  AND U951 ( .A(n804), .B(n803), .Z(n831) );
  NAND U952 ( .A(a[20]), .B(b[2]), .Z(n805) );
  XNOR U953 ( .A(n806), .B(n805), .Z(n823) );
  NAND U954 ( .A(b[1]), .B(a[21]), .Z(n824) );
  XNOR U955 ( .A(n823), .B(n824), .Z(n829) );
  NAND U956 ( .A(b[0]), .B(a[22]), .Z(n830) );
  XOR U957 ( .A(n829), .B(n830), .Z(n832) );
  XOR U958 ( .A(n831), .B(n832), .Z(n817) );
  NANDN U959 ( .A(n808), .B(n807), .Z(n812) );
  OR U960 ( .A(n810), .B(n809), .Z(n811) );
  AND U961 ( .A(n812), .B(n811), .Z(n816) );
  XOR U962 ( .A(n817), .B(n816), .Z(n819) );
  XNOR U963 ( .A(n818), .B(n819), .Z(n836) );
  XNOR U964 ( .A(sreg[146]), .B(n835), .Z(n815) );
  XNOR U965 ( .A(n836), .B(n815), .Z(c[146]) );
  NANDN U966 ( .A(n817), .B(n816), .Z(n821) );
  OR U967 ( .A(n819), .B(n818), .Z(n820) );
  AND U968 ( .A(n821), .B(n820), .Z(n841) );
  AND U969 ( .A(b[3]), .B(a[20]), .Z(n828) );
  AND U970 ( .A(b[2]), .B(a[19]), .Z(n822) );
  NAND U971 ( .A(n828), .B(n822), .Z(n826) );
  NANDN U972 ( .A(n824), .B(n823), .Z(n825) );
  AND U973 ( .A(n826), .B(n825), .Z(n853) );
  NAND U974 ( .A(a[21]), .B(b[2]), .Z(n827) );
  XNOR U975 ( .A(n828), .B(n827), .Z(n845) );
  NAND U976 ( .A(b[1]), .B(a[22]), .Z(n846) );
  XNOR U977 ( .A(n845), .B(n846), .Z(n851) );
  NAND U978 ( .A(b[0]), .B(a[23]), .Z(n852) );
  XOR U979 ( .A(n851), .B(n852), .Z(n854) );
  XOR U980 ( .A(n853), .B(n854), .Z(n839) );
  NANDN U981 ( .A(n830), .B(n829), .Z(n834) );
  OR U982 ( .A(n832), .B(n831), .Z(n833) );
  AND U983 ( .A(n834), .B(n833), .Z(n838) );
  XNOR U984 ( .A(n839), .B(n838), .Z(n840) );
  XNOR U985 ( .A(n841), .B(n840), .Z(n858) );
  XOR U986 ( .A(n857), .B(sreg[147]), .Z(n837) );
  XNOR U987 ( .A(n858), .B(n837), .Z(c[147]) );
  NANDN U988 ( .A(n839), .B(n838), .Z(n843) );
  NANDN U989 ( .A(n841), .B(n840), .Z(n842) );
  AND U990 ( .A(n843), .B(n842), .Z(n862) );
  AND U991 ( .A(b[3]), .B(a[21]), .Z(n850) );
  AND U992 ( .A(b[2]), .B(a[20]), .Z(n844) );
  NAND U993 ( .A(n850), .B(n844), .Z(n848) );
  NANDN U994 ( .A(n846), .B(n845), .Z(n847) );
  AND U995 ( .A(n848), .B(n847), .Z(n875) );
  NAND U996 ( .A(a[22]), .B(b[2]), .Z(n849) );
  XNOR U997 ( .A(n850), .B(n849), .Z(n867) );
  NAND U998 ( .A(b[1]), .B(a[23]), .Z(n868) );
  XNOR U999 ( .A(n867), .B(n868), .Z(n873) );
  NAND U1000 ( .A(b[0]), .B(a[24]), .Z(n874) );
  XOR U1001 ( .A(n873), .B(n874), .Z(n876) );
  XOR U1002 ( .A(n875), .B(n876), .Z(n861) );
  NANDN U1003 ( .A(n852), .B(n851), .Z(n856) );
  OR U1004 ( .A(n854), .B(n853), .Z(n855) );
  AND U1005 ( .A(n856), .B(n855), .Z(n860) );
  XOR U1006 ( .A(n861), .B(n860), .Z(n863) );
  XNOR U1007 ( .A(n862), .B(n863), .Z(n880) );
  XOR U1008 ( .A(sreg[148]), .B(n879), .Z(n859) );
  XNOR U1009 ( .A(n880), .B(n859), .Z(c[148]) );
  NANDN U1010 ( .A(n861), .B(n860), .Z(n865) );
  OR U1011 ( .A(n863), .B(n862), .Z(n864) );
  AND U1012 ( .A(n865), .B(n864), .Z(n885) );
  AND U1013 ( .A(b[3]), .B(a[22]), .Z(n872) );
  AND U1014 ( .A(b[2]), .B(a[21]), .Z(n866) );
  NAND U1015 ( .A(n872), .B(n866), .Z(n870) );
  NANDN U1016 ( .A(n868), .B(n867), .Z(n869) );
  AND U1017 ( .A(n870), .B(n869), .Z(n897) );
  NAND U1018 ( .A(a[23]), .B(b[2]), .Z(n871) );
  XNOR U1019 ( .A(n872), .B(n871), .Z(n889) );
  NAND U1020 ( .A(b[1]), .B(a[24]), .Z(n890) );
  XNOR U1021 ( .A(n889), .B(n890), .Z(n895) );
  NAND U1022 ( .A(b[0]), .B(a[25]), .Z(n896) );
  XOR U1023 ( .A(n895), .B(n896), .Z(n898) );
  XOR U1024 ( .A(n897), .B(n898), .Z(n883) );
  NANDN U1025 ( .A(n874), .B(n873), .Z(n878) );
  OR U1026 ( .A(n876), .B(n875), .Z(n877) );
  AND U1027 ( .A(n878), .B(n877), .Z(n882) );
  XNOR U1028 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U1029 ( .A(n885), .B(n884), .Z(n902) );
  XOR U1030 ( .A(n901), .B(sreg[149]), .Z(n881) );
  XNOR U1031 ( .A(n902), .B(n881), .Z(c[149]) );
  NANDN U1032 ( .A(n883), .B(n882), .Z(n887) );
  NANDN U1033 ( .A(n885), .B(n884), .Z(n886) );
  AND U1034 ( .A(n887), .B(n886), .Z(n906) );
  AND U1035 ( .A(b[3]), .B(a[23]), .Z(n894) );
  AND U1036 ( .A(b[2]), .B(a[22]), .Z(n888) );
  NAND U1037 ( .A(n894), .B(n888), .Z(n892) );
  NANDN U1038 ( .A(n890), .B(n889), .Z(n891) );
  AND U1039 ( .A(n892), .B(n891), .Z(n919) );
  NAND U1040 ( .A(a[24]), .B(b[2]), .Z(n893) );
  XNOR U1041 ( .A(n894), .B(n893), .Z(n911) );
  NAND U1042 ( .A(b[1]), .B(a[25]), .Z(n912) );
  XNOR U1043 ( .A(n911), .B(n912), .Z(n917) );
  NAND U1044 ( .A(b[0]), .B(a[26]), .Z(n918) );
  XOR U1045 ( .A(n917), .B(n918), .Z(n920) );
  XOR U1046 ( .A(n919), .B(n920), .Z(n905) );
  NANDN U1047 ( .A(n896), .B(n895), .Z(n900) );
  OR U1048 ( .A(n898), .B(n897), .Z(n899) );
  AND U1049 ( .A(n900), .B(n899), .Z(n904) );
  XOR U1050 ( .A(n905), .B(n904), .Z(n907) );
  XNOR U1051 ( .A(n906), .B(n907), .Z(n924) );
  XOR U1052 ( .A(sreg[150]), .B(n923), .Z(n903) );
  XNOR U1053 ( .A(n924), .B(n903), .Z(c[150]) );
  NANDN U1054 ( .A(n905), .B(n904), .Z(n909) );
  OR U1055 ( .A(n907), .B(n906), .Z(n908) );
  AND U1056 ( .A(n909), .B(n908), .Z(n928) );
  AND U1057 ( .A(b[3]), .B(a[24]), .Z(n916) );
  AND U1058 ( .A(b[2]), .B(a[23]), .Z(n910) );
  NAND U1059 ( .A(n916), .B(n910), .Z(n914) );
  NANDN U1060 ( .A(n912), .B(n911), .Z(n913) );
  AND U1061 ( .A(n914), .B(n913), .Z(n941) );
  NAND U1062 ( .A(a[25]), .B(b[2]), .Z(n915) );
  XNOR U1063 ( .A(n916), .B(n915), .Z(n933) );
  NAND U1064 ( .A(b[1]), .B(a[26]), .Z(n934) );
  XNOR U1065 ( .A(n933), .B(n934), .Z(n939) );
  NAND U1066 ( .A(b[0]), .B(a[27]), .Z(n940) );
  XOR U1067 ( .A(n939), .B(n940), .Z(n942) );
  XOR U1068 ( .A(n941), .B(n942), .Z(n927) );
  NANDN U1069 ( .A(n918), .B(n917), .Z(n922) );
  OR U1070 ( .A(n920), .B(n919), .Z(n921) );
  AND U1071 ( .A(n922), .B(n921), .Z(n926) );
  XOR U1072 ( .A(n927), .B(n926), .Z(n929) );
  XNOR U1073 ( .A(n928), .B(n929), .Z(n946) );
  XNOR U1074 ( .A(sreg[151]), .B(n945), .Z(n925) );
  XNOR U1075 ( .A(n946), .B(n925), .Z(c[151]) );
  NANDN U1076 ( .A(n927), .B(n926), .Z(n931) );
  OR U1077 ( .A(n929), .B(n928), .Z(n930) );
  AND U1078 ( .A(n931), .B(n930), .Z(n951) );
  AND U1079 ( .A(b[3]), .B(a[25]), .Z(n938) );
  AND U1080 ( .A(b[2]), .B(a[24]), .Z(n932) );
  NAND U1081 ( .A(n938), .B(n932), .Z(n936) );
  NANDN U1082 ( .A(n934), .B(n933), .Z(n935) );
  AND U1083 ( .A(n936), .B(n935), .Z(n963) );
  NAND U1084 ( .A(a[26]), .B(b[2]), .Z(n937) );
  XNOR U1085 ( .A(n938), .B(n937), .Z(n955) );
  NAND U1086 ( .A(b[1]), .B(a[27]), .Z(n956) );
  XNOR U1087 ( .A(n955), .B(n956), .Z(n961) );
  NAND U1088 ( .A(b[0]), .B(a[28]), .Z(n962) );
  XOR U1089 ( .A(n961), .B(n962), .Z(n964) );
  XOR U1090 ( .A(n963), .B(n964), .Z(n949) );
  NANDN U1091 ( .A(n940), .B(n939), .Z(n944) );
  OR U1092 ( .A(n942), .B(n941), .Z(n943) );
  AND U1093 ( .A(n944), .B(n943), .Z(n948) );
  XNOR U1094 ( .A(n949), .B(n948), .Z(n950) );
  XNOR U1095 ( .A(n951), .B(n950), .Z(n968) );
  XOR U1096 ( .A(n967), .B(sreg[152]), .Z(n947) );
  XNOR U1097 ( .A(n968), .B(n947), .Z(c[152]) );
  NANDN U1098 ( .A(n949), .B(n948), .Z(n953) );
  NANDN U1099 ( .A(n951), .B(n950), .Z(n952) );
  AND U1100 ( .A(n953), .B(n952), .Z(n973) );
  AND U1101 ( .A(b[3]), .B(a[26]), .Z(n960) );
  AND U1102 ( .A(b[2]), .B(a[25]), .Z(n954) );
  NAND U1103 ( .A(n960), .B(n954), .Z(n958) );
  NANDN U1104 ( .A(n956), .B(n955), .Z(n957) );
  AND U1105 ( .A(n958), .B(n957), .Z(n985) );
  NAND U1106 ( .A(a[27]), .B(b[2]), .Z(n959) );
  XNOR U1107 ( .A(n960), .B(n959), .Z(n977) );
  NAND U1108 ( .A(b[1]), .B(a[28]), .Z(n978) );
  XNOR U1109 ( .A(n977), .B(n978), .Z(n983) );
  NAND U1110 ( .A(b[0]), .B(a[29]), .Z(n984) );
  XOR U1111 ( .A(n983), .B(n984), .Z(n986) );
  XOR U1112 ( .A(n985), .B(n986), .Z(n971) );
  NANDN U1113 ( .A(n962), .B(n961), .Z(n966) );
  OR U1114 ( .A(n964), .B(n963), .Z(n965) );
  AND U1115 ( .A(n966), .B(n965), .Z(n970) );
  XNOR U1116 ( .A(n971), .B(n970), .Z(n972) );
  XNOR U1117 ( .A(n973), .B(n972), .Z(n990) );
  XNOR U1118 ( .A(n989), .B(sreg[153]), .Z(n969) );
  XNOR U1119 ( .A(n990), .B(n969), .Z(c[153]) );
  NANDN U1120 ( .A(n971), .B(n970), .Z(n975) );
  NANDN U1121 ( .A(n973), .B(n972), .Z(n974) );
  AND U1122 ( .A(n975), .B(n974), .Z(n994) );
  AND U1123 ( .A(b[3]), .B(a[27]), .Z(n982) );
  AND U1124 ( .A(b[2]), .B(a[26]), .Z(n976) );
  NAND U1125 ( .A(n982), .B(n976), .Z(n980) );
  NANDN U1126 ( .A(n978), .B(n977), .Z(n979) );
  AND U1127 ( .A(n980), .B(n979), .Z(n1007) );
  NAND U1128 ( .A(a[28]), .B(b[2]), .Z(n981) );
  XNOR U1129 ( .A(n982), .B(n981), .Z(n999) );
  NAND U1130 ( .A(b[1]), .B(a[29]), .Z(n1000) );
  XNOR U1131 ( .A(n999), .B(n1000), .Z(n1005) );
  NAND U1132 ( .A(b[0]), .B(a[30]), .Z(n1006) );
  XOR U1133 ( .A(n1005), .B(n1006), .Z(n1008) );
  XOR U1134 ( .A(n1007), .B(n1008), .Z(n993) );
  NANDN U1135 ( .A(n984), .B(n983), .Z(n988) );
  OR U1136 ( .A(n986), .B(n985), .Z(n987) );
  AND U1137 ( .A(n988), .B(n987), .Z(n992) );
  XOR U1138 ( .A(n993), .B(n992), .Z(n995) );
  XNOR U1139 ( .A(n994), .B(n995), .Z(n1012) );
  XOR U1140 ( .A(sreg[154]), .B(n1011), .Z(n991) );
  XNOR U1141 ( .A(n1012), .B(n991), .Z(c[154]) );
  NANDN U1142 ( .A(n993), .B(n992), .Z(n997) );
  OR U1143 ( .A(n995), .B(n994), .Z(n996) );
  AND U1144 ( .A(n997), .B(n996), .Z(n1016) );
  AND U1145 ( .A(b[3]), .B(a[28]), .Z(n1004) );
  AND U1146 ( .A(b[2]), .B(a[27]), .Z(n998) );
  NAND U1147 ( .A(n1004), .B(n998), .Z(n1002) );
  NANDN U1148 ( .A(n1000), .B(n999), .Z(n1001) );
  AND U1149 ( .A(n1002), .B(n1001), .Z(n1029) );
  NAND U1150 ( .A(a[29]), .B(b[2]), .Z(n1003) );
  XNOR U1151 ( .A(n1004), .B(n1003), .Z(n1021) );
  NAND U1152 ( .A(b[1]), .B(a[30]), .Z(n1022) );
  XNOR U1153 ( .A(n1021), .B(n1022), .Z(n1027) );
  NAND U1154 ( .A(b[0]), .B(a[31]), .Z(n1028) );
  XOR U1155 ( .A(n1027), .B(n1028), .Z(n1030) );
  XOR U1156 ( .A(n1029), .B(n1030), .Z(n1015) );
  NANDN U1157 ( .A(n1006), .B(n1005), .Z(n1010) );
  OR U1158 ( .A(n1008), .B(n1007), .Z(n1009) );
  AND U1159 ( .A(n1010), .B(n1009), .Z(n1014) );
  XOR U1160 ( .A(n1015), .B(n1014), .Z(n1017) );
  XNOR U1161 ( .A(n1016), .B(n1017), .Z(n1034) );
  XNOR U1162 ( .A(sreg[155]), .B(n1033), .Z(n1013) );
  XNOR U1163 ( .A(n1034), .B(n1013), .Z(c[155]) );
  NANDN U1164 ( .A(n1015), .B(n1014), .Z(n1019) );
  OR U1165 ( .A(n1017), .B(n1016), .Z(n1018) );
  AND U1166 ( .A(n1019), .B(n1018), .Z(n1039) );
  AND U1167 ( .A(b[3]), .B(a[29]), .Z(n1026) );
  AND U1168 ( .A(b[2]), .B(a[28]), .Z(n1020) );
  NAND U1169 ( .A(n1026), .B(n1020), .Z(n1024) );
  NANDN U1170 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1171 ( .A(n1024), .B(n1023), .Z(n1051) );
  NAND U1172 ( .A(a[30]), .B(b[2]), .Z(n1025) );
  XNOR U1173 ( .A(n1026), .B(n1025), .Z(n1043) );
  NAND U1174 ( .A(b[1]), .B(a[31]), .Z(n1044) );
  XNOR U1175 ( .A(n1043), .B(n1044), .Z(n1049) );
  NAND U1176 ( .A(b[0]), .B(a[32]), .Z(n1050) );
  XOR U1177 ( .A(n1049), .B(n1050), .Z(n1052) );
  XOR U1178 ( .A(n1051), .B(n1052), .Z(n1037) );
  NANDN U1179 ( .A(n1028), .B(n1027), .Z(n1032) );
  OR U1180 ( .A(n1030), .B(n1029), .Z(n1031) );
  AND U1181 ( .A(n1032), .B(n1031), .Z(n1036) );
  XNOR U1182 ( .A(n1037), .B(n1036), .Z(n1038) );
  XNOR U1183 ( .A(n1039), .B(n1038), .Z(n1056) );
  XOR U1184 ( .A(n1055), .B(sreg[156]), .Z(n1035) );
  XNOR U1185 ( .A(n1056), .B(n1035), .Z(c[156]) );
  NANDN U1186 ( .A(n1037), .B(n1036), .Z(n1041) );
  NANDN U1187 ( .A(n1039), .B(n1038), .Z(n1040) );
  AND U1188 ( .A(n1041), .B(n1040), .Z(n1060) );
  AND U1189 ( .A(b[3]), .B(a[30]), .Z(n1048) );
  AND U1190 ( .A(b[2]), .B(a[29]), .Z(n1042) );
  NAND U1191 ( .A(n1048), .B(n1042), .Z(n1046) );
  NANDN U1192 ( .A(n1044), .B(n1043), .Z(n1045) );
  AND U1193 ( .A(n1046), .B(n1045), .Z(n1073) );
  NAND U1194 ( .A(a[31]), .B(b[2]), .Z(n1047) );
  XNOR U1195 ( .A(n1048), .B(n1047), .Z(n1065) );
  NAND U1196 ( .A(b[1]), .B(a[32]), .Z(n1066) );
  XNOR U1197 ( .A(n1065), .B(n1066), .Z(n1071) );
  NAND U1198 ( .A(b[0]), .B(a[33]), .Z(n1072) );
  XOR U1199 ( .A(n1071), .B(n1072), .Z(n1074) );
  XOR U1200 ( .A(n1073), .B(n1074), .Z(n1059) );
  NANDN U1201 ( .A(n1050), .B(n1049), .Z(n1054) );
  OR U1202 ( .A(n1052), .B(n1051), .Z(n1053) );
  AND U1203 ( .A(n1054), .B(n1053), .Z(n1058) );
  XOR U1204 ( .A(n1059), .B(n1058), .Z(n1061) );
  XNOR U1205 ( .A(n1060), .B(n1061), .Z(n1078) );
  XOR U1206 ( .A(sreg[157]), .B(n1077), .Z(n1057) );
  XNOR U1207 ( .A(n1078), .B(n1057), .Z(c[157]) );
  NANDN U1208 ( .A(n1059), .B(n1058), .Z(n1063) );
  OR U1209 ( .A(n1061), .B(n1060), .Z(n1062) );
  AND U1210 ( .A(n1063), .B(n1062), .Z(n1082) );
  AND U1211 ( .A(b[3]), .B(a[31]), .Z(n1070) );
  AND U1212 ( .A(b[2]), .B(a[30]), .Z(n1064) );
  NAND U1213 ( .A(n1070), .B(n1064), .Z(n1068) );
  NANDN U1214 ( .A(n1066), .B(n1065), .Z(n1067) );
  AND U1215 ( .A(n1068), .B(n1067), .Z(n1095) );
  NAND U1216 ( .A(a[32]), .B(b[2]), .Z(n1069) );
  XNOR U1217 ( .A(n1070), .B(n1069), .Z(n1087) );
  NAND U1218 ( .A(b[1]), .B(a[33]), .Z(n1088) );
  XNOR U1219 ( .A(n1087), .B(n1088), .Z(n1093) );
  NAND U1220 ( .A(b[0]), .B(a[34]), .Z(n1094) );
  XOR U1221 ( .A(n1093), .B(n1094), .Z(n1096) );
  XOR U1222 ( .A(n1095), .B(n1096), .Z(n1081) );
  NANDN U1223 ( .A(n1072), .B(n1071), .Z(n1076) );
  OR U1224 ( .A(n1074), .B(n1073), .Z(n1075) );
  AND U1225 ( .A(n1076), .B(n1075), .Z(n1080) );
  XOR U1226 ( .A(n1081), .B(n1080), .Z(n1083) );
  XNOR U1227 ( .A(n1082), .B(n1083), .Z(n1100) );
  XNOR U1228 ( .A(sreg[158]), .B(n1099), .Z(n1079) );
  XNOR U1229 ( .A(n1100), .B(n1079), .Z(c[158]) );
  NANDN U1230 ( .A(n1081), .B(n1080), .Z(n1085) );
  OR U1231 ( .A(n1083), .B(n1082), .Z(n1084) );
  AND U1232 ( .A(n1085), .B(n1084), .Z(n1104) );
  AND U1233 ( .A(b[3]), .B(a[32]), .Z(n1092) );
  AND U1234 ( .A(b[2]), .B(a[31]), .Z(n1086) );
  NAND U1235 ( .A(n1092), .B(n1086), .Z(n1090) );
  NANDN U1236 ( .A(n1088), .B(n1087), .Z(n1089) );
  AND U1237 ( .A(n1090), .B(n1089), .Z(n1117) );
  NAND U1238 ( .A(a[33]), .B(b[2]), .Z(n1091) );
  XNOR U1239 ( .A(n1092), .B(n1091), .Z(n1109) );
  NAND U1240 ( .A(b[1]), .B(a[34]), .Z(n1110) );
  XNOR U1241 ( .A(n1109), .B(n1110), .Z(n1115) );
  NAND U1242 ( .A(b[0]), .B(a[35]), .Z(n1116) );
  XOR U1243 ( .A(n1115), .B(n1116), .Z(n1118) );
  XOR U1244 ( .A(n1117), .B(n1118), .Z(n1103) );
  NANDN U1245 ( .A(n1094), .B(n1093), .Z(n1098) );
  OR U1246 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1247 ( .A(n1098), .B(n1097), .Z(n1102) );
  XOR U1248 ( .A(n1103), .B(n1102), .Z(n1105) );
  XNOR U1249 ( .A(n1104), .B(n1105), .Z(n1122) );
  XNOR U1250 ( .A(sreg[159]), .B(n1121), .Z(n1101) );
  XNOR U1251 ( .A(n1122), .B(n1101), .Z(c[159]) );
  NANDN U1252 ( .A(n1103), .B(n1102), .Z(n1107) );
  OR U1253 ( .A(n1105), .B(n1104), .Z(n1106) );
  AND U1254 ( .A(n1107), .B(n1106), .Z(n1126) );
  AND U1255 ( .A(b[3]), .B(a[33]), .Z(n1114) );
  AND U1256 ( .A(b[2]), .B(a[32]), .Z(n1108) );
  NAND U1257 ( .A(n1114), .B(n1108), .Z(n1112) );
  NANDN U1258 ( .A(n1110), .B(n1109), .Z(n1111) );
  AND U1259 ( .A(n1112), .B(n1111), .Z(n1139) );
  NAND U1260 ( .A(a[34]), .B(b[2]), .Z(n1113) );
  XNOR U1261 ( .A(n1114), .B(n1113), .Z(n1131) );
  NAND U1262 ( .A(b[1]), .B(a[35]), .Z(n1132) );
  XNOR U1263 ( .A(n1131), .B(n1132), .Z(n1137) );
  NAND U1264 ( .A(b[0]), .B(a[36]), .Z(n1138) );
  XOR U1265 ( .A(n1137), .B(n1138), .Z(n1140) );
  XOR U1266 ( .A(n1139), .B(n1140), .Z(n1125) );
  NANDN U1267 ( .A(n1116), .B(n1115), .Z(n1120) );
  OR U1268 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U1269 ( .A(n1120), .B(n1119), .Z(n1124) );
  XOR U1270 ( .A(n1125), .B(n1124), .Z(n1127) );
  XNOR U1271 ( .A(n1126), .B(n1127), .Z(n1144) );
  XNOR U1272 ( .A(sreg[160]), .B(n1143), .Z(n1123) );
  XNOR U1273 ( .A(n1144), .B(n1123), .Z(c[160]) );
  NANDN U1274 ( .A(n1125), .B(n1124), .Z(n1129) );
  OR U1275 ( .A(n1127), .B(n1126), .Z(n1128) );
  AND U1276 ( .A(n1129), .B(n1128), .Z(n1148) );
  AND U1277 ( .A(b[3]), .B(a[34]), .Z(n1136) );
  AND U1278 ( .A(b[2]), .B(a[33]), .Z(n1130) );
  NAND U1279 ( .A(n1136), .B(n1130), .Z(n1134) );
  NANDN U1280 ( .A(n1132), .B(n1131), .Z(n1133) );
  AND U1281 ( .A(n1134), .B(n1133), .Z(n1161) );
  NAND U1282 ( .A(a[35]), .B(b[2]), .Z(n1135) );
  XNOR U1283 ( .A(n1136), .B(n1135), .Z(n1153) );
  NAND U1284 ( .A(b[1]), .B(a[36]), .Z(n1154) );
  XNOR U1285 ( .A(n1153), .B(n1154), .Z(n1159) );
  NAND U1286 ( .A(b[0]), .B(a[37]), .Z(n1160) );
  XOR U1287 ( .A(n1159), .B(n1160), .Z(n1162) );
  XOR U1288 ( .A(n1161), .B(n1162), .Z(n1147) );
  NANDN U1289 ( .A(n1138), .B(n1137), .Z(n1142) );
  OR U1290 ( .A(n1140), .B(n1139), .Z(n1141) );
  AND U1291 ( .A(n1142), .B(n1141), .Z(n1146) );
  XOR U1292 ( .A(n1147), .B(n1146), .Z(n1149) );
  XNOR U1293 ( .A(n1148), .B(n1149), .Z(n1166) );
  XNOR U1294 ( .A(sreg[161]), .B(n1165), .Z(n1145) );
  XNOR U1295 ( .A(n1166), .B(n1145), .Z(c[161]) );
  NANDN U1296 ( .A(n1147), .B(n1146), .Z(n1151) );
  OR U1297 ( .A(n1149), .B(n1148), .Z(n1150) );
  AND U1298 ( .A(n1151), .B(n1150), .Z(n1170) );
  AND U1299 ( .A(b[3]), .B(a[35]), .Z(n1158) );
  AND U1300 ( .A(b[2]), .B(a[34]), .Z(n1152) );
  NAND U1301 ( .A(n1158), .B(n1152), .Z(n1156) );
  NANDN U1302 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U1303 ( .A(n1156), .B(n1155), .Z(n1183) );
  NAND U1304 ( .A(a[36]), .B(b[2]), .Z(n1157) );
  XNOR U1305 ( .A(n1158), .B(n1157), .Z(n1175) );
  NAND U1306 ( .A(b[1]), .B(a[37]), .Z(n1176) );
  XNOR U1307 ( .A(n1175), .B(n1176), .Z(n1181) );
  NAND U1308 ( .A(b[0]), .B(a[38]), .Z(n1182) );
  XOR U1309 ( .A(n1181), .B(n1182), .Z(n1184) );
  XOR U1310 ( .A(n1183), .B(n1184), .Z(n1169) );
  NANDN U1311 ( .A(n1160), .B(n1159), .Z(n1164) );
  OR U1312 ( .A(n1162), .B(n1161), .Z(n1163) );
  AND U1313 ( .A(n1164), .B(n1163), .Z(n1168) );
  XOR U1314 ( .A(n1169), .B(n1168), .Z(n1171) );
  XNOR U1315 ( .A(n1170), .B(n1171), .Z(n1188) );
  XNOR U1316 ( .A(sreg[162]), .B(n1187), .Z(n1167) );
  XNOR U1317 ( .A(n1188), .B(n1167), .Z(c[162]) );
  NANDN U1318 ( .A(n1169), .B(n1168), .Z(n1173) );
  OR U1319 ( .A(n1171), .B(n1170), .Z(n1172) );
  AND U1320 ( .A(n1173), .B(n1172), .Z(n1193) );
  AND U1321 ( .A(b[3]), .B(a[36]), .Z(n1180) );
  AND U1322 ( .A(b[2]), .B(a[35]), .Z(n1174) );
  NAND U1323 ( .A(n1180), .B(n1174), .Z(n1178) );
  NANDN U1324 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1325 ( .A(n1178), .B(n1177), .Z(n1205) );
  NAND U1326 ( .A(a[37]), .B(b[2]), .Z(n1179) );
  XNOR U1327 ( .A(n1180), .B(n1179), .Z(n1197) );
  NAND U1328 ( .A(b[1]), .B(a[38]), .Z(n1198) );
  XNOR U1329 ( .A(n1197), .B(n1198), .Z(n1203) );
  NAND U1330 ( .A(b[0]), .B(a[39]), .Z(n1204) );
  XOR U1331 ( .A(n1203), .B(n1204), .Z(n1206) );
  XOR U1332 ( .A(n1205), .B(n1206), .Z(n1191) );
  NANDN U1333 ( .A(n1182), .B(n1181), .Z(n1186) );
  OR U1334 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U1335 ( .A(n1186), .B(n1185), .Z(n1190) );
  XNOR U1336 ( .A(n1191), .B(n1190), .Z(n1192) );
  XNOR U1337 ( .A(n1193), .B(n1192), .Z(n1210) );
  XOR U1338 ( .A(n1209), .B(sreg[163]), .Z(n1189) );
  XNOR U1339 ( .A(n1210), .B(n1189), .Z(c[163]) );
  NANDN U1340 ( .A(n1191), .B(n1190), .Z(n1195) );
  NANDN U1341 ( .A(n1193), .B(n1192), .Z(n1194) );
  AND U1342 ( .A(n1195), .B(n1194), .Z(n1214) );
  AND U1343 ( .A(b[3]), .B(a[37]), .Z(n1202) );
  AND U1344 ( .A(b[2]), .B(a[36]), .Z(n1196) );
  NAND U1345 ( .A(n1202), .B(n1196), .Z(n1200) );
  NANDN U1346 ( .A(n1198), .B(n1197), .Z(n1199) );
  AND U1347 ( .A(n1200), .B(n1199), .Z(n1227) );
  NAND U1348 ( .A(a[38]), .B(b[2]), .Z(n1201) );
  XNOR U1349 ( .A(n1202), .B(n1201), .Z(n1219) );
  NAND U1350 ( .A(b[1]), .B(a[39]), .Z(n1220) );
  XNOR U1351 ( .A(n1219), .B(n1220), .Z(n1225) );
  NAND U1352 ( .A(b[0]), .B(a[40]), .Z(n1226) );
  XOR U1353 ( .A(n1225), .B(n1226), .Z(n1228) );
  XOR U1354 ( .A(n1227), .B(n1228), .Z(n1213) );
  NANDN U1355 ( .A(n1204), .B(n1203), .Z(n1208) );
  OR U1356 ( .A(n1206), .B(n1205), .Z(n1207) );
  AND U1357 ( .A(n1208), .B(n1207), .Z(n1212) );
  XOR U1358 ( .A(n1213), .B(n1212), .Z(n1215) );
  XNOR U1359 ( .A(n1214), .B(n1215), .Z(n1232) );
  XOR U1360 ( .A(sreg[164]), .B(n1231), .Z(n1211) );
  XNOR U1361 ( .A(n1232), .B(n1211), .Z(c[164]) );
  NANDN U1362 ( .A(n1213), .B(n1212), .Z(n1217) );
  OR U1363 ( .A(n1215), .B(n1214), .Z(n1216) );
  AND U1364 ( .A(n1217), .B(n1216), .Z(n1237) );
  AND U1365 ( .A(b[3]), .B(a[38]), .Z(n1224) );
  AND U1366 ( .A(b[2]), .B(a[37]), .Z(n1218) );
  NAND U1367 ( .A(n1224), .B(n1218), .Z(n1222) );
  NANDN U1368 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U1369 ( .A(n1222), .B(n1221), .Z(n1249) );
  NAND U1370 ( .A(a[39]), .B(b[2]), .Z(n1223) );
  XNOR U1371 ( .A(n1224), .B(n1223), .Z(n1241) );
  NAND U1372 ( .A(b[1]), .B(a[40]), .Z(n1242) );
  XNOR U1373 ( .A(n1241), .B(n1242), .Z(n1247) );
  NAND U1374 ( .A(b[0]), .B(a[41]), .Z(n1248) );
  XOR U1375 ( .A(n1247), .B(n1248), .Z(n1250) );
  XOR U1376 ( .A(n1249), .B(n1250), .Z(n1235) );
  NANDN U1377 ( .A(n1226), .B(n1225), .Z(n1230) );
  OR U1378 ( .A(n1228), .B(n1227), .Z(n1229) );
  AND U1379 ( .A(n1230), .B(n1229), .Z(n1234) );
  XNOR U1380 ( .A(n1235), .B(n1234), .Z(n1236) );
  XNOR U1381 ( .A(n1237), .B(n1236), .Z(n1254) );
  XOR U1382 ( .A(n1253), .B(sreg[165]), .Z(n1233) );
  XNOR U1383 ( .A(n1254), .B(n1233), .Z(c[165]) );
  NANDN U1384 ( .A(n1235), .B(n1234), .Z(n1239) );
  NANDN U1385 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U1386 ( .A(n1239), .B(n1238), .Z(n1258) );
  AND U1387 ( .A(b[3]), .B(a[39]), .Z(n1246) );
  AND U1388 ( .A(b[2]), .B(a[38]), .Z(n1240) );
  NAND U1389 ( .A(n1246), .B(n1240), .Z(n1244) );
  NANDN U1390 ( .A(n1242), .B(n1241), .Z(n1243) );
  AND U1391 ( .A(n1244), .B(n1243), .Z(n1271) );
  NAND U1392 ( .A(a[40]), .B(b[2]), .Z(n1245) );
  XNOR U1393 ( .A(n1246), .B(n1245), .Z(n1263) );
  NAND U1394 ( .A(b[1]), .B(a[41]), .Z(n1264) );
  XNOR U1395 ( .A(n1263), .B(n1264), .Z(n1269) );
  NAND U1396 ( .A(b[0]), .B(a[42]), .Z(n1270) );
  XOR U1397 ( .A(n1269), .B(n1270), .Z(n1272) );
  XOR U1398 ( .A(n1271), .B(n1272), .Z(n1257) );
  NANDN U1399 ( .A(n1248), .B(n1247), .Z(n1252) );
  OR U1400 ( .A(n1250), .B(n1249), .Z(n1251) );
  AND U1401 ( .A(n1252), .B(n1251), .Z(n1256) );
  XOR U1402 ( .A(n1257), .B(n1256), .Z(n1259) );
  XNOR U1403 ( .A(n1258), .B(n1259), .Z(n1276) );
  XOR U1404 ( .A(sreg[166]), .B(n1275), .Z(n1255) );
  XNOR U1405 ( .A(n1276), .B(n1255), .Z(c[166]) );
  NANDN U1406 ( .A(n1257), .B(n1256), .Z(n1261) );
  OR U1407 ( .A(n1259), .B(n1258), .Z(n1260) );
  AND U1408 ( .A(n1261), .B(n1260), .Z(n1280) );
  AND U1409 ( .A(b[3]), .B(a[40]), .Z(n1268) );
  AND U1410 ( .A(b[2]), .B(a[39]), .Z(n1262) );
  NAND U1411 ( .A(n1268), .B(n1262), .Z(n1266) );
  NANDN U1412 ( .A(n1264), .B(n1263), .Z(n1265) );
  AND U1413 ( .A(n1266), .B(n1265), .Z(n1293) );
  NAND U1414 ( .A(a[41]), .B(b[2]), .Z(n1267) );
  XNOR U1415 ( .A(n1268), .B(n1267), .Z(n1285) );
  NAND U1416 ( .A(b[1]), .B(a[42]), .Z(n1286) );
  XNOR U1417 ( .A(n1285), .B(n1286), .Z(n1291) );
  NAND U1418 ( .A(b[0]), .B(a[43]), .Z(n1292) );
  XOR U1419 ( .A(n1291), .B(n1292), .Z(n1294) );
  XOR U1420 ( .A(n1293), .B(n1294), .Z(n1279) );
  NANDN U1421 ( .A(n1270), .B(n1269), .Z(n1274) );
  OR U1422 ( .A(n1272), .B(n1271), .Z(n1273) );
  AND U1423 ( .A(n1274), .B(n1273), .Z(n1278) );
  XOR U1424 ( .A(n1279), .B(n1278), .Z(n1281) );
  XNOR U1425 ( .A(n1280), .B(n1281), .Z(n1298) );
  XNOR U1426 ( .A(sreg[167]), .B(n1297), .Z(n1277) );
  XNOR U1427 ( .A(n1298), .B(n1277), .Z(c[167]) );
  NANDN U1428 ( .A(n1279), .B(n1278), .Z(n1283) );
  OR U1429 ( .A(n1281), .B(n1280), .Z(n1282) );
  AND U1430 ( .A(n1283), .B(n1282), .Z(n1302) );
  AND U1431 ( .A(b[3]), .B(a[41]), .Z(n1290) );
  AND U1432 ( .A(b[2]), .B(a[40]), .Z(n1284) );
  NAND U1433 ( .A(n1290), .B(n1284), .Z(n1288) );
  NANDN U1434 ( .A(n1286), .B(n1285), .Z(n1287) );
  AND U1435 ( .A(n1288), .B(n1287), .Z(n1315) );
  NAND U1436 ( .A(a[42]), .B(b[2]), .Z(n1289) );
  XNOR U1437 ( .A(n1290), .B(n1289), .Z(n1307) );
  NAND U1438 ( .A(b[1]), .B(a[43]), .Z(n1308) );
  XNOR U1439 ( .A(n1307), .B(n1308), .Z(n1313) );
  NAND U1440 ( .A(b[0]), .B(a[44]), .Z(n1314) );
  XOR U1441 ( .A(n1313), .B(n1314), .Z(n1316) );
  XOR U1442 ( .A(n1315), .B(n1316), .Z(n1301) );
  NANDN U1443 ( .A(n1292), .B(n1291), .Z(n1296) );
  OR U1444 ( .A(n1294), .B(n1293), .Z(n1295) );
  AND U1445 ( .A(n1296), .B(n1295), .Z(n1300) );
  XOR U1446 ( .A(n1301), .B(n1300), .Z(n1303) );
  XNOR U1447 ( .A(n1302), .B(n1303), .Z(n1320) );
  XNOR U1448 ( .A(sreg[168]), .B(n1319), .Z(n1299) );
  XNOR U1449 ( .A(n1320), .B(n1299), .Z(c[168]) );
  NANDN U1450 ( .A(n1301), .B(n1300), .Z(n1305) );
  OR U1451 ( .A(n1303), .B(n1302), .Z(n1304) );
  AND U1452 ( .A(n1305), .B(n1304), .Z(n1324) );
  AND U1453 ( .A(b[3]), .B(a[42]), .Z(n1312) );
  AND U1454 ( .A(b[2]), .B(a[41]), .Z(n1306) );
  NAND U1455 ( .A(n1312), .B(n1306), .Z(n1310) );
  NANDN U1456 ( .A(n1308), .B(n1307), .Z(n1309) );
  AND U1457 ( .A(n1310), .B(n1309), .Z(n1337) );
  NAND U1458 ( .A(a[43]), .B(b[2]), .Z(n1311) );
  XNOR U1459 ( .A(n1312), .B(n1311), .Z(n1329) );
  NAND U1460 ( .A(b[1]), .B(a[44]), .Z(n1330) );
  XNOR U1461 ( .A(n1329), .B(n1330), .Z(n1335) );
  NAND U1462 ( .A(b[0]), .B(a[45]), .Z(n1336) );
  XOR U1463 ( .A(n1335), .B(n1336), .Z(n1338) );
  XOR U1464 ( .A(n1337), .B(n1338), .Z(n1323) );
  NANDN U1465 ( .A(n1314), .B(n1313), .Z(n1318) );
  OR U1466 ( .A(n1316), .B(n1315), .Z(n1317) );
  AND U1467 ( .A(n1318), .B(n1317), .Z(n1322) );
  XOR U1468 ( .A(n1323), .B(n1322), .Z(n1325) );
  XNOR U1469 ( .A(n1324), .B(n1325), .Z(n1342) );
  XNOR U1470 ( .A(sreg[169]), .B(n1341), .Z(n1321) );
  XNOR U1471 ( .A(n1342), .B(n1321), .Z(c[169]) );
  NANDN U1472 ( .A(n1323), .B(n1322), .Z(n1327) );
  OR U1473 ( .A(n1325), .B(n1324), .Z(n1326) );
  AND U1474 ( .A(n1327), .B(n1326), .Z(n1346) );
  AND U1475 ( .A(b[3]), .B(a[43]), .Z(n1334) );
  AND U1476 ( .A(b[2]), .B(a[42]), .Z(n1328) );
  NAND U1477 ( .A(n1334), .B(n1328), .Z(n1332) );
  NANDN U1478 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U1479 ( .A(n1332), .B(n1331), .Z(n1359) );
  NAND U1480 ( .A(a[44]), .B(b[2]), .Z(n1333) );
  XNOR U1481 ( .A(n1334), .B(n1333), .Z(n1351) );
  NAND U1482 ( .A(b[1]), .B(a[45]), .Z(n1352) );
  XNOR U1483 ( .A(n1351), .B(n1352), .Z(n1357) );
  NAND U1484 ( .A(b[0]), .B(a[46]), .Z(n1358) );
  XOR U1485 ( .A(n1357), .B(n1358), .Z(n1360) );
  XOR U1486 ( .A(n1359), .B(n1360), .Z(n1345) );
  NANDN U1487 ( .A(n1336), .B(n1335), .Z(n1340) );
  OR U1488 ( .A(n1338), .B(n1337), .Z(n1339) );
  AND U1489 ( .A(n1340), .B(n1339), .Z(n1344) );
  XOR U1490 ( .A(n1345), .B(n1344), .Z(n1347) );
  XNOR U1491 ( .A(n1346), .B(n1347), .Z(n1364) );
  XNOR U1492 ( .A(sreg[170]), .B(n1363), .Z(n1343) );
  XNOR U1493 ( .A(n1364), .B(n1343), .Z(c[170]) );
  NANDN U1494 ( .A(n1345), .B(n1344), .Z(n1349) );
  OR U1495 ( .A(n1347), .B(n1346), .Z(n1348) );
  AND U1496 ( .A(n1349), .B(n1348), .Z(n1368) );
  AND U1497 ( .A(b[3]), .B(a[44]), .Z(n1356) );
  AND U1498 ( .A(b[2]), .B(a[43]), .Z(n1350) );
  NAND U1499 ( .A(n1356), .B(n1350), .Z(n1354) );
  NANDN U1500 ( .A(n1352), .B(n1351), .Z(n1353) );
  AND U1501 ( .A(n1354), .B(n1353), .Z(n1381) );
  NAND U1502 ( .A(a[45]), .B(b[2]), .Z(n1355) );
  XNOR U1503 ( .A(n1356), .B(n1355), .Z(n1373) );
  NAND U1504 ( .A(b[1]), .B(a[46]), .Z(n1374) );
  XNOR U1505 ( .A(n1373), .B(n1374), .Z(n1379) );
  NAND U1506 ( .A(b[0]), .B(a[47]), .Z(n1380) );
  XOR U1507 ( .A(n1379), .B(n1380), .Z(n1382) );
  XOR U1508 ( .A(n1381), .B(n1382), .Z(n1367) );
  NANDN U1509 ( .A(n1358), .B(n1357), .Z(n1362) );
  OR U1510 ( .A(n1360), .B(n1359), .Z(n1361) );
  AND U1511 ( .A(n1362), .B(n1361), .Z(n1366) );
  XOR U1512 ( .A(n1367), .B(n1366), .Z(n1369) );
  XNOR U1513 ( .A(n1368), .B(n1369), .Z(n1386) );
  XNOR U1514 ( .A(sreg[171]), .B(n1385), .Z(n1365) );
  XNOR U1515 ( .A(n1386), .B(n1365), .Z(c[171]) );
  NANDN U1516 ( .A(n1367), .B(n1366), .Z(n1371) );
  OR U1517 ( .A(n1369), .B(n1368), .Z(n1370) );
  AND U1518 ( .A(n1371), .B(n1370), .Z(n1390) );
  AND U1519 ( .A(b[3]), .B(a[45]), .Z(n1378) );
  AND U1520 ( .A(b[2]), .B(a[44]), .Z(n1372) );
  NAND U1521 ( .A(n1378), .B(n1372), .Z(n1376) );
  NANDN U1522 ( .A(n1374), .B(n1373), .Z(n1375) );
  AND U1523 ( .A(n1376), .B(n1375), .Z(n1403) );
  NAND U1524 ( .A(a[46]), .B(b[2]), .Z(n1377) );
  XNOR U1525 ( .A(n1378), .B(n1377), .Z(n1395) );
  NAND U1526 ( .A(b[1]), .B(a[47]), .Z(n1396) );
  XNOR U1527 ( .A(n1395), .B(n1396), .Z(n1401) );
  NAND U1528 ( .A(b[0]), .B(a[48]), .Z(n1402) );
  XOR U1529 ( .A(n1401), .B(n1402), .Z(n1404) );
  XOR U1530 ( .A(n1403), .B(n1404), .Z(n1389) );
  NANDN U1531 ( .A(n1380), .B(n1379), .Z(n1384) );
  OR U1532 ( .A(n1382), .B(n1381), .Z(n1383) );
  AND U1533 ( .A(n1384), .B(n1383), .Z(n1388) );
  XOR U1534 ( .A(n1389), .B(n1388), .Z(n1391) );
  XNOR U1535 ( .A(n1390), .B(n1391), .Z(n1408) );
  XNOR U1536 ( .A(sreg[172]), .B(n1407), .Z(n1387) );
  XNOR U1537 ( .A(n1408), .B(n1387), .Z(c[172]) );
  NANDN U1538 ( .A(n1389), .B(n1388), .Z(n1393) );
  OR U1539 ( .A(n1391), .B(n1390), .Z(n1392) );
  AND U1540 ( .A(n1393), .B(n1392), .Z(n1412) );
  AND U1541 ( .A(b[3]), .B(a[46]), .Z(n1400) );
  AND U1542 ( .A(b[2]), .B(a[45]), .Z(n1394) );
  NAND U1543 ( .A(n1400), .B(n1394), .Z(n1398) );
  NANDN U1544 ( .A(n1396), .B(n1395), .Z(n1397) );
  AND U1545 ( .A(n1398), .B(n1397), .Z(n1425) );
  NAND U1546 ( .A(a[47]), .B(b[2]), .Z(n1399) );
  XNOR U1547 ( .A(n1400), .B(n1399), .Z(n1417) );
  NAND U1548 ( .A(b[1]), .B(a[48]), .Z(n1418) );
  XNOR U1549 ( .A(n1417), .B(n1418), .Z(n1423) );
  NAND U1550 ( .A(b[0]), .B(a[49]), .Z(n1424) );
  XOR U1551 ( .A(n1423), .B(n1424), .Z(n1426) );
  XOR U1552 ( .A(n1425), .B(n1426), .Z(n1411) );
  NANDN U1553 ( .A(n1402), .B(n1401), .Z(n1406) );
  OR U1554 ( .A(n1404), .B(n1403), .Z(n1405) );
  AND U1555 ( .A(n1406), .B(n1405), .Z(n1410) );
  XOR U1556 ( .A(n1411), .B(n1410), .Z(n1413) );
  XNOR U1557 ( .A(n1412), .B(n1413), .Z(n1430) );
  XNOR U1558 ( .A(sreg[173]), .B(n1429), .Z(n1409) );
  XNOR U1559 ( .A(n1430), .B(n1409), .Z(c[173]) );
  NANDN U1560 ( .A(n1411), .B(n1410), .Z(n1415) );
  OR U1561 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U1562 ( .A(n1415), .B(n1414), .Z(n1435) );
  AND U1563 ( .A(b[3]), .B(a[47]), .Z(n1422) );
  AND U1564 ( .A(b[2]), .B(a[46]), .Z(n1416) );
  NAND U1565 ( .A(n1422), .B(n1416), .Z(n1420) );
  NANDN U1566 ( .A(n1418), .B(n1417), .Z(n1419) );
  AND U1567 ( .A(n1420), .B(n1419), .Z(n1447) );
  NAND U1568 ( .A(a[48]), .B(b[2]), .Z(n1421) );
  XNOR U1569 ( .A(n1422), .B(n1421), .Z(n1439) );
  NAND U1570 ( .A(b[1]), .B(a[49]), .Z(n1440) );
  XNOR U1571 ( .A(n1439), .B(n1440), .Z(n1445) );
  NAND U1572 ( .A(b[0]), .B(a[50]), .Z(n1446) );
  XOR U1573 ( .A(n1445), .B(n1446), .Z(n1448) );
  XOR U1574 ( .A(n1447), .B(n1448), .Z(n1433) );
  NANDN U1575 ( .A(n1424), .B(n1423), .Z(n1428) );
  OR U1576 ( .A(n1426), .B(n1425), .Z(n1427) );
  AND U1577 ( .A(n1428), .B(n1427), .Z(n1432) );
  XNOR U1578 ( .A(n1433), .B(n1432), .Z(n1434) );
  XNOR U1579 ( .A(n1435), .B(n1434), .Z(n1452) );
  XOR U1580 ( .A(n1451), .B(sreg[174]), .Z(n1431) );
  XNOR U1581 ( .A(n1452), .B(n1431), .Z(c[174]) );
  NANDN U1582 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U1583 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U1584 ( .A(n1437), .B(n1436), .Z(n1456) );
  AND U1585 ( .A(b[3]), .B(a[48]), .Z(n1444) );
  AND U1586 ( .A(b[2]), .B(a[47]), .Z(n1438) );
  NAND U1587 ( .A(n1444), .B(n1438), .Z(n1442) );
  NANDN U1588 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1589 ( .A(n1442), .B(n1441), .Z(n1469) );
  NAND U1590 ( .A(a[49]), .B(b[2]), .Z(n1443) );
  XNOR U1591 ( .A(n1444), .B(n1443), .Z(n1461) );
  NAND U1592 ( .A(b[1]), .B(a[50]), .Z(n1462) );
  XNOR U1593 ( .A(n1461), .B(n1462), .Z(n1467) );
  NAND U1594 ( .A(b[0]), .B(a[51]), .Z(n1468) );
  XOR U1595 ( .A(n1467), .B(n1468), .Z(n1470) );
  XOR U1596 ( .A(n1469), .B(n1470), .Z(n1455) );
  NANDN U1597 ( .A(n1446), .B(n1445), .Z(n1450) );
  OR U1598 ( .A(n1448), .B(n1447), .Z(n1449) );
  AND U1599 ( .A(n1450), .B(n1449), .Z(n1454) );
  XOR U1600 ( .A(n1455), .B(n1454), .Z(n1457) );
  XNOR U1601 ( .A(n1456), .B(n1457), .Z(n1474) );
  XOR U1602 ( .A(sreg[175]), .B(n1473), .Z(n1453) );
  XNOR U1603 ( .A(n1474), .B(n1453), .Z(c[175]) );
  NANDN U1604 ( .A(n1455), .B(n1454), .Z(n1459) );
  OR U1605 ( .A(n1457), .B(n1456), .Z(n1458) );
  AND U1606 ( .A(n1459), .B(n1458), .Z(n1478) );
  AND U1607 ( .A(b[3]), .B(a[49]), .Z(n1466) );
  AND U1608 ( .A(b[2]), .B(a[48]), .Z(n1460) );
  NAND U1609 ( .A(n1466), .B(n1460), .Z(n1464) );
  NANDN U1610 ( .A(n1462), .B(n1461), .Z(n1463) );
  AND U1611 ( .A(n1464), .B(n1463), .Z(n1491) );
  NAND U1612 ( .A(a[50]), .B(b[2]), .Z(n1465) );
  XNOR U1613 ( .A(n1466), .B(n1465), .Z(n1483) );
  NAND U1614 ( .A(b[1]), .B(a[51]), .Z(n1484) );
  XNOR U1615 ( .A(n1483), .B(n1484), .Z(n1489) );
  NAND U1616 ( .A(b[0]), .B(a[52]), .Z(n1490) );
  XOR U1617 ( .A(n1489), .B(n1490), .Z(n1492) );
  XOR U1618 ( .A(n1491), .B(n1492), .Z(n1477) );
  NANDN U1619 ( .A(n1468), .B(n1467), .Z(n1472) );
  OR U1620 ( .A(n1470), .B(n1469), .Z(n1471) );
  AND U1621 ( .A(n1472), .B(n1471), .Z(n1476) );
  XOR U1622 ( .A(n1477), .B(n1476), .Z(n1479) );
  XNOR U1623 ( .A(n1478), .B(n1479), .Z(n1496) );
  XNOR U1624 ( .A(sreg[176]), .B(n1495), .Z(n1475) );
  XNOR U1625 ( .A(n1496), .B(n1475), .Z(c[176]) );
  NANDN U1626 ( .A(n1477), .B(n1476), .Z(n1481) );
  OR U1627 ( .A(n1479), .B(n1478), .Z(n1480) );
  AND U1628 ( .A(n1481), .B(n1480), .Z(n1500) );
  AND U1629 ( .A(b[3]), .B(a[50]), .Z(n1488) );
  AND U1630 ( .A(b[2]), .B(a[49]), .Z(n1482) );
  NAND U1631 ( .A(n1488), .B(n1482), .Z(n1486) );
  NANDN U1632 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1633 ( .A(n1486), .B(n1485), .Z(n1513) );
  NAND U1634 ( .A(a[51]), .B(b[2]), .Z(n1487) );
  XNOR U1635 ( .A(n1488), .B(n1487), .Z(n1505) );
  NAND U1636 ( .A(b[1]), .B(a[52]), .Z(n1506) );
  XNOR U1637 ( .A(n1505), .B(n1506), .Z(n1511) );
  NAND U1638 ( .A(b[0]), .B(a[53]), .Z(n1512) );
  XOR U1639 ( .A(n1511), .B(n1512), .Z(n1514) );
  XOR U1640 ( .A(n1513), .B(n1514), .Z(n1499) );
  NANDN U1641 ( .A(n1490), .B(n1489), .Z(n1494) );
  OR U1642 ( .A(n1492), .B(n1491), .Z(n1493) );
  AND U1643 ( .A(n1494), .B(n1493), .Z(n1498) );
  XOR U1644 ( .A(n1499), .B(n1498), .Z(n1501) );
  XNOR U1645 ( .A(n1500), .B(n1501), .Z(n1518) );
  XNOR U1646 ( .A(sreg[177]), .B(n1517), .Z(n1497) );
  XNOR U1647 ( .A(n1518), .B(n1497), .Z(c[177]) );
  NANDN U1648 ( .A(n1499), .B(n1498), .Z(n1503) );
  OR U1649 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U1650 ( .A(n1503), .B(n1502), .Z(n1522) );
  AND U1651 ( .A(b[3]), .B(a[51]), .Z(n1510) );
  AND U1652 ( .A(b[2]), .B(a[50]), .Z(n1504) );
  NAND U1653 ( .A(n1510), .B(n1504), .Z(n1508) );
  NANDN U1654 ( .A(n1506), .B(n1505), .Z(n1507) );
  AND U1655 ( .A(n1508), .B(n1507), .Z(n1535) );
  NAND U1656 ( .A(a[52]), .B(b[2]), .Z(n1509) );
  XNOR U1657 ( .A(n1510), .B(n1509), .Z(n1527) );
  NAND U1658 ( .A(b[1]), .B(a[53]), .Z(n1528) );
  XNOR U1659 ( .A(n1527), .B(n1528), .Z(n1533) );
  NAND U1660 ( .A(b[0]), .B(a[54]), .Z(n1534) );
  XOR U1661 ( .A(n1533), .B(n1534), .Z(n1536) );
  XOR U1662 ( .A(n1535), .B(n1536), .Z(n1521) );
  NANDN U1663 ( .A(n1512), .B(n1511), .Z(n1516) );
  OR U1664 ( .A(n1514), .B(n1513), .Z(n1515) );
  AND U1665 ( .A(n1516), .B(n1515), .Z(n1520) );
  XOR U1666 ( .A(n1521), .B(n1520), .Z(n1523) );
  XNOR U1667 ( .A(n1522), .B(n1523), .Z(n1540) );
  XNOR U1668 ( .A(sreg[178]), .B(n1539), .Z(n1519) );
  XNOR U1669 ( .A(n1540), .B(n1519), .Z(c[178]) );
  NANDN U1670 ( .A(n1521), .B(n1520), .Z(n1525) );
  OR U1671 ( .A(n1523), .B(n1522), .Z(n1524) );
  AND U1672 ( .A(n1525), .B(n1524), .Z(n1545) );
  AND U1673 ( .A(b[3]), .B(a[52]), .Z(n1532) );
  AND U1674 ( .A(b[2]), .B(a[51]), .Z(n1526) );
  NAND U1675 ( .A(n1532), .B(n1526), .Z(n1530) );
  NANDN U1676 ( .A(n1528), .B(n1527), .Z(n1529) );
  AND U1677 ( .A(n1530), .B(n1529), .Z(n1557) );
  NAND U1678 ( .A(a[53]), .B(b[2]), .Z(n1531) );
  XNOR U1679 ( .A(n1532), .B(n1531), .Z(n1549) );
  NAND U1680 ( .A(b[1]), .B(a[54]), .Z(n1550) );
  XNOR U1681 ( .A(n1549), .B(n1550), .Z(n1555) );
  NAND U1682 ( .A(b[0]), .B(a[55]), .Z(n1556) );
  XOR U1683 ( .A(n1555), .B(n1556), .Z(n1558) );
  XOR U1684 ( .A(n1557), .B(n1558), .Z(n1543) );
  NANDN U1685 ( .A(n1534), .B(n1533), .Z(n1538) );
  OR U1686 ( .A(n1536), .B(n1535), .Z(n1537) );
  AND U1687 ( .A(n1538), .B(n1537), .Z(n1542) );
  XNOR U1688 ( .A(n1543), .B(n1542), .Z(n1544) );
  XNOR U1689 ( .A(n1545), .B(n1544), .Z(n1562) );
  XOR U1690 ( .A(n1561), .B(sreg[179]), .Z(n1541) );
  XNOR U1691 ( .A(n1562), .B(n1541), .Z(c[179]) );
  NANDN U1692 ( .A(n1543), .B(n1542), .Z(n1547) );
  NANDN U1693 ( .A(n1545), .B(n1544), .Z(n1546) );
  AND U1694 ( .A(n1547), .B(n1546), .Z(n1566) );
  AND U1695 ( .A(b[3]), .B(a[53]), .Z(n1554) );
  AND U1696 ( .A(b[2]), .B(a[52]), .Z(n1548) );
  NAND U1697 ( .A(n1554), .B(n1548), .Z(n1552) );
  NANDN U1698 ( .A(n1550), .B(n1549), .Z(n1551) );
  AND U1699 ( .A(n1552), .B(n1551), .Z(n1579) );
  NAND U1700 ( .A(a[54]), .B(b[2]), .Z(n1553) );
  XNOR U1701 ( .A(n1554), .B(n1553), .Z(n1571) );
  NAND U1702 ( .A(b[1]), .B(a[55]), .Z(n1572) );
  XNOR U1703 ( .A(n1571), .B(n1572), .Z(n1577) );
  NAND U1704 ( .A(b[0]), .B(a[56]), .Z(n1578) );
  XOR U1705 ( .A(n1577), .B(n1578), .Z(n1580) );
  XOR U1706 ( .A(n1579), .B(n1580), .Z(n1565) );
  NANDN U1707 ( .A(n1556), .B(n1555), .Z(n1560) );
  OR U1708 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U1709 ( .A(n1560), .B(n1559), .Z(n1564) );
  XOR U1710 ( .A(n1565), .B(n1564), .Z(n1567) );
  XNOR U1711 ( .A(n1566), .B(n1567), .Z(n1584) );
  XOR U1712 ( .A(sreg[180]), .B(n1583), .Z(n1563) );
  XNOR U1713 ( .A(n1584), .B(n1563), .Z(c[180]) );
  NANDN U1714 ( .A(n1565), .B(n1564), .Z(n1569) );
  OR U1715 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U1716 ( .A(n1569), .B(n1568), .Z(n1588) );
  AND U1717 ( .A(b[3]), .B(a[54]), .Z(n1576) );
  AND U1718 ( .A(b[2]), .B(a[53]), .Z(n1570) );
  NAND U1719 ( .A(n1576), .B(n1570), .Z(n1574) );
  NANDN U1720 ( .A(n1572), .B(n1571), .Z(n1573) );
  AND U1721 ( .A(n1574), .B(n1573), .Z(n1601) );
  NAND U1722 ( .A(a[55]), .B(b[2]), .Z(n1575) );
  XNOR U1723 ( .A(n1576), .B(n1575), .Z(n1593) );
  NAND U1724 ( .A(b[1]), .B(a[56]), .Z(n1594) );
  XNOR U1725 ( .A(n1593), .B(n1594), .Z(n1599) );
  NAND U1726 ( .A(b[0]), .B(a[57]), .Z(n1600) );
  XOR U1727 ( .A(n1599), .B(n1600), .Z(n1602) );
  XOR U1728 ( .A(n1601), .B(n1602), .Z(n1587) );
  NANDN U1729 ( .A(n1578), .B(n1577), .Z(n1582) );
  OR U1730 ( .A(n1580), .B(n1579), .Z(n1581) );
  AND U1731 ( .A(n1582), .B(n1581), .Z(n1586) );
  XOR U1732 ( .A(n1587), .B(n1586), .Z(n1589) );
  XNOR U1733 ( .A(n1588), .B(n1589), .Z(n1606) );
  XNOR U1734 ( .A(sreg[181]), .B(n1605), .Z(n1585) );
  XNOR U1735 ( .A(n1606), .B(n1585), .Z(c[181]) );
  NANDN U1736 ( .A(n1587), .B(n1586), .Z(n1591) );
  OR U1737 ( .A(n1589), .B(n1588), .Z(n1590) );
  AND U1738 ( .A(n1591), .B(n1590), .Z(n1610) );
  AND U1739 ( .A(b[3]), .B(a[55]), .Z(n1598) );
  AND U1740 ( .A(b[2]), .B(a[54]), .Z(n1592) );
  NAND U1741 ( .A(n1598), .B(n1592), .Z(n1596) );
  NANDN U1742 ( .A(n1594), .B(n1593), .Z(n1595) );
  AND U1743 ( .A(n1596), .B(n1595), .Z(n1623) );
  NAND U1744 ( .A(a[56]), .B(b[2]), .Z(n1597) );
  XNOR U1745 ( .A(n1598), .B(n1597), .Z(n1615) );
  NAND U1746 ( .A(b[1]), .B(a[57]), .Z(n1616) );
  XNOR U1747 ( .A(n1615), .B(n1616), .Z(n1621) );
  NAND U1748 ( .A(b[0]), .B(a[58]), .Z(n1622) );
  XOR U1749 ( .A(n1621), .B(n1622), .Z(n1624) );
  XOR U1750 ( .A(n1623), .B(n1624), .Z(n1609) );
  NANDN U1751 ( .A(n1600), .B(n1599), .Z(n1604) );
  OR U1752 ( .A(n1602), .B(n1601), .Z(n1603) );
  AND U1753 ( .A(n1604), .B(n1603), .Z(n1608) );
  XOR U1754 ( .A(n1609), .B(n1608), .Z(n1611) );
  XNOR U1755 ( .A(n1610), .B(n1611), .Z(n1628) );
  XNOR U1756 ( .A(sreg[182]), .B(n1627), .Z(n1607) );
  XNOR U1757 ( .A(n1628), .B(n1607), .Z(c[182]) );
  NANDN U1758 ( .A(n1609), .B(n1608), .Z(n1613) );
  OR U1759 ( .A(n1611), .B(n1610), .Z(n1612) );
  AND U1760 ( .A(n1613), .B(n1612), .Z(n1632) );
  AND U1761 ( .A(b[3]), .B(a[56]), .Z(n1620) );
  AND U1762 ( .A(b[2]), .B(a[55]), .Z(n1614) );
  NAND U1763 ( .A(n1620), .B(n1614), .Z(n1618) );
  NANDN U1764 ( .A(n1616), .B(n1615), .Z(n1617) );
  AND U1765 ( .A(n1618), .B(n1617), .Z(n1645) );
  NAND U1766 ( .A(a[57]), .B(b[2]), .Z(n1619) );
  XNOR U1767 ( .A(n1620), .B(n1619), .Z(n1637) );
  NAND U1768 ( .A(b[1]), .B(a[58]), .Z(n1638) );
  XNOR U1769 ( .A(n1637), .B(n1638), .Z(n1643) );
  NAND U1770 ( .A(b[0]), .B(a[59]), .Z(n1644) );
  XOR U1771 ( .A(n1643), .B(n1644), .Z(n1646) );
  XOR U1772 ( .A(n1645), .B(n1646), .Z(n1631) );
  NANDN U1773 ( .A(n1622), .B(n1621), .Z(n1626) );
  OR U1774 ( .A(n1624), .B(n1623), .Z(n1625) );
  AND U1775 ( .A(n1626), .B(n1625), .Z(n1630) );
  XOR U1776 ( .A(n1631), .B(n1630), .Z(n1633) );
  XNOR U1777 ( .A(n1632), .B(n1633), .Z(n1650) );
  XNOR U1778 ( .A(sreg[183]), .B(n1649), .Z(n1629) );
  XNOR U1779 ( .A(n1650), .B(n1629), .Z(c[183]) );
  NANDN U1780 ( .A(n1631), .B(n1630), .Z(n1635) );
  OR U1781 ( .A(n1633), .B(n1632), .Z(n1634) );
  AND U1782 ( .A(n1635), .B(n1634), .Z(n1654) );
  AND U1783 ( .A(b[3]), .B(a[57]), .Z(n1642) );
  AND U1784 ( .A(b[2]), .B(a[56]), .Z(n1636) );
  NAND U1785 ( .A(n1642), .B(n1636), .Z(n1640) );
  NANDN U1786 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U1787 ( .A(n1640), .B(n1639), .Z(n1667) );
  NAND U1788 ( .A(a[58]), .B(b[2]), .Z(n1641) );
  XNOR U1789 ( .A(n1642), .B(n1641), .Z(n1659) );
  NAND U1790 ( .A(b[1]), .B(a[59]), .Z(n1660) );
  XNOR U1791 ( .A(n1659), .B(n1660), .Z(n1665) );
  NAND U1792 ( .A(b[0]), .B(a[60]), .Z(n1666) );
  XOR U1793 ( .A(n1665), .B(n1666), .Z(n1668) );
  XOR U1794 ( .A(n1667), .B(n1668), .Z(n1653) );
  NANDN U1795 ( .A(n1644), .B(n1643), .Z(n1648) );
  OR U1796 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U1797 ( .A(n1648), .B(n1647), .Z(n1652) );
  XOR U1798 ( .A(n1653), .B(n1652), .Z(n1655) );
  XNOR U1799 ( .A(n1654), .B(n1655), .Z(n1672) );
  XNOR U1800 ( .A(sreg[184]), .B(n1671), .Z(n1651) );
  XNOR U1801 ( .A(n1672), .B(n1651), .Z(c[184]) );
  NANDN U1802 ( .A(n1653), .B(n1652), .Z(n1657) );
  OR U1803 ( .A(n1655), .B(n1654), .Z(n1656) );
  AND U1804 ( .A(n1657), .B(n1656), .Z(n1676) );
  AND U1805 ( .A(b[3]), .B(a[58]), .Z(n1664) );
  AND U1806 ( .A(b[2]), .B(a[57]), .Z(n1658) );
  NAND U1807 ( .A(n1664), .B(n1658), .Z(n1662) );
  NANDN U1808 ( .A(n1660), .B(n1659), .Z(n1661) );
  AND U1809 ( .A(n1662), .B(n1661), .Z(n1689) );
  NAND U1810 ( .A(a[59]), .B(b[2]), .Z(n1663) );
  XNOR U1811 ( .A(n1664), .B(n1663), .Z(n1681) );
  NAND U1812 ( .A(b[1]), .B(a[60]), .Z(n1682) );
  XNOR U1813 ( .A(n1681), .B(n1682), .Z(n1687) );
  NAND U1814 ( .A(b[0]), .B(a[61]), .Z(n1688) );
  XOR U1815 ( .A(n1687), .B(n1688), .Z(n1690) );
  XOR U1816 ( .A(n1689), .B(n1690), .Z(n1675) );
  NANDN U1817 ( .A(n1666), .B(n1665), .Z(n1670) );
  OR U1818 ( .A(n1668), .B(n1667), .Z(n1669) );
  AND U1819 ( .A(n1670), .B(n1669), .Z(n1674) );
  XOR U1820 ( .A(n1675), .B(n1674), .Z(n1677) );
  XNOR U1821 ( .A(n1676), .B(n1677), .Z(n1694) );
  XNOR U1822 ( .A(sreg[185]), .B(n1693), .Z(n1673) );
  XNOR U1823 ( .A(n1694), .B(n1673), .Z(c[185]) );
  NANDN U1824 ( .A(n1675), .B(n1674), .Z(n1679) );
  OR U1825 ( .A(n1677), .B(n1676), .Z(n1678) );
  AND U1826 ( .A(n1679), .B(n1678), .Z(n1698) );
  AND U1827 ( .A(b[3]), .B(a[59]), .Z(n1686) );
  AND U1828 ( .A(b[2]), .B(a[58]), .Z(n1680) );
  NAND U1829 ( .A(n1686), .B(n1680), .Z(n1684) );
  NANDN U1830 ( .A(n1682), .B(n1681), .Z(n1683) );
  AND U1831 ( .A(n1684), .B(n1683), .Z(n1711) );
  NAND U1832 ( .A(a[60]), .B(b[2]), .Z(n1685) );
  XNOR U1833 ( .A(n1686), .B(n1685), .Z(n1703) );
  NAND U1834 ( .A(b[1]), .B(a[61]), .Z(n1704) );
  XNOR U1835 ( .A(n1703), .B(n1704), .Z(n1709) );
  NAND U1836 ( .A(b[0]), .B(a[62]), .Z(n1710) );
  XOR U1837 ( .A(n1709), .B(n1710), .Z(n1712) );
  XOR U1838 ( .A(n1711), .B(n1712), .Z(n1697) );
  NANDN U1839 ( .A(n1688), .B(n1687), .Z(n1692) );
  OR U1840 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U1841 ( .A(n1692), .B(n1691), .Z(n1696) );
  XOR U1842 ( .A(n1697), .B(n1696), .Z(n1699) );
  XNOR U1843 ( .A(n1698), .B(n1699), .Z(n1716) );
  XNOR U1844 ( .A(sreg[186]), .B(n1715), .Z(n1695) );
  XNOR U1845 ( .A(n1716), .B(n1695), .Z(c[186]) );
  NANDN U1846 ( .A(n1697), .B(n1696), .Z(n1701) );
  OR U1847 ( .A(n1699), .B(n1698), .Z(n1700) );
  AND U1848 ( .A(n1701), .B(n1700), .Z(n1720) );
  AND U1849 ( .A(b[3]), .B(a[60]), .Z(n1708) );
  AND U1850 ( .A(b[2]), .B(a[59]), .Z(n1702) );
  NAND U1851 ( .A(n1708), .B(n1702), .Z(n1706) );
  NANDN U1852 ( .A(n1704), .B(n1703), .Z(n1705) );
  AND U1853 ( .A(n1706), .B(n1705), .Z(n1733) );
  NAND U1854 ( .A(a[61]), .B(b[2]), .Z(n1707) );
  XNOR U1855 ( .A(n1708), .B(n1707), .Z(n1725) );
  NAND U1856 ( .A(b[1]), .B(a[62]), .Z(n1726) );
  XNOR U1857 ( .A(n1725), .B(n1726), .Z(n1731) );
  NAND U1858 ( .A(b[0]), .B(a[63]), .Z(n1732) );
  XOR U1859 ( .A(n1731), .B(n1732), .Z(n1734) );
  XOR U1860 ( .A(n1733), .B(n1734), .Z(n1719) );
  NANDN U1861 ( .A(n1710), .B(n1709), .Z(n1714) );
  OR U1862 ( .A(n1712), .B(n1711), .Z(n1713) );
  AND U1863 ( .A(n1714), .B(n1713), .Z(n1718) );
  XOR U1864 ( .A(n1719), .B(n1718), .Z(n1721) );
  XNOR U1865 ( .A(n1720), .B(n1721), .Z(n1738) );
  XNOR U1866 ( .A(sreg[187]), .B(n1737), .Z(n1717) );
  XNOR U1867 ( .A(n1738), .B(n1717), .Z(c[187]) );
  NANDN U1868 ( .A(n1719), .B(n1718), .Z(n1723) );
  OR U1869 ( .A(n1721), .B(n1720), .Z(n1722) );
  AND U1870 ( .A(n1723), .B(n1722), .Z(n1742) );
  AND U1871 ( .A(b[3]), .B(a[61]), .Z(n1730) );
  AND U1872 ( .A(b[2]), .B(a[60]), .Z(n1724) );
  NAND U1873 ( .A(n1730), .B(n1724), .Z(n1728) );
  NANDN U1874 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U1875 ( .A(n1728), .B(n1727), .Z(n1755) );
  NAND U1876 ( .A(a[62]), .B(b[2]), .Z(n1729) );
  XNOR U1877 ( .A(n1730), .B(n1729), .Z(n1747) );
  NAND U1878 ( .A(b[1]), .B(a[63]), .Z(n1748) );
  XNOR U1879 ( .A(n1747), .B(n1748), .Z(n1753) );
  NAND U1880 ( .A(b[0]), .B(a[64]), .Z(n1754) );
  XOR U1881 ( .A(n1753), .B(n1754), .Z(n1756) );
  XOR U1882 ( .A(n1755), .B(n1756), .Z(n1741) );
  NANDN U1883 ( .A(n1732), .B(n1731), .Z(n1736) );
  OR U1884 ( .A(n1734), .B(n1733), .Z(n1735) );
  AND U1885 ( .A(n1736), .B(n1735), .Z(n1740) );
  XOR U1886 ( .A(n1741), .B(n1740), .Z(n1743) );
  XNOR U1887 ( .A(n1742), .B(n1743), .Z(n1760) );
  XNOR U1888 ( .A(sreg[188]), .B(n1759), .Z(n1739) );
  XNOR U1889 ( .A(n1760), .B(n1739), .Z(c[188]) );
  NANDN U1890 ( .A(n1741), .B(n1740), .Z(n1745) );
  OR U1891 ( .A(n1743), .B(n1742), .Z(n1744) );
  AND U1892 ( .A(n1745), .B(n1744), .Z(n1764) );
  AND U1893 ( .A(b[3]), .B(a[62]), .Z(n1752) );
  AND U1894 ( .A(b[2]), .B(a[61]), .Z(n1746) );
  NAND U1895 ( .A(n1752), .B(n1746), .Z(n1750) );
  NANDN U1896 ( .A(n1748), .B(n1747), .Z(n1749) );
  AND U1897 ( .A(n1750), .B(n1749), .Z(n1777) );
  NAND U1898 ( .A(a[63]), .B(b[2]), .Z(n1751) );
  XNOR U1899 ( .A(n1752), .B(n1751), .Z(n1769) );
  NAND U1900 ( .A(b[1]), .B(a[64]), .Z(n1770) );
  XNOR U1901 ( .A(n1769), .B(n1770), .Z(n1775) );
  NAND U1902 ( .A(b[0]), .B(a[65]), .Z(n1776) );
  XOR U1903 ( .A(n1775), .B(n1776), .Z(n1778) );
  XOR U1904 ( .A(n1777), .B(n1778), .Z(n1763) );
  NANDN U1905 ( .A(n1754), .B(n1753), .Z(n1758) );
  OR U1906 ( .A(n1756), .B(n1755), .Z(n1757) );
  AND U1907 ( .A(n1758), .B(n1757), .Z(n1762) );
  XOR U1908 ( .A(n1763), .B(n1762), .Z(n1765) );
  XNOR U1909 ( .A(n1764), .B(n1765), .Z(n1782) );
  XNOR U1910 ( .A(sreg[189]), .B(n1781), .Z(n1761) );
  XNOR U1911 ( .A(n1782), .B(n1761), .Z(c[189]) );
  NANDN U1912 ( .A(n1763), .B(n1762), .Z(n1767) );
  OR U1913 ( .A(n1765), .B(n1764), .Z(n1766) );
  AND U1914 ( .A(n1767), .B(n1766), .Z(n1787) );
  AND U1915 ( .A(b[3]), .B(a[63]), .Z(n1774) );
  AND U1916 ( .A(b[2]), .B(a[62]), .Z(n1768) );
  NAND U1917 ( .A(n1774), .B(n1768), .Z(n1772) );
  NANDN U1918 ( .A(n1770), .B(n1769), .Z(n1771) );
  AND U1919 ( .A(n1772), .B(n1771), .Z(n1799) );
  NAND U1920 ( .A(a[64]), .B(b[2]), .Z(n1773) );
  XNOR U1921 ( .A(n1774), .B(n1773), .Z(n1791) );
  NAND U1922 ( .A(b[1]), .B(a[65]), .Z(n1792) );
  XNOR U1923 ( .A(n1791), .B(n1792), .Z(n1797) );
  NAND U1924 ( .A(b[0]), .B(a[66]), .Z(n1798) );
  XOR U1925 ( .A(n1797), .B(n1798), .Z(n1800) );
  XOR U1926 ( .A(n1799), .B(n1800), .Z(n1785) );
  NANDN U1927 ( .A(n1776), .B(n1775), .Z(n1780) );
  OR U1928 ( .A(n1778), .B(n1777), .Z(n1779) );
  AND U1929 ( .A(n1780), .B(n1779), .Z(n1784) );
  XNOR U1930 ( .A(n1785), .B(n1784), .Z(n1786) );
  XNOR U1931 ( .A(n1787), .B(n1786), .Z(n1804) );
  XOR U1932 ( .A(n1803), .B(sreg[190]), .Z(n1783) );
  XNOR U1933 ( .A(n1804), .B(n1783), .Z(c[190]) );
  NANDN U1934 ( .A(n1785), .B(n1784), .Z(n1789) );
  NANDN U1935 ( .A(n1787), .B(n1786), .Z(n1788) );
  AND U1936 ( .A(n1789), .B(n1788), .Z(n1809) );
  AND U1937 ( .A(b[3]), .B(a[64]), .Z(n1796) );
  AND U1938 ( .A(b[2]), .B(a[63]), .Z(n1790) );
  NAND U1939 ( .A(n1796), .B(n1790), .Z(n1794) );
  NANDN U1940 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U1941 ( .A(n1794), .B(n1793), .Z(n1821) );
  NAND U1942 ( .A(a[65]), .B(b[2]), .Z(n1795) );
  XNOR U1943 ( .A(n1796), .B(n1795), .Z(n1813) );
  NAND U1944 ( .A(b[1]), .B(a[66]), .Z(n1814) );
  XNOR U1945 ( .A(n1813), .B(n1814), .Z(n1819) );
  NAND U1946 ( .A(b[0]), .B(a[67]), .Z(n1820) );
  XOR U1947 ( .A(n1819), .B(n1820), .Z(n1822) );
  XOR U1948 ( .A(n1821), .B(n1822), .Z(n1807) );
  NANDN U1949 ( .A(n1798), .B(n1797), .Z(n1802) );
  OR U1950 ( .A(n1800), .B(n1799), .Z(n1801) );
  AND U1951 ( .A(n1802), .B(n1801), .Z(n1806) );
  XNOR U1952 ( .A(n1807), .B(n1806), .Z(n1808) );
  XNOR U1953 ( .A(n1809), .B(n1808), .Z(n1826) );
  XNOR U1954 ( .A(n1825), .B(sreg[191]), .Z(n1805) );
  XNOR U1955 ( .A(n1826), .B(n1805), .Z(c[191]) );
  NANDN U1956 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U1957 ( .A(n1809), .B(n1808), .Z(n1810) );
  AND U1958 ( .A(n1811), .B(n1810), .Z(n1830) );
  AND U1959 ( .A(b[3]), .B(a[65]), .Z(n1818) );
  AND U1960 ( .A(b[2]), .B(a[64]), .Z(n1812) );
  NAND U1961 ( .A(n1818), .B(n1812), .Z(n1816) );
  NANDN U1962 ( .A(n1814), .B(n1813), .Z(n1815) );
  AND U1963 ( .A(n1816), .B(n1815), .Z(n1843) );
  NAND U1964 ( .A(a[66]), .B(b[2]), .Z(n1817) );
  XNOR U1965 ( .A(n1818), .B(n1817), .Z(n1835) );
  NAND U1966 ( .A(b[1]), .B(a[67]), .Z(n1836) );
  XNOR U1967 ( .A(n1835), .B(n1836), .Z(n1841) );
  NAND U1968 ( .A(b[0]), .B(a[68]), .Z(n1842) );
  XOR U1969 ( .A(n1841), .B(n1842), .Z(n1844) );
  XOR U1970 ( .A(n1843), .B(n1844), .Z(n1829) );
  NANDN U1971 ( .A(n1820), .B(n1819), .Z(n1824) );
  OR U1972 ( .A(n1822), .B(n1821), .Z(n1823) );
  AND U1973 ( .A(n1824), .B(n1823), .Z(n1828) );
  XOR U1974 ( .A(n1829), .B(n1828), .Z(n1831) );
  XNOR U1975 ( .A(n1830), .B(n1831), .Z(n1848) );
  XOR U1976 ( .A(sreg[192]), .B(n1847), .Z(n1827) );
  XNOR U1977 ( .A(n1848), .B(n1827), .Z(c[192]) );
  NANDN U1978 ( .A(n1829), .B(n1828), .Z(n1833) );
  OR U1979 ( .A(n1831), .B(n1830), .Z(n1832) );
  AND U1980 ( .A(n1833), .B(n1832), .Z(n1852) );
  AND U1981 ( .A(b[3]), .B(a[66]), .Z(n1840) );
  AND U1982 ( .A(b[2]), .B(a[65]), .Z(n1834) );
  NAND U1983 ( .A(n1840), .B(n1834), .Z(n1838) );
  NANDN U1984 ( .A(n1836), .B(n1835), .Z(n1837) );
  AND U1985 ( .A(n1838), .B(n1837), .Z(n1865) );
  NAND U1986 ( .A(a[67]), .B(b[2]), .Z(n1839) );
  XNOR U1987 ( .A(n1840), .B(n1839), .Z(n1857) );
  NAND U1988 ( .A(b[1]), .B(a[68]), .Z(n1858) );
  XNOR U1989 ( .A(n1857), .B(n1858), .Z(n1863) );
  NAND U1990 ( .A(b[0]), .B(a[69]), .Z(n1864) );
  XOR U1991 ( .A(n1863), .B(n1864), .Z(n1866) );
  XOR U1992 ( .A(n1865), .B(n1866), .Z(n1851) );
  NANDN U1993 ( .A(n1842), .B(n1841), .Z(n1846) );
  OR U1994 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U1995 ( .A(n1846), .B(n1845), .Z(n1850) );
  XOR U1996 ( .A(n1851), .B(n1850), .Z(n1853) );
  XNOR U1997 ( .A(n1852), .B(n1853), .Z(n1870) );
  XNOR U1998 ( .A(sreg[193]), .B(n1869), .Z(n1849) );
  XNOR U1999 ( .A(n1870), .B(n1849), .Z(c[193]) );
  NANDN U2000 ( .A(n1851), .B(n1850), .Z(n1855) );
  OR U2001 ( .A(n1853), .B(n1852), .Z(n1854) );
  AND U2002 ( .A(n1855), .B(n1854), .Z(n1874) );
  AND U2003 ( .A(b[3]), .B(a[67]), .Z(n1862) );
  AND U2004 ( .A(b[2]), .B(a[66]), .Z(n1856) );
  NAND U2005 ( .A(n1862), .B(n1856), .Z(n1860) );
  NANDN U2006 ( .A(n1858), .B(n1857), .Z(n1859) );
  AND U2007 ( .A(n1860), .B(n1859), .Z(n1887) );
  NAND U2008 ( .A(a[68]), .B(b[2]), .Z(n1861) );
  XNOR U2009 ( .A(n1862), .B(n1861), .Z(n1879) );
  NAND U2010 ( .A(b[1]), .B(a[69]), .Z(n1880) );
  XNOR U2011 ( .A(n1879), .B(n1880), .Z(n1885) );
  NAND U2012 ( .A(b[0]), .B(a[70]), .Z(n1886) );
  XOR U2013 ( .A(n1885), .B(n1886), .Z(n1888) );
  XOR U2014 ( .A(n1887), .B(n1888), .Z(n1873) );
  NANDN U2015 ( .A(n1864), .B(n1863), .Z(n1868) );
  OR U2016 ( .A(n1866), .B(n1865), .Z(n1867) );
  AND U2017 ( .A(n1868), .B(n1867), .Z(n1872) );
  XOR U2018 ( .A(n1873), .B(n1872), .Z(n1875) );
  XNOR U2019 ( .A(n1874), .B(n1875), .Z(n1892) );
  XNOR U2020 ( .A(sreg[194]), .B(n1891), .Z(n1871) );
  XNOR U2021 ( .A(n1892), .B(n1871), .Z(c[194]) );
  NANDN U2022 ( .A(n1873), .B(n1872), .Z(n1877) );
  OR U2023 ( .A(n1875), .B(n1874), .Z(n1876) );
  AND U2024 ( .A(n1877), .B(n1876), .Z(n1897) );
  AND U2025 ( .A(b[3]), .B(a[68]), .Z(n1884) );
  AND U2026 ( .A(b[2]), .B(a[67]), .Z(n1878) );
  NAND U2027 ( .A(n1884), .B(n1878), .Z(n1882) );
  NANDN U2028 ( .A(n1880), .B(n1879), .Z(n1881) );
  AND U2029 ( .A(n1882), .B(n1881), .Z(n1909) );
  NAND U2030 ( .A(a[69]), .B(b[2]), .Z(n1883) );
  XNOR U2031 ( .A(n1884), .B(n1883), .Z(n1901) );
  NAND U2032 ( .A(b[1]), .B(a[70]), .Z(n1902) );
  XNOR U2033 ( .A(n1901), .B(n1902), .Z(n1907) );
  NAND U2034 ( .A(b[0]), .B(a[71]), .Z(n1908) );
  XOR U2035 ( .A(n1907), .B(n1908), .Z(n1910) );
  XOR U2036 ( .A(n1909), .B(n1910), .Z(n1895) );
  NANDN U2037 ( .A(n1886), .B(n1885), .Z(n1890) );
  OR U2038 ( .A(n1888), .B(n1887), .Z(n1889) );
  AND U2039 ( .A(n1890), .B(n1889), .Z(n1894) );
  XNOR U2040 ( .A(n1895), .B(n1894), .Z(n1896) );
  XNOR U2041 ( .A(n1897), .B(n1896), .Z(n1914) );
  XOR U2042 ( .A(n1913), .B(sreg[195]), .Z(n1893) );
  XNOR U2043 ( .A(n1914), .B(n1893), .Z(c[195]) );
  NANDN U2044 ( .A(n1895), .B(n1894), .Z(n1899) );
  NANDN U2045 ( .A(n1897), .B(n1896), .Z(n1898) );
  AND U2046 ( .A(n1899), .B(n1898), .Z(n1918) );
  AND U2047 ( .A(b[3]), .B(a[69]), .Z(n1906) );
  AND U2048 ( .A(b[2]), .B(a[68]), .Z(n1900) );
  NAND U2049 ( .A(n1906), .B(n1900), .Z(n1904) );
  NANDN U2050 ( .A(n1902), .B(n1901), .Z(n1903) );
  AND U2051 ( .A(n1904), .B(n1903), .Z(n1931) );
  NAND U2052 ( .A(a[70]), .B(b[2]), .Z(n1905) );
  XNOR U2053 ( .A(n1906), .B(n1905), .Z(n1923) );
  NAND U2054 ( .A(b[1]), .B(a[71]), .Z(n1924) );
  XNOR U2055 ( .A(n1923), .B(n1924), .Z(n1929) );
  NAND U2056 ( .A(b[0]), .B(a[72]), .Z(n1930) );
  XOR U2057 ( .A(n1929), .B(n1930), .Z(n1932) );
  XOR U2058 ( .A(n1931), .B(n1932), .Z(n1917) );
  NANDN U2059 ( .A(n1908), .B(n1907), .Z(n1912) );
  OR U2060 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2061 ( .A(n1912), .B(n1911), .Z(n1916) );
  XOR U2062 ( .A(n1917), .B(n1916), .Z(n1919) );
  XNOR U2063 ( .A(n1918), .B(n1919), .Z(n1936) );
  XOR U2064 ( .A(sreg[196]), .B(n1935), .Z(n1915) );
  XNOR U2065 ( .A(n1936), .B(n1915), .Z(c[196]) );
  NANDN U2066 ( .A(n1917), .B(n1916), .Z(n1921) );
  OR U2067 ( .A(n1919), .B(n1918), .Z(n1920) );
  AND U2068 ( .A(n1921), .B(n1920), .Z(n1941) );
  AND U2069 ( .A(b[3]), .B(a[70]), .Z(n1928) );
  AND U2070 ( .A(b[2]), .B(a[69]), .Z(n1922) );
  NAND U2071 ( .A(n1928), .B(n1922), .Z(n1926) );
  NANDN U2072 ( .A(n1924), .B(n1923), .Z(n1925) );
  AND U2073 ( .A(n1926), .B(n1925), .Z(n1953) );
  NAND U2074 ( .A(a[71]), .B(b[2]), .Z(n1927) );
  XNOR U2075 ( .A(n1928), .B(n1927), .Z(n1945) );
  NAND U2076 ( .A(b[1]), .B(a[72]), .Z(n1946) );
  XNOR U2077 ( .A(n1945), .B(n1946), .Z(n1951) );
  NAND U2078 ( .A(b[0]), .B(a[73]), .Z(n1952) );
  XOR U2079 ( .A(n1951), .B(n1952), .Z(n1954) );
  XOR U2080 ( .A(n1953), .B(n1954), .Z(n1939) );
  NANDN U2081 ( .A(n1930), .B(n1929), .Z(n1934) );
  OR U2082 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2083 ( .A(n1934), .B(n1933), .Z(n1938) );
  XNOR U2084 ( .A(n1939), .B(n1938), .Z(n1940) );
  XNOR U2085 ( .A(n1941), .B(n1940), .Z(n1958) );
  XOR U2086 ( .A(n1957), .B(sreg[197]), .Z(n1937) );
  XNOR U2087 ( .A(n1958), .B(n1937), .Z(c[197]) );
  NANDN U2088 ( .A(n1939), .B(n1938), .Z(n1943) );
  NANDN U2089 ( .A(n1941), .B(n1940), .Z(n1942) );
  AND U2090 ( .A(n1943), .B(n1942), .Z(n1962) );
  AND U2091 ( .A(b[3]), .B(a[71]), .Z(n1950) );
  AND U2092 ( .A(b[2]), .B(a[70]), .Z(n1944) );
  NAND U2093 ( .A(n1950), .B(n1944), .Z(n1948) );
  NANDN U2094 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2095 ( .A(n1948), .B(n1947), .Z(n1975) );
  NAND U2096 ( .A(a[72]), .B(b[2]), .Z(n1949) );
  XNOR U2097 ( .A(n1950), .B(n1949), .Z(n1967) );
  NAND U2098 ( .A(b[1]), .B(a[73]), .Z(n1968) );
  XNOR U2099 ( .A(n1967), .B(n1968), .Z(n1973) );
  NAND U2100 ( .A(b[0]), .B(a[74]), .Z(n1974) );
  XOR U2101 ( .A(n1973), .B(n1974), .Z(n1976) );
  XOR U2102 ( .A(n1975), .B(n1976), .Z(n1961) );
  NANDN U2103 ( .A(n1952), .B(n1951), .Z(n1956) );
  OR U2104 ( .A(n1954), .B(n1953), .Z(n1955) );
  AND U2105 ( .A(n1956), .B(n1955), .Z(n1960) );
  XOR U2106 ( .A(n1961), .B(n1960), .Z(n1963) );
  XNOR U2107 ( .A(n1962), .B(n1963), .Z(n1980) );
  XOR U2108 ( .A(sreg[198]), .B(n1979), .Z(n1959) );
  XNOR U2109 ( .A(n1980), .B(n1959), .Z(c[198]) );
  NANDN U2110 ( .A(n1961), .B(n1960), .Z(n1965) );
  OR U2111 ( .A(n1963), .B(n1962), .Z(n1964) );
  AND U2112 ( .A(n1965), .B(n1964), .Z(n1984) );
  AND U2113 ( .A(b[3]), .B(a[72]), .Z(n1972) );
  AND U2114 ( .A(b[2]), .B(a[71]), .Z(n1966) );
  NAND U2115 ( .A(n1972), .B(n1966), .Z(n1970) );
  NANDN U2116 ( .A(n1968), .B(n1967), .Z(n1969) );
  AND U2117 ( .A(n1970), .B(n1969), .Z(n1997) );
  NAND U2118 ( .A(a[73]), .B(b[2]), .Z(n1971) );
  XNOR U2119 ( .A(n1972), .B(n1971), .Z(n1989) );
  NAND U2120 ( .A(b[1]), .B(a[74]), .Z(n1990) );
  XNOR U2121 ( .A(n1989), .B(n1990), .Z(n1995) );
  NAND U2122 ( .A(b[0]), .B(a[75]), .Z(n1996) );
  XOR U2123 ( .A(n1995), .B(n1996), .Z(n1998) );
  XOR U2124 ( .A(n1997), .B(n1998), .Z(n1983) );
  NANDN U2125 ( .A(n1974), .B(n1973), .Z(n1978) );
  OR U2126 ( .A(n1976), .B(n1975), .Z(n1977) );
  AND U2127 ( .A(n1978), .B(n1977), .Z(n1982) );
  XOR U2128 ( .A(n1983), .B(n1982), .Z(n1985) );
  XNOR U2129 ( .A(n1984), .B(n1985), .Z(n2002) );
  XNOR U2130 ( .A(sreg[199]), .B(n2001), .Z(n1981) );
  XNOR U2131 ( .A(n2002), .B(n1981), .Z(c[199]) );
  NANDN U2132 ( .A(n1983), .B(n1982), .Z(n1987) );
  OR U2133 ( .A(n1985), .B(n1984), .Z(n1986) );
  AND U2134 ( .A(n1987), .B(n1986), .Z(n2006) );
  AND U2135 ( .A(b[3]), .B(a[73]), .Z(n1994) );
  AND U2136 ( .A(b[2]), .B(a[72]), .Z(n1988) );
  NAND U2137 ( .A(n1994), .B(n1988), .Z(n1992) );
  NANDN U2138 ( .A(n1990), .B(n1989), .Z(n1991) );
  AND U2139 ( .A(n1992), .B(n1991), .Z(n2019) );
  NAND U2140 ( .A(a[74]), .B(b[2]), .Z(n1993) );
  XNOR U2141 ( .A(n1994), .B(n1993), .Z(n2011) );
  NAND U2142 ( .A(b[1]), .B(a[75]), .Z(n2012) );
  XNOR U2143 ( .A(n2011), .B(n2012), .Z(n2017) );
  NAND U2144 ( .A(b[0]), .B(a[76]), .Z(n2018) );
  XOR U2145 ( .A(n2017), .B(n2018), .Z(n2020) );
  XOR U2146 ( .A(n2019), .B(n2020), .Z(n2005) );
  NANDN U2147 ( .A(n1996), .B(n1995), .Z(n2000) );
  OR U2148 ( .A(n1998), .B(n1997), .Z(n1999) );
  AND U2149 ( .A(n2000), .B(n1999), .Z(n2004) );
  XOR U2150 ( .A(n2005), .B(n2004), .Z(n2007) );
  XNOR U2151 ( .A(n2006), .B(n2007), .Z(n2024) );
  XNOR U2152 ( .A(sreg[200]), .B(n2023), .Z(n2003) );
  XNOR U2153 ( .A(n2024), .B(n2003), .Z(c[200]) );
  NANDN U2154 ( .A(n2005), .B(n2004), .Z(n2009) );
  OR U2155 ( .A(n2007), .B(n2006), .Z(n2008) );
  AND U2156 ( .A(n2009), .B(n2008), .Z(n2028) );
  AND U2157 ( .A(b[3]), .B(a[74]), .Z(n2016) );
  AND U2158 ( .A(b[2]), .B(a[73]), .Z(n2010) );
  NAND U2159 ( .A(n2016), .B(n2010), .Z(n2014) );
  NANDN U2160 ( .A(n2012), .B(n2011), .Z(n2013) );
  AND U2161 ( .A(n2014), .B(n2013), .Z(n2041) );
  NAND U2162 ( .A(a[75]), .B(b[2]), .Z(n2015) );
  XNOR U2163 ( .A(n2016), .B(n2015), .Z(n2033) );
  NAND U2164 ( .A(b[1]), .B(a[76]), .Z(n2034) );
  XNOR U2165 ( .A(n2033), .B(n2034), .Z(n2039) );
  NAND U2166 ( .A(b[0]), .B(a[77]), .Z(n2040) );
  XOR U2167 ( .A(n2039), .B(n2040), .Z(n2042) );
  XOR U2168 ( .A(n2041), .B(n2042), .Z(n2027) );
  NANDN U2169 ( .A(n2018), .B(n2017), .Z(n2022) );
  OR U2170 ( .A(n2020), .B(n2019), .Z(n2021) );
  AND U2171 ( .A(n2022), .B(n2021), .Z(n2026) );
  XOR U2172 ( .A(n2027), .B(n2026), .Z(n2029) );
  XNOR U2173 ( .A(n2028), .B(n2029), .Z(n2046) );
  XNOR U2174 ( .A(sreg[201]), .B(n2045), .Z(n2025) );
  XNOR U2175 ( .A(n2046), .B(n2025), .Z(c[201]) );
  NANDN U2176 ( .A(n2027), .B(n2026), .Z(n2031) );
  OR U2177 ( .A(n2029), .B(n2028), .Z(n2030) );
  AND U2178 ( .A(n2031), .B(n2030), .Z(n2050) );
  AND U2179 ( .A(b[3]), .B(a[75]), .Z(n2038) );
  AND U2180 ( .A(b[2]), .B(a[74]), .Z(n2032) );
  NAND U2181 ( .A(n2038), .B(n2032), .Z(n2036) );
  NANDN U2182 ( .A(n2034), .B(n2033), .Z(n2035) );
  AND U2183 ( .A(n2036), .B(n2035), .Z(n2063) );
  NAND U2184 ( .A(a[76]), .B(b[2]), .Z(n2037) );
  XNOR U2185 ( .A(n2038), .B(n2037), .Z(n2055) );
  NAND U2186 ( .A(b[1]), .B(a[77]), .Z(n2056) );
  XNOR U2187 ( .A(n2055), .B(n2056), .Z(n2061) );
  NAND U2188 ( .A(b[0]), .B(a[78]), .Z(n2062) );
  XOR U2189 ( .A(n2061), .B(n2062), .Z(n2064) );
  XOR U2190 ( .A(n2063), .B(n2064), .Z(n2049) );
  NANDN U2191 ( .A(n2040), .B(n2039), .Z(n2044) );
  OR U2192 ( .A(n2042), .B(n2041), .Z(n2043) );
  AND U2193 ( .A(n2044), .B(n2043), .Z(n2048) );
  XOR U2194 ( .A(n2049), .B(n2048), .Z(n2051) );
  XNOR U2195 ( .A(n2050), .B(n2051), .Z(n2068) );
  XNOR U2196 ( .A(sreg[202]), .B(n2067), .Z(n2047) );
  XNOR U2197 ( .A(n2068), .B(n2047), .Z(c[202]) );
  NANDN U2198 ( .A(n2049), .B(n2048), .Z(n2053) );
  OR U2199 ( .A(n2051), .B(n2050), .Z(n2052) );
  AND U2200 ( .A(n2053), .B(n2052), .Z(n2072) );
  AND U2201 ( .A(b[3]), .B(a[76]), .Z(n2060) );
  AND U2202 ( .A(b[2]), .B(a[75]), .Z(n2054) );
  NAND U2203 ( .A(n2060), .B(n2054), .Z(n2058) );
  NANDN U2204 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U2205 ( .A(n2058), .B(n2057), .Z(n2085) );
  NAND U2206 ( .A(a[77]), .B(b[2]), .Z(n2059) );
  XNOR U2207 ( .A(n2060), .B(n2059), .Z(n2077) );
  NAND U2208 ( .A(b[1]), .B(a[78]), .Z(n2078) );
  XNOR U2209 ( .A(n2077), .B(n2078), .Z(n2083) );
  NAND U2210 ( .A(b[0]), .B(a[79]), .Z(n2084) );
  XOR U2211 ( .A(n2083), .B(n2084), .Z(n2086) );
  XOR U2212 ( .A(n2085), .B(n2086), .Z(n2071) );
  NANDN U2213 ( .A(n2062), .B(n2061), .Z(n2066) );
  OR U2214 ( .A(n2064), .B(n2063), .Z(n2065) );
  AND U2215 ( .A(n2066), .B(n2065), .Z(n2070) );
  XOR U2216 ( .A(n2071), .B(n2070), .Z(n2073) );
  XNOR U2217 ( .A(n2072), .B(n2073), .Z(n2090) );
  XNOR U2218 ( .A(sreg[203]), .B(n2089), .Z(n2069) );
  XNOR U2219 ( .A(n2090), .B(n2069), .Z(c[203]) );
  NANDN U2220 ( .A(n2071), .B(n2070), .Z(n2075) );
  OR U2221 ( .A(n2073), .B(n2072), .Z(n2074) );
  AND U2222 ( .A(n2075), .B(n2074), .Z(n2095) );
  AND U2223 ( .A(b[3]), .B(a[77]), .Z(n2082) );
  AND U2224 ( .A(b[2]), .B(a[76]), .Z(n2076) );
  NAND U2225 ( .A(n2082), .B(n2076), .Z(n2080) );
  NANDN U2226 ( .A(n2078), .B(n2077), .Z(n2079) );
  AND U2227 ( .A(n2080), .B(n2079), .Z(n2107) );
  NAND U2228 ( .A(a[78]), .B(b[2]), .Z(n2081) );
  XNOR U2229 ( .A(n2082), .B(n2081), .Z(n2099) );
  NAND U2230 ( .A(b[1]), .B(a[79]), .Z(n2100) );
  XNOR U2231 ( .A(n2099), .B(n2100), .Z(n2105) );
  NAND U2232 ( .A(b[0]), .B(a[80]), .Z(n2106) );
  XOR U2233 ( .A(n2105), .B(n2106), .Z(n2108) );
  XOR U2234 ( .A(n2107), .B(n2108), .Z(n2093) );
  NANDN U2235 ( .A(n2084), .B(n2083), .Z(n2088) );
  OR U2236 ( .A(n2086), .B(n2085), .Z(n2087) );
  AND U2237 ( .A(n2088), .B(n2087), .Z(n2092) );
  XNOR U2238 ( .A(n2093), .B(n2092), .Z(n2094) );
  XNOR U2239 ( .A(n2095), .B(n2094), .Z(n2112) );
  XOR U2240 ( .A(n2111), .B(sreg[204]), .Z(n2091) );
  XNOR U2241 ( .A(n2112), .B(n2091), .Z(c[204]) );
  NANDN U2242 ( .A(n2093), .B(n2092), .Z(n2097) );
  NANDN U2243 ( .A(n2095), .B(n2094), .Z(n2096) );
  AND U2244 ( .A(n2097), .B(n2096), .Z(n2116) );
  AND U2245 ( .A(b[3]), .B(a[78]), .Z(n2104) );
  AND U2246 ( .A(b[2]), .B(a[77]), .Z(n2098) );
  NAND U2247 ( .A(n2104), .B(n2098), .Z(n2102) );
  NANDN U2248 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2249 ( .A(n2102), .B(n2101), .Z(n2129) );
  NAND U2250 ( .A(a[79]), .B(b[2]), .Z(n2103) );
  XNOR U2251 ( .A(n2104), .B(n2103), .Z(n2121) );
  NAND U2252 ( .A(b[1]), .B(a[80]), .Z(n2122) );
  XNOR U2253 ( .A(n2121), .B(n2122), .Z(n2127) );
  NAND U2254 ( .A(b[0]), .B(a[81]), .Z(n2128) );
  XOR U2255 ( .A(n2127), .B(n2128), .Z(n2130) );
  XOR U2256 ( .A(n2129), .B(n2130), .Z(n2115) );
  NANDN U2257 ( .A(n2106), .B(n2105), .Z(n2110) );
  OR U2258 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U2259 ( .A(n2110), .B(n2109), .Z(n2114) );
  XOR U2260 ( .A(n2115), .B(n2114), .Z(n2117) );
  XNOR U2261 ( .A(n2116), .B(n2117), .Z(n2134) );
  XOR U2262 ( .A(sreg[205]), .B(n2133), .Z(n2113) );
  XNOR U2263 ( .A(n2134), .B(n2113), .Z(c[205]) );
  NANDN U2264 ( .A(n2115), .B(n2114), .Z(n2119) );
  OR U2265 ( .A(n2117), .B(n2116), .Z(n2118) );
  AND U2266 ( .A(n2119), .B(n2118), .Z(n2139) );
  AND U2267 ( .A(b[3]), .B(a[79]), .Z(n2126) );
  AND U2268 ( .A(b[2]), .B(a[78]), .Z(n2120) );
  NAND U2269 ( .A(n2126), .B(n2120), .Z(n2124) );
  NANDN U2270 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U2271 ( .A(n2124), .B(n2123), .Z(n2151) );
  NAND U2272 ( .A(a[80]), .B(b[2]), .Z(n2125) );
  XNOR U2273 ( .A(n2126), .B(n2125), .Z(n2143) );
  NAND U2274 ( .A(b[1]), .B(a[81]), .Z(n2144) );
  XNOR U2275 ( .A(n2143), .B(n2144), .Z(n2149) );
  NAND U2276 ( .A(b[0]), .B(a[82]), .Z(n2150) );
  XOR U2277 ( .A(n2149), .B(n2150), .Z(n2152) );
  XOR U2278 ( .A(n2151), .B(n2152), .Z(n2137) );
  NANDN U2279 ( .A(n2128), .B(n2127), .Z(n2132) );
  OR U2280 ( .A(n2130), .B(n2129), .Z(n2131) );
  AND U2281 ( .A(n2132), .B(n2131), .Z(n2136) );
  XNOR U2282 ( .A(n2137), .B(n2136), .Z(n2138) );
  XNOR U2283 ( .A(n2139), .B(n2138), .Z(n2156) );
  XOR U2284 ( .A(n2155), .B(sreg[206]), .Z(n2135) );
  XNOR U2285 ( .A(n2156), .B(n2135), .Z(c[206]) );
  NANDN U2286 ( .A(n2137), .B(n2136), .Z(n2141) );
  NANDN U2287 ( .A(n2139), .B(n2138), .Z(n2140) );
  AND U2288 ( .A(n2141), .B(n2140), .Z(n2160) );
  AND U2289 ( .A(b[3]), .B(a[80]), .Z(n2148) );
  AND U2290 ( .A(b[2]), .B(a[79]), .Z(n2142) );
  NAND U2291 ( .A(n2148), .B(n2142), .Z(n2146) );
  NANDN U2292 ( .A(n2144), .B(n2143), .Z(n2145) );
  AND U2293 ( .A(n2146), .B(n2145), .Z(n2173) );
  NAND U2294 ( .A(a[81]), .B(b[2]), .Z(n2147) );
  XNOR U2295 ( .A(n2148), .B(n2147), .Z(n2165) );
  NAND U2296 ( .A(b[1]), .B(a[82]), .Z(n2166) );
  XNOR U2297 ( .A(n2165), .B(n2166), .Z(n2171) );
  NAND U2298 ( .A(b[0]), .B(a[83]), .Z(n2172) );
  XOR U2299 ( .A(n2171), .B(n2172), .Z(n2174) );
  XOR U2300 ( .A(n2173), .B(n2174), .Z(n2159) );
  NANDN U2301 ( .A(n2150), .B(n2149), .Z(n2154) );
  OR U2302 ( .A(n2152), .B(n2151), .Z(n2153) );
  AND U2303 ( .A(n2154), .B(n2153), .Z(n2158) );
  XOR U2304 ( .A(n2159), .B(n2158), .Z(n2161) );
  XNOR U2305 ( .A(n2160), .B(n2161), .Z(n2178) );
  XOR U2306 ( .A(sreg[207]), .B(n2177), .Z(n2157) );
  XNOR U2307 ( .A(n2178), .B(n2157), .Z(c[207]) );
  NANDN U2308 ( .A(n2159), .B(n2158), .Z(n2163) );
  OR U2309 ( .A(n2161), .B(n2160), .Z(n2162) );
  AND U2310 ( .A(n2163), .B(n2162), .Z(n2182) );
  AND U2311 ( .A(b[3]), .B(a[81]), .Z(n2170) );
  AND U2312 ( .A(b[2]), .B(a[80]), .Z(n2164) );
  NAND U2313 ( .A(n2170), .B(n2164), .Z(n2168) );
  NANDN U2314 ( .A(n2166), .B(n2165), .Z(n2167) );
  AND U2315 ( .A(n2168), .B(n2167), .Z(n2195) );
  NAND U2316 ( .A(a[82]), .B(b[2]), .Z(n2169) );
  XNOR U2317 ( .A(n2170), .B(n2169), .Z(n2187) );
  NAND U2318 ( .A(b[1]), .B(a[83]), .Z(n2188) );
  XNOR U2319 ( .A(n2187), .B(n2188), .Z(n2193) );
  NAND U2320 ( .A(b[0]), .B(a[84]), .Z(n2194) );
  XOR U2321 ( .A(n2193), .B(n2194), .Z(n2196) );
  XOR U2322 ( .A(n2195), .B(n2196), .Z(n2181) );
  NANDN U2323 ( .A(n2172), .B(n2171), .Z(n2176) );
  OR U2324 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U2325 ( .A(n2176), .B(n2175), .Z(n2180) );
  XOR U2326 ( .A(n2181), .B(n2180), .Z(n2183) );
  XNOR U2327 ( .A(n2182), .B(n2183), .Z(n2200) );
  XNOR U2328 ( .A(sreg[208]), .B(n2199), .Z(n2179) );
  XNOR U2329 ( .A(n2200), .B(n2179), .Z(c[208]) );
  NANDN U2330 ( .A(n2181), .B(n2180), .Z(n2185) );
  OR U2331 ( .A(n2183), .B(n2182), .Z(n2184) );
  AND U2332 ( .A(n2185), .B(n2184), .Z(n2204) );
  AND U2333 ( .A(b[3]), .B(a[82]), .Z(n2192) );
  AND U2334 ( .A(b[2]), .B(a[81]), .Z(n2186) );
  NAND U2335 ( .A(n2192), .B(n2186), .Z(n2190) );
  NANDN U2336 ( .A(n2188), .B(n2187), .Z(n2189) );
  AND U2337 ( .A(n2190), .B(n2189), .Z(n2217) );
  NAND U2338 ( .A(a[83]), .B(b[2]), .Z(n2191) );
  XNOR U2339 ( .A(n2192), .B(n2191), .Z(n2209) );
  NAND U2340 ( .A(b[1]), .B(a[84]), .Z(n2210) );
  XNOR U2341 ( .A(n2209), .B(n2210), .Z(n2215) );
  NAND U2342 ( .A(b[0]), .B(a[85]), .Z(n2216) );
  XOR U2343 ( .A(n2215), .B(n2216), .Z(n2218) );
  XOR U2344 ( .A(n2217), .B(n2218), .Z(n2203) );
  NANDN U2345 ( .A(n2194), .B(n2193), .Z(n2198) );
  OR U2346 ( .A(n2196), .B(n2195), .Z(n2197) );
  AND U2347 ( .A(n2198), .B(n2197), .Z(n2202) );
  XOR U2348 ( .A(n2203), .B(n2202), .Z(n2205) );
  XNOR U2349 ( .A(n2204), .B(n2205), .Z(n2222) );
  XNOR U2350 ( .A(sreg[209]), .B(n2221), .Z(n2201) );
  XNOR U2351 ( .A(n2222), .B(n2201), .Z(c[209]) );
  NANDN U2352 ( .A(n2203), .B(n2202), .Z(n2207) );
  OR U2353 ( .A(n2205), .B(n2204), .Z(n2206) );
  AND U2354 ( .A(n2207), .B(n2206), .Z(n2226) );
  AND U2355 ( .A(b[3]), .B(a[83]), .Z(n2214) );
  AND U2356 ( .A(b[2]), .B(a[82]), .Z(n2208) );
  NAND U2357 ( .A(n2214), .B(n2208), .Z(n2212) );
  NANDN U2358 ( .A(n2210), .B(n2209), .Z(n2211) );
  AND U2359 ( .A(n2212), .B(n2211), .Z(n2239) );
  NAND U2360 ( .A(a[84]), .B(b[2]), .Z(n2213) );
  XNOR U2361 ( .A(n2214), .B(n2213), .Z(n2231) );
  NAND U2362 ( .A(b[1]), .B(a[85]), .Z(n2232) );
  XNOR U2363 ( .A(n2231), .B(n2232), .Z(n2237) );
  NAND U2364 ( .A(b[0]), .B(a[86]), .Z(n2238) );
  XOR U2365 ( .A(n2237), .B(n2238), .Z(n2240) );
  XOR U2366 ( .A(n2239), .B(n2240), .Z(n2225) );
  NANDN U2367 ( .A(n2216), .B(n2215), .Z(n2220) );
  OR U2368 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U2369 ( .A(n2220), .B(n2219), .Z(n2224) );
  XOR U2370 ( .A(n2225), .B(n2224), .Z(n2227) );
  XNOR U2371 ( .A(n2226), .B(n2227), .Z(n2244) );
  XNOR U2372 ( .A(sreg[210]), .B(n2243), .Z(n2223) );
  XNOR U2373 ( .A(n2244), .B(n2223), .Z(c[210]) );
  NANDN U2374 ( .A(n2225), .B(n2224), .Z(n2229) );
  OR U2375 ( .A(n2227), .B(n2226), .Z(n2228) );
  AND U2376 ( .A(n2229), .B(n2228), .Z(n2249) );
  AND U2377 ( .A(b[3]), .B(a[84]), .Z(n2236) );
  AND U2378 ( .A(b[2]), .B(a[83]), .Z(n2230) );
  NAND U2379 ( .A(n2236), .B(n2230), .Z(n2234) );
  NANDN U2380 ( .A(n2232), .B(n2231), .Z(n2233) );
  AND U2381 ( .A(n2234), .B(n2233), .Z(n2261) );
  NAND U2382 ( .A(a[85]), .B(b[2]), .Z(n2235) );
  XNOR U2383 ( .A(n2236), .B(n2235), .Z(n2253) );
  NAND U2384 ( .A(b[1]), .B(a[86]), .Z(n2254) );
  XNOR U2385 ( .A(n2253), .B(n2254), .Z(n2259) );
  NAND U2386 ( .A(b[0]), .B(a[87]), .Z(n2260) );
  XOR U2387 ( .A(n2259), .B(n2260), .Z(n2262) );
  XOR U2388 ( .A(n2261), .B(n2262), .Z(n2247) );
  NANDN U2389 ( .A(n2238), .B(n2237), .Z(n2242) );
  OR U2390 ( .A(n2240), .B(n2239), .Z(n2241) );
  AND U2391 ( .A(n2242), .B(n2241), .Z(n2246) );
  XNOR U2392 ( .A(n2247), .B(n2246), .Z(n2248) );
  XNOR U2393 ( .A(n2249), .B(n2248), .Z(n2266) );
  XOR U2394 ( .A(n2265), .B(sreg[211]), .Z(n2245) );
  XNOR U2395 ( .A(n2266), .B(n2245), .Z(c[211]) );
  NANDN U2396 ( .A(n2247), .B(n2246), .Z(n2251) );
  NANDN U2397 ( .A(n2249), .B(n2248), .Z(n2250) );
  AND U2398 ( .A(n2251), .B(n2250), .Z(n2270) );
  AND U2399 ( .A(b[3]), .B(a[85]), .Z(n2258) );
  AND U2400 ( .A(b[2]), .B(a[84]), .Z(n2252) );
  NAND U2401 ( .A(n2258), .B(n2252), .Z(n2256) );
  NANDN U2402 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2403 ( .A(n2256), .B(n2255), .Z(n2283) );
  NAND U2404 ( .A(a[86]), .B(b[2]), .Z(n2257) );
  XNOR U2405 ( .A(n2258), .B(n2257), .Z(n2275) );
  NAND U2406 ( .A(b[1]), .B(a[87]), .Z(n2276) );
  XNOR U2407 ( .A(n2275), .B(n2276), .Z(n2281) );
  NAND U2408 ( .A(b[0]), .B(a[88]), .Z(n2282) );
  XOR U2409 ( .A(n2281), .B(n2282), .Z(n2284) );
  XOR U2410 ( .A(n2283), .B(n2284), .Z(n2269) );
  NANDN U2411 ( .A(n2260), .B(n2259), .Z(n2264) );
  OR U2412 ( .A(n2262), .B(n2261), .Z(n2263) );
  AND U2413 ( .A(n2264), .B(n2263), .Z(n2268) );
  XOR U2414 ( .A(n2269), .B(n2268), .Z(n2271) );
  XNOR U2415 ( .A(n2270), .B(n2271), .Z(n2288) );
  XOR U2416 ( .A(sreg[212]), .B(n2287), .Z(n2267) );
  XNOR U2417 ( .A(n2288), .B(n2267), .Z(c[212]) );
  NANDN U2418 ( .A(n2269), .B(n2268), .Z(n2273) );
  OR U2419 ( .A(n2271), .B(n2270), .Z(n2272) );
  AND U2420 ( .A(n2273), .B(n2272), .Z(n2293) );
  AND U2421 ( .A(b[3]), .B(a[86]), .Z(n2280) );
  AND U2422 ( .A(b[2]), .B(a[85]), .Z(n2274) );
  NAND U2423 ( .A(n2280), .B(n2274), .Z(n2278) );
  NANDN U2424 ( .A(n2276), .B(n2275), .Z(n2277) );
  AND U2425 ( .A(n2278), .B(n2277), .Z(n2305) );
  NAND U2426 ( .A(a[87]), .B(b[2]), .Z(n2279) );
  XNOR U2427 ( .A(n2280), .B(n2279), .Z(n2297) );
  NAND U2428 ( .A(b[1]), .B(a[88]), .Z(n2298) );
  XNOR U2429 ( .A(n2297), .B(n2298), .Z(n2303) );
  NAND U2430 ( .A(b[0]), .B(a[89]), .Z(n2304) );
  XOR U2431 ( .A(n2303), .B(n2304), .Z(n2306) );
  XOR U2432 ( .A(n2305), .B(n2306), .Z(n2291) );
  NANDN U2433 ( .A(n2282), .B(n2281), .Z(n2286) );
  OR U2434 ( .A(n2284), .B(n2283), .Z(n2285) );
  AND U2435 ( .A(n2286), .B(n2285), .Z(n2290) );
  XNOR U2436 ( .A(n2291), .B(n2290), .Z(n2292) );
  XNOR U2437 ( .A(n2293), .B(n2292), .Z(n2310) );
  XOR U2438 ( .A(n2309), .B(sreg[213]), .Z(n2289) );
  XNOR U2439 ( .A(n2310), .B(n2289), .Z(c[213]) );
  NANDN U2440 ( .A(n2291), .B(n2290), .Z(n2295) );
  NANDN U2441 ( .A(n2293), .B(n2292), .Z(n2294) );
  AND U2442 ( .A(n2295), .B(n2294), .Z(n2315) );
  AND U2443 ( .A(b[3]), .B(a[87]), .Z(n2302) );
  AND U2444 ( .A(b[2]), .B(a[86]), .Z(n2296) );
  NAND U2445 ( .A(n2302), .B(n2296), .Z(n2300) );
  NANDN U2446 ( .A(n2298), .B(n2297), .Z(n2299) );
  AND U2447 ( .A(n2300), .B(n2299), .Z(n2327) );
  NAND U2448 ( .A(a[88]), .B(b[2]), .Z(n2301) );
  XNOR U2449 ( .A(n2302), .B(n2301), .Z(n2319) );
  NAND U2450 ( .A(b[1]), .B(a[89]), .Z(n2320) );
  XNOR U2451 ( .A(n2319), .B(n2320), .Z(n2325) );
  NAND U2452 ( .A(b[0]), .B(a[90]), .Z(n2326) );
  XOR U2453 ( .A(n2325), .B(n2326), .Z(n2328) );
  XOR U2454 ( .A(n2327), .B(n2328), .Z(n2313) );
  NANDN U2455 ( .A(n2304), .B(n2303), .Z(n2308) );
  OR U2456 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U2457 ( .A(n2308), .B(n2307), .Z(n2312) );
  XNOR U2458 ( .A(n2313), .B(n2312), .Z(n2314) );
  XNOR U2459 ( .A(n2315), .B(n2314), .Z(n2332) );
  XNOR U2460 ( .A(n2331), .B(sreg[214]), .Z(n2311) );
  XNOR U2461 ( .A(n2332), .B(n2311), .Z(c[214]) );
  NANDN U2462 ( .A(n2313), .B(n2312), .Z(n2317) );
  NANDN U2463 ( .A(n2315), .B(n2314), .Z(n2316) );
  AND U2464 ( .A(n2317), .B(n2316), .Z(n2336) );
  AND U2465 ( .A(b[3]), .B(a[88]), .Z(n2324) );
  AND U2466 ( .A(b[2]), .B(a[87]), .Z(n2318) );
  NAND U2467 ( .A(n2324), .B(n2318), .Z(n2322) );
  NANDN U2468 ( .A(n2320), .B(n2319), .Z(n2321) );
  AND U2469 ( .A(n2322), .B(n2321), .Z(n2349) );
  NAND U2470 ( .A(a[89]), .B(b[2]), .Z(n2323) );
  XNOR U2471 ( .A(n2324), .B(n2323), .Z(n2341) );
  NAND U2472 ( .A(b[1]), .B(a[90]), .Z(n2342) );
  XNOR U2473 ( .A(n2341), .B(n2342), .Z(n2347) );
  NAND U2474 ( .A(b[0]), .B(a[91]), .Z(n2348) );
  XOR U2475 ( .A(n2347), .B(n2348), .Z(n2350) );
  XOR U2476 ( .A(n2349), .B(n2350), .Z(n2335) );
  NANDN U2477 ( .A(n2326), .B(n2325), .Z(n2330) );
  OR U2478 ( .A(n2328), .B(n2327), .Z(n2329) );
  AND U2479 ( .A(n2330), .B(n2329), .Z(n2334) );
  XOR U2480 ( .A(n2335), .B(n2334), .Z(n2337) );
  XNOR U2481 ( .A(n2336), .B(n2337), .Z(n2354) );
  XOR U2482 ( .A(sreg[215]), .B(n2353), .Z(n2333) );
  XNOR U2483 ( .A(n2354), .B(n2333), .Z(c[215]) );
  NANDN U2484 ( .A(n2335), .B(n2334), .Z(n2339) );
  OR U2485 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U2486 ( .A(n2339), .B(n2338), .Z(n2358) );
  AND U2487 ( .A(b[3]), .B(a[89]), .Z(n2346) );
  AND U2488 ( .A(b[2]), .B(a[88]), .Z(n2340) );
  NAND U2489 ( .A(n2346), .B(n2340), .Z(n2344) );
  NANDN U2490 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U2491 ( .A(n2344), .B(n2343), .Z(n2371) );
  NAND U2492 ( .A(a[90]), .B(b[2]), .Z(n2345) );
  XNOR U2493 ( .A(n2346), .B(n2345), .Z(n2363) );
  NAND U2494 ( .A(b[1]), .B(a[91]), .Z(n2364) );
  XNOR U2495 ( .A(n2363), .B(n2364), .Z(n2369) );
  NAND U2496 ( .A(b[0]), .B(a[92]), .Z(n2370) );
  XOR U2497 ( .A(n2369), .B(n2370), .Z(n2372) );
  XOR U2498 ( .A(n2371), .B(n2372), .Z(n2357) );
  NANDN U2499 ( .A(n2348), .B(n2347), .Z(n2352) );
  OR U2500 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U2501 ( .A(n2352), .B(n2351), .Z(n2356) );
  XOR U2502 ( .A(n2357), .B(n2356), .Z(n2359) );
  XNOR U2503 ( .A(n2358), .B(n2359), .Z(n2376) );
  XNOR U2504 ( .A(sreg[216]), .B(n2375), .Z(n2355) );
  XNOR U2505 ( .A(n2376), .B(n2355), .Z(c[216]) );
  NANDN U2506 ( .A(n2357), .B(n2356), .Z(n2361) );
  OR U2507 ( .A(n2359), .B(n2358), .Z(n2360) );
  AND U2508 ( .A(n2361), .B(n2360), .Z(n2380) );
  AND U2509 ( .A(b[3]), .B(a[90]), .Z(n2368) );
  AND U2510 ( .A(b[2]), .B(a[89]), .Z(n2362) );
  NAND U2511 ( .A(n2368), .B(n2362), .Z(n2366) );
  NANDN U2512 ( .A(n2364), .B(n2363), .Z(n2365) );
  AND U2513 ( .A(n2366), .B(n2365), .Z(n2393) );
  NAND U2514 ( .A(a[91]), .B(b[2]), .Z(n2367) );
  XNOR U2515 ( .A(n2368), .B(n2367), .Z(n2385) );
  NAND U2516 ( .A(b[1]), .B(a[92]), .Z(n2386) );
  XNOR U2517 ( .A(n2385), .B(n2386), .Z(n2391) );
  NAND U2518 ( .A(b[0]), .B(a[93]), .Z(n2392) );
  XOR U2519 ( .A(n2391), .B(n2392), .Z(n2394) );
  XOR U2520 ( .A(n2393), .B(n2394), .Z(n2379) );
  NANDN U2521 ( .A(n2370), .B(n2369), .Z(n2374) );
  OR U2522 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U2523 ( .A(n2374), .B(n2373), .Z(n2378) );
  XOR U2524 ( .A(n2379), .B(n2378), .Z(n2381) );
  XNOR U2525 ( .A(n2380), .B(n2381), .Z(n2398) );
  XNOR U2526 ( .A(sreg[217]), .B(n2397), .Z(n2377) );
  XNOR U2527 ( .A(n2398), .B(n2377), .Z(c[217]) );
  NANDN U2528 ( .A(n2379), .B(n2378), .Z(n2383) );
  OR U2529 ( .A(n2381), .B(n2380), .Z(n2382) );
  AND U2530 ( .A(n2383), .B(n2382), .Z(n2402) );
  AND U2531 ( .A(b[3]), .B(a[91]), .Z(n2390) );
  AND U2532 ( .A(b[2]), .B(a[90]), .Z(n2384) );
  NAND U2533 ( .A(n2390), .B(n2384), .Z(n2388) );
  NANDN U2534 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U2535 ( .A(n2388), .B(n2387), .Z(n2415) );
  NAND U2536 ( .A(a[92]), .B(b[2]), .Z(n2389) );
  XNOR U2537 ( .A(n2390), .B(n2389), .Z(n2407) );
  NAND U2538 ( .A(b[1]), .B(a[93]), .Z(n2408) );
  XNOR U2539 ( .A(n2407), .B(n2408), .Z(n2413) );
  NAND U2540 ( .A(b[0]), .B(a[94]), .Z(n2414) );
  XOR U2541 ( .A(n2413), .B(n2414), .Z(n2416) );
  XOR U2542 ( .A(n2415), .B(n2416), .Z(n2401) );
  NANDN U2543 ( .A(n2392), .B(n2391), .Z(n2396) );
  OR U2544 ( .A(n2394), .B(n2393), .Z(n2395) );
  AND U2545 ( .A(n2396), .B(n2395), .Z(n2400) );
  XOR U2546 ( .A(n2401), .B(n2400), .Z(n2403) );
  XNOR U2547 ( .A(n2402), .B(n2403), .Z(n2420) );
  XNOR U2548 ( .A(sreg[218]), .B(n2419), .Z(n2399) );
  XNOR U2549 ( .A(n2420), .B(n2399), .Z(c[218]) );
  NANDN U2550 ( .A(n2401), .B(n2400), .Z(n2405) );
  OR U2551 ( .A(n2403), .B(n2402), .Z(n2404) );
  AND U2552 ( .A(n2405), .B(n2404), .Z(n2424) );
  AND U2553 ( .A(b[3]), .B(a[92]), .Z(n2412) );
  AND U2554 ( .A(b[2]), .B(a[91]), .Z(n2406) );
  NAND U2555 ( .A(n2412), .B(n2406), .Z(n2410) );
  NANDN U2556 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U2557 ( .A(n2410), .B(n2409), .Z(n2437) );
  NAND U2558 ( .A(a[93]), .B(b[2]), .Z(n2411) );
  XNOR U2559 ( .A(n2412), .B(n2411), .Z(n2429) );
  NAND U2560 ( .A(b[1]), .B(a[94]), .Z(n2430) );
  XNOR U2561 ( .A(n2429), .B(n2430), .Z(n2435) );
  NAND U2562 ( .A(b[0]), .B(a[95]), .Z(n2436) );
  XOR U2563 ( .A(n2435), .B(n2436), .Z(n2438) );
  XOR U2564 ( .A(n2437), .B(n2438), .Z(n2423) );
  NANDN U2565 ( .A(n2414), .B(n2413), .Z(n2418) );
  OR U2566 ( .A(n2416), .B(n2415), .Z(n2417) );
  AND U2567 ( .A(n2418), .B(n2417), .Z(n2422) );
  XOR U2568 ( .A(n2423), .B(n2422), .Z(n2425) );
  XNOR U2569 ( .A(n2424), .B(n2425), .Z(n2442) );
  XNOR U2570 ( .A(sreg[219]), .B(n2441), .Z(n2421) );
  XNOR U2571 ( .A(n2442), .B(n2421), .Z(c[219]) );
  NANDN U2572 ( .A(n2423), .B(n2422), .Z(n2427) );
  OR U2573 ( .A(n2425), .B(n2424), .Z(n2426) );
  AND U2574 ( .A(n2427), .B(n2426), .Z(n2447) );
  AND U2575 ( .A(b[3]), .B(a[93]), .Z(n2434) );
  AND U2576 ( .A(b[2]), .B(a[92]), .Z(n2428) );
  NAND U2577 ( .A(n2434), .B(n2428), .Z(n2432) );
  NANDN U2578 ( .A(n2430), .B(n2429), .Z(n2431) );
  AND U2579 ( .A(n2432), .B(n2431), .Z(n2459) );
  NAND U2580 ( .A(a[94]), .B(b[2]), .Z(n2433) );
  XNOR U2581 ( .A(n2434), .B(n2433), .Z(n2451) );
  NAND U2582 ( .A(b[1]), .B(a[95]), .Z(n2452) );
  XNOR U2583 ( .A(n2451), .B(n2452), .Z(n2457) );
  NAND U2584 ( .A(b[0]), .B(a[96]), .Z(n2458) );
  XOR U2585 ( .A(n2457), .B(n2458), .Z(n2460) );
  XOR U2586 ( .A(n2459), .B(n2460), .Z(n2445) );
  NANDN U2587 ( .A(n2436), .B(n2435), .Z(n2440) );
  OR U2588 ( .A(n2438), .B(n2437), .Z(n2439) );
  AND U2589 ( .A(n2440), .B(n2439), .Z(n2444) );
  XNOR U2590 ( .A(n2445), .B(n2444), .Z(n2446) );
  XNOR U2591 ( .A(n2447), .B(n2446), .Z(n2464) );
  XOR U2592 ( .A(n2463), .B(sreg[220]), .Z(n2443) );
  XNOR U2593 ( .A(n2464), .B(n2443), .Z(c[220]) );
  NANDN U2594 ( .A(n2445), .B(n2444), .Z(n2449) );
  NANDN U2595 ( .A(n2447), .B(n2446), .Z(n2448) );
  AND U2596 ( .A(n2449), .B(n2448), .Z(n2468) );
  AND U2597 ( .A(b[3]), .B(a[94]), .Z(n2456) );
  AND U2598 ( .A(b[2]), .B(a[93]), .Z(n2450) );
  NAND U2599 ( .A(n2456), .B(n2450), .Z(n2454) );
  NANDN U2600 ( .A(n2452), .B(n2451), .Z(n2453) );
  AND U2601 ( .A(n2454), .B(n2453), .Z(n2481) );
  NAND U2602 ( .A(a[95]), .B(b[2]), .Z(n2455) );
  XNOR U2603 ( .A(n2456), .B(n2455), .Z(n2473) );
  NAND U2604 ( .A(b[1]), .B(a[96]), .Z(n2474) );
  XNOR U2605 ( .A(n2473), .B(n2474), .Z(n2479) );
  NAND U2606 ( .A(b[0]), .B(a[97]), .Z(n2480) );
  XOR U2607 ( .A(n2479), .B(n2480), .Z(n2482) );
  XOR U2608 ( .A(n2481), .B(n2482), .Z(n2467) );
  NANDN U2609 ( .A(n2458), .B(n2457), .Z(n2462) );
  OR U2610 ( .A(n2460), .B(n2459), .Z(n2461) );
  AND U2611 ( .A(n2462), .B(n2461), .Z(n2466) );
  XOR U2612 ( .A(n2467), .B(n2466), .Z(n2469) );
  XNOR U2613 ( .A(n2468), .B(n2469), .Z(n2486) );
  XOR U2614 ( .A(sreg[221]), .B(n2485), .Z(n2465) );
  XNOR U2615 ( .A(n2486), .B(n2465), .Z(c[221]) );
  NANDN U2616 ( .A(n2467), .B(n2466), .Z(n2471) );
  OR U2617 ( .A(n2469), .B(n2468), .Z(n2470) );
  AND U2618 ( .A(n2471), .B(n2470), .Z(n2490) );
  AND U2619 ( .A(b[3]), .B(a[95]), .Z(n2478) );
  AND U2620 ( .A(b[2]), .B(a[94]), .Z(n2472) );
  NAND U2621 ( .A(n2478), .B(n2472), .Z(n2476) );
  NANDN U2622 ( .A(n2474), .B(n2473), .Z(n2475) );
  AND U2623 ( .A(n2476), .B(n2475), .Z(n2503) );
  NAND U2624 ( .A(a[96]), .B(b[2]), .Z(n2477) );
  XNOR U2625 ( .A(n2478), .B(n2477), .Z(n2495) );
  NAND U2626 ( .A(b[1]), .B(a[97]), .Z(n2496) );
  XNOR U2627 ( .A(n2495), .B(n2496), .Z(n2501) );
  NAND U2628 ( .A(b[0]), .B(a[98]), .Z(n2502) );
  XOR U2629 ( .A(n2501), .B(n2502), .Z(n2504) );
  XOR U2630 ( .A(n2503), .B(n2504), .Z(n2489) );
  NANDN U2631 ( .A(n2480), .B(n2479), .Z(n2484) );
  OR U2632 ( .A(n2482), .B(n2481), .Z(n2483) );
  AND U2633 ( .A(n2484), .B(n2483), .Z(n2488) );
  XOR U2634 ( .A(n2489), .B(n2488), .Z(n2491) );
  XNOR U2635 ( .A(n2490), .B(n2491), .Z(n2508) );
  XNOR U2636 ( .A(sreg[222]), .B(n2507), .Z(n2487) );
  XNOR U2637 ( .A(n2508), .B(n2487), .Z(c[222]) );
  NANDN U2638 ( .A(n2489), .B(n2488), .Z(n2493) );
  OR U2639 ( .A(n2491), .B(n2490), .Z(n2492) );
  AND U2640 ( .A(n2493), .B(n2492), .Z(n2512) );
  AND U2641 ( .A(b[3]), .B(a[96]), .Z(n2500) );
  AND U2642 ( .A(b[2]), .B(a[95]), .Z(n2494) );
  NAND U2643 ( .A(n2500), .B(n2494), .Z(n2498) );
  NANDN U2644 ( .A(n2496), .B(n2495), .Z(n2497) );
  AND U2645 ( .A(n2498), .B(n2497), .Z(n2525) );
  NAND U2646 ( .A(a[97]), .B(b[2]), .Z(n2499) );
  XNOR U2647 ( .A(n2500), .B(n2499), .Z(n2517) );
  NAND U2648 ( .A(b[1]), .B(a[98]), .Z(n2518) );
  XNOR U2649 ( .A(n2517), .B(n2518), .Z(n2523) );
  NAND U2650 ( .A(b[0]), .B(a[99]), .Z(n2524) );
  XOR U2651 ( .A(n2523), .B(n2524), .Z(n2526) );
  XOR U2652 ( .A(n2525), .B(n2526), .Z(n2511) );
  NANDN U2653 ( .A(n2502), .B(n2501), .Z(n2506) );
  OR U2654 ( .A(n2504), .B(n2503), .Z(n2505) );
  AND U2655 ( .A(n2506), .B(n2505), .Z(n2510) );
  XOR U2656 ( .A(n2511), .B(n2510), .Z(n2513) );
  XNOR U2657 ( .A(n2512), .B(n2513), .Z(n2530) );
  XNOR U2658 ( .A(sreg[223]), .B(n2529), .Z(n2509) );
  XNOR U2659 ( .A(n2530), .B(n2509), .Z(c[223]) );
  NANDN U2660 ( .A(n2511), .B(n2510), .Z(n2515) );
  OR U2661 ( .A(n2513), .B(n2512), .Z(n2514) );
  AND U2662 ( .A(n2515), .B(n2514), .Z(n2534) );
  AND U2663 ( .A(b[3]), .B(a[97]), .Z(n2522) );
  AND U2664 ( .A(b[2]), .B(a[96]), .Z(n2516) );
  NAND U2665 ( .A(n2522), .B(n2516), .Z(n2520) );
  NANDN U2666 ( .A(n2518), .B(n2517), .Z(n2519) );
  AND U2667 ( .A(n2520), .B(n2519), .Z(n2547) );
  NAND U2668 ( .A(a[98]), .B(b[2]), .Z(n2521) );
  XNOR U2669 ( .A(n2522), .B(n2521), .Z(n2539) );
  NAND U2670 ( .A(b[1]), .B(a[99]), .Z(n2540) );
  XNOR U2671 ( .A(n2539), .B(n2540), .Z(n2545) );
  NAND U2672 ( .A(b[0]), .B(a[100]), .Z(n2546) );
  XOR U2673 ( .A(n2545), .B(n2546), .Z(n2548) );
  XOR U2674 ( .A(n2547), .B(n2548), .Z(n2533) );
  NANDN U2675 ( .A(n2524), .B(n2523), .Z(n2528) );
  OR U2676 ( .A(n2526), .B(n2525), .Z(n2527) );
  AND U2677 ( .A(n2528), .B(n2527), .Z(n2532) );
  XOR U2678 ( .A(n2533), .B(n2532), .Z(n2535) );
  XNOR U2679 ( .A(n2534), .B(n2535), .Z(n2552) );
  XNOR U2680 ( .A(sreg[224]), .B(n2551), .Z(n2531) );
  XNOR U2681 ( .A(n2552), .B(n2531), .Z(c[224]) );
  NANDN U2682 ( .A(n2533), .B(n2532), .Z(n2537) );
  OR U2683 ( .A(n2535), .B(n2534), .Z(n2536) );
  AND U2684 ( .A(n2537), .B(n2536), .Z(n2556) );
  AND U2685 ( .A(b[3]), .B(a[98]), .Z(n2544) );
  AND U2686 ( .A(b[2]), .B(a[97]), .Z(n2538) );
  NAND U2687 ( .A(n2544), .B(n2538), .Z(n2542) );
  NANDN U2688 ( .A(n2540), .B(n2539), .Z(n2541) );
  AND U2689 ( .A(n2542), .B(n2541), .Z(n2569) );
  NAND U2690 ( .A(a[99]), .B(b[2]), .Z(n2543) );
  XNOR U2691 ( .A(n2544), .B(n2543), .Z(n2561) );
  NAND U2692 ( .A(b[1]), .B(a[100]), .Z(n2562) );
  XNOR U2693 ( .A(n2561), .B(n2562), .Z(n2567) );
  NAND U2694 ( .A(b[0]), .B(a[101]), .Z(n2568) );
  XOR U2695 ( .A(n2567), .B(n2568), .Z(n2570) );
  XOR U2696 ( .A(n2569), .B(n2570), .Z(n2555) );
  NANDN U2697 ( .A(n2546), .B(n2545), .Z(n2550) );
  OR U2698 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U2699 ( .A(n2550), .B(n2549), .Z(n2554) );
  XOR U2700 ( .A(n2555), .B(n2554), .Z(n2557) );
  XNOR U2701 ( .A(n2556), .B(n2557), .Z(n2574) );
  XNOR U2702 ( .A(sreg[225]), .B(n2573), .Z(n2553) );
  XNOR U2703 ( .A(n2574), .B(n2553), .Z(c[225]) );
  NANDN U2704 ( .A(n2555), .B(n2554), .Z(n2559) );
  OR U2705 ( .A(n2557), .B(n2556), .Z(n2558) );
  AND U2706 ( .A(n2559), .B(n2558), .Z(n2578) );
  AND U2707 ( .A(b[3]), .B(a[99]), .Z(n2566) );
  AND U2708 ( .A(b[2]), .B(a[98]), .Z(n2560) );
  NAND U2709 ( .A(n2566), .B(n2560), .Z(n2564) );
  NANDN U2710 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U2711 ( .A(n2564), .B(n2563), .Z(n2591) );
  NAND U2712 ( .A(a[100]), .B(b[2]), .Z(n2565) );
  XNOR U2713 ( .A(n2566), .B(n2565), .Z(n2583) );
  NAND U2714 ( .A(b[1]), .B(a[101]), .Z(n2584) );
  XNOR U2715 ( .A(n2583), .B(n2584), .Z(n2589) );
  NAND U2716 ( .A(b[0]), .B(a[102]), .Z(n2590) );
  XOR U2717 ( .A(n2589), .B(n2590), .Z(n2592) );
  XOR U2718 ( .A(n2591), .B(n2592), .Z(n2577) );
  NANDN U2719 ( .A(n2568), .B(n2567), .Z(n2572) );
  OR U2720 ( .A(n2570), .B(n2569), .Z(n2571) );
  AND U2721 ( .A(n2572), .B(n2571), .Z(n2576) );
  XOR U2722 ( .A(n2577), .B(n2576), .Z(n2579) );
  XNOR U2723 ( .A(n2578), .B(n2579), .Z(n2596) );
  XNOR U2724 ( .A(sreg[226]), .B(n2595), .Z(n2575) );
  XNOR U2725 ( .A(n2596), .B(n2575), .Z(c[226]) );
  NANDN U2726 ( .A(n2577), .B(n2576), .Z(n2581) );
  OR U2727 ( .A(n2579), .B(n2578), .Z(n2580) );
  AND U2728 ( .A(n2581), .B(n2580), .Z(n2600) );
  AND U2729 ( .A(b[3]), .B(a[100]), .Z(n2588) );
  AND U2730 ( .A(b[2]), .B(a[99]), .Z(n2582) );
  NAND U2731 ( .A(n2588), .B(n2582), .Z(n2586) );
  NANDN U2732 ( .A(n2584), .B(n2583), .Z(n2585) );
  AND U2733 ( .A(n2586), .B(n2585), .Z(n2613) );
  NAND U2734 ( .A(a[101]), .B(b[2]), .Z(n2587) );
  XNOR U2735 ( .A(n2588), .B(n2587), .Z(n2605) );
  NAND U2736 ( .A(b[1]), .B(a[102]), .Z(n2606) );
  XNOR U2737 ( .A(n2605), .B(n2606), .Z(n2611) );
  NAND U2738 ( .A(b[0]), .B(a[103]), .Z(n2612) );
  XOR U2739 ( .A(n2611), .B(n2612), .Z(n2614) );
  XOR U2740 ( .A(n2613), .B(n2614), .Z(n2599) );
  NANDN U2741 ( .A(n2590), .B(n2589), .Z(n2594) );
  OR U2742 ( .A(n2592), .B(n2591), .Z(n2593) );
  AND U2743 ( .A(n2594), .B(n2593), .Z(n2598) );
  XOR U2744 ( .A(n2599), .B(n2598), .Z(n2601) );
  XNOR U2745 ( .A(n2600), .B(n2601), .Z(n2618) );
  XNOR U2746 ( .A(sreg[227]), .B(n2617), .Z(n2597) );
  XNOR U2747 ( .A(n2618), .B(n2597), .Z(c[227]) );
  NANDN U2748 ( .A(n2599), .B(n2598), .Z(n2603) );
  OR U2749 ( .A(n2601), .B(n2600), .Z(n2602) );
  AND U2750 ( .A(n2603), .B(n2602), .Z(n2622) );
  AND U2751 ( .A(b[3]), .B(a[101]), .Z(n2610) );
  AND U2752 ( .A(b[2]), .B(a[100]), .Z(n2604) );
  NAND U2753 ( .A(n2610), .B(n2604), .Z(n2608) );
  NANDN U2754 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U2755 ( .A(n2608), .B(n2607), .Z(n2635) );
  NAND U2756 ( .A(a[102]), .B(b[2]), .Z(n2609) );
  XNOR U2757 ( .A(n2610), .B(n2609), .Z(n2627) );
  NAND U2758 ( .A(b[1]), .B(a[103]), .Z(n2628) );
  XNOR U2759 ( .A(n2627), .B(n2628), .Z(n2633) );
  NAND U2760 ( .A(b[0]), .B(a[104]), .Z(n2634) );
  XOR U2761 ( .A(n2633), .B(n2634), .Z(n2636) );
  XOR U2762 ( .A(n2635), .B(n2636), .Z(n2621) );
  NANDN U2763 ( .A(n2612), .B(n2611), .Z(n2616) );
  OR U2764 ( .A(n2614), .B(n2613), .Z(n2615) );
  AND U2765 ( .A(n2616), .B(n2615), .Z(n2620) );
  XOR U2766 ( .A(n2621), .B(n2620), .Z(n2623) );
  XNOR U2767 ( .A(n2622), .B(n2623), .Z(n2640) );
  XNOR U2768 ( .A(sreg[228]), .B(n2639), .Z(n2619) );
  XNOR U2769 ( .A(n2640), .B(n2619), .Z(c[228]) );
  NANDN U2770 ( .A(n2621), .B(n2620), .Z(n2625) );
  OR U2771 ( .A(n2623), .B(n2622), .Z(n2624) );
  AND U2772 ( .A(n2625), .B(n2624), .Z(n2644) );
  AND U2773 ( .A(b[3]), .B(a[102]), .Z(n2632) );
  AND U2774 ( .A(b[2]), .B(a[101]), .Z(n2626) );
  NAND U2775 ( .A(n2632), .B(n2626), .Z(n2630) );
  NANDN U2776 ( .A(n2628), .B(n2627), .Z(n2629) );
  AND U2777 ( .A(n2630), .B(n2629), .Z(n2657) );
  NAND U2778 ( .A(a[103]), .B(b[2]), .Z(n2631) );
  XNOR U2779 ( .A(n2632), .B(n2631), .Z(n2649) );
  NAND U2780 ( .A(b[1]), .B(a[104]), .Z(n2650) );
  XNOR U2781 ( .A(n2649), .B(n2650), .Z(n2655) );
  NAND U2782 ( .A(b[0]), .B(a[105]), .Z(n2656) );
  XOR U2783 ( .A(n2655), .B(n2656), .Z(n2658) );
  XOR U2784 ( .A(n2657), .B(n2658), .Z(n2643) );
  NANDN U2785 ( .A(n2634), .B(n2633), .Z(n2638) );
  OR U2786 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U2787 ( .A(n2638), .B(n2637), .Z(n2642) );
  XOR U2788 ( .A(n2643), .B(n2642), .Z(n2645) );
  XNOR U2789 ( .A(n2644), .B(n2645), .Z(n2662) );
  XNOR U2790 ( .A(sreg[229]), .B(n2661), .Z(n2641) );
  XNOR U2791 ( .A(n2662), .B(n2641), .Z(c[229]) );
  NANDN U2792 ( .A(n2643), .B(n2642), .Z(n2647) );
  OR U2793 ( .A(n2645), .B(n2644), .Z(n2646) );
  AND U2794 ( .A(n2647), .B(n2646), .Z(n2666) );
  AND U2795 ( .A(b[3]), .B(a[103]), .Z(n2654) );
  AND U2796 ( .A(b[2]), .B(a[102]), .Z(n2648) );
  NAND U2797 ( .A(n2654), .B(n2648), .Z(n2652) );
  NANDN U2798 ( .A(n2650), .B(n2649), .Z(n2651) );
  AND U2799 ( .A(n2652), .B(n2651), .Z(n2679) );
  NAND U2800 ( .A(a[104]), .B(b[2]), .Z(n2653) );
  XNOR U2801 ( .A(n2654), .B(n2653), .Z(n2671) );
  NAND U2802 ( .A(b[1]), .B(a[105]), .Z(n2672) );
  XNOR U2803 ( .A(n2671), .B(n2672), .Z(n2677) );
  NAND U2804 ( .A(b[0]), .B(a[106]), .Z(n2678) );
  XOR U2805 ( .A(n2677), .B(n2678), .Z(n2680) );
  XOR U2806 ( .A(n2679), .B(n2680), .Z(n2665) );
  NANDN U2807 ( .A(n2656), .B(n2655), .Z(n2660) );
  OR U2808 ( .A(n2658), .B(n2657), .Z(n2659) );
  AND U2809 ( .A(n2660), .B(n2659), .Z(n2664) );
  XOR U2810 ( .A(n2665), .B(n2664), .Z(n2667) );
  XNOR U2811 ( .A(n2666), .B(n2667), .Z(n2684) );
  XNOR U2812 ( .A(sreg[230]), .B(n2683), .Z(n2663) );
  XNOR U2813 ( .A(n2684), .B(n2663), .Z(c[230]) );
  NANDN U2814 ( .A(n2665), .B(n2664), .Z(n2669) );
  OR U2815 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U2816 ( .A(n2669), .B(n2668), .Z(n2688) );
  AND U2817 ( .A(b[3]), .B(a[104]), .Z(n2676) );
  AND U2818 ( .A(b[2]), .B(a[103]), .Z(n2670) );
  NAND U2819 ( .A(n2676), .B(n2670), .Z(n2674) );
  NANDN U2820 ( .A(n2672), .B(n2671), .Z(n2673) );
  AND U2821 ( .A(n2674), .B(n2673), .Z(n2701) );
  NAND U2822 ( .A(a[105]), .B(b[2]), .Z(n2675) );
  XNOR U2823 ( .A(n2676), .B(n2675), .Z(n2693) );
  NAND U2824 ( .A(b[1]), .B(a[106]), .Z(n2694) );
  XNOR U2825 ( .A(n2693), .B(n2694), .Z(n2699) );
  NAND U2826 ( .A(b[0]), .B(a[107]), .Z(n2700) );
  XOR U2827 ( .A(n2699), .B(n2700), .Z(n2702) );
  XOR U2828 ( .A(n2701), .B(n2702), .Z(n2687) );
  NANDN U2829 ( .A(n2678), .B(n2677), .Z(n2682) );
  OR U2830 ( .A(n2680), .B(n2679), .Z(n2681) );
  AND U2831 ( .A(n2682), .B(n2681), .Z(n2686) );
  XOR U2832 ( .A(n2687), .B(n2686), .Z(n2689) );
  XNOR U2833 ( .A(n2688), .B(n2689), .Z(n2706) );
  XNOR U2834 ( .A(sreg[231]), .B(n2705), .Z(n2685) );
  XNOR U2835 ( .A(n2706), .B(n2685), .Z(c[231]) );
  NANDN U2836 ( .A(n2687), .B(n2686), .Z(n2691) );
  OR U2837 ( .A(n2689), .B(n2688), .Z(n2690) );
  AND U2838 ( .A(n2691), .B(n2690), .Z(n2710) );
  AND U2839 ( .A(b[3]), .B(a[105]), .Z(n2698) );
  AND U2840 ( .A(b[2]), .B(a[104]), .Z(n2692) );
  NAND U2841 ( .A(n2698), .B(n2692), .Z(n2696) );
  NANDN U2842 ( .A(n2694), .B(n2693), .Z(n2695) );
  AND U2843 ( .A(n2696), .B(n2695), .Z(n2723) );
  NAND U2844 ( .A(a[106]), .B(b[2]), .Z(n2697) );
  XNOR U2845 ( .A(n2698), .B(n2697), .Z(n2715) );
  NAND U2846 ( .A(b[1]), .B(a[107]), .Z(n2716) );
  XNOR U2847 ( .A(n2715), .B(n2716), .Z(n2721) );
  NAND U2848 ( .A(b[0]), .B(a[108]), .Z(n2722) );
  XOR U2849 ( .A(n2721), .B(n2722), .Z(n2724) );
  XOR U2850 ( .A(n2723), .B(n2724), .Z(n2709) );
  NANDN U2851 ( .A(n2700), .B(n2699), .Z(n2704) );
  OR U2852 ( .A(n2702), .B(n2701), .Z(n2703) );
  AND U2853 ( .A(n2704), .B(n2703), .Z(n2708) );
  XOR U2854 ( .A(n2709), .B(n2708), .Z(n2711) );
  XNOR U2855 ( .A(n2710), .B(n2711), .Z(n2728) );
  XNOR U2856 ( .A(sreg[232]), .B(n2727), .Z(n2707) );
  XNOR U2857 ( .A(n2728), .B(n2707), .Z(c[232]) );
  NANDN U2858 ( .A(n2709), .B(n2708), .Z(n2713) );
  OR U2859 ( .A(n2711), .B(n2710), .Z(n2712) );
  AND U2860 ( .A(n2713), .B(n2712), .Z(n2732) );
  AND U2861 ( .A(b[3]), .B(a[106]), .Z(n2720) );
  AND U2862 ( .A(b[2]), .B(a[105]), .Z(n2714) );
  NAND U2863 ( .A(n2720), .B(n2714), .Z(n2718) );
  NANDN U2864 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U2865 ( .A(n2718), .B(n2717), .Z(n2745) );
  NAND U2866 ( .A(a[107]), .B(b[2]), .Z(n2719) );
  XNOR U2867 ( .A(n2720), .B(n2719), .Z(n2737) );
  NAND U2868 ( .A(b[1]), .B(a[108]), .Z(n2738) );
  XNOR U2869 ( .A(n2737), .B(n2738), .Z(n2743) );
  NAND U2870 ( .A(b[0]), .B(a[109]), .Z(n2744) );
  XOR U2871 ( .A(n2743), .B(n2744), .Z(n2746) );
  XOR U2872 ( .A(n2745), .B(n2746), .Z(n2731) );
  NANDN U2873 ( .A(n2722), .B(n2721), .Z(n2726) );
  OR U2874 ( .A(n2724), .B(n2723), .Z(n2725) );
  AND U2875 ( .A(n2726), .B(n2725), .Z(n2730) );
  XOR U2876 ( .A(n2731), .B(n2730), .Z(n2733) );
  XNOR U2877 ( .A(n2732), .B(n2733), .Z(n2750) );
  XNOR U2878 ( .A(sreg[233]), .B(n2749), .Z(n2729) );
  XNOR U2879 ( .A(n2750), .B(n2729), .Z(c[233]) );
  NANDN U2880 ( .A(n2731), .B(n2730), .Z(n2735) );
  OR U2881 ( .A(n2733), .B(n2732), .Z(n2734) );
  AND U2882 ( .A(n2735), .B(n2734), .Z(n2754) );
  AND U2883 ( .A(b[3]), .B(a[107]), .Z(n2742) );
  AND U2884 ( .A(b[2]), .B(a[106]), .Z(n2736) );
  NAND U2885 ( .A(n2742), .B(n2736), .Z(n2740) );
  NANDN U2886 ( .A(n2738), .B(n2737), .Z(n2739) );
  AND U2887 ( .A(n2740), .B(n2739), .Z(n2767) );
  NAND U2888 ( .A(a[108]), .B(b[2]), .Z(n2741) );
  XNOR U2889 ( .A(n2742), .B(n2741), .Z(n2759) );
  NAND U2890 ( .A(b[1]), .B(a[109]), .Z(n2760) );
  XNOR U2891 ( .A(n2759), .B(n2760), .Z(n2765) );
  NAND U2892 ( .A(b[0]), .B(a[110]), .Z(n2766) );
  XOR U2893 ( .A(n2765), .B(n2766), .Z(n2768) );
  XOR U2894 ( .A(n2767), .B(n2768), .Z(n2753) );
  NANDN U2895 ( .A(n2744), .B(n2743), .Z(n2748) );
  OR U2896 ( .A(n2746), .B(n2745), .Z(n2747) );
  AND U2897 ( .A(n2748), .B(n2747), .Z(n2752) );
  XOR U2898 ( .A(n2753), .B(n2752), .Z(n2755) );
  XNOR U2899 ( .A(n2754), .B(n2755), .Z(n2772) );
  XNOR U2900 ( .A(sreg[234]), .B(n2771), .Z(n2751) );
  XNOR U2901 ( .A(n2772), .B(n2751), .Z(c[234]) );
  NANDN U2902 ( .A(n2753), .B(n2752), .Z(n2757) );
  OR U2903 ( .A(n2755), .B(n2754), .Z(n2756) );
  AND U2904 ( .A(n2757), .B(n2756), .Z(n2776) );
  AND U2905 ( .A(b[3]), .B(a[108]), .Z(n2764) );
  AND U2906 ( .A(b[2]), .B(a[107]), .Z(n2758) );
  NAND U2907 ( .A(n2764), .B(n2758), .Z(n2762) );
  NANDN U2908 ( .A(n2760), .B(n2759), .Z(n2761) );
  AND U2909 ( .A(n2762), .B(n2761), .Z(n2789) );
  NAND U2910 ( .A(a[109]), .B(b[2]), .Z(n2763) );
  XNOR U2911 ( .A(n2764), .B(n2763), .Z(n2781) );
  NAND U2912 ( .A(b[1]), .B(a[110]), .Z(n2782) );
  XNOR U2913 ( .A(n2781), .B(n2782), .Z(n2787) );
  NAND U2914 ( .A(b[0]), .B(a[111]), .Z(n2788) );
  XOR U2915 ( .A(n2787), .B(n2788), .Z(n2790) );
  XOR U2916 ( .A(n2789), .B(n2790), .Z(n2775) );
  NANDN U2917 ( .A(n2766), .B(n2765), .Z(n2770) );
  OR U2918 ( .A(n2768), .B(n2767), .Z(n2769) );
  AND U2919 ( .A(n2770), .B(n2769), .Z(n2774) );
  XOR U2920 ( .A(n2775), .B(n2774), .Z(n2777) );
  XNOR U2921 ( .A(n2776), .B(n2777), .Z(n2794) );
  XNOR U2922 ( .A(sreg[235]), .B(n2793), .Z(n2773) );
  XNOR U2923 ( .A(n2794), .B(n2773), .Z(c[235]) );
  NANDN U2924 ( .A(n2775), .B(n2774), .Z(n2779) );
  OR U2925 ( .A(n2777), .B(n2776), .Z(n2778) );
  AND U2926 ( .A(n2779), .B(n2778), .Z(n2798) );
  AND U2927 ( .A(b[3]), .B(a[109]), .Z(n2786) );
  AND U2928 ( .A(b[2]), .B(a[108]), .Z(n2780) );
  NAND U2929 ( .A(n2786), .B(n2780), .Z(n2784) );
  NANDN U2930 ( .A(n2782), .B(n2781), .Z(n2783) );
  AND U2931 ( .A(n2784), .B(n2783), .Z(n2811) );
  NAND U2932 ( .A(a[110]), .B(b[2]), .Z(n2785) );
  XNOR U2933 ( .A(n2786), .B(n2785), .Z(n2803) );
  NAND U2934 ( .A(b[1]), .B(a[111]), .Z(n2804) );
  XNOR U2935 ( .A(n2803), .B(n2804), .Z(n2809) );
  NAND U2936 ( .A(b[0]), .B(a[112]), .Z(n2810) );
  XOR U2937 ( .A(n2809), .B(n2810), .Z(n2812) );
  XOR U2938 ( .A(n2811), .B(n2812), .Z(n2797) );
  NANDN U2939 ( .A(n2788), .B(n2787), .Z(n2792) );
  OR U2940 ( .A(n2790), .B(n2789), .Z(n2791) );
  AND U2941 ( .A(n2792), .B(n2791), .Z(n2796) );
  XOR U2942 ( .A(n2797), .B(n2796), .Z(n2799) );
  XNOR U2943 ( .A(n2798), .B(n2799), .Z(n2816) );
  XNOR U2944 ( .A(sreg[236]), .B(n2815), .Z(n2795) );
  XNOR U2945 ( .A(n2816), .B(n2795), .Z(c[236]) );
  NANDN U2946 ( .A(n2797), .B(n2796), .Z(n2801) );
  OR U2947 ( .A(n2799), .B(n2798), .Z(n2800) );
  AND U2948 ( .A(n2801), .B(n2800), .Z(n2820) );
  AND U2949 ( .A(b[3]), .B(a[110]), .Z(n2808) );
  AND U2950 ( .A(b[2]), .B(a[109]), .Z(n2802) );
  NAND U2951 ( .A(n2808), .B(n2802), .Z(n2806) );
  NANDN U2952 ( .A(n2804), .B(n2803), .Z(n2805) );
  AND U2953 ( .A(n2806), .B(n2805), .Z(n2833) );
  NAND U2954 ( .A(a[111]), .B(b[2]), .Z(n2807) );
  XNOR U2955 ( .A(n2808), .B(n2807), .Z(n2825) );
  NAND U2956 ( .A(b[1]), .B(a[112]), .Z(n2826) );
  XNOR U2957 ( .A(n2825), .B(n2826), .Z(n2831) );
  NAND U2958 ( .A(b[0]), .B(a[113]), .Z(n2832) );
  XOR U2959 ( .A(n2831), .B(n2832), .Z(n2834) );
  XOR U2960 ( .A(n2833), .B(n2834), .Z(n2819) );
  NANDN U2961 ( .A(n2810), .B(n2809), .Z(n2814) );
  OR U2962 ( .A(n2812), .B(n2811), .Z(n2813) );
  AND U2963 ( .A(n2814), .B(n2813), .Z(n2818) );
  XOR U2964 ( .A(n2819), .B(n2818), .Z(n2821) );
  XNOR U2965 ( .A(n2820), .B(n2821), .Z(n2838) );
  XNOR U2966 ( .A(sreg[237]), .B(n2837), .Z(n2817) );
  XNOR U2967 ( .A(n2838), .B(n2817), .Z(c[237]) );
  NANDN U2968 ( .A(n2819), .B(n2818), .Z(n2823) );
  OR U2969 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U2970 ( .A(n2823), .B(n2822), .Z(n2843) );
  AND U2971 ( .A(b[3]), .B(a[111]), .Z(n2830) );
  AND U2972 ( .A(b[2]), .B(a[110]), .Z(n2824) );
  NAND U2973 ( .A(n2830), .B(n2824), .Z(n2828) );
  NANDN U2974 ( .A(n2826), .B(n2825), .Z(n2827) );
  AND U2975 ( .A(n2828), .B(n2827), .Z(n2855) );
  NAND U2976 ( .A(a[112]), .B(b[2]), .Z(n2829) );
  XNOR U2977 ( .A(n2830), .B(n2829), .Z(n2847) );
  NAND U2978 ( .A(b[1]), .B(a[113]), .Z(n2848) );
  XNOR U2979 ( .A(n2847), .B(n2848), .Z(n2853) );
  NAND U2980 ( .A(b[0]), .B(a[114]), .Z(n2854) );
  XOR U2981 ( .A(n2853), .B(n2854), .Z(n2856) );
  XOR U2982 ( .A(n2855), .B(n2856), .Z(n2841) );
  NANDN U2983 ( .A(n2832), .B(n2831), .Z(n2836) );
  OR U2984 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U2985 ( .A(n2836), .B(n2835), .Z(n2840) );
  XNOR U2986 ( .A(n2841), .B(n2840), .Z(n2842) );
  XNOR U2987 ( .A(n2843), .B(n2842), .Z(n2860) );
  XOR U2988 ( .A(n2859), .B(sreg[238]), .Z(n2839) );
  XNOR U2989 ( .A(n2860), .B(n2839), .Z(c[238]) );
  NANDN U2990 ( .A(n2841), .B(n2840), .Z(n2845) );
  NANDN U2991 ( .A(n2843), .B(n2842), .Z(n2844) );
  AND U2992 ( .A(n2845), .B(n2844), .Z(n2864) );
  AND U2993 ( .A(b[3]), .B(a[112]), .Z(n2852) );
  AND U2994 ( .A(b[2]), .B(a[111]), .Z(n2846) );
  NAND U2995 ( .A(n2852), .B(n2846), .Z(n2850) );
  NANDN U2996 ( .A(n2848), .B(n2847), .Z(n2849) );
  AND U2997 ( .A(n2850), .B(n2849), .Z(n2877) );
  NAND U2998 ( .A(a[113]), .B(b[2]), .Z(n2851) );
  XNOR U2999 ( .A(n2852), .B(n2851), .Z(n2869) );
  NAND U3000 ( .A(b[1]), .B(a[114]), .Z(n2870) );
  XNOR U3001 ( .A(n2869), .B(n2870), .Z(n2875) );
  NAND U3002 ( .A(b[0]), .B(a[115]), .Z(n2876) );
  XOR U3003 ( .A(n2875), .B(n2876), .Z(n2878) );
  XOR U3004 ( .A(n2877), .B(n2878), .Z(n2863) );
  NANDN U3005 ( .A(n2854), .B(n2853), .Z(n2858) );
  OR U3006 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U3007 ( .A(n2858), .B(n2857), .Z(n2862) );
  XOR U3008 ( .A(n2863), .B(n2862), .Z(n2865) );
  XNOR U3009 ( .A(n2864), .B(n2865), .Z(n2882) );
  XOR U3010 ( .A(sreg[239]), .B(n2881), .Z(n2861) );
  XNOR U3011 ( .A(n2882), .B(n2861), .Z(c[239]) );
  NANDN U3012 ( .A(n2863), .B(n2862), .Z(n2867) );
  OR U3013 ( .A(n2865), .B(n2864), .Z(n2866) );
  AND U3014 ( .A(n2867), .B(n2866), .Z(n2886) );
  AND U3015 ( .A(b[3]), .B(a[113]), .Z(n2874) );
  AND U3016 ( .A(b[2]), .B(a[112]), .Z(n2868) );
  NAND U3017 ( .A(n2874), .B(n2868), .Z(n2872) );
  NANDN U3018 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3019 ( .A(n2872), .B(n2871), .Z(n2899) );
  NAND U3020 ( .A(a[114]), .B(b[2]), .Z(n2873) );
  XNOR U3021 ( .A(n2874), .B(n2873), .Z(n2891) );
  NAND U3022 ( .A(b[1]), .B(a[115]), .Z(n2892) );
  XNOR U3023 ( .A(n2891), .B(n2892), .Z(n2897) );
  NAND U3024 ( .A(b[0]), .B(a[116]), .Z(n2898) );
  XOR U3025 ( .A(n2897), .B(n2898), .Z(n2900) );
  XOR U3026 ( .A(n2899), .B(n2900), .Z(n2885) );
  NANDN U3027 ( .A(n2876), .B(n2875), .Z(n2880) );
  OR U3028 ( .A(n2878), .B(n2877), .Z(n2879) );
  AND U3029 ( .A(n2880), .B(n2879), .Z(n2884) );
  XOR U3030 ( .A(n2885), .B(n2884), .Z(n2887) );
  XNOR U3031 ( .A(n2886), .B(n2887), .Z(n2904) );
  XNOR U3032 ( .A(sreg[240]), .B(n2903), .Z(n2883) );
  XNOR U3033 ( .A(n2904), .B(n2883), .Z(c[240]) );
  NANDN U3034 ( .A(n2885), .B(n2884), .Z(n2889) );
  OR U3035 ( .A(n2887), .B(n2886), .Z(n2888) );
  AND U3036 ( .A(n2889), .B(n2888), .Z(n2908) );
  AND U3037 ( .A(b[3]), .B(a[114]), .Z(n2896) );
  AND U3038 ( .A(b[2]), .B(a[113]), .Z(n2890) );
  NAND U3039 ( .A(n2896), .B(n2890), .Z(n2894) );
  NANDN U3040 ( .A(n2892), .B(n2891), .Z(n2893) );
  AND U3041 ( .A(n2894), .B(n2893), .Z(n2921) );
  NAND U3042 ( .A(a[115]), .B(b[2]), .Z(n2895) );
  XNOR U3043 ( .A(n2896), .B(n2895), .Z(n2913) );
  NAND U3044 ( .A(b[1]), .B(a[116]), .Z(n2914) );
  XNOR U3045 ( .A(n2913), .B(n2914), .Z(n2919) );
  NAND U3046 ( .A(b[0]), .B(a[117]), .Z(n2920) );
  XOR U3047 ( .A(n2919), .B(n2920), .Z(n2922) );
  XOR U3048 ( .A(n2921), .B(n2922), .Z(n2907) );
  NANDN U3049 ( .A(n2898), .B(n2897), .Z(n2902) );
  OR U3050 ( .A(n2900), .B(n2899), .Z(n2901) );
  AND U3051 ( .A(n2902), .B(n2901), .Z(n2906) );
  XOR U3052 ( .A(n2907), .B(n2906), .Z(n2909) );
  XNOR U3053 ( .A(n2908), .B(n2909), .Z(n2926) );
  XNOR U3054 ( .A(sreg[241]), .B(n2925), .Z(n2905) );
  XNOR U3055 ( .A(n2926), .B(n2905), .Z(c[241]) );
  NANDN U3056 ( .A(n2907), .B(n2906), .Z(n2911) );
  OR U3057 ( .A(n2909), .B(n2908), .Z(n2910) );
  AND U3058 ( .A(n2911), .B(n2910), .Z(n2930) );
  AND U3059 ( .A(b[3]), .B(a[115]), .Z(n2918) );
  AND U3060 ( .A(b[2]), .B(a[114]), .Z(n2912) );
  NAND U3061 ( .A(n2918), .B(n2912), .Z(n2916) );
  NANDN U3062 ( .A(n2914), .B(n2913), .Z(n2915) );
  AND U3063 ( .A(n2916), .B(n2915), .Z(n2943) );
  NAND U3064 ( .A(a[116]), .B(b[2]), .Z(n2917) );
  XNOR U3065 ( .A(n2918), .B(n2917), .Z(n2935) );
  NAND U3066 ( .A(b[1]), .B(a[117]), .Z(n2936) );
  XNOR U3067 ( .A(n2935), .B(n2936), .Z(n2941) );
  NAND U3068 ( .A(b[0]), .B(a[118]), .Z(n2942) );
  XOR U3069 ( .A(n2941), .B(n2942), .Z(n2944) );
  XOR U3070 ( .A(n2943), .B(n2944), .Z(n2929) );
  NANDN U3071 ( .A(n2920), .B(n2919), .Z(n2924) );
  OR U3072 ( .A(n2922), .B(n2921), .Z(n2923) );
  AND U3073 ( .A(n2924), .B(n2923), .Z(n2928) );
  XOR U3074 ( .A(n2929), .B(n2928), .Z(n2931) );
  XNOR U3075 ( .A(n2930), .B(n2931), .Z(n2948) );
  XNOR U3076 ( .A(sreg[242]), .B(n2947), .Z(n2927) );
  XNOR U3077 ( .A(n2948), .B(n2927), .Z(c[242]) );
  NANDN U3078 ( .A(n2929), .B(n2928), .Z(n2933) );
  OR U3079 ( .A(n2931), .B(n2930), .Z(n2932) );
  AND U3080 ( .A(n2933), .B(n2932), .Z(n2953) );
  AND U3081 ( .A(b[3]), .B(a[116]), .Z(n2940) );
  AND U3082 ( .A(b[2]), .B(a[115]), .Z(n2934) );
  NAND U3083 ( .A(n2940), .B(n2934), .Z(n2938) );
  NANDN U3084 ( .A(n2936), .B(n2935), .Z(n2937) );
  AND U3085 ( .A(n2938), .B(n2937), .Z(n2965) );
  NAND U3086 ( .A(a[117]), .B(b[2]), .Z(n2939) );
  XNOR U3087 ( .A(n2940), .B(n2939), .Z(n2957) );
  NAND U3088 ( .A(b[1]), .B(a[118]), .Z(n2958) );
  XNOR U3089 ( .A(n2957), .B(n2958), .Z(n2963) );
  NAND U3090 ( .A(b[0]), .B(a[119]), .Z(n2964) );
  XOR U3091 ( .A(n2963), .B(n2964), .Z(n2966) );
  XOR U3092 ( .A(n2965), .B(n2966), .Z(n2951) );
  NANDN U3093 ( .A(n2942), .B(n2941), .Z(n2946) );
  OR U3094 ( .A(n2944), .B(n2943), .Z(n2945) );
  AND U3095 ( .A(n2946), .B(n2945), .Z(n2950) );
  XNOR U3096 ( .A(n2951), .B(n2950), .Z(n2952) );
  XNOR U3097 ( .A(n2953), .B(n2952), .Z(n2970) );
  XOR U3098 ( .A(n2969), .B(sreg[243]), .Z(n2949) );
  XNOR U3099 ( .A(n2970), .B(n2949), .Z(c[243]) );
  NANDN U3100 ( .A(n2951), .B(n2950), .Z(n2955) );
  NANDN U3101 ( .A(n2953), .B(n2952), .Z(n2954) );
  AND U3102 ( .A(n2955), .B(n2954), .Z(n2974) );
  AND U3103 ( .A(b[3]), .B(a[117]), .Z(n2962) );
  AND U3104 ( .A(b[2]), .B(a[116]), .Z(n2956) );
  NAND U3105 ( .A(n2962), .B(n2956), .Z(n2960) );
  NANDN U3106 ( .A(n2958), .B(n2957), .Z(n2959) );
  AND U3107 ( .A(n2960), .B(n2959), .Z(n2987) );
  NAND U3108 ( .A(a[118]), .B(b[2]), .Z(n2961) );
  XNOR U3109 ( .A(n2962), .B(n2961), .Z(n2979) );
  NAND U3110 ( .A(b[1]), .B(a[119]), .Z(n2980) );
  XNOR U3111 ( .A(n2979), .B(n2980), .Z(n2985) );
  NAND U3112 ( .A(b[0]), .B(a[120]), .Z(n2986) );
  XOR U3113 ( .A(n2985), .B(n2986), .Z(n2988) );
  XOR U3114 ( .A(n2987), .B(n2988), .Z(n2973) );
  NANDN U3115 ( .A(n2964), .B(n2963), .Z(n2968) );
  OR U3116 ( .A(n2966), .B(n2965), .Z(n2967) );
  AND U3117 ( .A(n2968), .B(n2967), .Z(n2972) );
  XOR U3118 ( .A(n2973), .B(n2972), .Z(n2975) );
  XNOR U3119 ( .A(n2974), .B(n2975), .Z(n2992) );
  XOR U3120 ( .A(sreg[244]), .B(n2991), .Z(n2971) );
  XNOR U3121 ( .A(n2992), .B(n2971), .Z(c[244]) );
  NANDN U3122 ( .A(n2973), .B(n2972), .Z(n2977) );
  OR U3123 ( .A(n2975), .B(n2974), .Z(n2976) );
  AND U3124 ( .A(n2977), .B(n2976), .Z(n2997) );
  AND U3125 ( .A(b[3]), .B(a[118]), .Z(n2984) );
  AND U3126 ( .A(b[2]), .B(a[117]), .Z(n2978) );
  NAND U3127 ( .A(n2984), .B(n2978), .Z(n2982) );
  NANDN U3128 ( .A(n2980), .B(n2979), .Z(n2981) );
  AND U3129 ( .A(n2982), .B(n2981), .Z(n3009) );
  NAND U3130 ( .A(a[119]), .B(b[2]), .Z(n2983) );
  XNOR U3131 ( .A(n2984), .B(n2983), .Z(n3001) );
  NAND U3132 ( .A(b[1]), .B(a[120]), .Z(n3002) );
  XNOR U3133 ( .A(n3001), .B(n3002), .Z(n3007) );
  NAND U3134 ( .A(b[0]), .B(a[121]), .Z(n3008) );
  XOR U3135 ( .A(n3007), .B(n3008), .Z(n3010) );
  XOR U3136 ( .A(n3009), .B(n3010), .Z(n2995) );
  NANDN U3137 ( .A(n2986), .B(n2985), .Z(n2990) );
  OR U3138 ( .A(n2988), .B(n2987), .Z(n2989) );
  AND U3139 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U3140 ( .A(n2995), .B(n2994), .Z(n2996) );
  XNOR U3141 ( .A(n2997), .B(n2996), .Z(n3014) );
  XOR U3142 ( .A(n3013), .B(sreg[245]), .Z(n2993) );
  XNOR U3143 ( .A(n3014), .B(n2993), .Z(c[245]) );
  NANDN U3144 ( .A(n2995), .B(n2994), .Z(n2999) );
  NANDN U3145 ( .A(n2997), .B(n2996), .Z(n2998) );
  AND U3146 ( .A(n2999), .B(n2998), .Z(n3018) );
  AND U3147 ( .A(b[3]), .B(a[119]), .Z(n3006) );
  AND U3148 ( .A(b[2]), .B(a[118]), .Z(n3000) );
  NAND U3149 ( .A(n3006), .B(n3000), .Z(n3004) );
  NANDN U3150 ( .A(n3002), .B(n3001), .Z(n3003) );
  AND U3151 ( .A(n3004), .B(n3003), .Z(n3031) );
  NAND U3152 ( .A(a[120]), .B(b[2]), .Z(n3005) );
  XNOR U3153 ( .A(n3006), .B(n3005), .Z(n3023) );
  NAND U3154 ( .A(b[1]), .B(a[121]), .Z(n3024) );
  XNOR U3155 ( .A(n3023), .B(n3024), .Z(n3029) );
  NAND U3156 ( .A(b[0]), .B(a[122]), .Z(n3030) );
  XOR U3157 ( .A(n3029), .B(n3030), .Z(n3032) );
  XOR U3158 ( .A(n3031), .B(n3032), .Z(n3017) );
  NANDN U3159 ( .A(n3008), .B(n3007), .Z(n3012) );
  OR U3160 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U3161 ( .A(n3012), .B(n3011), .Z(n3016) );
  XOR U3162 ( .A(n3017), .B(n3016), .Z(n3019) );
  XNOR U3163 ( .A(n3018), .B(n3019), .Z(n3036) );
  XOR U3164 ( .A(sreg[246]), .B(n3035), .Z(n3015) );
  XNOR U3165 ( .A(n3036), .B(n3015), .Z(c[246]) );
  NANDN U3166 ( .A(n3017), .B(n3016), .Z(n3021) );
  OR U3167 ( .A(n3019), .B(n3018), .Z(n3020) );
  AND U3168 ( .A(n3021), .B(n3020), .Z(n3040) );
  AND U3169 ( .A(b[3]), .B(a[120]), .Z(n3028) );
  AND U3170 ( .A(b[2]), .B(a[119]), .Z(n3022) );
  NAND U3171 ( .A(n3028), .B(n3022), .Z(n3026) );
  NANDN U3172 ( .A(n3024), .B(n3023), .Z(n3025) );
  AND U3173 ( .A(n3026), .B(n3025), .Z(n3053) );
  NAND U3174 ( .A(a[121]), .B(b[2]), .Z(n3027) );
  XNOR U3175 ( .A(n3028), .B(n3027), .Z(n3045) );
  NAND U3176 ( .A(b[1]), .B(a[122]), .Z(n3046) );
  XNOR U3177 ( .A(n3045), .B(n3046), .Z(n3051) );
  NAND U3178 ( .A(b[0]), .B(a[123]), .Z(n3052) );
  XOR U3179 ( .A(n3051), .B(n3052), .Z(n3054) );
  XOR U3180 ( .A(n3053), .B(n3054), .Z(n3039) );
  NANDN U3181 ( .A(n3030), .B(n3029), .Z(n3034) );
  OR U3182 ( .A(n3032), .B(n3031), .Z(n3033) );
  AND U3183 ( .A(n3034), .B(n3033), .Z(n3038) );
  XOR U3184 ( .A(n3039), .B(n3038), .Z(n3041) );
  XNOR U3185 ( .A(n3040), .B(n3041), .Z(n3058) );
  XNOR U3186 ( .A(sreg[247]), .B(n3057), .Z(n3037) );
  XNOR U3187 ( .A(n3058), .B(n3037), .Z(c[247]) );
  NANDN U3188 ( .A(n3039), .B(n3038), .Z(n3043) );
  OR U3189 ( .A(n3041), .B(n3040), .Z(n3042) );
  AND U3190 ( .A(n3043), .B(n3042), .Z(n3062) );
  AND U3191 ( .A(b[3]), .B(a[121]), .Z(n3050) );
  AND U3192 ( .A(b[2]), .B(a[120]), .Z(n3044) );
  NAND U3193 ( .A(n3050), .B(n3044), .Z(n3048) );
  NANDN U3194 ( .A(n3046), .B(n3045), .Z(n3047) );
  AND U3195 ( .A(n3048), .B(n3047), .Z(n3075) );
  NAND U3196 ( .A(a[122]), .B(b[2]), .Z(n3049) );
  XNOR U3197 ( .A(n3050), .B(n3049), .Z(n3067) );
  NAND U3198 ( .A(b[1]), .B(a[123]), .Z(n3068) );
  XNOR U3199 ( .A(n3067), .B(n3068), .Z(n3073) );
  NAND U3200 ( .A(a[124]), .B(b[0]), .Z(n3074) );
  XOR U3201 ( .A(n3073), .B(n3074), .Z(n3076) );
  XOR U3202 ( .A(n3075), .B(n3076), .Z(n3061) );
  NANDN U3203 ( .A(n3052), .B(n3051), .Z(n3056) );
  OR U3204 ( .A(n3054), .B(n3053), .Z(n3055) );
  AND U3205 ( .A(n3056), .B(n3055), .Z(n3060) );
  XOR U3206 ( .A(n3061), .B(n3060), .Z(n3063) );
  XNOR U3207 ( .A(n3062), .B(n3063), .Z(n3080) );
  XNOR U3208 ( .A(sreg[248]), .B(n3079), .Z(n3059) );
  XNOR U3209 ( .A(n3080), .B(n3059), .Z(c[248]) );
  NANDN U3210 ( .A(n3061), .B(n3060), .Z(n3065) );
  OR U3211 ( .A(n3063), .B(n3062), .Z(n3064) );
  AND U3212 ( .A(n3065), .B(n3064), .Z(n3084) );
  AND U3213 ( .A(b[3]), .B(a[122]), .Z(n3072) );
  AND U3214 ( .A(b[2]), .B(a[121]), .Z(n3066) );
  NAND U3215 ( .A(n3072), .B(n3066), .Z(n3070) );
  NANDN U3216 ( .A(n3068), .B(n3067), .Z(n3069) );
  AND U3217 ( .A(n3070), .B(n3069), .Z(n3097) );
  NAND U3218 ( .A(a[123]), .B(b[2]), .Z(n3071) );
  XNOR U3219 ( .A(n3072), .B(n3071), .Z(n3089) );
  NAND U3220 ( .A(b[1]), .B(a[124]), .Z(n3090) );
  XNOR U3221 ( .A(n3089), .B(n3090), .Z(n3095) );
  NAND U3222 ( .A(a[125]), .B(b[0]), .Z(n3096) );
  XOR U3223 ( .A(n3095), .B(n3096), .Z(n3098) );
  XOR U3224 ( .A(n3097), .B(n3098), .Z(n3083) );
  NANDN U3225 ( .A(n3074), .B(n3073), .Z(n3078) );
  OR U3226 ( .A(n3076), .B(n3075), .Z(n3077) );
  AND U3227 ( .A(n3078), .B(n3077), .Z(n3082) );
  XOR U3228 ( .A(n3083), .B(n3082), .Z(n3085) );
  XNOR U3229 ( .A(n3084), .B(n3085), .Z(n3102) );
  XNOR U3230 ( .A(sreg[249]), .B(n3101), .Z(n3081) );
  XNOR U3231 ( .A(n3102), .B(n3081), .Z(c[249]) );
  NANDN U3232 ( .A(n3083), .B(n3082), .Z(n3087) );
  OR U3233 ( .A(n3085), .B(n3084), .Z(n3086) );
  AND U3234 ( .A(n3087), .B(n3086), .Z(n3106) );
  AND U3235 ( .A(b[3]), .B(a[123]), .Z(n3094) );
  AND U3236 ( .A(b[2]), .B(a[122]), .Z(n3088) );
  NAND U3237 ( .A(n3094), .B(n3088), .Z(n3092) );
  NANDN U3238 ( .A(n3090), .B(n3089), .Z(n3091) );
  AND U3239 ( .A(n3092), .B(n3091), .Z(n3119) );
  NAND U3240 ( .A(a[124]), .B(b[2]), .Z(n3093) );
  XNOR U3241 ( .A(n3094), .B(n3093), .Z(n3111) );
  NAND U3242 ( .A(b[1]), .B(a[125]), .Z(n3112) );
  XNOR U3243 ( .A(n3111), .B(n3112), .Z(n3117) );
  NAND U3244 ( .A(a[126]), .B(b[0]), .Z(n3118) );
  XOR U3245 ( .A(n3117), .B(n3118), .Z(n3120) );
  XOR U3246 ( .A(n3119), .B(n3120), .Z(n3105) );
  NANDN U3247 ( .A(n3096), .B(n3095), .Z(n3100) );
  OR U3248 ( .A(n3098), .B(n3097), .Z(n3099) );
  AND U3249 ( .A(n3100), .B(n3099), .Z(n3104) );
  XOR U3250 ( .A(n3105), .B(n3104), .Z(n3107) );
  XNOR U3251 ( .A(n3106), .B(n3107), .Z(n3124) );
  XNOR U3252 ( .A(sreg[250]), .B(n3123), .Z(n3103) );
  XNOR U3253 ( .A(n3124), .B(n3103), .Z(c[250]) );
  NANDN U3254 ( .A(n3105), .B(n3104), .Z(n3109) );
  OR U3255 ( .A(n3107), .B(n3106), .Z(n3108) );
  AND U3256 ( .A(n3109), .B(n3108), .Z(n3130) );
  AND U3257 ( .A(b[3]), .B(a[124]), .Z(n3116) );
  AND U3258 ( .A(b[2]), .B(a[123]), .Z(n3110) );
  NAND U3259 ( .A(n3116), .B(n3110), .Z(n3114) );
  NANDN U3260 ( .A(n3112), .B(n3111), .Z(n3113) );
  AND U3261 ( .A(n3114), .B(n3113), .Z(n3142) );
  NAND U3262 ( .A(a[126]), .B(b[1]), .Z(n3159) );
  NAND U3263 ( .A(a[125]), .B(b[2]), .Z(n3115) );
  XOR U3264 ( .A(n3116), .B(n3115), .Z(n3135) );
  XOR U3265 ( .A(n3159), .B(n3135), .Z(n3140) );
  NAND U3266 ( .A(a[127]), .B(b[0]), .Z(n3141) );
  XOR U3267 ( .A(n3140), .B(n3141), .Z(n3143) );
  XOR U3268 ( .A(n3142), .B(n3143), .Z(n3129) );
  NANDN U3269 ( .A(n3118), .B(n3117), .Z(n3122) );
  OR U3270 ( .A(n3120), .B(n3119), .Z(n3121) );
  AND U3271 ( .A(n3122), .B(n3121), .Z(n3128) );
  XOR U3272 ( .A(n3129), .B(n3128), .Z(n3131) );
  XNOR U3273 ( .A(n3130), .B(n3131), .Z(n3127) );
  XNOR U3274 ( .A(sreg[251]), .B(n3126), .Z(n3125) );
  XNOR U3275 ( .A(n3127), .B(n3125), .Z(c[251]) );
  NANDN U3276 ( .A(n3129), .B(n3128), .Z(n3133) );
  OR U3277 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U3278 ( .A(n3133), .B(n3132), .Z(n3151) );
  AND U3279 ( .A(b[3]), .B(a[125]), .Z(n3154) );
  AND U3280 ( .A(b[2]), .B(a[124]), .Z(n3134) );
  NAND U3281 ( .A(n3154), .B(n3134), .Z(n3137) );
  IV U3282 ( .A(n3159), .Z(n3152) );
  NANDN U3283 ( .A(n3135), .B(n3152), .Z(n3136) );
  AND U3284 ( .A(n3137), .B(n3136), .Z(n3156) );
  AND U3285 ( .A(a[126]), .B(b[2]), .Z(n3139) );
  NAND U3286 ( .A(b[1]), .B(a[127]), .Z(n3138) );
  XNOR U3287 ( .A(n3139), .B(n3138), .Z(n3153) );
  XOR U3288 ( .A(n3153), .B(n3154), .Z(n3155) );
  XOR U3289 ( .A(n3156), .B(n3155), .Z(n3148) );
  NANDN U3290 ( .A(n3141), .B(n3140), .Z(n3145) );
  OR U3291 ( .A(n3143), .B(n3142), .Z(n3144) );
  AND U3292 ( .A(n3145), .B(n3144), .Z(n3149) );
  XOR U3293 ( .A(n3148), .B(n3149), .Z(n3150) );
  XOR U3294 ( .A(n3151), .B(n3150), .Z(n3146) );
  XOR U3295 ( .A(n3147), .B(n3146), .Z(c[252]) );
  AND U3296 ( .A(n3147), .B(n3146), .Z(n3168) );
  NAND U3297 ( .A(b[3]), .B(a[126]), .Z(n3160) );
  AND U3298 ( .A(a[127]), .B(b[2]), .Z(n3162) );
  NAND U3299 ( .A(n3154), .B(n3153), .Z(n3158) );
  NANDN U3300 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U3301 ( .A(n3158), .B(n3157), .Z(n3164) );
  XOR U3302 ( .A(n3163), .B(n3164), .Z(n3165) );
  XOR U3303 ( .A(n3166), .B(n3165), .Z(n3167) );
  XOR U3304 ( .A(n3168), .B(n3167), .Z(c[253]) );
  NAND U3305 ( .A(n3160), .B(n3159), .Z(n3161) );
  AND U3306 ( .A(n3162), .B(n3161), .Z(n3174) );
  AND U3307 ( .A(a[127]), .B(b[3]), .Z(n3171) );
  XNOR U3308 ( .A(n3171), .B(n3170), .Z(n3175) );
  XNOR U3309 ( .A(n3174), .B(n3175), .Z(n3169) );
  AND U3310 ( .A(n3168), .B(n3167), .Z(n3177) );
  XNOR U3311 ( .A(n3169), .B(n3177), .Z(c[254]) );
  NANDN U3312 ( .A(n3171), .B(n3170), .Z(n3173) );
  NANDN U3313 ( .A(n3174), .B(n3175), .Z(n3172) );
  NAND U3314 ( .A(n3173), .B(n3172), .Z(n3179) );
  XOR U3315 ( .A(n3175), .B(n3174), .Z(n3176) );
  NAND U3316 ( .A(n3177), .B(n3176), .Z(n3178) );
  NAND U3317 ( .A(n3179), .B(n3178), .Z(c[255]) );
endmodule

