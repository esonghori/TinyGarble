
module compare_N16384_CC16 ( clk, rst, x, y, g, e );
  input [1023:0] x;
  input [1023:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  NAND U10 ( .A(n7035), .B(n7036), .Z(n8) );
  NAND U11 ( .A(n7037), .B(n8), .Z(n9) );
  ANDN U12 ( .B(n9), .A(n7038), .Z(n10) );
  NANDN U13 ( .A(n10), .B(n7039), .Z(n11) );
  NANDN U14 ( .A(n7040), .B(n11), .Z(n12) );
  NAND U15 ( .A(n7041), .B(n12), .Z(n13) );
  ANDN U16 ( .B(n5424), .A(n5423), .Z(n14) );
  NAND U17 ( .A(n13), .B(n14), .Z(n15) );
  NAND U18 ( .A(n7042), .B(n15), .Z(n16) );
  NANDN U19 ( .A(n5422), .B(n16), .Z(n17) );
  NAND U20 ( .A(n7043), .B(n17), .Z(n18) );
  ANDN U21 ( .B(n18), .A(n7044), .Z(n19) );
  AND U22 ( .A(n7046), .B(n7047), .Z(n20) );
  NANDN U23 ( .A(n19), .B(n7045), .Z(n21) );
  AND U24 ( .A(n20), .B(n21), .Z(n22) );
  NANDN U25 ( .A(n22), .B(n7048), .Z(n23) );
  NAND U26 ( .A(n7049), .B(n23), .Z(n24) );
  NANDN U27 ( .A(n7050), .B(n24), .Z(n7051) );
  NANDN U28 ( .A(y[850]), .B(x[850]), .Z(n25) );
  NANDN U29 ( .A(y[849]), .B(x[849]), .Z(n26) );
  AND U30 ( .A(n25), .B(n26), .Z(n27) );
  NANDN U31 ( .A(n27), .B(n239), .Z(n28) );
  NANDN U32 ( .A(y[851]), .B(x[851]), .Z(n29) );
  AND U33 ( .A(n28), .B(n29), .Z(n5058) );
  ANDN U34 ( .B(n1702), .A(n1701), .Z(n7116) );
  NANDN U35 ( .A(n1684), .B(n1685), .Z(n7148) );
  NANDN U36 ( .A(n7204), .B(n7205), .Z(n30) );
  NANDN U37 ( .A(n7207), .B(n30), .Z(n31) );
  AND U38 ( .A(n7208), .B(n31), .Z(n32) );
  OR U39 ( .A(n7209), .B(n32), .Z(n33) );
  NAND U40 ( .A(n7210), .B(n33), .Z(n34) );
  NANDN U41 ( .A(n7211), .B(n34), .Z(n35) );
  NAND U42 ( .A(n7212), .B(n35), .Z(n36) );
  NAND U43 ( .A(n7213), .B(n36), .Z(n37) );
  ANDN U44 ( .B(n37), .A(n7214), .Z(n38) );
  NANDN U45 ( .A(n38), .B(n7215), .Z(n39) );
  NANDN U46 ( .A(n7216), .B(n39), .Z(n40) );
  NAND U47 ( .A(n7217), .B(n40), .Z(n41) );
  NAND U48 ( .A(n7218), .B(n41), .Z(n42) );
  NANDN U49 ( .A(n7219), .B(n42), .Z(n43) );
  AND U50 ( .A(n7220), .B(n43), .Z(n44) );
  NANDN U51 ( .A(n44), .B(n7221), .Z(n45) );
  NAND U52 ( .A(n7222), .B(n45), .Z(n46) );
  NAND U53 ( .A(n7223), .B(n46), .Z(n47) );
  AND U54 ( .A(n7224), .B(n47), .Z(n7226) );
  OR U55 ( .A(n7270), .B(n7271), .Z(n48) );
  NAND U56 ( .A(n7272), .B(n48), .Z(n49) );
  NAND U57 ( .A(n7273), .B(n49), .Z(n50) );
  NAND U58 ( .A(n7274), .B(n50), .Z(n51) );
  NAND U59 ( .A(n7275), .B(n51), .Z(n52) );
  AND U60 ( .A(n7276), .B(n52), .Z(n53) );
  OR U61 ( .A(n5397), .B(n53), .Z(n54) );
  NAND U62 ( .A(n5396), .B(n54), .Z(n55) );
  NANDN U63 ( .A(n7277), .B(n55), .Z(n56) );
  NAND U64 ( .A(n7278), .B(n56), .Z(n57) );
  NANDN U65 ( .A(n7279), .B(n57), .Z(n58) );
  ANDN U66 ( .B(n58), .A(n7280), .Z(n59) );
  NANDN U67 ( .A(n59), .B(n7281), .Z(n60) );
  AND U68 ( .A(n7282), .B(n60), .Z(n61) );
  NAND U69 ( .A(n7283), .B(n61), .Z(n62) );
  NAND U70 ( .A(n7284), .B(n62), .Z(n63) );
  NANDN U71 ( .A(n5395), .B(n63), .Z(n7285) );
  XNOR U72 ( .A(x[1007]), .B(y[1007]), .Z(n64) );
  NANDN U73 ( .A(n5370), .B(n64), .Z(n65) );
  NAND U74 ( .A(n5371), .B(n65), .Z(n5390) );
  NAND U75 ( .A(n7052), .B(n7051), .Z(n66) );
  NANDN U76 ( .A(n7053), .B(n66), .Z(n67) );
  NAND U77 ( .A(n7054), .B(n67), .Z(n68) );
  NANDN U78 ( .A(n7055), .B(n68), .Z(n69) );
  NAND U79 ( .A(n7056), .B(n69), .Z(n70) );
  ANDN U80 ( .B(n70), .A(n7057), .Z(n71) );
  NANDN U81 ( .A(n71), .B(n7058), .Z(n72) );
  NAND U82 ( .A(n7059), .B(n72), .Z(n73) );
  NAND U83 ( .A(n7060), .B(n73), .Z(n74) );
  NANDN U84 ( .A(n7061), .B(n74), .Z(n75) );
  NAND U85 ( .A(n7062), .B(n75), .Z(n76) );
  ANDN U86 ( .B(n76), .A(n7063), .Z(n77) );
  NOR U87 ( .A(n7065), .B(n7064), .Z(n78) );
  OR U88 ( .A(n5421), .B(n77), .Z(n79) );
  AND U89 ( .A(n78), .B(n79), .Z(n80) );
  NANDN U90 ( .A(n80), .B(n7066), .Z(n81) );
  NANDN U91 ( .A(n7067), .B(n81), .Z(n82) );
  NAND U92 ( .A(n7068), .B(n82), .Z(n83) );
  NAND U93 ( .A(n7069), .B(n83), .Z(n7072) );
  NANDN U94 ( .A(n1699), .B(n1700), .Z(n7118) );
  ANDN U95 ( .B(n1683), .A(n1682), .Z(n7150) );
  NANDN U96 ( .A(n1662), .B(n1663), .Z(n7189) );
  ANDN U97 ( .B(n1631), .A(n1630), .Z(n7222) );
  ANDN U98 ( .B(n5236), .A(n5235), .Z(n84) );
  AND U99 ( .A(n84), .B(n5241), .Z(n7235) );
  ANDN U100 ( .B(n1597), .A(n1596), .Z(n7276) );
  NAND U101 ( .A(n5311), .B(n5310), .Z(n85) );
  AND U102 ( .A(n5312), .B(n85), .Z(n7290) );
  NANDN U103 ( .A(n1538), .B(n1535), .Z(n86) );
  ANDN U104 ( .B(n86), .A(n1540), .Z(n7332) );
  ANDN U105 ( .B(n1762), .A(n1761), .Z(n7041) );
  NANDN U106 ( .A(n1745), .B(n1746), .Z(n7057) );
  ANDN U107 ( .B(n1728), .A(n1727), .Z(n7073) );
  ANDN U108 ( .B(n1698), .A(n1697), .Z(n7120) );
  NANDN U109 ( .A(n1680), .B(n1681), .Z(n7152) );
  NANDN U110 ( .A(n1658), .B(n1659), .Z(n7193) );
  OR U111 ( .A(n7225), .B(n7226), .Z(n87) );
  NANDN U112 ( .A(n7227), .B(n87), .Z(n88) );
  AND U113 ( .A(n7228), .B(n88), .Z(n89) );
  OR U114 ( .A(n7229), .B(n89), .Z(n90) );
  NAND U115 ( .A(n7230), .B(n90), .Z(n91) );
  NANDN U116 ( .A(n7231), .B(n91), .Z(n92) );
  NAND U117 ( .A(n7232), .B(n92), .Z(n93) );
  NANDN U118 ( .A(n7233), .B(n93), .Z(n94) );
  ANDN U119 ( .B(n94), .A(n7234), .Z(n95) );
  NANDN U120 ( .A(n95), .B(n7235), .Z(n96) );
  ANDN U121 ( .B(n96), .A(n5405), .Z(n97) );
  NANDN U122 ( .A(n97), .B(n7236), .Z(n98) );
  NANDN U123 ( .A(n5404), .B(n98), .Z(n99) );
  NAND U124 ( .A(n7237), .B(n99), .Z(n7238) );
  ANDN U125 ( .B(n1589), .A(n1588), .Z(n7281) );
  NAND U126 ( .A(n7320), .B(n7321), .Z(n100) );
  NANDN U127 ( .A(n7322), .B(n100), .Z(n101) );
  AND U128 ( .A(n5391), .B(n101), .Z(n102) );
  NANDN U129 ( .A(n102), .B(n7323), .Z(n103) );
  NAND U130 ( .A(n7324), .B(n103), .Z(n104) );
  NANDN U131 ( .A(n7325), .B(n104), .Z(n105) );
  NAND U132 ( .A(n7326), .B(n105), .Z(n106) );
  NANDN U133 ( .A(n7327), .B(n106), .Z(n107) );
  AND U134 ( .A(n7328), .B(n107), .Z(n108) );
  ANDN U135 ( .B(n7330), .A(n108), .Z(n109) );
  NAND U136 ( .A(n7329), .B(n109), .Z(n110) );
  AND U137 ( .A(n5390), .B(n110), .Z(n111) );
  NANDN U138 ( .A(n111), .B(n7331), .Z(n112) );
  NAND U139 ( .A(n7332), .B(n112), .Z(n113) );
  NAND U140 ( .A(n7333), .B(n113), .Z(n7334) );
  ANDN U141 ( .B(n1837), .A(n1836), .Z(n6708) );
  ANDN U142 ( .B(n1749), .A(n1748), .Z(n7045) );
  NANDN U143 ( .A(n1738), .B(n1739), .Z(n7061) );
  NANDN U144 ( .A(n5083), .B(n5084), .Z(n114) );
  NAND U145 ( .A(n5085), .B(n114), .Z(n7085) );
  NANDN U146 ( .A(n1695), .B(n1696), .Z(n7122) );
  ANDN U147 ( .B(n1677), .A(n1676), .Z(n7156) );
  NANDN U148 ( .A(n1656), .B(n1655), .Z(n115) );
  AND U149 ( .A(n1657), .B(n115), .Z(n7195) );
  ANDN U150 ( .B(n5212), .A(n5211), .Z(n7223) );
  ANDN U151 ( .B(n1623), .A(n1622), .Z(n7236) );
  ANDN U152 ( .B(n1613), .A(n1612), .Z(n7260) );
  ANDN U153 ( .B(n1591), .A(n1590), .Z(n7284) );
  NANDN U154 ( .A(y[984]), .B(x[984]), .Z(n116) );
  ANDN U155 ( .B(n116), .A(n1580), .Z(n7311) );
  NANDN U156 ( .A(n1550), .B(n1549), .Z(n117) );
  NAND U157 ( .A(n5359), .B(n117), .Z(n118) );
  ANDN U158 ( .B(n118), .A(n1548), .Z(n119) );
  XNOR U159 ( .A(x[1003]), .B(n1554), .Z(n120) );
  NAND U160 ( .A(y[1003]), .B(n120), .Z(n121) );
  NANDN U161 ( .A(x[1003]), .B(n1554), .Z(n122) );
  NAND U162 ( .A(n121), .B(n122), .Z(n123) );
  NAND U163 ( .A(n1553), .B(n119), .Z(n124) );
  NANDN U164 ( .A(n5358), .B(n124), .Z(n125) );
  AND U165 ( .A(n123), .B(n125), .Z(n7326) );
  NANDN U166 ( .A(n5384), .B(n5383), .Z(n5388) );
  NAND U167 ( .A(n2052), .B(n2053), .Z(n126) );
  AND U168 ( .A(n2051), .B(n126), .Z(n127) );
  NAND U169 ( .A(n127), .B(n2050), .Z(n128) );
  NAND U170 ( .A(n2054), .B(n128), .Z(n129) );
  NAND U171 ( .A(n2049), .B(n129), .Z(n130) );
  ANDN U172 ( .B(n130), .A(n2055), .Z(n131) );
  NANDN U173 ( .A(n131), .B(n2056), .Z(n132) );
  NANDN U174 ( .A(n2048), .B(n132), .Z(n133) );
  NAND U175 ( .A(n2047), .B(n133), .Z(n134) );
  NANDN U176 ( .A(n2046), .B(n134), .Z(n135) );
  NAND U177 ( .A(n2045), .B(n135), .Z(n136) );
  ANDN U178 ( .B(n136), .A(n2057), .Z(n5427) );
  NANDN U179 ( .A(n6697), .B(n6696), .Z(n137) );
  NAND U180 ( .A(n6698), .B(n137), .Z(n138) );
  ANDN U181 ( .B(n138), .A(n6699), .Z(n139) );
  NANDN U182 ( .A(n139), .B(n6700), .Z(n140) );
  NANDN U183 ( .A(n6701), .B(n140), .Z(n141) );
  NAND U184 ( .A(n6702), .B(n141), .Z(n142) );
  NANDN U185 ( .A(n6703), .B(n142), .Z(n143) );
  NAND U186 ( .A(n6704), .B(n143), .Z(n144) );
  ANDN U187 ( .B(n144), .A(n6705), .Z(n145) );
  OR U188 ( .A(n6706), .B(n145), .Z(n146) );
  NAND U189 ( .A(n6707), .B(n146), .Z(n147) );
  NANDN U190 ( .A(n5425), .B(n147), .Z(n148) );
  NAND U191 ( .A(n6708), .B(n148), .Z(n149) );
  NANDN U192 ( .A(n6709), .B(n149), .Z(n150) );
  AND U193 ( .A(n6710), .B(n150), .Z(n151) );
  NANDN U194 ( .A(n151), .B(n6711), .Z(n152) );
  NANDN U195 ( .A(n6712), .B(n152), .Z(n153) );
  NAND U196 ( .A(n6713), .B(n153), .Z(n154) );
  NANDN U197 ( .A(n6714), .B(n154), .Z(n6715) );
  NANDN U198 ( .A(y[834]), .B(x[834]), .Z(n155) );
  ANDN U199 ( .B(n155), .A(n1747), .Z(n7048) );
  NAND U200 ( .A(n1740), .B(n1741), .Z(n156) );
  ANDN U201 ( .B(n156), .A(n1742), .Z(n7059) );
  NOR U202 ( .A(n1723), .B(n1724), .Z(n7080) );
  ANDN U203 ( .B(n1707), .A(n1706), .Z(n7112) );
  NAND U204 ( .A(n5145), .B(n5146), .Z(n157) );
  ANDN U205 ( .B(n157), .A(n5147), .Z(n7161) );
  NANDN U206 ( .A(n1653), .B(n1652), .Z(n158) );
  AND U207 ( .A(n1654), .B(n158), .Z(n7199) );
  ANDN U208 ( .B(n5234), .A(n5233), .Z(n5241) );
  ANDN U209 ( .B(n1629), .A(n1628), .Z(n7224) );
  NANDN U210 ( .A(n5248), .B(n5249), .Z(n159) );
  NAND U211 ( .A(n5250), .B(n159), .Z(n5404) );
  ANDN U212 ( .B(n5278), .A(n5277), .Z(n7267) );
  NAND U213 ( .A(n1593), .B(n1592), .Z(n160) );
  NAND U214 ( .A(n1594), .B(n160), .Z(n161) );
  NANDN U215 ( .A(n1595), .B(n161), .Z(n5397) );
  NOR U216 ( .A(n1557), .B(n1558), .Z(n5352) );
  ANDN U217 ( .B(n1552), .A(n1551), .Z(n5359) );
  NANDN U218 ( .A(y[986]), .B(x[986]), .Z(n162) );
  ANDN U219 ( .B(n162), .A(n1579), .Z(n7317) );
  AND U220 ( .A(e), .B(n7341), .Z(n163) );
  AND U221 ( .A(n5380), .B(n5379), .Z(n164) );
  NANDN U222 ( .A(n5382), .B(n5381), .Z(n165) );
  NAND U223 ( .A(n164), .B(n165), .Z(n166) );
  AND U224 ( .A(n5387), .B(n5388), .Z(n167) );
  NANDN U225 ( .A(n7335), .B(n7334), .Z(n168) );
  AND U226 ( .A(n167), .B(n168), .Z(n169) );
  NAND U227 ( .A(n7336), .B(n169), .Z(n170) );
  NAND U228 ( .A(n7337), .B(n170), .Z(n171) );
  AND U229 ( .A(n7338), .B(n171), .Z(n172) );
  OR U230 ( .A(n166), .B(n172), .Z(n173) );
  NAND U231 ( .A(n5378), .B(n173), .Z(n174) );
  NAND U232 ( .A(n7339), .B(n174), .Z(n175) );
  NANDN U233 ( .A(n163), .B(g), .Z(n176) );
  AND U234 ( .A(n7340), .B(n175), .Z(n177) );
  NAND U235 ( .A(n163), .B(n177), .Z(n178) );
  NAND U236 ( .A(n176), .B(n178), .Z(n4) );
  IV U237 ( .A(ebreg), .Z(e) );
  NANDN U238 ( .A(x[1013]), .B(y[1013]), .Z(n180) );
  NANDN U239 ( .A(x[1012]), .B(y[1012]), .Z(n179) );
  AND U240 ( .A(n180), .B(n179), .Z(n5386) );
  NANDN U241 ( .A(x[1011]), .B(y[1011]), .Z(n182) );
  NANDN U242 ( .A(x[1010]), .B(y[1010]), .Z(n181) );
  AND U243 ( .A(n182), .B(n181), .Z(n7333) );
  AND U244 ( .A(n5386), .B(n7333), .Z(n188) );
  NANDN U245 ( .A(y[1018]), .B(x[1018]), .Z(n184) );
  NANDN U246 ( .A(y[1019]), .B(x[1019]), .Z(n183) );
  AND U247 ( .A(n184), .B(n183), .Z(n5382) );
  NANDN U248 ( .A(y[1017]), .B(x[1017]), .Z(n186) );
  NANDN U249 ( .A(y[1016]), .B(x[1016]), .Z(n185) );
  AND U250 ( .A(n186), .B(n185), .Z(n7337) );
  AND U251 ( .A(n5382), .B(n7337), .Z(n187) );
  AND U252 ( .A(n188), .B(n187), .Z(n189) );
  NANDN U253 ( .A(x[1023]), .B(y[1023]), .Z(n7340) );
  AND U254 ( .A(n189), .B(n7340), .Z(n193) );
  NANDN U255 ( .A(x[1015]), .B(y[1015]), .Z(n191) );
  NANDN U256 ( .A(x[1014]), .B(y[1014]), .Z(n190) );
  AND U257 ( .A(n191), .B(n190), .Z(n5384) );
  NANDN U258 ( .A(y[1020]), .B(x[1020]), .Z(n5379) );
  AND U259 ( .A(n5384), .B(n5379), .Z(n192) );
  AND U260 ( .A(n193), .B(n192), .Z(n203) );
  NANDN U261 ( .A(y[1014]), .B(x[1014]), .Z(n195) );
  NANDN U262 ( .A(y[1013]), .B(x[1013]), .Z(n194) );
  AND U263 ( .A(n195), .B(n194), .Z(n196) );
  NANDN U264 ( .A(y[1015]), .B(x[1015]), .Z(n5383) );
  AND U265 ( .A(n196), .B(n5383), .Z(n5385) );
  NANDN U266 ( .A(y[1010]), .B(x[1010]), .Z(n1541) );
  NANDN U267 ( .A(x[1011]), .B(n1541), .Z(n199) );
  XNOR U268 ( .A(x[1011]), .B(n1541), .Z(n197) );
  NAND U269 ( .A(n197), .B(y[1011]), .Z(n198) );
  NAND U270 ( .A(n199), .B(n198), .Z(n200) );
  AND U271 ( .A(n5385), .B(n200), .Z(n202) );
  NANDN U272 ( .A(y[1012]), .B(x[1012]), .Z(n201) );
  AND U273 ( .A(n202), .B(n201), .Z(n5389) );
  AND U274 ( .A(n203), .B(n5389), .Z(n204) );
  ANDN U275 ( .B(y[1009]), .A(x[1009]), .Z(n1538) );
  ANDN U276 ( .B(x[1008]), .A(y[1008]), .Z(n1535) );
  ANDN U277 ( .B(x[1009]), .A(y[1009]), .Z(n1540) );
  AND U278 ( .A(n204), .B(n7332), .Z(n218) );
  NANDN U279 ( .A(y[1023]), .B(x[1023]), .Z(n206) );
  NANDN U280 ( .A(y[1022]), .B(x[1022]), .Z(n205) );
  AND U281 ( .A(n206), .B(n205), .Z(n7339) );
  NANDN U282 ( .A(x[1016]), .B(y[1016]), .Z(n7336) );
  AND U283 ( .A(n7339), .B(n7336), .Z(n210) );
  NANDN U284 ( .A(y[1021]), .B(x[1021]), .Z(n5380) );
  NANDN U285 ( .A(x[1022]), .B(y[1022]), .Z(n208) );
  NANDN U286 ( .A(x[1021]), .B(y[1021]), .Z(n207) );
  AND U287 ( .A(n208), .B(n207), .Z(n5378) );
  AND U288 ( .A(n5380), .B(n5378), .Z(n209) );
  AND U289 ( .A(n210), .B(n209), .Z(n216) );
  NANDN U290 ( .A(x[1018]), .B(y[1018]), .Z(n212) );
  NANDN U291 ( .A(x[1017]), .B(y[1017]), .Z(n211) );
  AND U292 ( .A(n212), .B(n211), .Z(n215) );
  NANDN U293 ( .A(x[1020]), .B(y[1020]), .Z(n214) );
  NANDN U294 ( .A(x[1019]), .B(y[1019]), .Z(n213) );
  AND U295 ( .A(n214), .B(n213), .Z(n5381) );
  AND U296 ( .A(n215), .B(n5381), .Z(n7338) );
  AND U297 ( .A(n216), .B(n7338), .Z(n217) );
  AND U298 ( .A(n218), .B(n217), .Z(n1545) );
  NANDN U299 ( .A(x[1007]), .B(y[1007]), .Z(n5371) );
  NANDN U300 ( .A(x[1006]), .B(y[1006]), .Z(n219) );
  AND U301 ( .A(n5371), .B(n219), .Z(n7329) );
  NANDN U302 ( .A(x[1005]), .B(y[1005]), .Z(n7330) );
  ANDN U303 ( .B(y[1004]), .A(x[1004]), .Z(n7327) );
  ANDN U304 ( .B(n7330), .A(n7327), .Z(n1531) );
  NANDN U305 ( .A(x[1003]), .B(y[1003]), .Z(n221) );
  NANDN U306 ( .A(x[1002]), .B(y[1002]), .Z(n220) );
  AND U307 ( .A(n221), .B(n220), .Z(n1547) );
  NANDN U308 ( .A(y[1002]), .B(x[1002]), .Z(n1554) );
  NANDN U309 ( .A(x[1001]), .B(y[1001]), .Z(n1546) );
  NANDN U310 ( .A(x[1000]), .B(y[1000]), .Z(n1552) );
  AND U311 ( .A(n1546), .B(n1552), .Z(n1525) );
  ANDN U312 ( .B(x[999]), .A(y[999]), .Z(n1550) );
  NANDN U313 ( .A(y[1000]), .B(x[1000]), .Z(n1553) );
  ANDN U314 ( .B(y[998]), .A(x[998]), .Z(n5363) );
  NANDN U315 ( .A(y[998]), .B(x[998]), .Z(n1549) );
  ANDN U316 ( .B(y[996]), .A(x[996]), .Z(n1557) );
  NANDN U317 ( .A(y[995]), .B(x[995]), .Z(n5349) );
  NANDN U318 ( .A(y[996]), .B(x[996]), .Z(n5354) );
  AND U319 ( .A(n5349), .B(n5354), .Z(n1516) );
  ANDN U320 ( .B(y[995]), .A(x[995]), .Z(n1558) );
  NANDN U321 ( .A(x[994]), .B(y[994]), .Z(n1556) );
  NANDN U322 ( .A(y[993]), .B(x[993]), .Z(n1562) );
  NANDN U323 ( .A(x[993]), .B(y[993]), .Z(n1555) );
  ANDN U324 ( .B(x[992]), .A(y[992]), .Z(n1560) );
  NANDN U325 ( .A(x[991]), .B(y[991]), .Z(n1566) );
  ANDN U326 ( .B(x[990]), .A(y[990]), .Z(n1563) );
  NANDN U327 ( .A(x[989]), .B(y[989]), .Z(n1573) );
  NANDN U328 ( .A(x[988]), .B(y[988]), .Z(n5341) );
  AND U329 ( .A(n1573), .B(n5341), .Z(n1504) );
  ANDN U330 ( .B(x[987]), .A(y[987]), .Z(n1579) );
  NANDN U331 ( .A(x[987]), .B(y[987]), .Z(n5342) );
  XNOR U332 ( .A(x[986]), .B(y[986]), .Z(n5337) );
  ANDN U333 ( .B(y[984]), .A(x[984]), .Z(n7309) );
  NANDN U334 ( .A(x[985]), .B(y[985]), .Z(n7315) );
  ANDN U335 ( .B(x[983]), .A(y[983]), .Z(n7306) );
  NANDN U336 ( .A(x[982]), .B(y[982]), .Z(n222) );
  NANDN U337 ( .A(x[983]), .B(y[983]), .Z(n5334) );
  NAND U338 ( .A(n222), .B(n5334), .Z(n7303) );
  XNOR U339 ( .A(x[982]), .B(y[982]), .Z(n5327) );
  ANDN U340 ( .B(x[981]), .A(y[981]), .Z(n1582) );
  ANDN U341 ( .B(n5327), .A(n1582), .Z(n7302) );
  ANDN U342 ( .B(y[980]), .A(x[980]), .Z(n5321) );
  NANDN U343 ( .A(x[981]), .B(y[981]), .Z(n5326) );
  NANDN U344 ( .A(n5321), .B(n5326), .Z(n7300) );
  NANDN U345 ( .A(y[979]), .B(x[979]), .Z(n5317) );
  ANDN U346 ( .B(x[980]), .A(y[980]), .Z(n1581) );
  ANDN U347 ( .B(n5317), .A(n1581), .Z(n7298) );
  NANDN U348 ( .A(x[977]), .B(y[977]), .Z(n5309) );
  NANDN U349 ( .A(x[976]), .B(y[976]), .Z(n223) );
  AND U350 ( .A(n5309), .B(n223), .Z(n7291) );
  ANDN U351 ( .B(y[978]), .A(x[978]), .Z(n5316) );
  ANDN U352 ( .B(y[979]), .A(x[979]), .Z(n5322) );
  NOR U353 ( .A(n5316), .B(n5322), .Z(n7295) );
  NAND U354 ( .A(n7291), .B(n7295), .Z(n1489) );
  NANDN U355 ( .A(y[976]), .B(x[976]), .Z(n5306) );
  NANDN U356 ( .A(x[974]), .B(y[974]), .Z(n224) );
  NANDN U357 ( .A(x[975]), .B(y[975]), .Z(n5310) );
  AND U358 ( .A(n224), .B(n5310), .Z(n1584) );
  ANDN U359 ( .B(x[974]), .A(y[974]), .Z(n5311) );
  NANDN U360 ( .A(x[973]), .B(y[973]), .Z(n1583) );
  NANDN U361 ( .A(y[971]), .B(x[971]), .Z(n1591) );
  NANDN U362 ( .A(x[970]), .B(y[970]), .Z(n7282) );
  ANDN U363 ( .B(x[970]), .A(y[970]), .Z(n1590) );
  ANDN U364 ( .B(y[968]), .A(x[968]), .Z(n7280) );
  NANDN U365 ( .A(x[969]), .B(y[969]), .Z(n7283) );
  ANDN U366 ( .B(x[968]), .A(y[968]), .Z(n1588) );
  NANDN U367 ( .A(x[966]), .B(y[966]), .Z(n5290) );
  NANDN U368 ( .A(x[967]), .B(y[967]), .Z(n5297) );
  AND U369 ( .A(n5290), .B(n5297), .Z(n7278) );
  ANDN U370 ( .B(x[965]), .A(y[965]), .Z(n5286) );
  ANDN U371 ( .B(x[966]), .A(y[966]), .Z(n5294) );
  OR U372 ( .A(n5286), .B(n5294), .Z(n7277) );
  NANDN U373 ( .A(x[965]), .B(y[965]), .Z(n5289) );
  NANDN U374 ( .A(x[964]), .B(y[964]), .Z(n225) );
  AND U375 ( .A(n5289), .B(n225), .Z(n5396) );
  NANDN U376 ( .A(x[963]), .B(y[963]), .Z(n1594) );
  NANDN U377 ( .A(x[962]), .B(y[962]), .Z(n226) );
  AND U378 ( .A(n1594), .B(n226), .Z(n1597) );
  ANDN U379 ( .B(x[961]), .A(y[961]), .Z(n1598) );
  ANDN U380 ( .B(y[960]), .A(x[960]), .Z(n1601) );
  NANDN U381 ( .A(y[960]), .B(x[960]), .Z(n1600) );
  NANDN U382 ( .A(x[959]), .B(y[959]), .Z(n1603) );
  NANDN U383 ( .A(x[958]), .B(y[958]), .Z(n1609) );
  AND U384 ( .A(n1603), .B(n1609), .Z(n1458) );
  ANDN U385 ( .B(x[958]), .A(y[958]), .Z(n1604) );
  NANDN U386 ( .A(y[957]), .B(x[957]), .Z(n1611) );
  ANDN U387 ( .B(y[956]), .A(x[956]), .Z(n5277) );
  NANDN U388 ( .A(y[956]), .B(x[956]), .Z(n1610) );
  NANDN U389 ( .A(x[955]), .B(y[955]), .Z(n5278) );
  NANDN U390 ( .A(x[954]), .B(y[954]), .Z(n7262) );
  AND U391 ( .A(n5278), .B(n7262), .Z(n1450) );
  NANDN U392 ( .A(y[953]), .B(x[953]), .Z(n1613) );
  NANDN U393 ( .A(y[954]), .B(x[954]), .Z(n1614) );
  ANDN U394 ( .B(y[953]), .A(x[953]), .Z(n5399) );
  NANDN U395 ( .A(x[950]), .B(y[950]), .Z(n5266) );
  NANDN U396 ( .A(x[951]), .B(y[951]), .Z(n5273) );
  AND U397 ( .A(n5266), .B(n5273), .Z(n7254) );
  ANDN U398 ( .B(x[949]), .A(y[949]), .Z(n5262) );
  ANDN U399 ( .B(x[950]), .A(y[950]), .Z(n5270) );
  OR U400 ( .A(n5262), .B(n5270), .Z(n7252) );
  NANDN U401 ( .A(x[948]), .B(y[948]), .Z(n5260) );
  NANDN U402 ( .A(x[949]), .B(y[949]), .Z(n5265) );
  NAND U403 ( .A(n5260), .B(n5265), .Z(n5401) );
  NANDN U404 ( .A(y[948]), .B(x[948]), .Z(n1616) );
  NANDN U405 ( .A(x[946]), .B(y[946]), .Z(n227) );
  NANDN U406 ( .A(x[947]), .B(y[947]), .Z(n5403) );
  NAND U407 ( .A(n227), .B(n5403), .Z(n7240) );
  NANDN U408 ( .A(y[945]), .B(x[945]), .Z(n1619) );
  XNOR U409 ( .A(x[946]), .B(y[946]), .Z(n1618) );
  ANDN U410 ( .B(y[944]), .A(x[944]), .Z(n1621) );
  NANDN U411 ( .A(y[943]), .B(x[943]), .Z(n5250) );
  NANDN U412 ( .A(x[943]), .B(y[943]), .Z(n5249) );
  NANDN U413 ( .A(x[942]), .B(y[942]), .Z(n228) );
  NAND U414 ( .A(n5249), .B(n228), .Z(n1622) );
  NANDN U415 ( .A(y[942]), .B(x[942]), .Z(n5248) );
  NANDN U416 ( .A(y[941]), .B(x[941]), .Z(n5243) );
  NANDN U417 ( .A(y[940]), .B(x[940]), .Z(n5244) );
  NANDN U418 ( .A(y[939]), .B(x[939]), .Z(n5238) );
  AND U419 ( .A(n5244), .B(n5238), .Z(n1425) );
  ANDN U420 ( .B(y[938]), .A(x[938]), .Z(n5235) );
  NANDN U421 ( .A(y[938]), .B(x[938]), .Z(n5239) );
  ANDN U422 ( .B(y[936]), .A(x[936]), .Z(n7233) );
  NANDN U423 ( .A(y[935]), .B(x[935]), .Z(n7232) );
  NANDN U424 ( .A(y[933]), .B(x[933]), .Z(n5220) );
  XOR U425 ( .A(x[934]), .B(y[934]), .Z(n5225) );
  ANDN U426 ( .B(n5220), .A(n5225), .Z(n7230) );
  ANDN U427 ( .B(y[932]), .A(x[932]), .Z(n5216) );
  ANDN U428 ( .B(y[933]), .A(x[933]), .Z(n5222) );
  OR U429 ( .A(n5216), .B(n5222), .Z(n7229) );
  NANDN U430 ( .A(y[932]), .B(x[932]), .Z(n7228) );
  NANDN U431 ( .A(y[931]), .B(x[931]), .Z(n1626) );
  ANDN U432 ( .B(y[931]), .A(x[931]), .Z(n7227) );
  NANDN U433 ( .A(y[930]), .B(x[930]), .Z(n1627) );
  NANDN U434 ( .A(x[929]), .B(y[929]), .Z(n1629) );
  ANDN U435 ( .B(y[928]), .A(x[928]), .Z(n1630) );
  ANDN U436 ( .B(n1629), .A(n1630), .Z(n1405) );
  ANDN U437 ( .B(x[927]), .A(y[927]), .Z(n1633) );
  NANDN U438 ( .A(x[927]), .B(y[927]), .Z(n1631) );
  ANDN U439 ( .B(x[925]), .A(y[925]), .Z(n1637) );
  NANDN U440 ( .A(x[925]), .B(y[925]), .Z(n1636) );
  ANDN U441 ( .B(x[923]), .A(y[923]), .Z(n1642) );
  NANDN U442 ( .A(x[922]), .B(y[922]), .Z(n229) );
  ANDN U443 ( .B(y[923]), .A(x[923]), .Z(n1641) );
  ANDN U444 ( .B(n229), .A(n1641), .Z(n1646) );
  ANDN U445 ( .B(x[921]), .A(y[921]), .Z(n1647) );
  NANDN U446 ( .A(x[921]), .B(y[921]), .Z(n1645) );
  NANDN U447 ( .A(y[919]), .B(x[919]), .Z(n7213) );
  ANDN U448 ( .B(y[918]), .A(x[918]), .Z(n5193) );
  ANDN U449 ( .B(y[919]), .A(x[919]), .Z(n5201) );
  NOR U450 ( .A(n5193), .B(n5201), .Z(n7212) );
  NANDN U451 ( .A(y[917]), .B(x[917]), .Z(n5190) );
  XNOR U452 ( .A(y[918]), .B(x[918]), .Z(n230) );
  NAND U453 ( .A(n5190), .B(n230), .Z(n7211) );
  ANDN U454 ( .B(y[916]), .A(x[916]), .Z(n5186) );
  ANDN U455 ( .B(y[917]), .A(x[917]), .Z(n5196) );
  NOR U456 ( .A(n5186), .B(n5196), .Z(n7210) );
  NANDN U457 ( .A(y[915]), .B(x[915]), .Z(n5182) );
  NANDN U458 ( .A(y[916]), .B(x[916]), .Z(n5191) );
  NAND U459 ( .A(n5182), .B(n5191), .Z(n7209) );
  ANDN U460 ( .B(y[914]), .A(x[914]), .Z(n5181) );
  ANDN U461 ( .B(y[915]), .A(x[915]), .Z(n5188) );
  NOR U462 ( .A(n5181), .B(n5188), .Z(n7208) );
  ANDN U463 ( .B(y[912]), .A(x[912]), .Z(n7201) );
  ANDN U464 ( .B(y[913]), .A(x[913]), .Z(n7204) );
  OR U465 ( .A(n7201), .B(n7204), .Z(n1379) );
  NANDN U466 ( .A(y[911]), .B(x[911]), .Z(n1654) );
  NANDN U467 ( .A(x[910]), .B(y[910]), .Z(n231) );
  NANDN U468 ( .A(x[911]), .B(y[911]), .Z(n1652) );
  AND U469 ( .A(n231), .B(n1652), .Z(n7197) );
  NANDN U470 ( .A(y[909]), .B(x[909]), .Z(n1657) );
  NANDN U471 ( .A(x[908]), .B(y[908]), .Z(n232) );
  NANDN U472 ( .A(x[909]), .B(y[909]), .Z(n1655) );
  AND U473 ( .A(n232), .B(n1655), .Z(n1659) );
  NANDN U474 ( .A(y[907]), .B(x[907]), .Z(n1660) );
  ANDN U475 ( .B(y[906]), .A(x[906]), .Z(n1662) );
  NANDN U476 ( .A(y[905]), .B(x[905]), .Z(n1666) );
  NANDN U477 ( .A(x[902]), .B(y[902]), .Z(n233) );
  ANDN U478 ( .B(y[903]), .A(x[903]), .Z(n5168) );
  ANDN U479 ( .B(n233), .A(n5168), .Z(n7181) );
  ANDN U480 ( .B(x[901]), .A(y[901]), .Z(n5159) );
  XNOR U481 ( .A(x[902]), .B(y[902]), .Z(n1667) );
  NANDN U482 ( .A(n5159), .B(n1667), .Z(n7178) );
  NANDN U483 ( .A(x[900]), .B(y[900]), .Z(n5155) );
  NANDN U484 ( .A(x[901]), .B(y[901]), .Z(n1668) );
  NAND U485 ( .A(n5155), .B(n1668), .Z(n7175) );
  NANDN U486 ( .A(y[900]), .B(x[900]), .Z(n5160) );
  NANDN U487 ( .A(x[898]), .B(y[898]), .Z(n5151) );
  NANDN U488 ( .A(x[899]), .B(y[899]), .Z(n5408) );
  NAND U489 ( .A(n5151), .B(n5408), .Z(n7166) );
  NANDN U490 ( .A(x[897]), .B(y[897]), .Z(n7169) );
  NANDN U491 ( .A(x[896]), .B(y[896]), .Z(n7162) );
  AND U492 ( .A(n7169), .B(n7162), .Z(n1353) );
  ANDN U493 ( .B(x[895]), .A(y[895]), .Z(n5147) );
  NANDN U494 ( .A(x[894]), .B(y[894]), .Z(n234) );
  NANDN U495 ( .A(x[895]), .B(y[895]), .Z(n5145) );
  AND U496 ( .A(n234), .B(n5145), .Z(n1675) );
  NANDN U497 ( .A(y[893]), .B(x[893]), .Z(n1677) );
  NANDN U498 ( .A(x[892]), .B(y[892]), .Z(n1678) );
  ANDN U499 ( .B(x[891]), .A(y[891]), .Z(n1680) );
  NANDN U500 ( .A(x[891]), .B(y[891]), .Z(n1679) );
  NANDN U501 ( .A(y[890]), .B(x[890]), .Z(n1681) );
  ANDN U502 ( .B(x[889]), .A(y[889]), .Z(n1684) );
  ANDN U503 ( .B(n1681), .A(n1684), .Z(n1340) );
  ANDN U504 ( .B(y[888]), .A(x[888]), .Z(n1686) );
  NANDN U505 ( .A(y[888]), .B(x[888]), .Z(n1685) );
  ANDN U506 ( .B(y[886]), .A(x[886]), .Z(n5133) );
  NANDN U507 ( .A(x[887]), .B(y[887]), .Z(n1687) );
  NANDN U508 ( .A(n5133), .B(n1687), .Z(n7140) );
  NANDN U509 ( .A(y[885]), .B(x[885]), .Z(n1689) );
  XNOR U510 ( .A(y[886]), .B(x[886]), .Z(n235) );
  AND U511 ( .A(n1689), .B(n235), .Z(n5409) );
  NANDN U512 ( .A(y[884]), .B(x[884]), .Z(n1690) );
  ANDN U513 ( .B(x[883]), .A(y[883]), .Z(n5123) );
  ANDN U514 ( .B(n1690), .A(n5123), .Z(n7135) );
  ANDN U515 ( .B(y[883]), .A(x[883]), .Z(n5127) );
  NANDN U516 ( .A(x[882]), .B(y[882]), .Z(n5118) );
  NANDN U517 ( .A(n5127), .B(n5118), .Z(n5411) );
  NANDN U518 ( .A(y[882]), .B(x[882]), .Z(n1691) );
  NANDN U519 ( .A(y[881]), .B(x[881]), .Z(n1692) );
  XNOR U520 ( .A(x[880]), .B(y[880]), .Z(n1694) );
  NANDN U521 ( .A(y[879]), .B(x[879]), .Z(n1696) );
  AND U522 ( .A(n1694), .B(n1696), .Z(n1325) );
  ANDN U523 ( .B(y[878]), .A(x[878]), .Z(n1697) );
  NANDN U524 ( .A(x[879]), .B(y[879]), .Z(n7126) );
  ANDN U525 ( .B(x[877]), .A(y[877]), .Z(n1699) );
  NANDN U526 ( .A(x[877]), .B(y[877]), .Z(n1698) );
  NANDN U527 ( .A(y[876]), .B(x[876]), .Z(n1700) );
  ANDN U528 ( .B(x[875]), .A(y[875]), .Z(n1703) );
  ANDN U529 ( .B(n1700), .A(n1703), .Z(n1317) );
  ANDN U530 ( .B(y[874]), .A(x[874]), .Z(n1706) );
  NANDN U531 ( .A(y[874]), .B(x[874]), .Z(n1704) );
  ANDN U532 ( .B(y[872]), .A(x[872]), .Z(n1710) );
  NANDN U533 ( .A(x[870]), .B(y[870]), .Z(n1712) );
  NANDN U534 ( .A(x[871]), .B(y[871]), .Z(n1711) );
  NAND U535 ( .A(n1712), .B(n1711), .Z(n7102) );
  ANDN U536 ( .B(x[869]), .A(y[869]), .Z(n5097) );
  ANDN U537 ( .B(x[870]), .A(y[870]), .Z(n5103) );
  NOR U538 ( .A(n5097), .B(n5103), .Z(n7101) );
  NANDN U539 ( .A(x[868]), .B(y[868]), .Z(n5093) );
  NANDN U540 ( .A(x[869]), .B(y[869]), .Z(n1713) );
  NAND U541 ( .A(n5093), .B(n1713), .Z(n5414) );
  NANDN U542 ( .A(y[868]), .B(x[868]), .Z(n5098) );
  NANDN U543 ( .A(x[866]), .B(y[866]), .Z(n5089) );
  NANDN U544 ( .A(x[867]), .B(y[867]), .Z(n5416) );
  NAND U545 ( .A(n5089), .B(n5416), .Z(n5417) );
  NANDN U546 ( .A(y[865]), .B(x[865]), .Z(n1716) );
  ANDN U547 ( .B(y[864]), .A(x[864]), .Z(n1718) );
  NANDN U548 ( .A(y[863]), .B(x[863]), .Z(n5085) );
  NANDN U549 ( .A(x[863]), .B(y[863]), .Z(n5084) );
  NANDN U550 ( .A(x[862]), .B(y[862]), .Z(n236) );
  AND U551 ( .A(n5084), .B(n236), .Z(n1720) );
  NANDN U552 ( .A(y[862]), .B(x[862]), .Z(n5083) );
  NANDN U553 ( .A(y[861]), .B(x[861]), .Z(n1722) );
  NANDN U554 ( .A(y[860]), .B(x[860]), .Z(n1721) );
  NANDN U555 ( .A(y[859]), .B(x[859]), .Z(n1726) );
  AND U556 ( .A(n1721), .B(n1726), .Z(n1290) );
  ANDN U557 ( .B(y[858]), .A(x[858]), .Z(n5076) );
  NANDN U558 ( .A(y[858]), .B(x[858]), .Z(n1725) );
  NANDN U559 ( .A(x[857]), .B(y[857]), .Z(n5077) );
  ANDN U560 ( .B(y[856]), .A(x[856]), .Z(n7070) );
  ANDN U561 ( .B(n5077), .A(n7070), .Z(n1284) );
  NANDN U562 ( .A(y[855]), .B(x[855]), .Z(n7069) );
  NANDN U563 ( .A(x[854]), .B(y[854]), .Z(n5067) );
  ANDN U564 ( .B(y[855]), .A(x[855]), .Z(n5074) );
  ANDN U565 ( .B(n5067), .A(n5074), .Z(n7068) );
  ANDN U566 ( .B(x[853]), .A(y[853]), .Z(n5063) );
  NANDN U567 ( .A(y[854]), .B(x[854]), .Z(n1729) );
  NANDN U568 ( .A(n5063), .B(n1729), .Z(n7067) );
  NANDN U569 ( .A(x[852]), .B(y[852]), .Z(n5061) );
  ANDN U570 ( .B(y[853]), .A(x[853]), .Z(n5069) );
  ANDN U571 ( .B(n5061), .A(n5069), .Z(n7066) );
  ANDN U572 ( .B(x[852]), .A(y[852]), .Z(n5065) );
  NANDN U573 ( .A(x[851]), .B(y[851]), .Z(n238) );
  NANDN U574 ( .A(x[850]), .B(y[850]), .Z(n237) );
  AND U575 ( .A(n238), .B(n237), .Z(n239) );
  NANDN U576 ( .A(n5065), .B(n5058), .Z(n7064) );
  NANDN U577 ( .A(x[849]), .B(y[849]), .Z(n240) );
  AND U578 ( .A(n240), .B(n239), .Z(n1731) );
  NANDN U579 ( .A(x[848]), .B(y[848]), .Z(n241) );
  AND U580 ( .A(n1731), .B(n241), .Z(n1733) );
  NANDN U581 ( .A(y[847]), .B(x[847]), .Z(n1734) );
  NANDN U582 ( .A(x[846]), .B(y[846]), .Z(n1736) );
  NANDN U583 ( .A(x[845]), .B(y[845]), .Z(n1737) );
  NANDN U584 ( .A(x[844]), .B(y[844]), .Z(n7060) );
  AND U585 ( .A(n1737), .B(n7060), .Z(n1269) );
  ANDN U586 ( .B(x[843]), .A(y[843]), .Z(n1742) );
  NANDN U587 ( .A(x[842]), .B(y[842]), .Z(n242) );
  NANDN U588 ( .A(x[843]), .B(y[843]), .Z(n1740) );
  AND U589 ( .A(n242), .B(n1740), .Z(n1744) );
  NANDN U590 ( .A(y[841]), .B(x[841]), .Z(n1746) );
  NANDN U591 ( .A(x[841]), .B(y[841]), .Z(n1743) );
  ANDN U592 ( .B(x[839]), .A(y[839]), .Z(n7055) );
  NANDN U593 ( .A(x[838]), .B(y[838]), .Z(n243) );
  NANDN U594 ( .A(x[839]), .B(y[839]), .Z(n5046) );
  AND U595 ( .A(n243), .B(n5046), .Z(n7054) );
  ANDN U596 ( .B(x[837]), .A(y[837]), .Z(n5037) );
  XNOR U597 ( .A(x[838]), .B(y[838]), .Z(n5040) );
  NANDN U598 ( .A(n5037), .B(n5040), .Z(n7053) );
  NANDN U599 ( .A(x[836]), .B(y[836]), .Z(n5034) );
  NANDN U600 ( .A(x[837]), .B(y[837]), .Z(n5041) );
  AND U601 ( .A(n5034), .B(n5041), .Z(n7052) );
  ANDN U602 ( .B(x[836]), .A(y[836]), .Z(n7050) );
  NANDN U603 ( .A(x[834]), .B(y[834]), .Z(n7047) );
  NANDN U604 ( .A(x[835]), .B(y[835]), .Z(n7049) );
  AND U605 ( .A(n7047), .B(n7049), .Z(n1253) );
  XNOR U606 ( .A(x[834]), .B(y[834]), .Z(n5029) );
  NANDN U607 ( .A(x[833]), .B(y[833]), .Z(n7046) );
  ANDN U608 ( .B(x[831]), .A(y[831]), .Z(n1753) );
  NANDN U609 ( .A(x[830]), .B(y[830]), .Z(n244) );
  NANDN U610 ( .A(x[831]), .B(y[831]), .Z(n1750) );
  AND U611 ( .A(n244), .B(n1750), .Z(n1757) );
  ANDN U612 ( .B(x[829]), .A(y[829]), .Z(n1758) );
  NANDN U613 ( .A(x[828]), .B(y[828]), .Z(n5424) );
  XOR U614 ( .A(x[828]), .B(y[828]), .Z(n5023) );
  ANDN U615 ( .B(y[827]), .A(x[827]), .Z(n5423) );
  NANDN U616 ( .A(y[825]), .B(x[825]), .Z(n1767) );
  ANDN U617 ( .B(y[822]), .A(x[822]), .Z(n1769) );
  ANDN U618 ( .B(y[823]), .A(x[823]), .Z(n5016) );
  NOR U619 ( .A(n1769), .B(n5016), .Z(n7036) );
  ANDN U620 ( .B(x[821]), .A(y[821]), .Z(n5007) );
  NANDN U621 ( .A(y[822]), .B(x[822]), .Z(n5012) );
  NANDN U622 ( .A(n5007), .B(n5012), .Z(n7034) );
  NANDN U623 ( .A(x[820]), .B(y[820]), .Z(n5003) );
  ANDN U624 ( .B(y[821]), .A(x[821]), .Z(n1768) );
  ANDN U625 ( .B(n5003), .A(n1768), .Z(n7032) );
  ANDN U626 ( .B(x[819]), .A(y[819]), .Z(n4998) );
  ANDN U627 ( .B(x[820]), .A(y[820]), .Z(n5008) );
  OR U628 ( .A(n4998), .B(n5008), .Z(n7030) );
  NANDN U629 ( .A(x[818]), .B(y[818]), .Z(n4995) );
  NANDN U630 ( .A(x[819]), .B(y[819]), .Z(n5002) );
  AND U631 ( .A(n4995), .B(n5002), .Z(n7028) );
  ANDN U632 ( .B(x[817]), .A(y[817]), .Z(n4991) );
  XNOR U633 ( .A(y[818]), .B(x[818]), .Z(n245) );
  NANDN U634 ( .A(n4991), .B(n245), .Z(n7026) );
  NANDN U635 ( .A(x[816]), .B(y[816]), .Z(n246) );
  NANDN U636 ( .A(x[817]), .B(y[817]), .Z(n4996) );
  AND U637 ( .A(n246), .B(n4996), .Z(n7024) );
  ANDN U638 ( .B(x[815]), .A(y[815]), .Z(n1770) );
  XNOR U639 ( .A(x[816]), .B(y[816]), .Z(n4987) );
  NANDN U640 ( .A(n1770), .B(n4987), .Z(n7022) );
  NANDN U641 ( .A(x[814]), .B(y[814]), .Z(n247) );
  NANDN U642 ( .A(x[815]), .B(y[815]), .Z(n4986) );
  AND U643 ( .A(n247), .B(n4986), .Z(n7020) );
  XNOR U644 ( .A(x[814]), .B(y[814]), .Z(n4981) );
  NANDN U645 ( .A(y[813]), .B(x[813]), .Z(n4977) );
  NAND U646 ( .A(n4981), .B(n4977), .Z(n7018) );
  NANDN U647 ( .A(x[813]), .B(y[813]), .Z(n4980) );
  ANDN U648 ( .B(y[812]), .A(x[812]), .Z(n4975) );
  ANDN U649 ( .B(n4980), .A(n4975), .Z(n7016) );
  NANDN U650 ( .A(y[811]), .B(x[811]), .Z(n1772) );
  NANDN U651 ( .A(y[812]), .B(x[812]), .Z(n4978) );
  NAND U652 ( .A(n1772), .B(n4978), .Z(n7014) );
  NANDN U653 ( .A(x[810]), .B(y[810]), .Z(n248) );
  ANDN U654 ( .B(y[811]), .A(x[811]), .Z(n4972) );
  ANDN U655 ( .B(n248), .A(n4972), .Z(n7012) );
  XOR U656 ( .A(x[810]), .B(y[810]), .Z(n4968) );
  NANDN U657 ( .A(y[809]), .B(x[809]), .Z(n4963) );
  NANDN U658 ( .A(n4968), .B(n4963), .Z(n7010) );
  ANDN U659 ( .B(y[808]), .A(x[808]), .Z(n4958) );
  ANDN U660 ( .B(y[809]), .A(x[809]), .Z(n4967) );
  NOR U661 ( .A(n4958), .B(n4967), .Z(n7008) );
  NANDN U662 ( .A(y[807]), .B(x[807]), .Z(n4955) );
  XNOR U663 ( .A(y[808]), .B(x[808]), .Z(n249) );
  NAND U664 ( .A(n4955), .B(n249), .Z(n7006) );
  ANDN U665 ( .B(y[806]), .A(x[806]), .Z(n4951) );
  ANDN U666 ( .B(y[807]), .A(x[807]), .Z(n4961) );
  NOR U667 ( .A(n4951), .B(n4961), .Z(n7004) );
  NANDN U668 ( .A(y[805]), .B(x[805]), .Z(n4947) );
  XNOR U669 ( .A(y[806]), .B(x[806]), .Z(n250) );
  NAND U670 ( .A(n4947), .B(n250), .Z(n7002) );
  ANDN U671 ( .B(y[804]), .A(x[804]), .Z(n1775) );
  ANDN U672 ( .B(y[805]), .A(x[805]), .Z(n4953) );
  NOR U673 ( .A(n1775), .B(n4953), .Z(n7000) );
  ANDN U674 ( .B(x[803]), .A(y[803]), .Z(n4942) );
  XNOR U675 ( .A(y[804]), .B(x[804]), .Z(n251) );
  NANDN U676 ( .A(n4942), .B(n251), .Z(n6998) );
  NANDN U677 ( .A(x[802]), .B(y[802]), .Z(n252) );
  ANDN U678 ( .B(y[803]), .A(x[803]), .Z(n1774) );
  ANDN U679 ( .B(n252), .A(n1774), .Z(n6996) );
  ANDN U680 ( .B(x[801]), .A(y[801]), .Z(n4935) );
  XNOR U681 ( .A(x[802]), .B(y[802]), .Z(n4937) );
  NANDN U682 ( .A(n4935), .B(n4937), .Z(n6994) );
  NANDN U683 ( .A(x[800]), .B(y[800]), .Z(n253) );
  NANDN U684 ( .A(x[801]), .B(y[801]), .Z(n4936) );
  AND U685 ( .A(n253), .B(n4936), .Z(n6992) );
  XNOR U686 ( .A(x[800]), .B(y[800]), .Z(n4929) );
  NANDN U687 ( .A(y[799]), .B(x[799]), .Z(n4925) );
  NAND U688 ( .A(n4929), .B(n4925), .Z(n6990) );
  NANDN U689 ( .A(x[799]), .B(y[799]), .Z(n4930) );
  ANDN U690 ( .B(y[798]), .A(x[798]), .Z(n4921) );
  ANDN U691 ( .B(n4930), .A(n4921), .Z(n6988) );
  ANDN U692 ( .B(x[798]), .A(y[798]), .Z(n4927) );
  NANDN U693 ( .A(y[797]), .B(x[797]), .Z(n4917) );
  NANDN U694 ( .A(n4927), .B(n4917), .Z(n6986) );
  NANDN U695 ( .A(x[796]), .B(y[796]), .Z(n254) );
  ANDN U696 ( .B(y[797]), .A(x[797]), .Z(n4923) );
  ANDN U697 ( .B(n254), .A(n4923), .Z(n6984) );
  XOR U698 ( .A(x[796]), .B(y[796]), .Z(n1776) );
  ANDN U699 ( .B(x[795]), .A(y[795]), .Z(n4911) );
  OR U700 ( .A(n1776), .B(n4911), .Z(n6982) );
  NANDN U701 ( .A(x[794]), .B(y[794]), .Z(n4907) );
  ANDN U702 ( .B(y[795]), .A(x[795]), .Z(n1777) );
  ANDN U703 ( .B(n4907), .A(n1777), .Z(n6980) );
  ANDN U704 ( .B(x[793]), .A(y[793]), .Z(n4902) );
  ANDN U705 ( .B(x[794]), .A(y[794]), .Z(n4912) );
  OR U706 ( .A(n4902), .B(n4912), .Z(n6978) );
  NANDN U707 ( .A(x[792]), .B(y[792]), .Z(n4899) );
  NANDN U708 ( .A(x[793]), .B(y[793]), .Z(n4906) );
  AND U709 ( .A(n4899), .B(n4906), .Z(n6976) );
  ANDN U710 ( .B(x[792]), .A(y[792]), .Z(n4905) );
  NANDN U711 ( .A(y[791]), .B(x[791]), .Z(n4895) );
  NANDN U712 ( .A(n4905), .B(n4895), .Z(n6974) );
  NANDN U713 ( .A(x[791]), .B(y[791]), .Z(n4900) );
  ANDN U714 ( .B(y[790]), .A(x[790]), .Z(n4891) );
  ANDN U715 ( .B(n4900), .A(n4891), .Z(n6972) );
  ANDN U716 ( .B(x[790]), .A(y[790]), .Z(n4897) );
  NANDN U717 ( .A(y[789]), .B(x[789]), .Z(n4887) );
  NANDN U718 ( .A(n4897), .B(n4887), .Z(n6970) );
  NANDN U719 ( .A(x[788]), .B(y[788]), .Z(n255) );
  ANDN U720 ( .B(y[789]), .A(x[789]), .Z(n4893) );
  ANDN U721 ( .B(n255), .A(n4893), .Z(n6968) );
  XOR U722 ( .A(x[788]), .B(y[788]), .Z(n1778) );
  ANDN U723 ( .B(x[787]), .A(y[787]), .Z(n4881) );
  OR U724 ( .A(n1778), .B(n4881), .Z(n6966) );
  NANDN U725 ( .A(x[786]), .B(y[786]), .Z(n4877) );
  ANDN U726 ( .B(y[787]), .A(x[787]), .Z(n1779) );
  ANDN U727 ( .B(n4877), .A(n1779), .Z(n6964) );
  ANDN U728 ( .B(x[785]), .A(y[785]), .Z(n4872) );
  ANDN U729 ( .B(x[786]), .A(y[786]), .Z(n4882) );
  OR U730 ( .A(n4872), .B(n4882), .Z(n6962) );
  NANDN U731 ( .A(x[784]), .B(y[784]), .Z(n4869) );
  NANDN U732 ( .A(x[785]), .B(y[785]), .Z(n4876) );
  AND U733 ( .A(n4869), .B(n4876), .Z(n6960) );
  ANDN U734 ( .B(x[784]), .A(y[784]), .Z(n4875) );
  NANDN U735 ( .A(y[783]), .B(x[783]), .Z(n4865) );
  NANDN U736 ( .A(n4875), .B(n4865), .Z(n6958) );
  NANDN U737 ( .A(x[783]), .B(y[783]), .Z(n4870) );
  ANDN U738 ( .B(y[782]), .A(x[782]), .Z(n4861) );
  ANDN U739 ( .B(n4870), .A(n4861), .Z(n6956) );
  ANDN U740 ( .B(x[782]), .A(y[782]), .Z(n4867) );
  NANDN U741 ( .A(y[781]), .B(x[781]), .Z(n4857) );
  NANDN U742 ( .A(n4867), .B(n4857), .Z(n6954) );
  NANDN U743 ( .A(x[780]), .B(y[780]), .Z(n256) );
  ANDN U744 ( .B(y[781]), .A(x[781]), .Z(n4863) );
  ANDN U745 ( .B(n256), .A(n4863), .Z(n6952) );
  XOR U746 ( .A(x[780]), .B(y[780]), .Z(n1780) );
  ANDN U747 ( .B(x[779]), .A(y[779]), .Z(n4852) );
  OR U748 ( .A(n1780), .B(n4852), .Z(n6950) );
  NANDN U749 ( .A(x[778]), .B(y[778]), .Z(n257) );
  ANDN U750 ( .B(y[779]), .A(x[779]), .Z(n1781) );
  ANDN U751 ( .B(n257), .A(n1781), .Z(n6948) );
  ANDN U752 ( .B(x[777]), .A(y[777]), .Z(n4842) );
  XNOR U753 ( .A(x[778]), .B(y[778]), .Z(n4847) );
  NANDN U754 ( .A(n4842), .B(n4847), .Z(n6946) );
  NANDN U755 ( .A(x[776]), .B(y[776]), .Z(n4839) );
  NANDN U756 ( .A(x[777]), .B(y[777]), .Z(n4846) );
  AND U757 ( .A(n4839), .B(n4846), .Z(n6944) );
  ANDN U758 ( .B(x[775]), .A(y[775]), .Z(n4835) );
  ANDN U759 ( .B(x[776]), .A(y[776]), .Z(n4845) );
  OR U760 ( .A(n4835), .B(n4845), .Z(n6942) );
  NANDN U761 ( .A(x[774]), .B(y[774]), .Z(n4831) );
  NANDN U762 ( .A(x[775]), .B(y[775]), .Z(n4840) );
  AND U763 ( .A(n4831), .B(n4840), .Z(n6940) );
  ANDN U764 ( .B(x[773]), .A(y[773]), .Z(n1782) );
  XNOR U765 ( .A(y[774]), .B(x[774]), .Z(n258) );
  NANDN U766 ( .A(n1782), .B(n258), .Z(n6938) );
  NANDN U767 ( .A(x[772]), .B(y[772]), .Z(n259) );
  NANDN U768 ( .A(x[773]), .B(y[773]), .Z(n4830) );
  AND U769 ( .A(n259), .B(n4830), .Z(n6936) );
  XNOR U770 ( .A(x[772]), .B(y[772]), .Z(n4825) );
  NANDN U771 ( .A(y[771]), .B(x[771]), .Z(n4821) );
  NAND U772 ( .A(n4825), .B(n4821), .Z(n6934) );
  NANDN U773 ( .A(x[771]), .B(y[771]), .Z(n4824) );
  ANDN U774 ( .B(y[770]), .A(x[770]), .Z(n4819) );
  ANDN U775 ( .B(n4824), .A(n4819), .Z(n6932) );
  NANDN U776 ( .A(y[769]), .B(x[769]), .Z(n1784) );
  NANDN U777 ( .A(y[770]), .B(x[770]), .Z(n4822) );
  NAND U778 ( .A(n1784), .B(n4822), .Z(n6930) );
  NANDN U779 ( .A(x[768]), .B(y[768]), .Z(n4811) );
  ANDN U780 ( .B(y[769]), .A(x[769]), .Z(n4816) );
  ANDN U781 ( .B(n4811), .A(n4816), .Z(n6928) );
  ANDN U782 ( .B(x[767]), .A(y[767]), .Z(n4807) );
  NANDN U783 ( .A(y[768]), .B(x[768]), .Z(n1785) );
  NANDN U784 ( .A(n4807), .B(n1785), .Z(n6926) );
  NANDN U785 ( .A(x[766]), .B(y[766]), .Z(n4803) );
  ANDN U786 ( .B(y[767]), .A(x[767]), .Z(n4813) );
  ANDN U787 ( .B(n4803), .A(n4813), .Z(n6924) );
  ANDN U788 ( .B(x[765]), .A(y[765]), .Z(n1787) );
  ANDN U789 ( .B(x[766]), .A(y[766]), .Z(n4809) );
  OR U790 ( .A(n1787), .B(n4809), .Z(n6922) );
  NANDN U791 ( .A(x[765]), .B(y[765]), .Z(n4802) );
  ANDN U792 ( .B(y[764]), .A(x[764]), .Z(n4797) );
  ANDN U793 ( .B(n4802), .A(n4797), .Z(n6920) );
  NANDN U794 ( .A(y[763]), .B(x[763]), .Z(n4793) );
  XNOR U795 ( .A(x[764]), .B(y[764]), .Z(n260) );
  NAND U796 ( .A(n4793), .B(n260), .Z(n6918) );
  NANDN U797 ( .A(x[762]), .B(y[762]), .Z(n261) );
  ANDN U798 ( .B(y[763]), .A(x[763]), .Z(n4798) );
  ANDN U799 ( .B(n261), .A(n4798), .Z(n6916) );
  XOR U800 ( .A(x[762]), .B(y[762]), .Z(n4791) );
  NANDN U801 ( .A(y[761]), .B(x[761]), .Z(n4785) );
  NANDN U802 ( .A(n4791), .B(n4785), .Z(n6914) );
  NANDN U803 ( .A(x[760]), .B(y[760]), .Z(n1788) );
  ANDN U804 ( .B(y[761]), .A(x[761]), .Z(n4788) );
  ANDN U805 ( .B(n1788), .A(n4788), .Z(n6912) );
  NANDN U806 ( .A(y[759]), .B(x[759]), .Z(n4778) );
  XNOR U807 ( .A(y[760]), .B(x[760]), .Z(n262) );
  NAND U808 ( .A(n4778), .B(n262), .Z(n6910) );
  NANDN U809 ( .A(x[758]), .B(y[758]), .Z(n4775) );
  NANDN U810 ( .A(x[759]), .B(y[759]), .Z(n1789) );
  AND U811 ( .A(n4775), .B(n1789), .Z(n6908) );
  ANDN U812 ( .B(x[757]), .A(y[757]), .Z(n4773) );
  NANDN U813 ( .A(y[758]), .B(x[758]), .Z(n4779) );
  NANDN U814 ( .A(n4773), .B(n4779), .Z(n6906) );
  NANDN U815 ( .A(x[756]), .B(y[756]), .Z(n1790) );
  NANDN U816 ( .A(x[757]), .B(y[757]), .Z(n4776) );
  AND U817 ( .A(n1790), .B(n4776), .Z(n6904) );
  ANDN U818 ( .B(x[756]), .A(y[756]), .Z(n4770) );
  NANDN U819 ( .A(y[755]), .B(x[755]), .Z(n4765) );
  NANDN U820 ( .A(n4770), .B(n4765), .Z(n6902) );
  NANDN U821 ( .A(x[754]), .B(y[754]), .Z(n263) );
  NANDN U822 ( .A(x[755]), .B(y[755]), .Z(n1791) );
  AND U823 ( .A(n263), .B(n1791), .Z(n6900) );
  XOR U824 ( .A(x[754]), .B(y[754]), .Z(n4761) );
  NANDN U825 ( .A(y[753]), .B(x[753]), .Z(n4757) );
  NANDN U826 ( .A(n4761), .B(n4757), .Z(n6898) );
  NANDN U827 ( .A(x[752]), .B(y[752]), .Z(n264) );
  ANDN U828 ( .B(y[753]), .A(x[753]), .Z(n4763) );
  ANDN U829 ( .B(n264), .A(n4763), .Z(n6896) );
  XNOR U830 ( .A(x[752]), .B(y[752]), .Z(n1793) );
  NANDN U831 ( .A(y[751]), .B(x[751]), .Z(n4751) );
  NAND U832 ( .A(n1793), .B(n4751), .Z(n6894) );
  NANDN U833 ( .A(x[750]), .B(y[750]), .Z(n265) );
  NANDN U834 ( .A(x[751]), .B(y[751]), .Z(n1792) );
  AND U835 ( .A(n265), .B(n1792), .Z(n6892) );
  XOR U836 ( .A(x[750]), .B(y[750]), .Z(n4747) );
  NANDN U837 ( .A(y[749]), .B(x[749]), .Z(n4743) );
  NANDN U838 ( .A(n4747), .B(n4743), .Z(n6890) );
  NANDN U839 ( .A(x[748]), .B(y[748]), .Z(n266) );
  ANDN U840 ( .B(y[749]), .A(x[749]), .Z(n4749) );
  ANDN U841 ( .B(n266), .A(n4749), .Z(n6888) );
  XOR U842 ( .A(x[748]), .B(y[748]), .Z(n1794) );
  ANDN U843 ( .B(x[747]), .A(y[747]), .Z(n4737) );
  OR U844 ( .A(n1794), .B(n4737), .Z(n6886) );
  NANDN U845 ( .A(x[746]), .B(y[746]), .Z(n4733) );
  ANDN U846 ( .B(y[747]), .A(x[747]), .Z(n1795) );
  ANDN U847 ( .B(n4733), .A(n1795), .Z(n6884) );
  ANDN U848 ( .B(x[745]), .A(y[745]), .Z(n4728) );
  XNOR U849 ( .A(y[746]), .B(x[746]), .Z(n267) );
  NANDN U850 ( .A(n4728), .B(n267), .Z(n6882) );
  NANDN U851 ( .A(x[744]), .B(y[744]), .Z(n4725) );
  NANDN U852 ( .A(x[745]), .B(y[745]), .Z(n4732) );
  AND U853 ( .A(n4725), .B(n4732), .Z(n6880) );
  ANDN U854 ( .B(x[743]), .A(y[743]), .Z(n4721) );
  XNOR U855 ( .A(x[744]), .B(y[744]), .Z(n268) );
  NANDN U856 ( .A(n4721), .B(n268), .Z(n6878) );
  NANDN U857 ( .A(x[742]), .B(y[742]), .Z(n4717) );
  NANDN U858 ( .A(x[743]), .B(y[743]), .Z(n4726) );
  AND U859 ( .A(n4717), .B(n4726), .Z(n6876) );
  ANDN U860 ( .B(x[742]), .A(y[742]), .Z(n4723) );
  NANDN U861 ( .A(y[741]), .B(x[741]), .Z(n1796) );
  NANDN U862 ( .A(n4723), .B(n1796), .Z(n6874) );
  NANDN U863 ( .A(x[740]), .B(y[740]), .Z(n1798) );
  NANDN U864 ( .A(x[741]), .B(y[741]), .Z(n4716) );
  AND U865 ( .A(n1798), .B(n4716), .Z(n6872) );
  ANDN U866 ( .B(x[739]), .A(y[739]), .Z(n4709) );
  NANDN U867 ( .A(y[740]), .B(x[740]), .Z(n1797) );
  NANDN U868 ( .A(n4709), .B(n1797), .Z(n6870) );
  NANDN U869 ( .A(x[738]), .B(y[738]), .Z(n4705) );
  NANDN U870 ( .A(x[739]), .B(y[739]), .Z(n1799) );
  AND U871 ( .A(n4705), .B(n1799), .Z(n6868) );
  ANDN U872 ( .B(x[738]), .A(y[738]), .Z(n4710) );
  NANDN U873 ( .A(y[737]), .B(x[737]), .Z(n1800) );
  NANDN U874 ( .A(n4710), .B(n1800), .Z(n6866) );
  NANDN U875 ( .A(x[736]), .B(y[736]), .Z(n1802) );
  NANDN U876 ( .A(x[737]), .B(y[737]), .Z(n4704) );
  AND U877 ( .A(n1802), .B(n4704), .Z(n6864) );
  ANDN U878 ( .B(x[735]), .A(y[735]), .Z(n4697) );
  NANDN U879 ( .A(y[736]), .B(x[736]), .Z(n1801) );
  NANDN U880 ( .A(n4697), .B(n1801), .Z(n6862) );
  NANDN U881 ( .A(x[734]), .B(y[734]), .Z(n4693) );
  NANDN U882 ( .A(x[735]), .B(y[735]), .Z(n1803) );
  AND U883 ( .A(n4693), .B(n1803), .Z(n6860) );
  ANDN U884 ( .B(x[734]), .A(y[734]), .Z(n4698) );
  NANDN U885 ( .A(y[733]), .B(x[733]), .Z(n1805) );
  NANDN U886 ( .A(n4698), .B(n1805), .Z(n6858) );
  NANDN U887 ( .A(x[733]), .B(y[733]), .Z(n4692) );
  ANDN U888 ( .B(y[732]), .A(x[732]), .Z(n4687) );
  ANDN U889 ( .B(n4692), .A(n4687), .Z(n6856) );
  NANDN U890 ( .A(y[731]), .B(x[731]), .Z(n4683) );
  NANDN U891 ( .A(y[732]), .B(x[732]), .Z(n1804) );
  NAND U892 ( .A(n4683), .B(n1804), .Z(n6854) );
  NANDN U893 ( .A(x[730]), .B(y[730]), .Z(n269) );
  ANDN U894 ( .B(y[731]), .A(x[731]), .Z(n4688) );
  ANDN U895 ( .B(n269), .A(n4688), .Z(n6852) );
  XOR U896 ( .A(x[730]), .B(y[730]), .Z(n4681) );
  NANDN U897 ( .A(y[729]), .B(x[729]), .Z(n4675) );
  NANDN U898 ( .A(n4681), .B(n4675), .Z(n6850) );
  NANDN U899 ( .A(x[728]), .B(y[728]), .Z(n270) );
  ANDN U900 ( .B(y[729]), .A(x[729]), .Z(n4678) );
  ANDN U901 ( .B(n270), .A(n4678), .Z(n6848) );
  XOR U902 ( .A(x[728]), .B(y[728]), .Z(n4671) );
  NANDN U903 ( .A(y[727]), .B(x[727]), .Z(n1806) );
  NANDN U904 ( .A(n4671), .B(n1806), .Z(n6846) );
  ANDN U905 ( .B(y[726]), .A(x[726]), .Z(n4667) );
  ANDN U906 ( .B(y[727]), .A(x[727]), .Z(n4673) );
  NOR U907 ( .A(n4667), .B(n4673), .Z(n6844) );
  ANDN U908 ( .B(x[725]), .A(y[725]), .Z(n4660) );
  NANDN U909 ( .A(y[726]), .B(x[726]), .Z(n1807) );
  NANDN U910 ( .A(n4660), .B(n1807), .Z(n6842) );
  NANDN U911 ( .A(x[725]), .B(y[725]), .Z(n4663) );
  NANDN U912 ( .A(x[724]), .B(y[724]), .Z(n271) );
  NAND U913 ( .A(n4663), .B(n271), .Z(n6839) );
  ANDN U914 ( .B(x[724]), .A(y[724]), .Z(n4661) );
  NANDN U915 ( .A(y[723]), .B(x[723]), .Z(n4654) );
  NANDN U916 ( .A(n4661), .B(n4654), .Z(n6838) );
  NANDN U917 ( .A(x[722]), .B(y[722]), .Z(n4652) );
  ANDN U918 ( .B(y[723]), .A(x[723]), .Z(n4658) );
  ANDN U919 ( .B(n4652), .A(n4658), .Z(n6836) );
  ANDN U920 ( .B(x[721]), .A(y[721]), .Z(n4650) );
  XNOR U921 ( .A(x[722]), .B(y[722]), .Z(n272) );
  NANDN U922 ( .A(n4650), .B(n272), .Z(n6834) );
  NANDN U923 ( .A(x[721]), .B(y[721]), .Z(n4644) );
  NANDN U924 ( .A(x[720]), .B(y[720]), .Z(n273) );
  AND U925 ( .A(n4644), .B(n273), .Z(n6832) );
  NANDN U926 ( .A(y[719]), .B(x[719]), .Z(n4638) );
  NANDN U927 ( .A(y[720]), .B(x[720]), .Z(n274) );
  NAND U928 ( .A(n4638), .B(n274), .Z(n6830) );
  ANDN U929 ( .B(y[718]), .A(x[718]), .Z(n4633) );
  ANDN U930 ( .B(y[719]), .A(x[719]), .Z(n4642) );
  NOR U931 ( .A(n4633), .B(n4642), .Z(n6828) );
  NANDN U932 ( .A(y[717]), .B(x[717]), .Z(n4630) );
  XNOR U933 ( .A(x[718]), .B(y[718]), .Z(n275) );
  NAND U934 ( .A(n4630), .B(n275), .Z(n6826) );
  NANDN U935 ( .A(x[716]), .B(y[716]), .Z(n1808) );
  ANDN U936 ( .B(y[717]), .A(x[717]), .Z(n4636) );
  ANDN U937 ( .B(n1808), .A(n4636), .Z(n6824) );
  NANDN U938 ( .A(y[715]), .B(x[715]), .Z(n4623) );
  NANDN U939 ( .A(y[716]), .B(x[716]), .Z(n4631) );
  NAND U940 ( .A(n4623), .B(n4631), .Z(n6822) );
  NANDN U941 ( .A(x[714]), .B(y[714]), .Z(n276) );
  NANDN U942 ( .A(x[715]), .B(y[715]), .Z(n1809) );
  AND U943 ( .A(n276), .B(n1809), .Z(n6820) );
  ANDN U944 ( .B(x[713]), .A(y[713]), .Z(n4616) );
  XNOR U945 ( .A(x[714]), .B(y[714]), .Z(n4620) );
  NANDN U946 ( .A(n4616), .B(n4620), .Z(n6818) );
  NANDN U947 ( .A(x[712]), .B(y[712]), .Z(n277) );
  NANDN U948 ( .A(x[713]), .B(y[713]), .Z(n4621) );
  AND U949 ( .A(n277), .B(n4621), .Z(n6816) );
  ANDN U950 ( .B(x[711]), .A(y[711]), .Z(n1811) );
  XNOR U951 ( .A(x[712]), .B(y[712]), .Z(n4612) );
  NANDN U952 ( .A(n1811), .B(n4612), .Z(n6814) );
  NANDN U953 ( .A(x[711]), .B(y[711]), .Z(n4611) );
  ANDN U954 ( .B(y[710]), .A(x[710]), .Z(n4606) );
  ANDN U955 ( .B(n4611), .A(n4606), .Z(n6812) );
  ANDN U956 ( .B(x[710]), .A(y[710]), .Z(n1810) );
  NANDN U957 ( .A(y[709]), .B(x[709]), .Z(n4602) );
  NANDN U958 ( .A(n1810), .B(n4602), .Z(n6810) );
  ANDN U959 ( .B(y[708]), .A(x[708]), .Z(n4597) );
  ANDN U960 ( .B(y[709]), .A(x[709]), .Z(n4607) );
  NOR U961 ( .A(n4597), .B(n4607), .Z(n6808) );
  NANDN U962 ( .A(y[707]), .B(x[707]), .Z(n4594) );
  XNOR U963 ( .A(x[708]), .B(y[708]), .Z(n278) );
  NAND U964 ( .A(n4594), .B(n278), .Z(n6806) );
  ANDN U965 ( .B(y[706]), .A(x[706]), .Z(n4590) );
  ANDN U966 ( .B(y[707]), .A(x[707]), .Z(n4600) );
  NOR U967 ( .A(n4590), .B(n4600), .Z(n6804) );
  NANDN U968 ( .A(y[705]), .B(x[705]), .Z(n4586) );
  XNOR U969 ( .A(y[706]), .B(x[706]), .Z(n279) );
  NAND U970 ( .A(n4586), .B(n279), .Z(n6802) );
  NANDN U971 ( .A(x[704]), .B(y[704]), .Z(n1812) );
  ANDN U972 ( .B(y[705]), .A(x[705]), .Z(n4592) );
  ANDN U973 ( .B(n1812), .A(n4592), .Z(n6800) );
  NANDN U974 ( .A(y[703]), .B(x[703]), .Z(n4580) );
  NANDN U975 ( .A(y[704]), .B(x[704]), .Z(n4588) );
  NAND U976 ( .A(n4580), .B(n4588), .Z(n6798) );
  NANDN U977 ( .A(x[702]), .B(y[702]), .Z(n280) );
  NANDN U978 ( .A(x[703]), .B(y[703]), .Z(n1813) );
  AND U979 ( .A(n280), .B(n1813), .Z(n6796) );
  XOR U980 ( .A(x[702]), .B(y[702]), .Z(n4576) );
  NANDN U981 ( .A(y[701]), .B(x[701]), .Z(n4572) );
  NANDN U982 ( .A(n4576), .B(n4572), .Z(n6794) );
  NANDN U983 ( .A(x[700]), .B(y[700]), .Z(n1814) );
  ANDN U984 ( .B(y[701]), .A(x[701]), .Z(n4578) );
  ANDN U985 ( .B(n1814), .A(n4578), .Z(n6792) );
  NANDN U986 ( .A(y[699]), .B(x[699]), .Z(n1816) );
  NANDN U987 ( .A(y[700]), .B(x[700]), .Z(n4574) );
  NAND U988 ( .A(n1816), .B(n4574), .Z(n6790) );
  NANDN U989 ( .A(x[699]), .B(y[699]), .Z(n1815) );
  ANDN U990 ( .B(y[698]), .A(x[698]), .Z(n4564) );
  ANDN U991 ( .B(n1815), .A(n4564), .Z(n6788) );
  NANDN U992 ( .A(y[697]), .B(x[697]), .Z(n4560) );
  NANDN U993 ( .A(y[698]), .B(x[698]), .Z(n1817) );
  NAND U994 ( .A(n4560), .B(n1817), .Z(n6786) );
  NANDN U995 ( .A(x[696]), .B(y[696]), .Z(n1818) );
  ANDN U996 ( .B(y[697]), .A(x[697]), .Z(n4565) );
  ANDN U997 ( .B(n1818), .A(n4565), .Z(n6784) );
  NANDN U998 ( .A(y[695]), .B(x[695]), .Z(n1820) );
  NANDN U999 ( .A(y[696]), .B(x[696]), .Z(n4559) );
  NAND U1000 ( .A(n1820), .B(n4559), .Z(n6782) );
  NANDN U1001 ( .A(x[695]), .B(y[695]), .Z(n1819) );
  ANDN U1002 ( .B(y[694]), .A(x[694]), .Z(n4552) );
  ANDN U1003 ( .B(n1819), .A(n4552), .Z(n6780) );
  NANDN U1004 ( .A(y[693]), .B(x[693]), .Z(n4548) );
  NANDN U1005 ( .A(y[694]), .B(x[694]), .Z(n1821) );
  NAND U1006 ( .A(n4548), .B(n1821), .Z(n6778) );
  NANDN U1007 ( .A(x[692]), .B(y[692]), .Z(n4546) );
  ANDN U1008 ( .B(y[693]), .A(x[693]), .Z(n4553) );
  ANDN U1009 ( .B(n4546), .A(n4553), .Z(n6776) );
  ANDN U1010 ( .B(x[691]), .A(y[691]), .Z(n4544) );
  NANDN U1011 ( .A(y[692]), .B(x[692]), .Z(n4550) );
  NANDN U1012 ( .A(n4544), .B(n4550), .Z(n6774) );
  NANDN U1013 ( .A(x[691]), .B(y[691]), .Z(n4542) );
  NANDN U1014 ( .A(x[690]), .B(y[690]), .Z(n281) );
  AND U1015 ( .A(n4542), .B(n281), .Z(n6772) );
  ANDN U1016 ( .B(x[689]), .A(y[689]), .Z(n4534) );
  NANDN U1017 ( .A(y[690]), .B(x[690]), .Z(n4540) );
  NANDN U1018 ( .A(n4534), .B(n4540), .Z(n6770) );
  NANDN U1019 ( .A(x[688]), .B(y[688]), .Z(n1823) );
  NANDN U1020 ( .A(x[689]), .B(y[689]), .Z(n4536) );
  AND U1021 ( .A(n1823), .B(n4536), .Z(n6768) );
  ANDN U1022 ( .B(x[687]), .A(y[687]), .Z(n4526) );
  XNOR U1023 ( .A(y[688]), .B(x[688]), .Z(n282) );
  NANDN U1024 ( .A(n4526), .B(n282), .Z(n6766) );
  NANDN U1025 ( .A(x[686]), .B(y[686]), .Z(n4522) );
  NANDN U1026 ( .A(x[687]), .B(y[687]), .Z(n1822) );
  AND U1027 ( .A(n4522), .B(n1822), .Z(n6764) );
  ANDN U1028 ( .B(x[685]), .A(y[685]), .Z(n4520) );
  ANDN U1029 ( .B(x[686]), .A(y[686]), .Z(n4527) );
  OR U1030 ( .A(n4520), .B(n4527), .Z(n6762) );
  NANDN U1031 ( .A(x[684]), .B(y[684]), .Z(n283) );
  NANDN U1032 ( .A(x[685]), .B(y[685]), .Z(n4521) );
  AND U1033 ( .A(n283), .B(n4521), .Z(n6760) );
  XNOR U1034 ( .A(x[684]), .B(y[684]), .Z(n4514) );
  NANDN U1035 ( .A(y[683]), .B(x[683]), .Z(n4510) );
  NAND U1036 ( .A(n4514), .B(n4510), .Z(n6758) );
  NANDN U1037 ( .A(x[682]), .B(y[682]), .Z(n284) );
  NANDN U1038 ( .A(x[683]), .B(y[683]), .Z(n4515) );
  AND U1039 ( .A(n284), .B(n4515), .Z(n6756) );
  XNOR U1040 ( .A(x[682]), .B(y[682]), .Z(n4506) );
  NANDN U1041 ( .A(y[681]), .B(x[681]), .Z(n1824) );
  NAND U1042 ( .A(n4506), .B(n1824), .Z(n6754) );
  NANDN U1043 ( .A(x[680]), .B(y[680]), .Z(n285) );
  NANDN U1044 ( .A(x[681]), .B(y[681]), .Z(n4505) );
  AND U1045 ( .A(n285), .B(n4505), .Z(n6752) );
  XNOR U1046 ( .A(x[680]), .B(y[680]), .Z(n4500) );
  NANDN U1047 ( .A(y[679]), .B(x[679]), .Z(n4495) );
  NAND U1048 ( .A(n4500), .B(n4495), .Z(n6750) );
  NANDN U1049 ( .A(x[678]), .B(y[678]), .Z(n286) );
  ANDN U1050 ( .B(y[679]), .A(x[679]), .Z(n4501) );
  ANDN U1051 ( .B(n286), .A(n4501), .Z(n6748) );
  ANDN U1052 ( .B(x[677]), .A(y[677]), .Z(n4488) );
  XNOR U1053 ( .A(x[678]), .B(y[678]), .Z(n4492) );
  NANDN U1054 ( .A(n4488), .B(n4492), .Z(n6746) );
  NANDN U1055 ( .A(x[676]), .B(y[676]), .Z(n287) );
  NANDN U1056 ( .A(x[677]), .B(y[677]), .Z(n4493) );
  AND U1057 ( .A(n287), .B(n4493), .Z(n6744) );
  XNOR U1058 ( .A(x[676]), .B(y[676]), .Z(n4484) );
  NANDN U1059 ( .A(y[675]), .B(x[675]), .Z(n1826) );
  NAND U1060 ( .A(n4484), .B(n1826), .Z(n6742) );
  NANDN U1061 ( .A(x[674]), .B(y[674]), .Z(n288) );
  NANDN U1062 ( .A(x[675]), .B(y[675]), .Z(n4483) );
  AND U1063 ( .A(n288), .B(n4483), .Z(n6740) );
  ANDN U1064 ( .B(x[673]), .A(y[673]), .Z(n4474) );
  XNOR U1065 ( .A(x[674]), .B(y[674]), .Z(n4478) );
  NANDN U1066 ( .A(n4474), .B(n4478), .Z(n6738) );
  NANDN U1067 ( .A(x[672]), .B(y[672]), .Z(n289) );
  ANDN U1068 ( .B(y[673]), .A(x[673]), .Z(n4480) );
  ANDN U1069 ( .B(n289), .A(n4480), .Z(n6736) );
  XNOR U1070 ( .A(x[672]), .B(y[672]), .Z(n4470) );
  NANDN U1071 ( .A(y[671]), .B(x[671]), .Z(n1828) );
  NAND U1072 ( .A(n4470), .B(n1828), .Z(n6734) );
  NANDN U1073 ( .A(x[670]), .B(y[670]), .Z(n1830) );
  NANDN U1074 ( .A(x[671]), .B(y[671]), .Z(n4469) );
  AND U1075 ( .A(n1830), .B(n4469), .Z(n6732) );
  ANDN U1076 ( .B(x[669]), .A(y[669]), .Z(n4462) );
  NANDN U1077 ( .A(y[670]), .B(x[670]), .Z(n1829) );
  NANDN U1078 ( .A(n4462), .B(n1829), .Z(n6730) );
  NANDN U1079 ( .A(x[668]), .B(y[668]), .Z(n4458) );
  NANDN U1080 ( .A(x[669]), .B(y[669]), .Z(n1831) );
  AND U1081 ( .A(n4458), .B(n1831), .Z(n6728) );
  ANDN U1082 ( .B(x[667]), .A(y[667]), .Z(n1832) );
  ANDN U1083 ( .B(x[668]), .A(y[668]), .Z(n4463) );
  OR U1084 ( .A(n1832), .B(n4463), .Z(n6726) );
  NANDN U1085 ( .A(x[666]), .B(y[666]), .Z(n290) );
  NANDN U1086 ( .A(x[667]), .B(y[667]), .Z(n4457) );
  AND U1087 ( .A(n290), .B(n4457), .Z(n6724) );
  XNOR U1088 ( .A(x[666]), .B(y[666]), .Z(n4452) );
  NANDN U1089 ( .A(y[665]), .B(x[665]), .Z(n4448) );
  NAND U1090 ( .A(n4452), .B(n4448), .Z(n6722) );
  NANDN U1091 ( .A(x[665]), .B(y[665]), .Z(n4451) );
  ANDN U1092 ( .B(y[664]), .A(x[664]), .Z(n4446) );
  ANDN U1093 ( .B(n4451), .A(n4446), .Z(n6720) );
  NANDN U1094 ( .A(y[663]), .B(x[663]), .Z(n1835) );
  NANDN U1095 ( .A(y[664]), .B(x[664]), .Z(n4449) );
  NAND U1096 ( .A(n1835), .B(n4449), .Z(n6718) );
  ANDN U1097 ( .B(y[662]), .A(x[662]), .Z(n4438) );
  ANDN U1098 ( .B(y[663]), .A(x[663]), .Z(n4443) );
  NOR U1099 ( .A(n4438), .B(n4443), .Z(n6716) );
  NANDN U1100 ( .A(y[661]), .B(x[661]), .Z(n4434) );
  NANDN U1101 ( .A(y[662]), .B(x[662]), .Z(n1834) );
  NAND U1102 ( .A(n4434), .B(n1834), .Z(n6714) );
  ANDN U1103 ( .B(y[660]), .A(x[660]), .Z(n4429) );
  ANDN U1104 ( .B(y[661]), .A(x[661]), .Z(n4439) );
  NOR U1105 ( .A(n4429), .B(n4439), .Z(n6713) );
  NANDN U1106 ( .A(y[659]), .B(x[659]), .Z(n4427) );
  NANDN U1107 ( .A(y[660]), .B(x[660]), .Z(n4433) );
  NAND U1108 ( .A(n4427), .B(n4433), .Z(n6712) );
  ANDN U1109 ( .B(y[658]), .A(x[658]), .Z(n4424) );
  ANDN U1110 ( .B(y[659]), .A(x[659]), .Z(n4432) );
  NOR U1111 ( .A(n4424), .B(n4432), .Z(n6711) );
  NANDN U1112 ( .A(y[658]), .B(x[658]), .Z(n6710) );
  NANDN U1113 ( .A(x[655]), .B(y[655]), .Z(n4420) );
  ANDN U1114 ( .B(y[654]), .A(x[654]), .Z(n6706) );
  ANDN U1115 ( .B(n4420), .A(n6706), .Z(n1059) );
  NANDN U1116 ( .A(y[653]), .B(x[653]), .Z(n4411) );
  NANDN U1117 ( .A(y[654]), .B(x[654]), .Z(n1838) );
  NAND U1118 ( .A(n4411), .B(n1838), .Z(n6705) );
  ANDN U1119 ( .B(y[652]), .A(x[652]), .Z(n4406) );
  ANDN U1120 ( .B(y[653]), .A(x[653]), .Z(n4415) );
  NOR U1121 ( .A(n4406), .B(n4415), .Z(n6704) );
  NANDN U1122 ( .A(y[651]), .B(x[651]), .Z(n4403) );
  NANDN U1123 ( .A(y[652]), .B(x[652]), .Z(n4410) );
  NAND U1124 ( .A(n4403), .B(n4410), .Z(n6703) );
  NANDN U1125 ( .A(x[650]), .B(y[650]), .Z(n291) );
  ANDN U1126 ( .B(y[651]), .A(x[651]), .Z(n4409) );
  ANDN U1127 ( .B(n291), .A(n4409), .Z(n6702) );
  XOR U1128 ( .A(x[650]), .B(y[650]), .Z(n4399) );
  NANDN U1129 ( .A(y[649]), .B(x[649]), .Z(n4395) );
  NANDN U1130 ( .A(n4399), .B(n4395), .Z(n6701) );
  NANDN U1131 ( .A(x[648]), .B(y[648]), .Z(n292) );
  ANDN U1132 ( .B(y[649]), .A(x[649]), .Z(n4401) );
  ANDN U1133 ( .B(n292), .A(n4401), .Z(n6700) );
  XOR U1134 ( .A(x[648]), .B(y[648]), .Z(n4393) );
  NANDN U1135 ( .A(y[647]), .B(x[647]), .Z(n4387) );
  NANDN U1136 ( .A(n4393), .B(n4387), .Z(n6699) );
  NANDN U1137 ( .A(x[646]), .B(y[646]), .Z(n293) );
  ANDN U1138 ( .B(y[647]), .A(x[647]), .Z(n4390) );
  ANDN U1139 ( .B(n293), .A(n4390), .Z(n6698) );
  XOR U1140 ( .A(x[646]), .B(y[646]), .Z(n4383) );
  NANDN U1141 ( .A(y[645]), .B(x[645]), .Z(n1840) );
  NANDN U1142 ( .A(n4383), .B(n1840), .Z(n6697) );
  ANDN U1143 ( .B(y[644]), .A(x[644]), .Z(n4377) );
  ANDN U1144 ( .B(y[645]), .A(x[645]), .Z(n4385) );
  NOR U1145 ( .A(n4377), .B(n4385), .Z(n6695) );
  NANDN U1146 ( .A(y[643]), .B(x[643]), .Z(n4373) );
  NANDN U1147 ( .A(y[644]), .B(x[644]), .Z(n1839) );
  NAND U1148 ( .A(n4373), .B(n1839), .Z(n6693) );
  ANDN U1149 ( .B(y[642]), .A(x[642]), .Z(n4368) );
  ANDN U1150 ( .B(y[643]), .A(x[643]), .Z(n4378) );
  NOR U1151 ( .A(n4368), .B(n4378), .Z(n6691) );
  NANDN U1152 ( .A(y[641]), .B(x[641]), .Z(n4365) );
  NANDN U1153 ( .A(y[642]), .B(x[642]), .Z(n4372) );
  NAND U1154 ( .A(n4365), .B(n4372), .Z(n6689) );
  ANDN U1155 ( .B(y[640]), .A(x[640]), .Z(n4363) );
  ANDN U1156 ( .B(y[641]), .A(x[641]), .Z(n4371) );
  NOR U1157 ( .A(n4363), .B(n4371), .Z(n6687) );
  NANDN U1158 ( .A(y[639]), .B(x[639]), .Z(n1842) );
  NANDN U1159 ( .A(y[640]), .B(x[640]), .Z(n4366) );
  NAND U1160 ( .A(n1842), .B(n4366), .Z(n6685) );
  ANDN U1161 ( .B(y[638]), .A(x[638]), .Z(n4355) );
  ANDN U1162 ( .B(y[639]), .A(x[639]), .Z(n4360) );
  NOR U1163 ( .A(n4355), .B(n4360), .Z(n6683) );
  NANDN U1164 ( .A(y[637]), .B(x[637]), .Z(n4351) );
  NANDN U1165 ( .A(y[638]), .B(x[638]), .Z(n1841) );
  NAND U1166 ( .A(n4351), .B(n1841), .Z(n6681) );
  ANDN U1167 ( .B(y[636]), .A(x[636]), .Z(n4346) );
  ANDN U1168 ( .B(y[637]), .A(x[637]), .Z(n4356) );
  NOR U1169 ( .A(n4346), .B(n4356), .Z(n6679) );
  NANDN U1170 ( .A(y[635]), .B(x[635]), .Z(n4343) );
  NANDN U1171 ( .A(y[636]), .B(x[636]), .Z(n4350) );
  NAND U1172 ( .A(n4343), .B(n4350), .Z(n6677) );
  ANDN U1173 ( .B(y[634]), .A(x[634]), .Z(n4341) );
  ANDN U1174 ( .B(y[635]), .A(x[635]), .Z(n4349) );
  NOR U1175 ( .A(n4341), .B(n4349), .Z(n6675) );
  NANDN U1176 ( .A(y[633]), .B(x[633]), .Z(n1844) );
  NANDN U1177 ( .A(y[634]), .B(x[634]), .Z(n4344) );
  NAND U1178 ( .A(n1844), .B(n4344), .Z(n6673) );
  ANDN U1179 ( .B(y[632]), .A(x[632]), .Z(n4333) );
  ANDN U1180 ( .B(y[633]), .A(x[633]), .Z(n4338) );
  NOR U1181 ( .A(n4333), .B(n4338), .Z(n6671) );
  NANDN U1182 ( .A(y[631]), .B(x[631]), .Z(n4329) );
  NANDN U1183 ( .A(y[632]), .B(x[632]), .Z(n1843) );
  NAND U1184 ( .A(n4329), .B(n1843), .Z(n6669) );
  NANDN U1185 ( .A(x[630]), .B(y[630]), .Z(n294) );
  ANDN U1186 ( .B(y[631]), .A(x[631]), .Z(n4334) );
  ANDN U1187 ( .B(n294), .A(n4334), .Z(n6667) );
  XOR U1188 ( .A(x[630]), .B(y[630]), .Z(n4327) );
  NANDN U1189 ( .A(y[629]), .B(x[629]), .Z(n4321) );
  NANDN U1190 ( .A(n4327), .B(n4321), .Z(n6665) );
  ANDN U1191 ( .B(y[628]), .A(x[628]), .Z(n4319) );
  ANDN U1192 ( .B(y[629]), .A(x[629]), .Z(n4324) );
  NOR U1193 ( .A(n4319), .B(n4324), .Z(n6663) );
  NANDN U1194 ( .A(y[627]), .B(x[627]), .Z(n1845) );
  NANDN U1195 ( .A(y[628]), .B(x[628]), .Z(n4322) );
  NAND U1196 ( .A(n1845), .B(n4322), .Z(n6661) );
  NANDN U1197 ( .A(x[626]), .B(y[626]), .Z(n295) );
  ANDN U1198 ( .B(y[627]), .A(x[627]), .Z(n4316) );
  ANDN U1199 ( .B(n295), .A(n4316), .Z(n6659) );
  XOR U1200 ( .A(x[626]), .B(y[626]), .Z(n4311) );
  NANDN U1201 ( .A(y[625]), .B(x[625]), .Z(n4307) );
  NANDN U1202 ( .A(n4311), .B(n4307), .Z(n6657) );
  ANDN U1203 ( .B(y[624]), .A(x[624]), .Z(n4302) );
  ANDN U1204 ( .B(y[625]), .A(x[625]), .Z(n4312) );
  NOR U1205 ( .A(n4302), .B(n4312), .Z(n6655) );
  NANDN U1206 ( .A(y[623]), .B(x[623]), .Z(n4299) );
  NANDN U1207 ( .A(y[624]), .B(x[624]), .Z(n4309) );
  NAND U1208 ( .A(n4299), .B(n4309), .Z(n6653) );
  ANDN U1209 ( .B(y[622]), .A(x[622]), .Z(n4297) );
  ANDN U1210 ( .B(y[623]), .A(x[623]), .Z(n4305) );
  NOR U1211 ( .A(n4297), .B(n4305), .Z(n6651) );
  NANDN U1212 ( .A(y[621]), .B(x[621]), .Z(n1848) );
  NANDN U1213 ( .A(y[622]), .B(x[622]), .Z(n4300) );
  NAND U1214 ( .A(n1848), .B(n4300), .Z(n6649) );
  ANDN U1215 ( .B(y[620]), .A(x[620]), .Z(n4289) );
  ANDN U1216 ( .B(y[621]), .A(x[621]), .Z(n4294) );
  NOR U1217 ( .A(n4289), .B(n4294), .Z(n6647) );
  NANDN U1218 ( .A(y[619]), .B(x[619]), .Z(n4285) );
  NANDN U1219 ( .A(y[620]), .B(x[620]), .Z(n1847) );
  NAND U1220 ( .A(n4285), .B(n1847), .Z(n6645) );
  ANDN U1221 ( .B(y[618]), .A(x[618]), .Z(n4280) );
  ANDN U1222 ( .B(y[619]), .A(x[619]), .Z(n4290) );
  NOR U1223 ( .A(n4280), .B(n4290), .Z(n6643) );
  NANDN U1224 ( .A(y[617]), .B(x[617]), .Z(n4277) );
  NANDN U1225 ( .A(y[618]), .B(x[618]), .Z(n4284) );
  NAND U1226 ( .A(n4277), .B(n4284), .Z(n6641) );
  NANDN U1227 ( .A(x[616]), .B(y[616]), .Z(n296) );
  ANDN U1228 ( .B(y[617]), .A(x[617]), .Z(n4283) );
  ANDN U1229 ( .B(n296), .A(n4283), .Z(n6639) );
  XOR U1230 ( .A(x[616]), .B(y[616]), .Z(n4273) );
  NANDN U1231 ( .A(y[615]), .B(x[615]), .Z(n1850) );
  NANDN U1232 ( .A(n4273), .B(n1850), .Z(n6637) );
  ANDN U1233 ( .B(y[614]), .A(x[614]), .Z(n4267) );
  ANDN U1234 ( .B(y[615]), .A(x[615]), .Z(n4275) );
  NOR U1235 ( .A(n4267), .B(n4275), .Z(n6635) );
  NANDN U1236 ( .A(y[613]), .B(x[613]), .Z(n4263) );
  NANDN U1237 ( .A(y[614]), .B(x[614]), .Z(n1849) );
  NAND U1238 ( .A(n4263), .B(n1849), .Z(n6633) );
  ANDN U1239 ( .B(y[612]), .A(x[612]), .Z(n4258) );
  ANDN U1240 ( .B(y[613]), .A(x[613]), .Z(n4268) );
  NOR U1241 ( .A(n4258), .B(n4268), .Z(n6631) );
  NANDN U1242 ( .A(y[611]), .B(x[611]), .Z(n4255) );
  NANDN U1243 ( .A(y[612]), .B(x[612]), .Z(n4262) );
  NAND U1244 ( .A(n4255), .B(n4262), .Z(n6629) );
  NANDN U1245 ( .A(x[610]), .B(y[610]), .Z(n297) );
  ANDN U1246 ( .B(y[611]), .A(x[611]), .Z(n4261) );
  ANDN U1247 ( .B(n297), .A(n4261), .Z(n6627) );
  XOR U1248 ( .A(x[610]), .B(y[610]), .Z(n4251) );
  NANDN U1249 ( .A(y[609]), .B(x[609]), .Z(n1851) );
  NANDN U1250 ( .A(n4251), .B(n1851), .Z(n6625) );
  NANDN U1251 ( .A(x[608]), .B(y[608]), .Z(n298) );
  ANDN U1252 ( .B(y[609]), .A(x[609]), .Z(n4253) );
  ANDN U1253 ( .B(n298), .A(n4253), .Z(n6623) );
  XOR U1254 ( .A(x[608]), .B(y[608]), .Z(n4245) );
  NANDN U1255 ( .A(y[607]), .B(x[607]), .Z(n4241) );
  NANDN U1256 ( .A(n4245), .B(n4241), .Z(n6621) );
  ANDN U1257 ( .B(y[606]), .A(x[606]), .Z(n4236) );
  ANDN U1258 ( .B(y[607]), .A(x[607]), .Z(n4246) );
  NOR U1259 ( .A(n4236), .B(n4246), .Z(n6619) );
  NANDN U1260 ( .A(y[605]), .B(x[605]), .Z(n4233) );
  NANDN U1261 ( .A(y[606]), .B(x[606]), .Z(n4243) );
  NAND U1262 ( .A(n4233), .B(n4243), .Z(n6617) );
  ANDN U1263 ( .B(y[604]), .A(x[604]), .Z(n4231) );
  ANDN U1264 ( .B(y[605]), .A(x[605]), .Z(n4239) );
  NOR U1265 ( .A(n4231), .B(n4239), .Z(n6615) );
  NANDN U1266 ( .A(y[603]), .B(x[603]), .Z(n1854) );
  NANDN U1267 ( .A(y[604]), .B(x[604]), .Z(n4234) );
  NAND U1268 ( .A(n1854), .B(n4234), .Z(n6613) );
  ANDN U1269 ( .B(y[602]), .A(x[602]), .Z(n4223) );
  ANDN U1270 ( .B(y[603]), .A(x[603]), .Z(n4228) );
  NOR U1271 ( .A(n4223), .B(n4228), .Z(n6611) );
  NANDN U1272 ( .A(y[601]), .B(x[601]), .Z(n4219) );
  NANDN U1273 ( .A(y[602]), .B(x[602]), .Z(n1853) );
  NAND U1274 ( .A(n4219), .B(n1853), .Z(n6609) );
  ANDN U1275 ( .B(y[600]), .A(x[600]), .Z(n4214) );
  ANDN U1276 ( .B(y[601]), .A(x[601]), .Z(n4224) );
  NOR U1277 ( .A(n4214), .B(n4224), .Z(n6607) );
  NANDN U1278 ( .A(y[599]), .B(x[599]), .Z(n4211) );
  NANDN U1279 ( .A(y[600]), .B(x[600]), .Z(n4218) );
  NAND U1280 ( .A(n4211), .B(n4218), .Z(n6605) );
  ANDN U1281 ( .B(y[598]), .A(x[598]), .Z(n4209) );
  ANDN U1282 ( .B(y[599]), .A(x[599]), .Z(n4217) );
  NOR U1283 ( .A(n4209), .B(n4217), .Z(n6603) );
  NANDN U1284 ( .A(y[597]), .B(x[597]), .Z(n1856) );
  NANDN U1285 ( .A(y[598]), .B(x[598]), .Z(n4212) );
  NAND U1286 ( .A(n1856), .B(n4212), .Z(n6601) );
  ANDN U1287 ( .B(y[596]), .A(x[596]), .Z(n4201) );
  ANDN U1288 ( .B(y[597]), .A(x[597]), .Z(n4206) );
  NOR U1289 ( .A(n4201), .B(n4206), .Z(n6599) );
  NANDN U1290 ( .A(y[595]), .B(x[595]), .Z(n4197) );
  NANDN U1291 ( .A(y[596]), .B(x[596]), .Z(n1855) );
  NAND U1292 ( .A(n4197), .B(n1855), .Z(n6597) );
  ANDN U1293 ( .B(y[594]), .A(x[594]), .Z(n4192) );
  ANDN U1294 ( .B(y[595]), .A(x[595]), .Z(n4202) );
  NOR U1295 ( .A(n4192), .B(n4202), .Z(n6595) );
  NANDN U1296 ( .A(y[593]), .B(x[593]), .Z(n4189) );
  NANDN U1297 ( .A(y[594]), .B(x[594]), .Z(n4196) );
  NAND U1298 ( .A(n4189), .B(n4196), .Z(n6593) );
  ANDN U1299 ( .B(y[592]), .A(x[592]), .Z(n4187) );
  ANDN U1300 ( .B(y[593]), .A(x[593]), .Z(n4195) );
  NOR U1301 ( .A(n4187), .B(n4195), .Z(n6591) );
  NANDN U1302 ( .A(y[591]), .B(x[591]), .Z(n1858) );
  NANDN U1303 ( .A(y[592]), .B(x[592]), .Z(n4190) );
  NAND U1304 ( .A(n1858), .B(n4190), .Z(n6589) );
  ANDN U1305 ( .B(y[590]), .A(x[590]), .Z(n4179) );
  ANDN U1306 ( .B(y[591]), .A(x[591]), .Z(n4184) );
  NOR U1307 ( .A(n4179), .B(n4184), .Z(n6587) );
  NANDN U1308 ( .A(y[589]), .B(x[589]), .Z(n4175) );
  NANDN U1309 ( .A(y[590]), .B(x[590]), .Z(n1857) );
  NAND U1310 ( .A(n4175), .B(n1857), .Z(n6585) );
  ANDN U1311 ( .B(y[588]), .A(x[588]), .Z(n4170) );
  ANDN U1312 ( .B(y[589]), .A(x[589]), .Z(n4180) );
  NOR U1313 ( .A(n4170), .B(n4180), .Z(n6583) );
  NANDN U1314 ( .A(y[587]), .B(x[587]), .Z(n4167) );
  NANDN U1315 ( .A(y[588]), .B(x[588]), .Z(n4174) );
  NAND U1316 ( .A(n4167), .B(n4174), .Z(n6581) );
  NANDN U1317 ( .A(x[586]), .B(y[586]), .Z(n299) );
  ANDN U1318 ( .B(y[587]), .A(x[587]), .Z(n4173) );
  ANDN U1319 ( .B(n299), .A(n4173), .Z(n6579) );
  XOR U1320 ( .A(x[586]), .B(y[586]), .Z(n4163) );
  NANDN U1321 ( .A(y[585]), .B(x[585]), .Z(n1859) );
  NANDN U1322 ( .A(n4163), .B(n1859), .Z(n6577) );
  NANDN U1323 ( .A(x[584]), .B(y[584]), .Z(n300) );
  ANDN U1324 ( .B(y[585]), .A(x[585]), .Z(n4165) );
  ANDN U1325 ( .B(n300), .A(n4165), .Z(n6575) );
  XOR U1326 ( .A(x[584]), .B(y[584]), .Z(n4157) );
  NANDN U1327 ( .A(y[583]), .B(x[583]), .Z(n4153) );
  NANDN U1328 ( .A(n4157), .B(n4153), .Z(n6573) );
  NANDN U1329 ( .A(x[582]), .B(y[582]), .Z(n301) );
  ANDN U1330 ( .B(y[583]), .A(x[583]), .Z(n4158) );
  ANDN U1331 ( .B(n301), .A(n4158), .Z(n6571) );
  XOR U1332 ( .A(x[582]), .B(y[582]), .Z(n4151) );
  NANDN U1333 ( .A(y[581]), .B(x[581]), .Z(n4145) );
  NANDN U1334 ( .A(n4151), .B(n4145), .Z(n6569) );
  NANDN U1335 ( .A(x[580]), .B(y[580]), .Z(n302) );
  ANDN U1336 ( .B(y[581]), .A(x[581]), .Z(n4148) );
  ANDN U1337 ( .B(n302), .A(n4148), .Z(n6567) );
  XOR U1338 ( .A(x[580]), .B(y[580]), .Z(n4141) );
  NANDN U1339 ( .A(y[579]), .B(x[579]), .Z(n1862) );
  NANDN U1340 ( .A(n4141), .B(n1862), .Z(n6565) );
  ANDN U1341 ( .B(y[578]), .A(x[578]), .Z(n4137) );
  ANDN U1342 ( .B(y[579]), .A(x[579]), .Z(n4143) );
  NOR U1343 ( .A(n4137), .B(n4143), .Z(n6563) );
  NANDN U1344 ( .A(y[577]), .B(x[577]), .Z(n4135) );
  NANDN U1345 ( .A(y[578]), .B(x[578]), .Z(n1861) );
  NAND U1346 ( .A(n4135), .B(n1861), .Z(n6561) );
  NANDN U1347 ( .A(x[577]), .B(y[577]), .Z(n304) );
  NANDN U1348 ( .A(x[576]), .B(y[576]), .Z(n303) );
  NAND U1349 ( .A(n304), .B(n303), .Z(n6558) );
  NANDN U1350 ( .A(x[574]), .B(y[574]), .Z(n305) );
  ANDN U1351 ( .B(y[575]), .A(x[575]), .Z(n4126) );
  ANDN U1352 ( .B(n305), .A(n4126), .Z(n6555) );
  NANDN U1353 ( .A(y[573]), .B(x[573]), .Z(n4121) );
  NANDN U1354 ( .A(y[574]), .B(x[574]), .Z(n306) );
  NAND U1355 ( .A(n4121), .B(n306), .Z(n6553) );
  ANDN U1356 ( .B(y[572]), .A(x[572]), .Z(n4116) );
  ANDN U1357 ( .B(y[573]), .A(x[573]), .Z(n4125) );
  NOR U1358 ( .A(n4116), .B(n4125), .Z(n6551) );
  NANDN U1359 ( .A(y[571]), .B(x[571]), .Z(n4113) );
  NANDN U1360 ( .A(y[572]), .B(x[572]), .Z(n4120) );
  NAND U1361 ( .A(n4113), .B(n4120), .Z(n6549) );
  ANDN U1362 ( .B(y[570]), .A(x[570]), .Z(n4109) );
  ANDN U1363 ( .B(y[571]), .A(x[571]), .Z(n4119) );
  NOR U1364 ( .A(n4109), .B(n4119), .Z(n6547) );
  NANDN U1365 ( .A(y[569]), .B(x[569]), .Z(n4105) );
  NANDN U1366 ( .A(y[570]), .B(x[570]), .Z(n4114) );
  NAND U1367 ( .A(n4105), .B(n4114), .Z(n6545) );
  ANDN U1368 ( .B(y[568]), .A(x[568]), .Z(n4100) );
  ANDN U1369 ( .B(y[569]), .A(x[569]), .Z(n4111) );
  NOR U1370 ( .A(n4100), .B(n4111), .Z(n6543) );
  NANDN U1371 ( .A(y[567]), .B(x[567]), .Z(n4097) );
  NANDN U1372 ( .A(y[568]), .B(x[568]), .Z(n4104) );
  NAND U1373 ( .A(n4097), .B(n4104), .Z(n6541) );
  ANDN U1374 ( .B(y[566]), .A(x[566]), .Z(n4095) );
  ANDN U1375 ( .B(y[567]), .A(x[567]), .Z(n4103) );
  NOR U1376 ( .A(n4095), .B(n4103), .Z(n6539) );
  NANDN U1377 ( .A(y[565]), .B(x[565]), .Z(n1864) );
  NANDN U1378 ( .A(y[566]), .B(x[566]), .Z(n4098) );
  NAND U1379 ( .A(n1864), .B(n4098), .Z(n6537) );
  ANDN U1380 ( .B(y[564]), .A(x[564]), .Z(n4087) );
  ANDN U1381 ( .B(y[565]), .A(x[565]), .Z(n4092) );
  NOR U1382 ( .A(n4087), .B(n4092), .Z(n6535) );
  NANDN U1383 ( .A(y[563]), .B(x[563]), .Z(n4083) );
  NANDN U1384 ( .A(y[564]), .B(x[564]), .Z(n1863) );
  NAND U1385 ( .A(n4083), .B(n1863), .Z(n6533) );
  NANDN U1386 ( .A(x[562]), .B(y[562]), .Z(n307) );
  ANDN U1387 ( .B(y[563]), .A(x[563]), .Z(n4088) );
  ANDN U1388 ( .B(n307), .A(n4088), .Z(n6531) );
  XOR U1389 ( .A(x[562]), .B(y[562]), .Z(n4081) );
  NANDN U1390 ( .A(y[561]), .B(x[561]), .Z(n4075) );
  NANDN U1391 ( .A(n4081), .B(n4075), .Z(n6529) );
  NANDN U1392 ( .A(x[560]), .B(y[560]), .Z(n308) );
  ANDN U1393 ( .B(y[561]), .A(x[561]), .Z(n4078) );
  ANDN U1394 ( .B(n308), .A(n4078), .Z(n6527) );
  XOR U1395 ( .A(x[560]), .B(y[560]), .Z(n4071) );
  NANDN U1396 ( .A(y[559]), .B(x[559]), .Z(n1866) );
  NANDN U1397 ( .A(n4071), .B(n1866), .Z(n6525) );
  ANDN U1398 ( .B(y[558]), .A(x[558]), .Z(n4065) );
  ANDN U1399 ( .B(y[559]), .A(x[559]), .Z(n4073) );
  NOR U1400 ( .A(n4065), .B(n4073), .Z(n6523) );
  NANDN U1401 ( .A(y[557]), .B(x[557]), .Z(n4061) );
  NANDN U1402 ( .A(y[558]), .B(x[558]), .Z(n1865) );
  NAND U1403 ( .A(n4061), .B(n1865), .Z(n6521) );
  ANDN U1404 ( .B(y[556]), .A(x[556]), .Z(n4056) );
  ANDN U1405 ( .B(y[557]), .A(x[557]), .Z(n4066) );
  NOR U1406 ( .A(n4056), .B(n4066), .Z(n6519) );
  NANDN U1407 ( .A(y[555]), .B(x[555]), .Z(n4053) );
  NANDN U1408 ( .A(y[556]), .B(x[556]), .Z(n4060) );
  NAND U1409 ( .A(n4053), .B(n4060), .Z(n6517) );
  ANDN U1410 ( .B(y[554]), .A(x[554]), .Z(n4051) );
  ANDN U1411 ( .B(y[555]), .A(x[555]), .Z(n4059) );
  NOR U1412 ( .A(n4051), .B(n4059), .Z(n6515) );
  NANDN U1413 ( .A(y[553]), .B(x[553]), .Z(n1868) );
  NANDN U1414 ( .A(y[554]), .B(x[554]), .Z(n4054) );
  NAND U1415 ( .A(n1868), .B(n4054), .Z(n6513) );
  ANDN U1416 ( .B(y[552]), .A(x[552]), .Z(n4043) );
  ANDN U1417 ( .B(y[553]), .A(x[553]), .Z(n4048) );
  NOR U1418 ( .A(n4043), .B(n4048), .Z(n6511) );
  NANDN U1419 ( .A(y[551]), .B(x[551]), .Z(n4039) );
  NANDN U1420 ( .A(y[552]), .B(x[552]), .Z(n1867) );
  NAND U1421 ( .A(n4039), .B(n1867), .Z(n6509) );
  NANDN U1422 ( .A(x[550]), .B(y[550]), .Z(n309) );
  ANDN U1423 ( .B(y[551]), .A(x[551]), .Z(n4044) );
  ANDN U1424 ( .B(n309), .A(n4044), .Z(n6507) );
  XOR U1425 ( .A(x[550]), .B(y[550]), .Z(n4037) );
  NANDN U1426 ( .A(y[549]), .B(x[549]), .Z(n4031) );
  NANDN U1427 ( .A(n4037), .B(n4031), .Z(n6505) );
  ANDN U1428 ( .B(y[548]), .A(x[548]), .Z(n4029) );
  ANDN U1429 ( .B(y[549]), .A(x[549]), .Z(n4034) );
  NOR U1430 ( .A(n4029), .B(n4034), .Z(n6503) );
  NANDN U1431 ( .A(y[547]), .B(x[547]), .Z(n1870) );
  NANDN U1432 ( .A(y[548]), .B(x[548]), .Z(n4032) );
  NAND U1433 ( .A(n1870), .B(n4032), .Z(n6501) );
  ANDN U1434 ( .B(y[546]), .A(x[546]), .Z(n4021) );
  ANDN U1435 ( .B(y[547]), .A(x[547]), .Z(n4026) );
  NOR U1436 ( .A(n4021), .B(n4026), .Z(n6499) );
  NANDN U1437 ( .A(y[545]), .B(x[545]), .Z(n4017) );
  NANDN U1438 ( .A(y[546]), .B(x[546]), .Z(n1869) );
  NAND U1439 ( .A(n4017), .B(n1869), .Z(n6497) );
  ANDN U1440 ( .B(y[544]), .A(x[544]), .Z(n4012) );
  ANDN U1441 ( .B(y[545]), .A(x[545]), .Z(n4022) );
  NOR U1442 ( .A(n4012), .B(n4022), .Z(n6495) );
  NANDN U1443 ( .A(y[543]), .B(x[543]), .Z(n4009) );
  NANDN U1444 ( .A(y[544]), .B(x[544]), .Z(n4016) );
  NAND U1445 ( .A(n4009), .B(n4016), .Z(n6493) );
  ANDN U1446 ( .B(y[542]), .A(x[542]), .Z(n4007) );
  ANDN U1447 ( .B(y[543]), .A(x[543]), .Z(n4015) );
  NOR U1448 ( .A(n4007), .B(n4015), .Z(n6491) );
  NANDN U1449 ( .A(y[541]), .B(x[541]), .Z(n1872) );
  NANDN U1450 ( .A(y[542]), .B(x[542]), .Z(n4010) );
  NAND U1451 ( .A(n1872), .B(n4010), .Z(n6489) );
  ANDN U1452 ( .B(y[540]), .A(x[540]), .Z(n3999) );
  ANDN U1453 ( .B(y[541]), .A(x[541]), .Z(n4004) );
  NOR U1454 ( .A(n3999), .B(n4004), .Z(n6487) );
  NANDN U1455 ( .A(y[539]), .B(x[539]), .Z(n3995) );
  NANDN U1456 ( .A(y[540]), .B(x[540]), .Z(n1871) );
  NAND U1457 ( .A(n3995), .B(n1871), .Z(n6485) );
  NANDN U1458 ( .A(x[538]), .B(y[538]), .Z(n310) );
  ANDN U1459 ( .B(y[539]), .A(x[539]), .Z(n4000) );
  ANDN U1460 ( .B(n310), .A(n4000), .Z(n6483) );
  XOR U1461 ( .A(x[538]), .B(y[538]), .Z(n3993) );
  NANDN U1462 ( .A(y[537]), .B(x[537]), .Z(n3987) );
  NANDN U1463 ( .A(n3993), .B(n3987), .Z(n6481) );
  ANDN U1464 ( .B(y[536]), .A(x[536]), .Z(n3985) );
  ANDN U1465 ( .B(y[537]), .A(x[537]), .Z(n3990) );
  NOR U1466 ( .A(n3985), .B(n3990), .Z(n6479) );
  NANDN U1467 ( .A(y[535]), .B(x[535]), .Z(n1874) );
  NANDN U1468 ( .A(y[536]), .B(x[536]), .Z(n3988) );
  NAND U1469 ( .A(n1874), .B(n3988), .Z(n6477) );
  ANDN U1470 ( .B(y[534]), .A(x[534]), .Z(n3977) );
  ANDN U1471 ( .B(y[535]), .A(x[535]), .Z(n3982) );
  NOR U1472 ( .A(n3977), .B(n3982), .Z(n6475) );
  NANDN U1473 ( .A(y[533]), .B(x[533]), .Z(n3973) );
  NANDN U1474 ( .A(y[534]), .B(x[534]), .Z(n1873) );
  NAND U1475 ( .A(n3973), .B(n1873), .Z(n6473) );
  NANDN U1476 ( .A(x[532]), .B(y[532]), .Z(n311) );
  ANDN U1477 ( .B(y[533]), .A(x[533]), .Z(n3978) );
  ANDN U1478 ( .B(n311), .A(n3978), .Z(n6471) );
  XOR U1479 ( .A(x[532]), .B(y[532]), .Z(n3971) );
  NANDN U1480 ( .A(y[531]), .B(x[531]), .Z(n3965) );
  NANDN U1481 ( .A(n3971), .B(n3965), .Z(n6469) );
  NANDN U1482 ( .A(x[530]), .B(y[530]), .Z(n312) );
  ANDN U1483 ( .B(y[531]), .A(x[531]), .Z(n3968) );
  ANDN U1484 ( .B(n312), .A(n3968), .Z(n6467) );
  XOR U1485 ( .A(x[530]), .B(y[530]), .Z(n3961) );
  NANDN U1486 ( .A(y[529]), .B(x[529]), .Z(n1875) );
  NANDN U1487 ( .A(n3961), .B(n1875), .Z(n6465) );
  NANDN U1488 ( .A(x[528]), .B(y[528]), .Z(n313) );
  ANDN U1489 ( .B(y[529]), .A(x[529]), .Z(n3963) );
  ANDN U1490 ( .B(n313), .A(n3963), .Z(n6463) );
  XOR U1491 ( .A(x[528]), .B(y[528]), .Z(n3955) );
  NANDN U1492 ( .A(y[527]), .B(x[527]), .Z(n3951) );
  NANDN U1493 ( .A(n3955), .B(n3951), .Z(n6461) );
  NANDN U1494 ( .A(x[526]), .B(y[526]), .Z(n314) );
  ANDN U1495 ( .B(y[527]), .A(x[527]), .Z(n3956) );
  ANDN U1496 ( .B(n314), .A(n3956), .Z(n6459) );
  XOR U1497 ( .A(x[526]), .B(y[526]), .Z(n3949) );
  NANDN U1498 ( .A(y[525]), .B(x[525]), .Z(n3943) );
  NANDN U1499 ( .A(n3949), .B(n3943), .Z(n6457) );
  ANDN U1500 ( .B(y[524]), .A(x[524]), .Z(n3941) );
  ANDN U1501 ( .B(y[525]), .A(x[525]), .Z(n3946) );
  NOR U1502 ( .A(n3941), .B(n3946), .Z(n6455) );
  NANDN U1503 ( .A(y[523]), .B(x[523]), .Z(n1878) );
  NANDN U1504 ( .A(y[524]), .B(x[524]), .Z(n3944) );
  NAND U1505 ( .A(n1878), .B(n3944), .Z(n6453) );
  ANDN U1506 ( .B(y[522]), .A(x[522]), .Z(n3933) );
  ANDN U1507 ( .B(y[523]), .A(x[523]), .Z(n3938) );
  NOR U1508 ( .A(n3933), .B(n3938), .Z(n6451) );
  NANDN U1509 ( .A(y[521]), .B(x[521]), .Z(n3929) );
  NANDN U1510 ( .A(y[522]), .B(x[522]), .Z(n1877) );
  NAND U1511 ( .A(n3929), .B(n1877), .Z(n6449) );
  ANDN U1512 ( .B(y[520]), .A(x[520]), .Z(n3924) );
  ANDN U1513 ( .B(y[521]), .A(x[521]), .Z(n3934) );
  NOR U1514 ( .A(n3924), .B(n3934), .Z(n6447) );
  NANDN U1515 ( .A(y[519]), .B(x[519]), .Z(n3921) );
  NANDN U1516 ( .A(y[520]), .B(x[520]), .Z(n3928) );
  NAND U1517 ( .A(n3921), .B(n3928), .Z(n6445) );
  ANDN U1518 ( .B(y[518]), .A(x[518]), .Z(n3919) );
  ANDN U1519 ( .B(y[519]), .A(x[519]), .Z(n3927) );
  NOR U1520 ( .A(n3919), .B(n3927), .Z(n6443) );
  NANDN U1521 ( .A(y[517]), .B(x[517]), .Z(n1880) );
  NANDN U1522 ( .A(y[518]), .B(x[518]), .Z(n3922) );
  NAND U1523 ( .A(n1880), .B(n3922), .Z(n6441) );
  ANDN U1524 ( .B(y[516]), .A(x[516]), .Z(n3911) );
  ANDN U1525 ( .B(y[517]), .A(x[517]), .Z(n3916) );
  NOR U1526 ( .A(n3911), .B(n3916), .Z(n6439) );
  NANDN U1527 ( .A(y[515]), .B(x[515]), .Z(n3907) );
  NANDN U1528 ( .A(y[516]), .B(x[516]), .Z(n1879) );
  NAND U1529 ( .A(n3907), .B(n1879), .Z(n6437) );
  NANDN U1530 ( .A(x[514]), .B(y[514]), .Z(n315) );
  ANDN U1531 ( .B(y[515]), .A(x[515]), .Z(n3912) );
  ANDN U1532 ( .B(n315), .A(n3912), .Z(n6435) );
  XOR U1533 ( .A(x[514]), .B(y[514]), .Z(n3905) );
  NANDN U1534 ( .A(y[513]), .B(x[513]), .Z(n3899) );
  NANDN U1535 ( .A(n3905), .B(n3899), .Z(n6433) );
  ANDN U1536 ( .B(y[512]), .A(x[512]), .Z(n3897) );
  ANDN U1537 ( .B(y[513]), .A(x[513]), .Z(n3902) );
  NOR U1538 ( .A(n3897), .B(n3902), .Z(n6431) );
  NANDN U1539 ( .A(y[511]), .B(x[511]), .Z(n1882) );
  NANDN U1540 ( .A(y[512]), .B(x[512]), .Z(n3900) );
  NAND U1541 ( .A(n1882), .B(n3900), .Z(n6429) );
  ANDN U1542 ( .B(y[510]), .A(x[510]), .Z(n3889) );
  ANDN U1543 ( .B(y[511]), .A(x[511]), .Z(n3894) );
  NOR U1544 ( .A(n3889), .B(n3894), .Z(n6427) );
  NANDN U1545 ( .A(y[509]), .B(x[509]), .Z(n3885) );
  NANDN U1546 ( .A(y[510]), .B(x[510]), .Z(n1881) );
  NAND U1547 ( .A(n3885), .B(n1881), .Z(n6425) );
  NANDN U1548 ( .A(x[508]), .B(y[508]), .Z(n316) );
  ANDN U1549 ( .B(y[509]), .A(x[509]), .Z(n3890) );
  ANDN U1550 ( .B(n316), .A(n3890), .Z(n6423) );
  XOR U1551 ( .A(x[508]), .B(y[508]), .Z(n3883) );
  NANDN U1552 ( .A(y[507]), .B(x[507]), .Z(n3877) );
  NANDN U1553 ( .A(n3883), .B(n3877), .Z(n6421) );
  ANDN U1554 ( .B(y[506]), .A(x[506]), .Z(n3875) );
  ANDN U1555 ( .B(y[507]), .A(x[507]), .Z(n3880) );
  NOR U1556 ( .A(n3875), .B(n3880), .Z(n6419) );
  NANDN U1557 ( .A(y[505]), .B(x[505]), .Z(n1884) );
  NANDN U1558 ( .A(y[506]), .B(x[506]), .Z(n3878) );
  NAND U1559 ( .A(n1884), .B(n3878), .Z(n6417) );
  ANDN U1560 ( .B(y[504]), .A(x[504]), .Z(n3867) );
  ANDN U1561 ( .B(y[505]), .A(x[505]), .Z(n3872) );
  NOR U1562 ( .A(n3867), .B(n3872), .Z(n6415) );
  NANDN U1563 ( .A(y[503]), .B(x[503]), .Z(n3863) );
  NANDN U1564 ( .A(y[504]), .B(x[504]), .Z(n1883) );
  NAND U1565 ( .A(n3863), .B(n1883), .Z(n6413) );
  ANDN U1566 ( .B(y[502]), .A(x[502]), .Z(n3858) );
  ANDN U1567 ( .B(y[503]), .A(x[503]), .Z(n3868) );
  NOR U1568 ( .A(n3858), .B(n3868), .Z(n6411) );
  NANDN U1569 ( .A(y[501]), .B(x[501]), .Z(n3855) );
  NANDN U1570 ( .A(y[502]), .B(x[502]), .Z(n3862) );
  NAND U1571 ( .A(n3855), .B(n3862), .Z(n6409) );
  ANDN U1572 ( .B(y[500]), .A(x[500]), .Z(n3853) );
  ANDN U1573 ( .B(y[501]), .A(x[501]), .Z(n3861) );
  NOR U1574 ( .A(n3853), .B(n3861), .Z(n6407) );
  NANDN U1575 ( .A(y[499]), .B(x[499]), .Z(n1886) );
  NANDN U1576 ( .A(y[500]), .B(x[500]), .Z(n3856) );
  NAND U1577 ( .A(n1886), .B(n3856), .Z(n6405) );
  ANDN U1578 ( .B(y[498]), .A(x[498]), .Z(n3845) );
  ANDN U1579 ( .B(y[499]), .A(x[499]), .Z(n3850) );
  NOR U1580 ( .A(n3845), .B(n3850), .Z(n6403) );
  NANDN U1581 ( .A(y[497]), .B(x[497]), .Z(n3841) );
  NANDN U1582 ( .A(y[498]), .B(x[498]), .Z(n1885) );
  NAND U1583 ( .A(n3841), .B(n1885), .Z(n6401) );
  NANDN U1584 ( .A(x[496]), .B(y[496]), .Z(n317) );
  ANDN U1585 ( .B(y[497]), .A(x[497]), .Z(n3846) );
  ANDN U1586 ( .B(n317), .A(n3846), .Z(n6399) );
  XOR U1587 ( .A(x[496]), .B(y[496]), .Z(n3839) );
  NANDN U1588 ( .A(y[495]), .B(x[495]), .Z(n3833) );
  NANDN U1589 ( .A(n3839), .B(n3833), .Z(n6397) );
  ANDN U1590 ( .B(y[494]), .A(x[494]), .Z(n3831) );
  ANDN U1591 ( .B(y[495]), .A(x[495]), .Z(n3836) );
  NOR U1592 ( .A(n3831), .B(n3836), .Z(n6395) );
  NANDN U1593 ( .A(y[493]), .B(x[493]), .Z(n1888) );
  NANDN U1594 ( .A(y[494]), .B(x[494]), .Z(n3834) );
  NAND U1595 ( .A(n1888), .B(n3834), .Z(n6393) );
  ANDN U1596 ( .B(y[492]), .A(x[492]), .Z(n3823) );
  ANDN U1597 ( .B(y[493]), .A(x[493]), .Z(n3828) );
  NOR U1598 ( .A(n3823), .B(n3828), .Z(n6391) );
  NANDN U1599 ( .A(y[491]), .B(x[491]), .Z(n3819) );
  NANDN U1600 ( .A(y[492]), .B(x[492]), .Z(n1887) );
  NAND U1601 ( .A(n3819), .B(n1887), .Z(n6389) );
  NANDN U1602 ( .A(x[490]), .B(y[490]), .Z(n318) );
  ANDN U1603 ( .B(y[491]), .A(x[491]), .Z(n3824) );
  ANDN U1604 ( .B(n318), .A(n3824), .Z(n6387) );
  XOR U1605 ( .A(x[490]), .B(y[490]), .Z(n3817) );
  NANDN U1606 ( .A(y[489]), .B(x[489]), .Z(n3811) );
  NANDN U1607 ( .A(n3817), .B(n3811), .Z(n6385) );
  NANDN U1608 ( .A(x[488]), .B(y[488]), .Z(n319) );
  ANDN U1609 ( .B(y[489]), .A(x[489]), .Z(n3814) );
  ANDN U1610 ( .B(n319), .A(n3814), .Z(n6383) );
  XOR U1611 ( .A(x[488]), .B(y[488]), .Z(n3807) );
  NANDN U1612 ( .A(y[487]), .B(x[487]), .Z(n1889) );
  NANDN U1613 ( .A(n3807), .B(n1889), .Z(n6381) );
  NANDN U1614 ( .A(x[486]), .B(y[486]), .Z(n320) );
  ANDN U1615 ( .B(y[487]), .A(x[487]), .Z(n3809) );
  ANDN U1616 ( .B(n320), .A(n3809), .Z(n6379) );
  XOR U1617 ( .A(x[486]), .B(y[486]), .Z(n3801) );
  NANDN U1618 ( .A(y[485]), .B(x[485]), .Z(n3797) );
  NANDN U1619 ( .A(n3801), .B(n3797), .Z(n6377) );
  NANDN U1620 ( .A(x[484]), .B(y[484]), .Z(n321) );
  ANDN U1621 ( .B(y[485]), .A(x[485]), .Z(n3802) );
  ANDN U1622 ( .B(n321), .A(n3802), .Z(n6375) );
  XOR U1623 ( .A(x[484]), .B(y[484]), .Z(n3795) );
  NANDN U1624 ( .A(y[483]), .B(x[483]), .Z(n3789) );
  NANDN U1625 ( .A(n3795), .B(n3789), .Z(n6373) );
  ANDN U1626 ( .B(y[482]), .A(x[482]), .Z(n3787) );
  ANDN U1627 ( .B(y[483]), .A(x[483]), .Z(n3792) );
  NOR U1628 ( .A(n3787), .B(n3792), .Z(n6371) );
  NANDN U1629 ( .A(y[481]), .B(x[481]), .Z(n1891) );
  NANDN U1630 ( .A(y[482]), .B(x[482]), .Z(n3790) );
  NAND U1631 ( .A(n1891), .B(n3790), .Z(n6369) );
  NANDN U1632 ( .A(x[480]), .B(y[480]), .Z(n322) );
  ANDN U1633 ( .B(y[481]), .A(x[481]), .Z(n3784) );
  ANDN U1634 ( .B(n322), .A(n3784), .Z(n6367) );
  XOR U1635 ( .A(x[480]), .B(y[480]), .Z(n3779) );
  NANDN U1636 ( .A(y[479]), .B(x[479]), .Z(n3775) );
  NANDN U1637 ( .A(n3779), .B(n3775), .Z(n6365) );
  ANDN U1638 ( .B(y[478]), .A(x[478]), .Z(n3770) );
  ANDN U1639 ( .B(y[479]), .A(x[479]), .Z(n3780) );
  NOR U1640 ( .A(n3770), .B(n3780), .Z(n6363) );
  NANDN U1641 ( .A(y[477]), .B(x[477]), .Z(n3767) );
  NANDN U1642 ( .A(y[478]), .B(x[478]), .Z(n3777) );
  NAND U1643 ( .A(n3767), .B(n3777), .Z(n6361) );
  ANDN U1644 ( .B(y[476]), .A(x[476]), .Z(n3765) );
  ANDN U1645 ( .B(y[477]), .A(x[477]), .Z(n3773) );
  NOR U1646 ( .A(n3765), .B(n3773), .Z(n6359) );
  NANDN U1647 ( .A(y[475]), .B(x[475]), .Z(n1893) );
  NANDN U1648 ( .A(y[476]), .B(x[476]), .Z(n3768) );
  NAND U1649 ( .A(n1893), .B(n3768), .Z(n6357) );
  NANDN U1650 ( .A(x[474]), .B(y[474]), .Z(n323) );
  ANDN U1651 ( .B(y[475]), .A(x[475]), .Z(n3762) );
  ANDN U1652 ( .B(n323), .A(n3762), .Z(n6355) );
  XOR U1653 ( .A(x[474]), .B(y[474]), .Z(n3757) );
  NANDN U1654 ( .A(y[473]), .B(x[473]), .Z(n3753) );
  NANDN U1655 ( .A(n3757), .B(n3753), .Z(n6353) );
  NANDN U1656 ( .A(x[472]), .B(y[472]), .Z(n324) );
  ANDN U1657 ( .B(y[473]), .A(x[473]), .Z(n3758) );
  ANDN U1658 ( .B(n324), .A(n3758), .Z(n6351) );
  XOR U1659 ( .A(x[472]), .B(y[472]), .Z(n3751) );
  NANDN U1660 ( .A(y[471]), .B(x[471]), .Z(n3745) );
  NANDN U1661 ( .A(n3751), .B(n3745), .Z(n6349) );
  ANDN U1662 ( .B(y[470]), .A(x[470]), .Z(n3743) );
  ANDN U1663 ( .B(y[471]), .A(x[471]), .Z(n3748) );
  NOR U1664 ( .A(n3743), .B(n3748), .Z(n6347) );
  NANDN U1665 ( .A(y[469]), .B(x[469]), .Z(n1895) );
  NANDN U1666 ( .A(y[470]), .B(x[470]), .Z(n3746) );
  NAND U1667 ( .A(n1895), .B(n3746), .Z(n6345) );
  NANDN U1668 ( .A(x[468]), .B(y[468]), .Z(n325) );
  ANDN U1669 ( .B(y[469]), .A(x[469]), .Z(n3740) );
  ANDN U1670 ( .B(n325), .A(n3740), .Z(n6343) );
  XOR U1671 ( .A(x[468]), .B(y[468]), .Z(n3735) );
  NANDN U1672 ( .A(y[467]), .B(x[467]), .Z(n3731) );
  NANDN U1673 ( .A(n3735), .B(n3731), .Z(n6341) );
  NANDN U1674 ( .A(x[466]), .B(y[466]), .Z(n326) );
  ANDN U1675 ( .B(y[467]), .A(x[467]), .Z(n3736) );
  ANDN U1676 ( .B(n326), .A(n3736), .Z(n6339) );
  XOR U1677 ( .A(x[466]), .B(y[466]), .Z(n3729) );
  NANDN U1678 ( .A(y[465]), .B(x[465]), .Z(n3723) );
  NANDN U1679 ( .A(n3729), .B(n3723), .Z(n6337) );
  NANDN U1680 ( .A(x[464]), .B(y[464]), .Z(n327) );
  ANDN U1681 ( .B(y[465]), .A(x[465]), .Z(n3726) );
  ANDN U1682 ( .B(n327), .A(n3726), .Z(n6335) );
  XOR U1683 ( .A(x[464]), .B(y[464]), .Z(n3719) );
  NANDN U1684 ( .A(y[463]), .B(x[463]), .Z(n1897) );
  NANDN U1685 ( .A(n3719), .B(n1897), .Z(n6333) );
  NANDN U1686 ( .A(x[462]), .B(y[462]), .Z(n328) );
  ANDN U1687 ( .B(y[463]), .A(x[463]), .Z(n3721) );
  ANDN U1688 ( .B(n328), .A(n3721), .Z(n6331) );
  XOR U1689 ( .A(x[462]), .B(y[462]), .Z(n3713) );
  NANDN U1690 ( .A(y[461]), .B(x[461]), .Z(n3709) );
  NANDN U1691 ( .A(n3713), .B(n3709), .Z(n6329) );
  ANDN U1692 ( .B(y[460]), .A(x[460]), .Z(n3704) );
  ANDN U1693 ( .B(y[461]), .A(x[461]), .Z(n3714) );
  NOR U1694 ( .A(n3704), .B(n3714), .Z(n6327) );
  NANDN U1695 ( .A(y[459]), .B(x[459]), .Z(n3701) );
  NANDN U1696 ( .A(y[460]), .B(x[460]), .Z(n3711) );
  NAND U1697 ( .A(n3701), .B(n3711), .Z(n6325) );
  ANDN U1698 ( .B(y[458]), .A(x[458]), .Z(n3699) );
  ANDN U1699 ( .B(y[459]), .A(x[459]), .Z(n3707) );
  NOR U1700 ( .A(n3699), .B(n3707), .Z(n6323) );
  NANDN U1701 ( .A(y[457]), .B(x[457]), .Z(n1900) );
  NANDN U1702 ( .A(y[458]), .B(x[458]), .Z(n3702) );
  NAND U1703 ( .A(n1900), .B(n3702), .Z(n6321) );
  ANDN U1704 ( .B(y[456]), .A(x[456]), .Z(n3691) );
  ANDN U1705 ( .B(y[457]), .A(x[457]), .Z(n3696) );
  NOR U1706 ( .A(n3691), .B(n3696), .Z(n6319) );
  NANDN U1707 ( .A(y[455]), .B(x[455]), .Z(n3687) );
  NANDN U1708 ( .A(y[456]), .B(x[456]), .Z(n1899) );
  NAND U1709 ( .A(n3687), .B(n1899), .Z(n6317) );
  ANDN U1710 ( .B(y[454]), .A(x[454]), .Z(n3682) );
  ANDN U1711 ( .B(y[455]), .A(x[455]), .Z(n3692) );
  NOR U1712 ( .A(n3682), .B(n3692), .Z(n6315) );
  NANDN U1713 ( .A(y[453]), .B(x[453]), .Z(n3679) );
  NANDN U1714 ( .A(y[454]), .B(x[454]), .Z(n3686) );
  NAND U1715 ( .A(n3679), .B(n3686), .Z(n6313) );
  ANDN U1716 ( .B(y[452]), .A(x[452]), .Z(n3677) );
  ANDN U1717 ( .B(y[453]), .A(x[453]), .Z(n3685) );
  NOR U1718 ( .A(n3677), .B(n3685), .Z(n6311) );
  NANDN U1719 ( .A(y[451]), .B(x[451]), .Z(n1902) );
  NANDN U1720 ( .A(y[452]), .B(x[452]), .Z(n3680) );
  NAND U1721 ( .A(n1902), .B(n3680), .Z(n6309) );
  ANDN U1722 ( .B(y[450]), .A(x[450]), .Z(n3669) );
  ANDN U1723 ( .B(y[451]), .A(x[451]), .Z(n3674) );
  NOR U1724 ( .A(n3669), .B(n3674), .Z(n6307) );
  NANDN U1725 ( .A(y[449]), .B(x[449]), .Z(n3665) );
  NANDN U1726 ( .A(y[450]), .B(x[450]), .Z(n1901) );
  NAND U1727 ( .A(n3665), .B(n1901), .Z(n6305) );
  ANDN U1728 ( .B(y[448]), .A(x[448]), .Z(n3660) );
  ANDN U1729 ( .B(y[449]), .A(x[449]), .Z(n3670) );
  NOR U1730 ( .A(n3660), .B(n3670), .Z(n6303) );
  NANDN U1731 ( .A(y[447]), .B(x[447]), .Z(n3657) );
  NANDN U1732 ( .A(y[448]), .B(x[448]), .Z(n3664) );
  NAND U1733 ( .A(n3657), .B(n3664), .Z(n6301) );
  ANDN U1734 ( .B(y[446]), .A(x[446]), .Z(n3655) );
  ANDN U1735 ( .B(y[447]), .A(x[447]), .Z(n3663) );
  NOR U1736 ( .A(n3655), .B(n3663), .Z(n6299) );
  NANDN U1737 ( .A(y[445]), .B(x[445]), .Z(n1904) );
  NANDN U1738 ( .A(y[446]), .B(x[446]), .Z(n3658) );
  NAND U1739 ( .A(n1904), .B(n3658), .Z(n6297) );
  ANDN U1740 ( .B(y[444]), .A(x[444]), .Z(n3647) );
  ANDN U1741 ( .B(y[445]), .A(x[445]), .Z(n3652) );
  NOR U1742 ( .A(n3647), .B(n3652), .Z(n6295) );
  NANDN U1743 ( .A(y[443]), .B(x[443]), .Z(n3643) );
  NANDN U1744 ( .A(y[444]), .B(x[444]), .Z(n1903) );
  NAND U1745 ( .A(n3643), .B(n1903), .Z(n6293) );
  NANDN U1746 ( .A(x[442]), .B(y[442]), .Z(n329) );
  ANDN U1747 ( .B(y[443]), .A(x[443]), .Z(n3648) );
  ANDN U1748 ( .B(n329), .A(n3648), .Z(n6291) );
  XOR U1749 ( .A(x[442]), .B(y[442]), .Z(n3641) );
  NANDN U1750 ( .A(y[441]), .B(x[441]), .Z(n3635) );
  NANDN U1751 ( .A(n3641), .B(n3635), .Z(n6289) );
  ANDN U1752 ( .B(y[440]), .A(x[440]), .Z(n3633) );
  ANDN U1753 ( .B(y[441]), .A(x[441]), .Z(n3638) );
  NOR U1754 ( .A(n3633), .B(n3638), .Z(n6287) );
  NANDN U1755 ( .A(y[439]), .B(x[439]), .Z(n1906) );
  NANDN U1756 ( .A(y[440]), .B(x[440]), .Z(n3636) );
  NAND U1757 ( .A(n1906), .B(n3636), .Z(n6285) );
  ANDN U1758 ( .B(y[438]), .A(x[438]), .Z(n3625) );
  ANDN U1759 ( .B(y[439]), .A(x[439]), .Z(n3630) );
  NOR U1760 ( .A(n3625), .B(n3630), .Z(n6283) );
  NANDN U1761 ( .A(y[437]), .B(x[437]), .Z(n3621) );
  NANDN U1762 ( .A(y[438]), .B(x[438]), .Z(n1905) );
  NAND U1763 ( .A(n3621), .B(n1905), .Z(n6281) );
  NANDN U1764 ( .A(x[436]), .B(y[436]), .Z(n330) );
  ANDN U1765 ( .B(y[437]), .A(x[437]), .Z(n3626) );
  ANDN U1766 ( .B(n330), .A(n3626), .Z(n6279) );
  XOR U1767 ( .A(x[436]), .B(y[436]), .Z(n3619) );
  NANDN U1768 ( .A(y[435]), .B(x[435]), .Z(n3613) );
  NANDN U1769 ( .A(n3619), .B(n3613), .Z(n6277) );
  NANDN U1770 ( .A(x[434]), .B(y[434]), .Z(n331) );
  ANDN U1771 ( .B(y[435]), .A(x[435]), .Z(n3616) );
  ANDN U1772 ( .B(n331), .A(n3616), .Z(n6275) );
  XOR U1773 ( .A(x[434]), .B(y[434]), .Z(n3609) );
  NANDN U1774 ( .A(y[433]), .B(x[433]), .Z(n1908) );
  NANDN U1775 ( .A(n3609), .B(n1908), .Z(n6273) );
  ANDN U1776 ( .B(y[432]), .A(x[432]), .Z(n3603) );
  ANDN U1777 ( .B(y[433]), .A(x[433]), .Z(n3611) );
  NOR U1778 ( .A(n3603), .B(n3611), .Z(n6271) );
  NANDN U1779 ( .A(y[431]), .B(x[431]), .Z(n3599) );
  NANDN U1780 ( .A(y[432]), .B(x[432]), .Z(n1907) );
  NAND U1781 ( .A(n3599), .B(n1907), .Z(n6269) );
  ANDN U1782 ( .B(y[430]), .A(x[430]), .Z(n3594) );
  ANDN U1783 ( .B(y[431]), .A(x[431]), .Z(n3604) );
  NOR U1784 ( .A(n3594), .B(n3604), .Z(n6267) );
  NANDN U1785 ( .A(y[429]), .B(x[429]), .Z(n3591) );
  NANDN U1786 ( .A(y[430]), .B(x[430]), .Z(n3598) );
  NAND U1787 ( .A(n3591), .B(n3598), .Z(n6265) );
  ANDN U1788 ( .B(y[428]), .A(x[428]), .Z(n3589) );
  ANDN U1789 ( .B(y[429]), .A(x[429]), .Z(n3597) );
  NOR U1790 ( .A(n3589), .B(n3597), .Z(n6263) );
  NANDN U1791 ( .A(y[427]), .B(x[427]), .Z(n1910) );
  NANDN U1792 ( .A(y[428]), .B(x[428]), .Z(n3592) );
  NAND U1793 ( .A(n1910), .B(n3592), .Z(n6261) );
  ANDN U1794 ( .B(y[426]), .A(x[426]), .Z(n3581) );
  ANDN U1795 ( .B(y[427]), .A(x[427]), .Z(n3586) );
  NOR U1796 ( .A(n3581), .B(n3586), .Z(n6259) );
  NANDN U1797 ( .A(y[425]), .B(x[425]), .Z(n3577) );
  NANDN U1798 ( .A(y[426]), .B(x[426]), .Z(n1909) );
  NAND U1799 ( .A(n3577), .B(n1909), .Z(n6257) );
  ANDN U1800 ( .B(y[424]), .A(x[424]), .Z(n3572) );
  ANDN U1801 ( .B(y[425]), .A(x[425]), .Z(n3582) );
  NOR U1802 ( .A(n3572), .B(n3582), .Z(n6255) );
  NANDN U1803 ( .A(y[423]), .B(x[423]), .Z(n3569) );
  NANDN U1804 ( .A(y[424]), .B(x[424]), .Z(n3576) );
  NAND U1805 ( .A(n3569), .B(n3576), .Z(n6253) );
  ANDN U1806 ( .B(y[422]), .A(x[422]), .Z(n3567) );
  ANDN U1807 ( .B(y[423]), .A(x[423]), .Z(n3575) );
  NOR U1808 ( .A(n3567), .B(n3575), .Z(n6251) );
  NANDN U1809 ( .A(y[421]), .B(x[421]), .Z(n1912) );
  NANDN U1810 ( .A(y[422]), .B(x[422]), .Z(n3570) );
  NAND U1811 ( .A(n1912), .B(n3570), .Z(n6249) );
  ANDN U1812 ( .B(y[420]), .A(x[420]), .Z(n3559) );
  ANDN U1813 ( .B(y[421]), .A(x[421]), .Z(n3564) );
  NOR U1814 ( .A(n3559), .B(n3564), .Z(n6247) );
  NANDN U1815 ( .A(y[419]), .B(x[419]), .Z(n3555) );
  NANDN U1816 ( .A(y[420]), .B(x[420]), .Z(n1911) );
  NAND U1817 ( .A(n3555), .B(n1911), .Z(n6245) );
  NANDN U1818 ( .A(x[418]), .B(y[418]), .Z(n332) );
  ANDN U1819 ( .B(y[419]), .A(x[419]), .Z(n3560) );
  ANDN U1820 ( .B(n332), .A(n3560), .Z(n6243) );
  XOR U1821 ( .A(x[418]), .B(y[418]), .Z(n3553) );
  NANDN U1822 ( .A(y[417]), .B(x[417]), .Z(n3547) );
  NANDN U1823 ( .A(n3553), .B(n3547), .Z(n6241) );
  ANDN U1824 ( .B(y[416]), .A(x[416]), .Z(n3545) );
  ANDN U1825 ( .B(y[417]), .A(x[417]), .Z(n3550) );
  NOR U1826 ( .A(n3545), .B(n3550), .Z(n6239) );
  NANDN U1827 ( .A(y[415]), .B(x[415]), .Z(n1914) );
  NANDN U1828 ( .A(y[416]), .B(x[416]), .Z(n3548) );
  NAND U1829 ( .A(n1914), .B(n3548), .Z(n6237) );
  ANDN U1830 ( .B(y[414]), .A(x[414]), .Z(n3537) );
  ANDN U1831 ( .B(y[415]), .A(x[415]), .Z(n3542) );
  NOR U1832 ( .A(n3537), .B(n3542), .Z(n6235) );
  NANDN U1833 ( .A(y[413]), .B(x[413]), .Z(n3533) );
  NANDN U1834 ( .A(y[414]), .B(x[414]), .Z(n1913) );
  NAND U1835 ( .A(n3533), .B(n1913), .Z(n6233) );
  ANDN U1836 ( .B(y[412]), .A(x[412]), .Z(n3528) );
  ANDN U1837 ( .B(y[413]), .A(x[413]), .Z(n3538) );
  NOR U1838 ( .A(n3528), .B(n3538), .Z(n6231) );
  NANDN U1839 ( .A(y[411]), .B(x[411]), .Z(n3525) );
  NANDN U1840 ( .A(y[412]), .B(x[412]), .Z(n3532) );
  NAND U1841 ( .A(n3525), .B(n3532), .Z(n6229) );
  ANDN U1842 ( .B(y[410]), .A(x[410]), .Z(n3523) );
  ANDN U1843 ( .B(y[411]), .A(x[411]), .Z(n3531) );
  NOR U1844 ( .A(n3523), .B(n3531), .Z(n6227) );
  NANDN U1845 ( .A(y[409]), .B(x[409]), .Z(n1916) );
  NANDN U1846 ( .A(y[410]), .B(x[410]), .Z(n3526) );
  NAND U1847 ( .A(n1916), .B(n3526), .Z(n6225) );
  ANDN U1848 ( .B(y[408]), .A(x[408]), .Z(n3515) );
  ANDN U1849 ( .B(y[409]), .A(x[409]), .Z(n3520) );
  NOR U1850 ( .A(n3515), .B(n3520), .Z(n6223) );
  NANDN U1851 ( .A(y[407]), .B(x[407]), .Z(n3511) );
  NANDN U1852 ( .A(y[408]), .B(x[408]), .Z(n1915) );
  NAND U1853 ( .A(n3511), .B(n1915), .Z(n6221) );
  NANDN U1854 ( .A(x[406]), .B(y[406]), .Z(n333) );
  ANDN U1855 ( .B(y[407]), .A(x[407]), .Z(n3516) );
  ANDN U1856 ( .B(n333), .A(n3516), .Z(n6219) );
  XOR U1857 ( .A(x[406]), .B(y[406]), .Z(n3509) );
  NANDN U1858 ( .A(y[405]), .B(x[405]), .Z(n3503) );
  NANDN U1859 ( .A(n3509), .B(n3503), .Z(n6217) );
  ANDN U1860 ( .B(y[404]), .A(x[404]), .Z(n3501) );
  ANDN U1861 ( .B(y[405]), .A(x[405]), .Z(n3506) );
  NOR U1862 ( .A(n3501), .B(n3506), .Z(n6215) );
  NANDN U1863 ( .A(y[403]), .B(x[403]), .Z(n1917) );
  NANDN U1864 ( .A(y[404]), .B(x[404]), .Z(n3504) );
  NAND U1865 ( .A(n1917), .B(n3504), .Z(n6213) );
  NANDN U1866 ( .A(x[402]), .B(y[402]), .Z(n334) );
  ANDN U1867 ( .B(y[403]), .A(x[403]), .Z(n3498) );
  ANDN U1868 ( .B(n334), .A(n3498), .Z(n6211) );
  XOR U1869 ( .A(x[402]), .B(y[402]), .Z(n3493) );
  NANDN U1870 ( .A(y[401]), .B(x[401]), .Z(n3489) );
  NANDN U1871 ( .A(n3493), .B(n3489), .Z(n6209) );
  NANDN U1872 ( .A(x[400]), .B(y[400]), .Z(n335) );
  ANDN U1873 ( .B(y[401]), .A(x[401]), .Z(n3494) );
  ANDN U1874 ( .B(n335), .A(n3494), .Z(n6207) );
  XOR U1875 ( .A(x[400]), .B(y[400]), .Z(n3487) );
  NANDN U1876 ( .A(y[399]), .B(x[399]), .Z(n3481) );
  NANDN U1877 ( .A(n3487), .B(n3481), .Z(n6205) );
  NANDN U1878 ( .A(x[398]), .B(y[398]), .Z(n336) );
  ANDN U1879 ( .B(y[399]), .A(x[399]), .Z(n3484) );
  ANDN U1880 ( .B(n336), .A(n3484), .Z(n6203) );
  XOR U1881 ( .A(x[398]), .B(y[398]), .Z(n3477) );
  NANDN U1882 ( .A(y[397]), .B(x[397]), .Z(n1920) );
  NANDN U1883 ( .A(n3477), .B(n1920), .Z(n6201) );
  ANDN U1884 ( .B(y[396]), .A(x[396]), .Z(n3471) );
  ANDN U1885 ( .B(y[397]), .A(x[397]), .Z(n3479) );
  NOR U1886 ( .A(n3471), .B(n3479), .Z(n6199) );
  NANDN U1887 ( .A(y[395]), .B(x[395]), .Z(n3467) );
  NANDN U1888 ( .A(y[396]), .B(x[396]), .Z(n1919) );
  NAND U1889 ( .A(n3467), .B(n1919), .Z(n6197) );
  NANDN U1890 ( .A(x[394]), .B(y[394]), .Z(n337) );
  ANDN U1891 ( .B(y[395]), .A(x[395]), .Z(n3472) );
  ANDN U1892 ( .B(n337), .A(n3472), .Z(n6195) );
  XOR U1893 ( .A(x[394]), .B(y[394]), .Z(n3465) );
  NANDN U1894 ( .A(y[393]), .B(x[393]), .Z(n3459) );
  NANDN U1895 ( .A(n3465), .B(n3459), .Z(n6193) );
  NANDN U1896 ( .A(x[392]), .B(y[392]), .Z(n338) );
  ANDN U1897 ( .B(y[393]), .A(x[393]), .Z(n3462) );
  ANDN U1898 ( .B(n338), .A(n3462), .Z(n6191) );
  XOR U1899 ( .A(x[392]), .B(y[392]), .Z(n3455) );
  NANDN U1900 ( .A(y[391]), .B(x[391]), .Z(n1922) );
  NANDN U1901 ( .A(n3455), .B(n1922), .Z(n6189) );
  ANDN U1902 ( .B(y[390]), .A(x[390]), .Z(n3449) );
  ANDN U1903 ( .B(y[391]), .A(x[391]), .Z(n3457) );
  NOR U1904 ( .A(n3449), .B(n3457), .Z(n6187) );
  NANDN U1905 ( .A(y[389]), .B(x[389]), .Z(n3445) );
  NANDN U1906 ( .A(y[390]), .B(x[390]), .Z(n1921) );
  NAND U1907 ( .A(n3445), .B(n1921), .Z(n6185) );
  ANDN U1908 ( .B(y[388]), .A(x[388]), .Z(n3440) );
  ANDN U1909 ( .B(y[389]), .A(x[389]), .Z(n3450) );
  NOR U1910 ( .A(n3440), .B(n3450), .Z(n6183) );
  NANDN U1911 ( .A(y[387]), .B(x[387]), .Z(n3437) );
  NANDN U1912 ( .A(y[388]), .B(x[388]), .Z(n3444) );
  NAND U1913 ( .A(n3437), .B(n3444), .Z(n6181) );
  ANDN U1914 ( .B(y[386]), .A(x[386]), .Z(n3435) );
  ANDN U1915 ( .B(y[387]), .A(x[387]), .Z(n3443) );
  NOR U1916 ( .A(n3435), .B(n3443), .Z(n6179) );
  NANDN U1917 ( .A(y[385]), .B(x[385]), .Z(n1924) );
  NANDN U1918 ( .A(y[386]), .B(x[386]), .Z(n3438) );
  NAND U1919 ( .A(n1924), .B(n3438), .Z(n6177) );
  ANDN U1920 ( .B(y[384]), .A(x[384]), .Z(n3427) );
  ANDN U1921 ( .B(y[385]), .A(x[385]), .Z(n3432) );
  NOR U1922 ( .A(n3427), .B(n3432), .Z(n6175) );
  NANDN U1923 ( .A(y[383]), .B(x[383]), .Z(n3423) );
  NANDN U1924 ( .A(y[384]), .B(x[384]), .Z(n1923) );
  NAND U1925 ( .A(n3423), .B(n1923), .Z(n6173) );
  NANDN U1926 ( .A(x[382]), .B(y[382]), .Z(n339) );
  ANDN U1927 ( .B(y[383]), .A(x[383]), .Z(n3428) );
  ANDN U1928 ( .B(n339), .A(n3428), .Z(n6171) );
  XOR U1929 ( .A(x[382]), .B(y[382]), .Z(n3421) );
  NANDN U1930 ( .A(y[381]), .B(x[381]), .Z(n3415) );
  NANDN U1931 ( .A(n3421), .B(n3415), .Z(n6169) );
  ANDN U1932 ( .B(y[380]), .A(x[380]), .Z(n3413) );
  ANDN U1933 ( .B(y[381]), .A(x[381]), .Z(n3418) );
  NOR U1934 ( .A(n3413), .B(n3418), .Z(n6167) );
  NANDN U1935 ( .A(y[379]), .B(x[379]), .Z(n1925) );
  NANDN U1936 ( .A(y[380]), .B(x[380]), .Z(n3416) );
  NAND U1937 ( .A(n1925), .B(n3416), .Z(n6165) );
  NANDN U1938 ( .A(x[378]), .B(y[378]), .Z(n340) );
  ANDN U1939 ( .B(y[379]), .A(x[379]), .Z(n3410) );
  ANDN U1940 ( .B(n340), .A(n3410), .Z(n6163) );
  XOR U1941 ( .A(x[378]), .B(y[378]), .Z(n3405) );
  NANDN U1942 ( .A(y[377]), .B(x[377]), .Z(n3401) );
  NANDN U1943 ( .A(n3405), .B(n3401), .Z(n6161) );
  NANDN U1944 ( .A(x[376]), .B(y[376]), .Z(n341) );
  ANDN U1945 ( .B(y[377]), .A(x[377]), .Z(n3406) );
  ANDN U1946 ( .B(n341), .A(n3406), .Z(n6159) );
  XOR U1947 ( .A(x[376]), .B(y[376]), .Z(n3399) );
  NANDN U1948 ( .A(y[375]), .B(x[375]), .Z(n3393) );
  NANDN U1949 ( .A(n3399), .B(n3393), .Z(n6157) );
  ANDN U1950 ( .B(y[374]), .A(x[374]), .Z(n3391) );
  ANDN U1951 ( .B(y[375]), .A(x[375]), .Z(n3396) );
  NOR U1952 ( .A(n3391), .B(n3396), .Z(n6155) );
  NANDN U1953 ( .A(y[373]), .B(x[373]), .Z(n1927) );
  NANDN U1954 ( .A(y[374]), .B(x[374]), .Z(n3394) );
  NAND U1955 ( .A(n1927), .B(n3394), .Z(n6153) );
  NANDN U1956 ( .A(x[372]), .B(y[372]), .Z(n342) );
  ANDN U1957 ( .B(y[373]), .A(x[373]), .Z(n3388) );
  ANDN U1958 ( .B(n342), .A(n3388), .Z(n6151) );
  XOR U1959 ( .A(x[372]), .B(y[372]), .Z(n3383) );
  NANDN U1960 ( .A(y[371]), .B(x[371]), .Z(n3379) );
  NANDN U1961 ( .A(n3383), .B(n3379), .Z(n6149) );
  NANDN U1962 ( .A(x[370]), .B(y[370]), .Z(n343) );
  ANDN U1963 ( .B(y[371]), .A(x[371]), .Z(n3384) );
  ANDN U1964 ( .B(n343), .A(n3384), .Z(n6147) );
  XOR U1965 ( .A(x[370]), .B(y[370]), .Z(n3377) );
  NANDN U1966 ( .A(y[369]), .B(x[369]), .Z(n3371) );
  NANDN U1967 ( .A(n3377), .B(n3371), .Z(n6145) );
  ANDN U1968 ( .B(y[368]), .A(x[368]), .Z(n3369) );
  ANDN U1969 ( .B(y[369]), .A(x[369]), .Z(n3374) );
  NOR U1970 ( .A(n3369), .B(n3374), .Z(n6143) );
  NANDN U1971 ( .A(y[367]), .B(x[367]), .Z(n1930) );
  NANDN U1972 ( .A(y[368]), .B(x[368]), .Z(n3372) );
  NAND U1973 ( .A(n1930), .B(n3372), .Z(n6141) );
  ANDN U1974 ( .B(y[366]), .A(x[366]), .Z(n3361) );
  ANDN U1975 ( .B(y[367]), .A(x[367]), .Z(n3366) );
  NOR U1976 ( .A(n3361), .B(n3366), .Z(n6139) );
  NANDN U1977 ( .A(y[365]), .B(x[365]), .Z(n3357) );
  NANDN U1978 ( .A(y[366]), .B(x[366]), .Z(n1929) );
  NAND U1979 ( .A(n3357), .B(n1929), .Z(n6137) );
  NANDN U1980 ( .A(x[364]), .B(y[364]), .Z(n344) );
  ANDN U1981 ( .B(y[365]), .A(x[365]), .Z(n3362) );
  ANDN U1982 ( .B(n344), .A(n3362), .Z(n6135) );
  XOR U1983 ( .A(x[364]), .B(y[364]), .Z(n3355) );
  NANDN U1984 ( .A(y[363]), .B(x[363]), .Z(n3349) );
  NANDN U1985 ( .A(n3355), .B(n3349), .Z(n6133) );
  NANDN U1986 ( .A(x[362]), .B(y[362]), .Z(n345) );
  ANDN U1987 ( .B(y[363]), .A(x[363]), .Z(n3352) );
  ANDN U1988 ( .B(n345), .A(n3352), .Z(n6131) );
  XOR U1989 ( .A(x[362]), .B(y[362]), .Z(n3345) );
  NANDN U1990 ( .A(y[361]), .B(x[361]), .Z(n1932) );
  NANDN U1991 ( .A(n3345), .B(n1932), .Z(n6129) );
  ANDN U1992 ( .B(y[360]), .A(x[360]), .Z(n3339) );
  ANDN U1993 ( .B(y[361]), .A(x[361]), .Z(n3347) );
  NOR U1994 ( .A(n3339), .B(n3347), .Z(n6127) );
  NANDN U1995 ( .A(y[359]), .B(x[359]), .Z(n3335) );
  NANDN U1996 ( .A(y[360]), .B(x[360]), .Z(n1931) );
  NAND U1997 ( .A(n3335), .B(n1931), .Z(n6125) );
  NANDN U1998 ( .A(x[358]), .B(y[358]), .Z(n346) );
  ANDN U1999 ( .B(y[359]), .A(x[359]), .Z(n3340) );
  ANDN U2000 ( .B(n346), .A(n3340), .Z(n6123) );
  XOR U2001 ( .A(x[358]), .B(y[358]), .Z(n3333) );
  NANDN U2002 ( .A(y[357]), .B(x[357]), .Z(n3327) );
  NANDN U2003 ( .A(n3333), .B(n3327), .Z(n6121) );
  NANDN U2004 ( .A(x[356]), .B(y[356]), .Z(n347) );
  ANDN U2005 ( .B(y[357]), .A(x[357]), .Z(n3330) );
  ANDN U2006 ( .B(n347), .A(n3330), .Z(n6119) );
  XOR U2007 ( .A(x[356]), .B(y[356]), .Z(n3323) );
  NANDN U2008 ( .A(y[355]), .B(x[355]), .Z(n1933) );
  NANDN U2009 ( .A(n3323), .B(n1933), .Z(n6117) );
  NANDN U2010 ( .A(x[354]), .B(y[354]), .Z(n348) );
  ANDN U2011 ( .B(y[355]), .A(x[355]), .Z(n3325) );
  ANDN U2012 ( .B(n348), .A(n3325), .Z(n6115) );
  XOR U2013 ( .A(x[354]), .B(y[354]), .Z(n3317) );
  NANDN U2014 ( .A(y[353]), .B(x[353]), .Z(n3313) );
  NANDN U2015 ( .A(n3317), .B(n3313), .Z(n6113) );
  NANDN U2016 ( .A(x[352]), .B(y[352]), .Z(n349) );
  ANDN U2017 ( .B(y[353]), .A(x[353]), .Z(n3318) );
  ANDN U2018 ( .B(n349), .A(n3318), .Z(n6111) );
  XOR U2019 ( .A(x[352]), .B(y[352]), .Z(n3311) );
  NANDN U2020 ( .A(y[351]), .B(x[351]), .Z(n3305) );
  NANDN U2021 ( .A(n3311), .B(n3305), .Z(n6109) );
  ANDN U2022 ( .B(y[350]), .A(x[350]), .Z(n3303) );
  ANDN U2023 ( .B(y[351]), .A(x[351]), .Z(n3308) );
  NOR U2024 ( .A(n3303), .B(n3308), .Z(n6107) );
  NANDN U2025 ( .A(y[349]), .B(x[349]), .Z(n1935) );
  NANDN U2026 ( .A(y[350]), .B(x[350]), .Z(n3306) );
  NAND U2027 ( .A(n1935), .B(n3306), .Z(n6105) );
  NANDN U2028 ( .A(x[348]), .B(y[348]), .Z(n350) );
  ANDN U2029 ( .B(y[349]), .A(x[349]), .Z(n3300) );
  ANDN U2030 ( .B(n350), .A(n3300), .Z(n6103) );
  XOR U2031 ( .A(x[348]), .B(y[348]), .Z(n3295) );
  NANDN U2032 ( .A(y[347]), .B(x[347]), .Z(n3291) );
  NANDN U2033 ( .A(n3295), .B(n3291), .Z(n6101) );
  ANDN U2034 ( .B(y[346]), .A(x[346]), .Z(n3286) );
  ANDN U2035 ( .B(y[347]), .A(x[347]), .Z(n3296) );
  NOR U2036 ( .A(n3286), .B(n3296), .Z(n6099) );
  NANDN U2037 ( .A(y[345]), .B(x[345]), .Z(n3283) );
  NANDN U2038 ( .A(y[346]), .B(x[346]), .Z(n3293) );
  NAND U2039 ( .A(n3283), .B(n3293), .Z(n6097) );
  NANDN U2040 ( .A(x[344]), .B(y[344]), .Z(n351) );
  ANDN U2041 ( .B(y[345]), .A(x[345]), .Z(n3289) );
  ANDN U2042 ( .B(n351), .A(n3289), .Z(n6095) );
  XOR U2043 ( .A(x[344]), .B(y[344]), .Z(n3279) );
  NANDN U2044 ( .A(y[343]), .B(x[343]), .Z(n1938) );
  NANDN U2045 ( .A(n3279), .B(n1938), .Z(n6093) );
  ANDN U2046 ( .B(y[342]), .A(x[342]), .Z(n3273) );
  ANDN U2047 ( .B(y[343]), .A(x[343]), .Z(n3281) );
  NOR U2048 ( .A(n3273), .B(n3281), .Z(n6091) );
  NANDN U2049 ( .A(y[341]), .B(x[341]), .Z(n3269) );
  NANDN U2050 ( .A(y[342]), .B(x[342]), .Z(n1937) );
  NAND U2051 ( .A(n3269), .B(n1937), .Z(n6089) );
  ANDN U2052 ( .B(y[340]), .A(x[340]), .Z(n3264) );
  ANDN U2053 ( .B(y[341]), .A(x[341]), .Z(n3274) );
  NOR U2054 ( .A(n3264), .B(n3274), .Z(n6087) );
  NANDN U2055 ( .A(y[339]), .B(x[339]), .Z(n3261) );
  NANDN U2056 ( .A(y[340]), .B(x[340]), .Z(n3268) );
  NAND U2057 ( .A(n3261), .B(n3268), .Z(n6085) );
  NANDN U2058 ( .A(x[338]), .B(y[338]), .Z(n352) );
  ANDN U2059 ( .B(y[339]), .A(x[339]), .Z(n3267) );
  ANDN U2060 ( .B(n352), .A(n3267), .Z(n6083) );
  XOR U2061 ( .A(x[338]), .B(y[338]), .Z(n3257) );
  NANDN U2062 ( .A(y[337]), .B(x[337]), .Z(n1940) );
  NANDN U2063 ( .A(n3257), .B(n1940), .Z(n6081) );
  ANDN U2064 ( .B(y[336]), .A(x[336]), .Z(n3251) );
  ANDN U2065 ( .B(y[337]), .A(x[337]), .Z(n3259) );
  NOR U2066 ( .A(n3251), .B(n3259), .Z(n6079) );
  NANDN U2067 ( .A(y[335]), .B(x[335]), .Z(n3247) );
  NANDN U2068 ( .A(y[336]), .B(x[336]), .Z(n1939) );
  NAND U2069 ( .A(n3247), .B(n1939), .Z(n6077) );
  ANDN U2070 ( .B(y[334]), .A(x[334]), .Z(n3242) );
  ANDN U2071 ( .B(y[335]), .A(x[335]), .Z(n3252) );
  NOR U2072 ( .A(n3242), .B(n3252), .Z(n6075) );
  NANDN U2073 ( .A(y[333]), .B(x[333]), .Z(n3239) );
  NANDN U2074 ( .A(y[334]), .B(x[334]), .Z(n3246) );
  NAND U2075 ( .A(n3239), .B(n3246), .Z(n6073) );
  ANDN U2076 ( .B(y[332]), .A(x[332]), .Z(n3237) );
  ANDN U2077 ( .B(y[333]), .A(x[333]), .Z(n3245) );
  NOR U2078 ( .A(n3237), .B(n3245), .Z(n6071) );
  NANDN U2079 ( .A(y[331]), .B(x[331]), .Z(n1941) );
  NANDN U2080 ( .A(y[332]), .B(x[332]), .Z(n3240) );
  NAND U2081 ( .A(n1941), .B(n3240), .Z(n6069) );
  NANDN U2082 ( .A(x[330]), .B(y[330]), .Z(n353) );
  ANDN U2083 ( .B(y[331]), .A(x[331]), .Z(n3234) );
  ANDN U2084 ( .B(n353), .A(n3234), .Z(n6067) );
  XOR U2085 ( .A(x[330]), .B(y[330]), .Z(n3229) );
  NANDN U2086 ( .A(y[329]), .B(x[329]), .Z(n3225) );
  NANDN U2087 ( .A(n3229), .B(n3225), .Z(n6065) );
  ANDN U2088 ( .B(y[328]), .A(x[328]), .Z(n3220) );
  ANDN U2089 ( .B(y[329]), .A(x[329]), .Z(n3230) );
  NOR U2090 ( .A(n3220), .B(n3230), .Z(n6063) );
  NANDN U2091 ( .A(y[327]), .B(x[327]), .Z(n3217) );
  NANDN U2092 ( .A(y[328]), .B(x[328]), .Z(n3227) );
  NAND U2093 ( .A(n3217), .B(n3227), .Z(n6061) );
  ANDN U2094 ( .B(y[326]), .A(x[326]), .Z(n3215) );
  ANDN U2095 ( .B(y[327]), .A(x[327]), .Z(n3223) );
  NOR U2096 ( .A(n3215), .B(n3223), .Z(n6059) );
  NANDN U2097 ( .A(y[325]), .B(x[325]), .Z(n1944) );
  NANDN U2098 ( .A(y[326]), .B(x[326]), .Z(n3218) );
  NAND U2099 ( .A(n1944), .B(n3218), .Z(n6057) );
  ANDN U2100 ( .B(y[324]), .A(x[324]), .Z(n3207) );
  ANDN U2101 ( .B(y[325]), .A(x[325]), .Z(n3212) );
  NOR U2102 ( .A(n3207), .B(n3212), .Z(n6055) );
  NANDN U2103 ( .A(y[323]), .B(x[323]), .Z(n3203) );
  NANDN U2104 ( .A(y[324]), .B(x[324]), .Z(n1943) );
  NAND U2105 ( .A(n3203), .B(n1943), .Z(n6053) );
  ANDN U2106 ( .B(y[322]), .A(x[322]), .Z(n3198) );
  ANDN U2107 ( .B(y[323]), .A(x[323]), .Z(n3208) );
  NOR U2108 ( .A(n3198), .B(n3208), .Z(n6051) );
  NANDN U2109 ( .A(y[321]), .B(x[321]), .Z(n3195) );
  NANDN U2110 ( .A(y[322]), .B(x[322]), .Z(n3202) );
  NAND U2111 ( .A(n3195), .B(n3202), .Z(n6049) );
  ANDN U2112 ( .B(y[320]), .A(x[320]), .Z(n3193) );
  ANDN U2113 ( .B(y[321]), .A(x[321]), .Z(n3201) );
  NOR U2114 ( .A(n3193), .B(n3201), .Z(n6047) );
  NANDN U2115 ( .A(y[319]), .B(x[319]), .Z(n1946) );
  NANDN U2116 ( .A(y[320]), .B(x[320]), .Z(n3196) );
  NAND U2117 ( .A(n1946), .B(n3196), .Z(n6045) );
  ANDN U2118 ( .B(y[318]), .A(x[318]), .Z(n3185) );
  ANDN U2119 ( .B(y[319]), .A(x[319]), .Z(n3190) );
  NOR U2120 ( .A(n3185), .B(n3190), .Z(n6043) );
  NANDN U2121 ( .A(y[317]), .B(x[317]), .Z(n3181) );
  NANDN U2122 ( .A(y[318]), .B(x[318]), .Z(n1945) );
  NAND U2123 ( .A(n3181), .B(n1945), .Z(n6041) );
  ANDN U2124 ( .B(y[316]), .A(x[316]), .Z(n3176) );
  ANDN U2125 ( .B(y[317]), .A(x[317]), .Z(n3186) );
  NOR U2126 ( .A(n3176), .B(n3186), .Z(n6039) );
  NANDN U2127 ( .A(y[315]), .B(x[315]), .Z(n3173) );
  NANDN U2128 ( .A(y[316]), .B(x[316]), .Z(n3180) );
  NAND U2129 ( .A(n3173), .B(n3180), .Z(n6037) );
  NANDN U2130 ( .A(x[314]), .B(y[314]), .Z(n354) );
  ANDN U2131 ( .B(y[315]), .A(x[315]), .Z(n3179) );
  ANDN U2132 ( .B(n354), .A(n3179), .Z(n6035) );
  XOR U2133 ( .A(x[314]), .B(y[314]), .Z(n3169) );
  NANDN U2134 ( .A(y[313]), .B(x[313]), .Z(n1947) );
  NANDN U2135 ( .A(n3169), .B(n1947), .Z(n6033) );
  NANDN U2136 ( .A(x[312]), .B(y[312]), .Z(n355) );
  ANDN U2137 ( .B(y[313]), .A(x[313]), .Z(n3171) );
  ANDN U2138 ( .B(n355), .A(n3171), .Z(n6031) );
  XOR U2139 ( .A(x[312]), .B(y[312]), .Z(n3163) );
  NANDN U2140 ( .A(y[311]), .B(x[311]), .Z(n3159) );
  NANDN U2141 ( .A(n3163), .B(n3159), .Z(n6029) );
  ANDN U2142 ( .B(y[310]), .A(x[310]), .Z(n3154) );
  ANDN U2143 ( .B(y[311]), .A(x[311]), .Z(n3164) );
  NOR U2144 ( .A(n3154), .B(n3164), .Z(n6027) );
  NANDN U2145 ( .A(y[309]), .B(x[309]), .Z(n3151) );
  NANDN U2146 ( .A(y[310]), .B(x[310]), .Z(n3161) );
  NAND U2147 ( .A(n3151), .B(n3161), .Z(n6025) );
  ANDN U2148 ( .B(y[308]), .A(x[308]), .Z(n3149) );
  ANDN U2149 ( .B(y[309]), .A(x[309]), .Z(n3157) );
  NOR U2150 ( .A(n3149), .B(n3157), .Z(n6023) );
  NANDN U2151 ( .A(y[307]), .B(x[307]), .Z(n1950) );
  NANDN U2152 ( .A(y[308]), .B(x[308]), .Z(n3152) );
  NAND U2153 ( .A(n1950), .B(n3152), .Z(n6021) );
  ANDN U2154 ( .B(y[306]), .A(x[306]), .Z(n3141) );
  ANDN U2155 ( .B(y[307]), .A(x[307]), .Z(n3146) );
  NOR U2156 ( .A(n3141), .B(n3146), .Z(n6019) );
  NANDN U2157 ( .A(y[305]), .B(x[305]), .Z(n3137) );
  NANDN U2158 ( .A(y[306]), .B(x[306]), .Z(n1949) );
  NAND U2159 ( .A(n3137), .B(n1949), .Z(n6017) );
  ANDN U2160 ( .B(y[304]), .A(x[304]), .Z(n3132) );
  ANDN U2161 ( .B(y[305]), .A(x[305]), .Z(n3142) );
  NOR U2162 ( .A(n3132), .B(n3142), .Z(n6015) );
  NANDN U2163 ( .A(y[303]), .B(x[303]), .Z(n3129) );
  NANDN U2164 ( .A(y[304]), .B(x[304]), .Z(n3136) );
  NAND U2165 ( .A(n3129), .B(n3136), .Z(n6013) );
  ANDN U2166 ( .B(y[302]), .A(x[302]), .Z(n3127) );
  ANDN U2167 ( .B(y[303]), .A(x[303]), .Z(n3135) );
  NOR U2168 ( .A(n3127), .B(n3135), .Z(n6011) );
  NANDN U2169 ( .A(y[301]), .B(x[301]), .Z(n3123) );
  NANDN U2170 ( .A(y[302]), .B(x[302]), .Z(n3130) );
  NAND U2171 ( .A(n3123), .B(n3130), .Z(n6009) );
  ANDN U2172 ( .B(y[300]), .A(x[300]), .Z(n3121) );
  ANDN U2173 ( .B(y[301]), .A(x[301]), .Z(n3124) );
  NOR U2174 ( .A(n3121), .B(n3124), .Z(n6007) );
  NANDN U2175 ( .A(x[298]), .B(y[298]), .Z(n356) );
  ANDN U2176 ( .B(y[299]), .A(x[299]), .Z(n3113) );
  ANDN U2177 ( .B(n356), .A(n3113), .Z(n6003) );
  NANDN U2178 ( .A(y[297]), .B(x[297]), .Z(n3108) );
  NANDN U2179 ( .A(y[298]), .B(x[298]), .Z(n357) );
  NAND U2180 ( .A(n3108), .B(n357), .Z(n6001) );
  ANDN U2181 ( .B(y[296]), .A(x[296]), .Z(n3103) );
  ANDN U2182 ( .B(y[297]), .A(x[297]), .Z(n3112) );
  NOR U2183 ( .A(n3103), .B(n3112), .Z(n5999) );
  NANDN U2184 ( .A(y[295]), .B(x[295]), .Z(n3100) );
  NANDN U2185 ( .A(y[296]), .B(x[296]), .Z(n3107) );
  NAND U2186 ( .A(n3100), .B(n3107), .Z(n5997) );
  ANDN U2187 ( .B(y[294]), .A(x[294]), .Z(n3096) );
  ANDN U2188 ( .B(y[295]), .A(x[295]), .Z(n3106) );
  NOR U2189 ( .A(n3096), .B(n3106), .Z(n5995) );
  NANDN U2190 ( .A(y[293]), .B(x[293]), .Z(n3092) );
  NANDN U2191 ( .A(y[294]), .B(x[294]), .Z(n3101) );
  NAND U2192 ( .A(n3092), .B(n3101), .Z(n5993) );
  ANDN U2193 ( .B(y[292]), .A(x[292]), .Z(n3087) );
  ANDN U2194 ( .B(y[293]), .A(x[293]), .Z(n3098) );
  NOR U2195 ( .A(n3087), .B(n3098), .Z(n5991) );
  NANDN U2196 ( .A(y[291]), .B(x[291]), .Z(n3084) );
  NANDN U2197 ( .A(y[292]), .B(x[292]), .Z(n3091) );
  NAND U2198 ( .A(n3084), .B(n3091), .Z(n5989) );
  ANDN U2199 ( .B(y[290]), .A(x[290]), .Z(n3082) );
  ANDN U2200 ( .B(y[291]), .A(x[291]), .Z(n3090) );
  NOR U2201 ( .A(n3082), .B(n3090), .Z(n5987) );
  NANDN U2202 ( .A(y[289]), .B(x[289]), .Z(n1951) );
  NANDN U2203 ( .A(y[290]), .B(x[290]), .Z(n3085) );
  NAND U2204 ( .A(n1951), .B(n3085), .Z(n5985) );
  NANDN U2205 ( .A(x[288]), .B(y[288]), .Z(n358) );
  ANDN U2206 ( .B(y[289]), .A(x[289]), .Z(n3079) );
  ANDN U2207 ( .B(n358), .A(n3079), .Z(n5983) );
  XOR U2208 ( .A(x[288]), .B(y[288]), .Z(n3074) );
  NANDN U2209 ( .A(y[287]), .B(x[287]), .Z(n3070) );
  NANDN U2210 ( .A(n3074), .B(n3070), .Z(n5981) );
  ANDN U2211 ( .B(y[286]), .A(x[286]), .Z(n3065) );
  ANDN U2212 ( .B(y[287]), .A(x[287]), .Z(n3075) );
  NOR U2213 ( .A(n3065), .B(n3075), .Z(n5979) );
  NANDN U2214 ( .A(y[285]), .B(x[285]), .Z(n3062) );
  NANDN U2215 ( .A(y[286]), .B(x[286]), .Z(n3072) );
  NAND U2216 ( .A(n3062), .B(n3072), .Z(n5977) );
  ANDN U2217 ( .B(y[284]), .A(x[284]), .Z(n3060) );
  ANDN U2218 ( .B(y[285]), .A(x[285]), .Z(n3068) );
  NOR U2219 ( .A(n3060), .B(n3068), .Z(n5975) );
  NANDN U2220 ( .A(y[283]), .B(x[283]), .Z(n1954) );
  NANDN U2221 ( .A(y[284]), .B(x[284]), .Z(n3063) );
  NAND U2222 ( .A(n1954), .B(n3063), .Z(n5973) );
  ANDN U2223 ( .B(y[282]), .A(x[282]), .Z(n3052) );
  ANDN U2224 ( .B(y[283]), .A(x[283]), .Z(n3057) );
  NOR U2225 ( .A(n3052), .B(n3057), .Z(n5971) );
  NANDN U2226 ( .A(y[281]), .B(x[281]), .Z(n3048) );
  NANDN U2227 ( .A(y[282]), .B(x[282]), .Z(n1953) );
  NAND U2228 ( .A(n3048), .B(n1953), .Z(n5969) );
  ANDN U2229 ( .B(y[280]), .A(x[280]), .Z(n3043) );
  ANDN U2230 ( .B(y[281]), .A(x[281]), .Z(n3053) );
  NOR U2231 ( .A(n3043), .B(n3053), .Z(n5967) );
  NANDN U2232 ( .A(y[279]), .B(x[279]), .Z(n3040) );
  NANDN U2233 ( .A(y[280]), .B(x[280]), .Z(n3047) );
  NAND U2234 ( .A(n3040), .B(n3047), .Z(n5965) );
  NANDN U2235 ( .A(x[278]), .B(y[278]), .Z(n359) );
  ANDN U2236 ( .B(y[279]), .A(x[279]), .Z(n3046) );
  ANDN U2237 ( .B(n359), .A(n3046), .Z(n5963) );
  XOR U2238 ( .A(x[278]), .B(y[278]), .Z(n3036) );
  NANDN U2239 ( .A(y[277]), .B(x[277]), .Z(n1956) );
  NANDN U2240 ( .A(n3036), .B(n1956), .Z(n5961) );
  ANDN U2241 ( .B(y[276]), .A(x[276]), .Z(n3030) );
  ANDN U2242 ( .B(y[277]), .A(x[277]), .Z(n3038) );
  NOR U2243 ( .A(n3030), .B(n3038), .Z(n5959) );
  NANDN U2244 ( .A(y[275]), .B(x[275]), .Z(n3026) );
  NANDN U2245 ( .A(y[276]), .B(x[276]), .Z(n1955) );
  NAND U2246 ( .A(n3026), .B(n1955), .Z(n5957) );
  ANDN U2247 ( .B(y[274]), .A(x[274]), .Z(n3021) );
  ANDN U2248 ( .B(y[275]), .A(x[275]), .Z(n3031) );
  NOR U2249 ( .A(n3021), .B(n3031), .Z(n5955) );
  NANDN U2250 ( .A(y[273]), .B(x[273]), .Z(n3018) );
  NANDN U2251 ( .A(y[274]), .B(x[274]), .Z(n3025) );
  NAND U2252 ( .A(n3018), .B(n3025), .Z(n5953) );
  NANDN U2253 ( .A(x[272]), .B(y[272]), .Z(n360) );
  ANDN U2254 ( .B(y[273]), .A(x[273]), .Z(n3024) );
  ANDN U2255 ( .B(n360), .A(n3024), .Z(n5951) );
  XOR U2256 ( .A(x[272]), .B(y[272]), .Z(n3014) );
  NANDN U2257 ( .A(y[271]), .B(x[271]), .Z(n1958) );
  NANDN U2258 ( .A(n3014), .B(n1958), .Z(n5949) );
  ANDN U2259 ( .B(y[270]), .A(x[270]), .Z(n3008) );
  ANDN U2260 ( .B(y[271]), .A(x[271]), .Z(n3016) );
  NOR U2261 ( .A(n3008), .B(n3016), .Z(n5947) );
  NANDN U2262 ( .A(y[269]), .B(x[269]), .Z(n3004) );
  NANDN U2263 ( .A(y[270]), .B(x[270]), .Z(n1957) );
  NAND U2264 ( .A(n3004), .B(n1957), .Z(n5945) );
  ANDN U2265 ( .B(y[268]), .A(x[268]), .Z(n2999) );
  ANDN U2266 ( .B(y[269]), .A(x[269]), .Z(n3009) );
  NOR U2267 ( .A(n2999), .B(n3009), .Z(n5943) );
  NANDN U2268 ( .A(y[267]), .B(x[267]), .Z(n2996) );
  NANDN U2269 ( .A(y[268]), .B(x[268]), .Z(n3003) );
  NAND U2270 ( .A(n2996), .B(n3003), .Z(n5941) );
  NANDN U2271 ( .A(x[266]), .B(y[266]), .Z(n361) );
  ANDN U2272 ( .B(y[267]), .A(x[267]), .Z(n3002) );
  ANDN U2273 ( .B(n361), .A(n3002), .Z(n5939) );
  XOR U2274 ( .A(x[266]), .B(y[266]), .Z(n2992) );
  NANDN U2275 ( .A(y[265]), .B(x[265]), .Z(n1960) );
  NANDN U2276 ( .A(n2992), .B(n1960), .Z(n5937) );
  ANDN U2277 ( .B(y[264]), .A(x[264]), .Z(n2986) );
  ANDN U2278 ( .B(y[265]), .A(x[265]), .Z(n2994) );
  NOR U2279 ( .A(n2986), .B(n2994), .Z(n5935) );
  NANDN U2280 ( .A(y[263]), .B(x[263]), .Z(n2982) );
  NANDN U2281 ( .A(y[264]), .B(x[264]), .Z(n1959) );
  NAND U2282 ( .A(n2982), .B(n1959), .Z(n5933) );
  ANDN U2283 ( .B(y[262]), .A(x[262]), .Z(n2977) );
  ANDN U2284 ( .B(y[263]), .A(x[263]), .Z(n2987) );
  NOR U2285 ( .A(n2977), .B(n2987), .Z(n5931) );
  NANDN U2286 ( .A(y[261]), .B(x[261]), .Z(n2974) );
  NANDN U2287 ( .A(y[262]), .B(x[262]), .Z(n2981) );
  NAND U2288 ( .A(n2974), .B(n2981), .Z(n5929) );
  ANDN U2289 ( .B(y[260]), .A(x[260]), .Z(n2972) );
  ANDN U2290 ( .B(y[261]), .A(x[261]), .Z(n2980) );
  NOR U2291 ( .A(n2972), .B(n2980), .Z(n5927) );
  NANDN U2292 ( .A(y[259]), .B(x[259]), .Z(n1962) );
  NANDN U2293 ( .A(y[260]), .B(x[260]), .Z(n2975) );
  NAND U2294 ( .A(n1962), .B(n2975), .Z(n5925) );
  ANDN U2295 ( .B(y[258]), .A(x[258]), .Z(n2964) );
  ANDN U2296 ( .B(y[259]), .A(x[259]), .Z(n2969) );
  NOR U2297 ( .A(n2964), .B(n2969), .Z(n5923) );
  NANDN U2298 ( .A(y[257]), .B(x[257]), .Z(n2960) );
  NANDN U2299 ( .A(y[258]), .B(x[258]), .Z(n1961) );
  NAND U2300 ( .A(n2960), .B(n1961), .Z(n5921) );
  ANDN U2301 ( .B(y[256]), .A(x[256]), .Z(n2955) );
  ANDN U2302 ( .B(y[257]), .A(x[257]), .Z(n2965) );
  NOR U2303 ( .A(n2955), .B(n2965), .Z(n5919) );
  NANDN U2304 ( .A(y[255]), .B(x[255]), .Z(n2952) );
  NANDN U2305 ( .A(y[256]), .B(x[256]), .Z(n2959) );
  NAND U2306 ( .A(n2952), .B(n2959), .Z(n5917) );
  NANDN U2307 ( .A(x[254]), .B(y[254]), .Z(n362) );
  ANDN U2308 ( .B(y[255]), .A(x[255]), .Z(n2958) );
  ANDN U2309 ( .B(n362), .A(n2958), .Z(n5915) );
  XOR U2310 ( .A(x[254]), .B(y[254]), .Z(n2948) );
  NANDN U2311 ( .A(y[253]), .B(x[253]), .Z(n1964) );
  NANDN U2312 ( .A(n2948), .B(n1964), .Z(n5913) );
  ANDN U2313 ( .B(y[252]), .A(x[252]), .Z(n2942) );
  ANDN U2314 ( .B(y[253]), .A(x[253]), .Z(n2950) );
  NOR U2315 ( .A(n2942), .B(n2950), .Z(n5911) );
  NANDN U2316 ( .A(y[251]), .B(x[251]), .Z(n2938) );
  NANDN U2317 ( .A(y[252]), .B(x[252]), .Z(n1963) );
  NAND U2318 ( .A(n2938), .B(n1963), .Z(n5909) );
  NANDN U2319 ( .A(x[250]), .B(y[250]), .Z(n363) );
  ANDN U2320 ( .B(y[251]), .A(x[251]), .Z(n2943) );
  ANDN U2321 ( .B(n363), .A(n2943), .Z(n5907) );
  XOR U2322 ( .A(x[250]), .B(y[250]), .Z(n2936) );
  NANDN U2323 ( .A(y[249]), .B(x[249]), .Z(n2930) );
  NANDN U2324 ( .A(n2936), .B(n2930), .Z(n5905) );
  ANDN U2325 ( .B(y[248]), .A(x[248]), .Z(n2928) );
  ANDN U2326 ( .B(y[249]), .A(x[249]), .Z(n2933) );
  NOR U2327 ( .A(n2928), .B(n2933), .Z(n5903) );
  NANDN U2328 ( .A(y[247]), .B(x[247]), .Z(n1966) );
  NANDN U2329 ( .A(y[248]), .B(x[248]), .Z(n2931) );
  NAND U2330 ( .A(n1966), .B(n2931), .Z(n5901) );
  ANDN U2331 ( .B(y[246]), .A(x[246]), .Z(n2920) );
  ANDN U2332 ( .B(y[247]), .A(x[247]), .Z(n2925) );
  NOR U2333 ( .A(n2920), .B(n2925), .Z(n5899) );
  NANDN U2334 ( .A(y[245]), .B(x[245]), .Z(n2916) );
  NANDN U2335 ( .A(y[246]), .B(x[246]), .Z(n1965) );
  NAND U2336 ( .A(n2916), .B(n1965), .Z(n5897) );
  ANDN U2337 ( .B(y[244]), .A(x[244]), .Z(n2911) );
  ANDN U2338 ( .B(y[245]), .A(x[245]), .Z(n2921) );
  NOR U2339 ( .A(n2911), .B(n2921), .Z(n5895) );
  NANDN U2340 ( .A(y[243]), .B(x[243]), .Z(n2908) );
  NANDN U2341 ( .A(y[244]), .B(x[244]), .Z(n2915) );
  NAND U2342 ( .A(n2908), .B(n2915), .Z(n5893) );
  ANDN U2343 ( .B(y[242]), .A(x[242]), .Z(n2906) );
  ANDN U2344 ( .B(y[243]), .A(x[243]), .Z(n2914) );
  NOR U2345 ( .A(n2906), .B(n2914), .Z(n5891) );
  NANDN U2346 ( .A(y[241]), .B(x[241]), .Z(n1968) );
  NANDN U2347 ( .A(y[242]), .B(x[242]), .Z(n2909) );
  NAND U2348 ( .A(n1968), .B(n2909), .Z(n5889) );
  ANDN U2349 ( .B(y[240]), .A(x[240]), .Z(n2898) );
  ANDN U2350 ( .B(y[241]), .A(x[241]), .Z(n2903) );
  NOR U2351 ( .A(n2898), .B(n2903), .Z(n5887) );
  NANDN U2352 ( .A(y[239]), .B(x[239]), .Z(n2894) );
  NANDN U2353 ( .A(y[240]), .B(x[240]), .Z(n1967) );
  NAND U2354 ( .A(n2894), .B(n1967), .Z(n5885) );
  ANDN U2355 ( .B(y[238]), .A(x[238]), .Z(n2889) );
  ANDN U2356 ( .B(y[239]), .A(x[239]), .Z(n2899) );
  NOR U2357 ( .A(n2889), .B(n2899), .Z(n5883) );
  NANDN U2358 ( .A(y[237]), .B(x[237]), .Z(n2886) );
  NANDN U2359 ( .A(y[238]), .B(x[238]), .Z(n2893) );
  NAND U2360 ( .A(n2886), .B(n2893), .Z(n5881) );
  ANDN U2361 ( .B(y[236]), .A(x[236]), .Z(n2884) );
  ANDN U2362 ( .B(y[237]), .A(x[237]), .Z(n2892) );
  NOR U2363 ( .A(n2884), .B(n2892), .Z(n5879) );
  NANDN U2364 ( .A(y[235]), .B(x[235]), .Z(n1970) );
  NANDN U2365 ( .A(y[236]), .B(x[236]), .Z(n2887) );
  NAND U2366 ( .A(n1970), .B(n2887), .Z(n5877) );
  ANDN U2367 ( .B(y[234]), .A(x[234]), .Z(n2876) );
  ANDN U2368 ( .B(y[235]), .A(x[235]), .Z(n2881) );
  NOR U2369 ( .A(n2876), .B(n2881), .Z(n5875) );
  NANDN U2370 ( .A(y[233]), .B(x[233]), .Z(n2872) );
  NANDN U2371 ( .A(y[234]), .B(x[234]), .Z(n1969) );
  NAND U2372 ( .A(n2872), .B(n1969), .Z(n5873) );
  ANDN U2373 ( .B(y[232]), .A(x[232]), .Z(n2867) );
  ANDN U2374 ( .B(y[233]), .A(x[233]), .Z(n2877) );
  NOR U2375 ( .A(n2867), .B(n2877), .Z(n5871) );
  NANDN U2376 ( .A(y[231]), .B(x[231]), .Z(n2864) );
  NANDN U2377 ( .A(y[232]), .B(x[232]), .Z(n2871) );
  NAND U2378 ( .A(n2864), .B(n2871), .Z(n5869) );
  ANDN U2379 ( .B(y[230]), .A(x[230]), .Z(n2862) );
  ANDN U2380 ( .B(y[231]), .A(x[231]), .Z(n2870) );
  NOR U2381 ( .A(n2862), .B(n2870), .Z(n5867) );
  NANDN U2382 ( .A(y[229]), .B(x[229]), .Z(n1971) );
  NANDN U2383 ( .A(y[230]), .B(x[230]), .Z(n2865) );
  NAND U2384 ( .A(n1971), .B(n2865), .Z(n5865) );
  NANDN U2385 ( .A(x[228]), .B(y[228]), .Z(n364) );
  ANDN U2386 ( .B(y[229]), .A(x[229]), .Z(n2859) );
  ANDN U2387 ( .B(n364), .A(n2859), .Z(n5863) );
  XOR U2388 ( .A(x[228]), .B(y[228]), .Z(n2854) );
  NANDN U2389 ( .A(y[227]), .B(x[227]), .Z(n2850) );
  NANDN U2390 ( .A(n2854), .B(n2850), .Z(n5861) );
  ANDN U2391 ( .B(y[226]), .A(x[226]), .Z(n2845) );
  ANDN U2392 ( .B(y[227]), .A(x[227]), .Z(n2855) );
  NOR U2393 ( .A(n2845), .B(n2855), .Z(n5859) );
  NANDN U2394 ( .A(y[225]), .B(x[225]), .Z(n2842) );
  NANDN U2395 ( .A(y[226]), .B(x[226]), .Z(n2852) );
  NAND U2396 ( .A(n2842), .B(n2852), .Z(n5857) );
  NANDN U2397 ( .A(x[224]), .B(y[224]), .Z(n365) );
  ANDN U2398 ( .B(y[225]), .A(x[225]), .Z(n2848) );
  ANDN U2399 ( .B(n365), .A(n2848), .Z(n5855) );
  XOR U2400 ( .A(x[224]), .B(y[224]), .Z(n2838) );
  NANDN U2401 ( .A(y[223]), .B(x[223]), .Z(n1974) );
  NANDN U2402 ( .A(n2838), .B(n1974), .Z(n5853) );
  ANDN U2403 ( .B(y[222]), .A(x[222]), .Z(n2832) );
  ANDN U2404 ( .B(y[223]), .A(x[223]), .Z(n2840) );
  NOR U2405 ( .A(n2832), .B(n2840), .Z(n5851) );
  NANDN U2406 ( .A(y[221]), .B(x[221]), .Z(n2828) );
  NANDN U2407 ( .A(y[222]), .B(x[222]), .Z(n1973) );
  NAND U2408 ( .A(n2828), .B(n1973), .Z(n5849) );
  NANDN U2409 ( .A(x[220]), .B(y[220]), .Z(n366) );
  ANDN U2410 ( .B(y[221]), .A(x[221]), .Z(n2833) );
  ANDN U2411 ( .B(n366), .A(n2833), .Z(n5847) );
  XOR U2412 ( .A(x[220]), .B(y[220]), .Z(n2826) );
  NANDN U2413 ( .A(y[219]), .B(x[219]), .Z(n2820) );
  NANDN U2414 ( .A(n2826), .B(n2820), .Z(n5845) );
  NANDN U2415 ( .A(x[218]), .B(y[218]), .Z(n367) );
  ANDN U2416 ( .B(y[219]), .A(x[219]), .Z(n2823) );
  ANDN U2417 ( .B(n367), .A(n2823), .Z(n5843) );
  XOR U2418 ( .A(x[218]), .B(y[218]), .Z(n2816) );
  NANDN U2419 ( .A(y[217]), .B(x[217]), .Z(n1976) );
  NANDN U2420 ( .A(n2816), .B(n1976), .Z(n5841) );
  ANDN U2421 ( .B(y[216]), .A(x[216]), .Z(n2810) );
  ANDN U2422 ( .B(y[217]), .A(x[217]), .Z(n2818) );
  NOR U2423 ( .A(n2810), .B(n2818), .Z(n5839) );
  NANDN U2424 ( .A(y[215]), .B(x[215]), .Z(n2806) );
  NANDN U2425 ( .A(y[216]), .B(x[216]), .Z(n1975) );
  NAND U2426 ( .A(n2806), .B(n1975), .Z(n5837) );
  ANDN U2427 ( .B(y[214]), .A(x[214]), .Z(n2801) );
  ANDN U2428 ( .B(y[215]), .A(x[215]), .Z(n2811) );
  NOR U2429 ( .A(n2801), .B(n2811), .Z(n5835) );
  NANDN U2430 ( .A(y[213]), .B(x[213]), .Z(n2798) );
  NANDN U2431 ( .A(y[214]), .B(x[214]), .Z(n2805) );
  NAND U2432 ( .A(n2798), .B(n2805), .Z(n5833) );
  ANDN U2433 ( .B(y[212]), .A(x[212]), .Z(n2796) );
  ANDN U2434 ( .B(y[213]), .A(x[213]), .Z(n2804) );
  NOR U2435 ( .A(n2796), .B(n2804), .Z(n5831) );
  NANDN U2436 ( .A(y[211]), .B(x[211]), .Z(n1978) );
  NANDN U2437 ( .A(y[212]), .B(x[212]), .Z(n2799) );
  NAND U2438 ( .A(n1978), .B(n2799), .Z(n5829) );
  ANDN U2439 ( .B(y[210]), .A(x[210]), .Z(n2788) );
  ANDN U2440 ( .B(y[211]), .A(x[211]), .Z(n2793) );
  NOR U2441 ( .A(n2788), .B(n2793), .Z(n5827) );
  NANDN U2442 ( .A(y[209]), .B(x[209]), .Z(n2784) );
  NANDN U2443 ( .A(y[210]), .B(x[210]), .Z(n1977) );
  NAND U2444 ( .A(n2784), .B(n1977), .Z(n5825) );
  NANDN U2445 ( .A(x[208]), .B(y[208]), .Z(n368) );
  ANDN U2446 ( .B(y[209]), .A(x[209]), .Z(n2789) );
  ANDN U2447 ( .B(n368), .A(n2789), .Z(n5823) );
  XOR U2448 ( .A(x[208]), .B(y[208]), .Z(n2782) );
  NANDN U2449 ( .A(y[207]), .B(x[207]), .Z(n2776) );
  NANDN U2450 ( .A(n2782), .B(n2776), .Z(n5821) );
  ANDN U2451 ( .B(y[206]), .A(x[206]), .Z(n2774) );
  ANDN U2452 ( .B(y[207]), .A(x[207]), .Z(n2779) );
  NOR U2453 ( .A(n2774), .B(n2779), .Z(n5819) );
  NANDN U2454 ( .A(y[205]), .B(x[205]), .Z(n1980) );
  NANDN U2455 ( .A(y[206]), .B(x[206]), .Z(n2777) );
  NAND U2456 ( .A(n1980), .B(n2777), .Z(n5817) );
  ANDN U2457 ( .B(y[204]), .A(x[204]), .Z(n2766) );
  ANDN U2458 ( .B(y[205]), .A(x[205]), .Z(n2771) );
  NOR U2459 ( .A(n2766), .B(n2771), .Z(n5815) );
  NANDN U2460 ( .A(y[203]), .B(x[203]), .Z(n2762) );
  NANDN U2461 ( .A(y[204]), .B(x[204]), .Z(n1979) );
  NAND U2462 ( .A(n2762), .B(n1979), .Z(n5813) );
  ANDN U2463 ( .B(y[202]), .A(x[202]), .Z(n2757) );
  ANDN U2464 ( .B(y[203]), .A(x[203]), .Z(n2767) );
  NOR U2465 ( .A(n2757), .B(n2767), .Z(n5811) );
  NANDN U2466 ( .A(y[201]), .B(x[201]), .Z(n2754) );
  NANDN U2467 ( .A(y[202]), .B(x[202]), .Z(n2761) );
  NAND U2468 ( .A(n2754), .B(n2761), .Z(n5809) );
  ANDN U2469 ( .B(y[200]), .A(x[200]), .Z(n2752) );
  ANDN U2470 ( .B(y[201]), .A(x[201]), .Z(n2760) );
  NOR U2471 ( .A(n2752), .B(n2760), .Z(n5807) );
  NANDN U2472 ( .A(y[199]), .B(x[199]), .Z(n1982) );
  NANDN U2473 ( .A(y[200]), .B(x[200]), .Z(n2755) );
  NAND U2474 ( .A(n1982), .B(n2755), .Z(n5805) );
  ANDN U2475 ( .B(y[198]), .A(x[198]), .Z(n2744) );
  ANDN U2476 ( .B(y[199]), .A(x[199]), .Z(n2749) );
  NOR U2477 ( .A(n2744), .B(n2749), .Z(n5803) );
  NANDN U2478 ( .A(y[197]), .B(x[197]), .Z(n2740) );
  NANDN U2479 ( .A(y[198]), .B(x[198]), .Z(n1981) );
  NAND U2480 ( .A(n2740), .B(n1981), .Z(n5801) );
  ANDN U2481 ( .B(y[196]), .A(x[196]), .Z(n2735) );
  ANDN U2482 ( .B(y[197]), .A(x[197]), .Z(n2745) );
  NOR U2483 ( .A(n2735), .B(n2745), .Z(n5799) );
  NANDN U2484 ( .A(y[195]), .B(x[195]), .Z(n2732) );
  NANDN U2485 ( .A(y[196]), .B(x[196]), .Z(n2739) );
  NAND U2486 ( .A(n2732), .B(n2739), .Z(n5797) );
  ANDN U2487 ( .B(y[194]), .A(x[194]), .Z(n2730) );
  ANDN U2488 ( .B(y[195]), .A(x[195]), .Z(n2738) );
  NOR U2489 ( .A(n2730), .B(n2738), .Z(n5795) );
  NANDN U2490 ( .A(y[193]), .B(x[193]), .Z(n1984) );
  NANDN U2491 ( .A(y[194]), .B(x[194]), .Z(n2733) );
  NAND U2492 ( .A(n1984), .B(n2733), .Z(n5793) );
  ANDN U2493 ( .B(y[192]), .A(x[192]), .Z(n2722) );
  ANDN U2494 ( .B(y[193]), .A(x[193]), .Z(n2727) );
  NOR U2495 ( .A(n2722), .B(n2727), .Z(n5791) );
  NANDN U2496 ( .A(y[191]), .B(x[191]), .Z(n2718) );
  NANDN U2497 ( .A(y[192]), .B(x[192]), .Z(n1983) );
  NAND U2498 ( .A(n2718), .B(n1983), .Z(n5789) );
  ANDN U2499 ( .B(y[190]), .A(x[190]), .Z(n2713) );
  ANDN U2500 ( .B(y[191]), .A(x[191]), .Z(n2723) );
  NOR U2501 ( .A(n2713), .B(n2723), .Z(n5787) );
  NANDN U2502 ( .A(y[189]), .B(x[189]), .Z(n2710) );
  NANDN U2503 ( .A(y[190]), .B(x[190]), .Z(n2717) );
  NAND U2504 ( .A(n2710), .B(n2717), .Z(n5785) );
  ANDN U2505 ( .B(y[188]), .A(x[188]), .Z(n2708) );
  ANDN U2506 ( .B(y[189]), .A(x[189]), .Z(n2716) );
  NOR U2507 ( .A(n2708), .B(n2716), .Z(n5783) );
  NANDN U2508 ( .A(y[187]), .B(x[187]), .Z(n1986) );
  NANDN U2509 ( .A(y[188]), .B(x[188]), .Z(n2711) );
  NAND U2510 ( .A(n1986), .B(n2711), .Z(n5781) );
  ANDN U2511 ( .B(y[186]), .A(x[186]), .Z(n2700) );
  ANDN U2512 ( .B(y[187]), .A(x[187]), .Z(n2705) );
  NOR U2513 ( .A(n2700), .B(n2705), .Z(n5779) );
  NANDN U2514 ( .A(y[185]), .B(x[185]), .Z(n2696) );
  NANDN U2515 ( .A(y[186]), .B(x[186]), .Z(n1985) );
  NAND U2516 ( .A(n2696), .B(n1985), .Z(n5777) );
  NANDN U2517 ( .A(x[184]), .B(y[184]), .Z(n369) );
  ANDN U2518 ( .B(y[185]), .A(x[185]), .Z(n2701) );
  ANDN U2519 ( .B(n369), .A(n2701), .Z(n5775) );
  XOR U2520 ( .A(x[184]), .B(y[184]), .Z(n2694) );
  NANDN U2521 ( .A(y[183]), .B(x[183]), .Z(n2688) );
  NANDN U2522 ( .A(n2694), .B(n2688), .Z(n5773) );
  ANDN U2523 ( .B(y[182]), .A(x[182]), .Z(n2686) );
  ANDN U2524 ( .B(y[183]), .A(x[183]), .Z(n2691) );
  NOR U2525 ( .A(n2686), .B(n2691), .Z(n5771) );
  NANDN U2526 ( .A(y[181]), .B(x[181]), .Z(n1988) );
  NANDN U2527 ( .A(y[182]), .B(x[182]), .Z(n2689) );
  NAND U2528 ( .A(n1988), .B(n2689), .Z(n5769) );
  ANDN U2529 ( .B(y[180]), .A(x[180]), .Z(n2678) );
  ANDN U2530 ( .B(y[181]), .A(x[181]), .Z(n2683) );
  NOR U2531 ( .A(n2678), .B(n2683), .Z(n5767) );
  NANDN U2532 ( .A(y[179]), .B(x[179]), .Z(n2674) );
  NANDN U2533 ( .A(y[180]), .B(x[180]), .Z(n1987) );
  NAND U2534 ( .A(n2674), .B(n1987), .Z(n5765) );
  ANDN U2535 ( .B(y[178]), .A(x[178]), .Z(n2669) );
  ANDN U2536 ( .B(y[179]), .A(x[179]), .Z(n2679) );
  NOR U2537 ( .A(n2669), .B(n2679), .Z(n5763) );
  NANDN U2538 ( .A(y[177]), .B(x[177]), .Z(n2666) );
  NANDN U2539 ( .A(y[178]), .B(x[178]), .Z(n2673) );
  NAND U2540 ( .A(n2666), .B(n2673), .Z(n5761) );
  NANDN U2541 ( .A(x[176]), .B(y[176]), .Z(n370) );
  ANDN U2542 ( .B(y[177]), .A(x[177]), .Z(n2672) );
  ANDN U2543 ( .B(n370), .A(n2672), .Z(n5759) );
  XOR U2544 ( .A(x[176]), .B(y[176]), .Z(n2662) );
  NANDN U2545 ( .A(y[175]), .B(x[175]), .Z(n1990) );
  NANDN U2546 ( .A(n2662), .B(n1990), .Z(n5757) );
  ANDN U2547 ( .B(y[174]), .A(x[174]), .Z(n2656) );
  ANDN U2548 ( .B(y[175]), .A(x[175]), .Z(n2664) );
  NOR U2549 ( .A(n2656), .B(n2664), .Z(n5755) );
  NANDN U2550 ( .A(y[173]), .B(x[173]), .Z(n2652) );
  NANDN U2551 ( .A(y[174]), .B(x[174]), .Z(n1989) );
  NAND U2552 ( .A(n2652), .B(n1989), .Z(n5753) );
  ANDN U2553 ( .B(y[172]), .A(x[172]), .Z(n2647) );
  ANDN U2554 ( .B(y[173]), .A(x[173]), .Z(n2657) );
  NOR U2555 ( .A(n2647), .B(n2657), .Z(n5751) );
  NANDN U2556 ( .A(y[171]), .B(x[171]), .Z(n2644) );
  NANDN U2557 ( .A(y[172]), .B(x[172]), .Z(n2651) );
  NAND U2558 ( .A(n2644), .B(n2651), .Z(n5749) );
  NANDN U2559 ( .A(x[170]), .B(y[170]), .Z(n371) );
  ANDN U2560 ( .B(y[171]), .A(x[171]), .Z(n2650) );
  ANDN U2561 ( .B(n371), .A(n2650), .Z(n5747) );
  XOR U2562 ( .A(x[170]), .B(y[170]), .Z(n2640) );
  NANDN U2563 ( .A(y[169]), .B(x[169]), .Z(n1991) );
  NANDN U2564 ( .A(n2640), .B(n1991), .Z(n5745) );
  NANDN U2565 ( .A(x[168]), .B(y[168]), .Z(n372) );
  ANDN U2566 ( .B(y[169]), .A(x[169]), .Z(n2642) );
  ANDN U2567 ( .B(n372), .A(n2642), .Z(n5743) );
  XOR U2568 ( .A(x[168]), .B(y[168]), .Z(n2634) );
  NANDN U2569 ( .A(y[167]), .B(x[167]), .Z(n2630) );
  NANDN U2570 ( .A(n2634), .B(n2630), .Z(n5741) );
  NANDN U2571 ( .A(x[166]), .B(y[166]), .Z(n373) );
  ANDN U2572 ( .B(y[167]), .A(x[167]), .Z(n2635) );
  ANDN U2573 ( .B(n373), .A(n2635), .Z(n5739) );
  XOR U2574 ( .A(x[166]), .B(y[166]), .Z(n2628) );
  NANDN U2575 ( .A(y[165]), .B(x[165]), .Z(n2622) );
  NANDN U2576 ( .A(n2628), .B(n2622), .Z(n5737) );
  ANDN U2577 ( .B(y[164]), .A(x[164]), .Z(n2620) );
  ANDN U2578 ( .B(y[165]), .A(x[165]), .Z(n2625) );
  NOR U2579 ( .A(n2620), .B(n2625), .Z(n5735) );
  NANDN U2580 ( .A(y[163]), .B(x[163]), .Z(n1993) );
  NANDN U2581 ( .A(y[164]), .B(x[164]), .Z(n2623) );
  NAND U2582 ( .A(n1993), .B(n2623), .Z(n5733) );
  NANDN U2583 ( .A(x[162]), .B(y[162]), .Z(n374) );
  ANDN U2584 ( .B(y[163]), .A(x[163]), .Z(n2617) );
  ANDN U2585 ( .B(n374), .A(n2617), .Z(n5731) );
  XOR U2586 ( .A(x[162]), .B(y[162]), .Z(n2612) );
  NANDN U2587 ( .A(y[161]), .B(x[161]), .Z(n2608) );
  NANDN U2588 ( .A(n2612), .B(n2608), .Z(n5729) );
  ANDN U2589 ( .B(y[160]), .A(x[160]), .Z(n2603) );
  ANDN U2590 ( .B(y[161]), .A(x[161]), .Z(n2613) );
  NOR U2591 ( .A(n2603), .B(n2613), .Z(n5727) );
  NANDN U2592 ( .A(y[159]), .B(x[159]), .Z(n2600) );
  NANDN U2593 ( .A(y[160]), .B(x[160]), .Z(n2610) );
  NAND U2594 ( .A(n2600), .B(n2610), .Z(n5725) );
  ANDN U2595 ( .B(y[158]), .A(x[158]), .Z(n2598) );
  ANDN U2596 ( .B(y[159]), .A(x[159]), .Z(n2606) );
  NOR U2597 ( .A(n2598), .B(n2606), .Z(n5723) );
  NANDN U2598 ( .A(y[157]), .B(x[157]), .Z(n1996) );
  NANDN U2599 ( .A(y[158]), .B(x[158]), .Z(n2601) );
  NAND U2600 ( .A(n1996), .B(n2601), .Z(n5721) );
  ANDN U2601 ( .B(y[156]), .A(x[156]), .Z(n2590) );
  ANDN U2602 ( .B(y[157]), .A(x[157]), .Z(n2595) );
  NOR U2603 ( .A(n2590), .B(n2595), .Z(n5719) );
  NANDN U2604 ( .A(y[155]), .B(x[155]), .Z(n2586) );
  NANDN U2605 ( .A(y[156]), .B(x[156]), .Z(n1995) );
  NAND U2606 ( .A(n2586), .B(n1995), .Z(n5717) );
  ANDN U2607 ( .B(y[154]), .A(x[154]), .Z(n2581) );
  ANDN U2608 ( .B(y[155]), .A(x[155]), .Z(n2591) );
  NOR U2609 ( .A(n2581), .B(n2591), .Z(n5715) );
  NANDN U2610 ( .A(y[153]), .B(x[153]), .Z(n2578) );
  NANDN U2611 ( .A(y[154]), .B(x[154]), .Z(n2585) );
  NAND U2612 ( .A(n2578), .B(n2585), .Z(n5713) );
  ANDN U2613 ( .B(y[152]), .A(x[152]), .Z(n2576) );
  ANDN U2614 ( .B(y[153]), .A(x[153]), .Z(n2584) );
  NOR U2615 ( .A(n2576), .B(n2584), .Z(n5711) );
  NANDN U2616 ( .A(y[151]), .B(x[151]), .Z(n1998) );
  NANDN U2617 ( .A(y[152]), .B(x[152]), .Z(n2579) );
  NAND U2618 ( .A(n1998), .B(n2579), .Z(n5709) );
  ANDN U2619 ( .B(y[150]), .A(x[150]), .Z(n2568) );
  ANDN U2620 ( .B(y[151]), .A(x[151]), .Z(n2573) );
  NOR U2621 ( .A(n2568), .B(n2573), .Z(n5707) );
  NANDN U2622 ( .A(y[149]), .B(x[149]), .Z(n2564) );
  NANDN U2623 ( .A(y[150]), .B(x[150]), .Z(n1997) );
  NAND U2624 ( .A(n2564), .B(n1997), .Z(n5705) );
  ANDN U2625 ( .B(y[148]), .A(x[148]), .Z(n2559) );
  ANDN U2626 ( .B(y[149]), .A(x[149]), .Z(n2569) );
  NOR U2627 ( .A(n2559), .B(n2569), .Z(n5703) );
  NANDN U2628 ( .A(y[147]), .B(x[147]), .Z(n2556) );
  NANDN U2629 ( .A(y[148]), .B(x[148]), .Z(n2563) );
  NAND U2630 ( .A(n2556), .B(n2563), .Z(n5701) );
  NANDN U2631 ( .A(x[146]), .B(y[146]), .Z(n375) );
  ANDN U2632 ( .B(y[147]), .A(x[147]), .Z(n2562) );
  ANDN U2633 ( .B(n375), .A(n2562), .Z(n5699) );
  XOR U2634 ( .A(x[146]), .B(y[146]), .Z(n2552) );
  NANDN U2635 ( .A(y[145]), .B(x[145]), .Z(n2000) );
  NANDN U2636 ( .A(n2552), .B(n2000), .Z(n5697) );
  ANDN U2637 ( .B(y[144]), .A(x[144]), .Z(n2546) );
  ANDN U2638 ( .B(y[145]), .A(x[145]), .Z(n2554) );
  NOR U2639 ( .A(n2546), .B(n2554), .Z(n5695) );
  NANDN U2640 ( .A(y[143]), .B(x[143]), .Z(n2542) );
  NANDN U2641 ( .A(y[144]), .B(x[144]), .Z(n1999) );
  NAND U2642 ( .A(n2542), .B(n1999), .Z(n5693) );
  ANDN U2643 ( .B(y[142]), .A(x[142]), .Z(n2537) );
  ANDN U2644 ( .B(y[143]), .A(x[143]), .Z(n2547) );
  NOR U2645 ( .A(n2537), .B(n2547), .Z(n5691) );
  NANDN U2646 ( .A(y[141]), .B(x[141]), .Z(n2534) );
  NANDN U2647 ( .A(y[142]), .B(x[142]), .Z(n2541) );
  NAND U2648 ( .A(n2534), .B(n2541), .Z(n5689) );
  ANDN U2649 ( .B(y[140]), .A(x[140]), .Z(n2532) );
  ANDN U2650 ( .B(y[141]), .A(x[141]), .Z(n2540) );
  NOR U2651 ( .A(n2532), .B(n2540), .Z(n5687) );
  NANDN U2652 ( .A(y[139]), .B(x[139]), .Z(n2002) );
  NANDN U2653 ( .A(y[140]), .B(x[140]), .Z(n2535) );
  NAND U2654 ( .A(n2002), .B(n2535), .Z(n5685) );
  ANDN U2655 ( .B(y[138]), .A(x[138]), .Z(n2524) );
  ANDN U2656 ( .B(y[139]), .A(x[139]), .Z(n2529) );
  NOR U2657 ( .A(n2524), .B(n2529), .Z(n5683) );
  NANDN U2658 ( .A(y[137]), .B(x[137]), .Z(n2520) );
  NANDN U2659 ( .A(y[138]), .B(x[138]), .Z(n2001) );
  NAND U2660 ( .A(n2520), .B(n2001), .Z(n5681) );
  ANDN U2661 ( .B(y[136]), .A(x[136]), .Z(n2515) );
  ANDN U2662 ( .B(y[137]), .A(x[137]), .Z(n2525) );
  NOR U2663 ( .A(n2515), .B(n2525), .Z(n5679) );
  NANDN U2664 ( .A(y[135]), .B(x[135]), .Z(n2512) );
  NANDN U2665 ( .A(y[136]), .B(x[136]), .Z(n2519) );
  NAND U2666 ( .A(n2512), .B(n2519), .Z(n5677) );
  ANDN U2667 ( .B(y[134]), .A(x[134]), .Z(n2510) );
  ANDN U2668 ( .B(y[135]), .A(x[135]), .Z(n2518) );
  NOR U2669 ( .A(n2510), .B(n2518), .Z(n5675) );
  NANDN U2670 ( .A(y[133]), .B(x[133]), .Z(n2004) );
  NANDN U2671 ( .A(y[134]), .B(x[134]), .Z(n2513) );
  NAND U2672 ( .A(n2004), .B(n2513), .Z(n5673) );
  ANDN U2673 ( .B(y[132]), .A(x[132]), .Z(n2502) );
  ANDN U2674 ( .B(y[133]), .A(x[133]), .Z(n2507) );
  NOR U2675 ( .A(n2502), .B(n2507), .Z(n5671) );
  NANDN U2676 ( .A(y[131]), .B(x[131]), .Z(n2498) );
  NANDN U2677 ( .A(y[132]), .B(x[132]), .Z(n2003) );
  NAND U2678 ( .A(n2498), .B(n2003), .Z(n5669) );
  ANDN U2679 ( .B(y[130]), .A(x[130]), .Z(n2493) );
  ANDN U2680 ( .B(y[131]), .A(x[131]), .Z(n2503) );
  NOR U2681 ( .A(n2493), .B(n2503), .Z(n5667) );
  NANDN U2682 ( .A(y[129]), .B(x[129]), .Z(n2490) );
  NANDN U2683 ( .A(y[130]), .B(x[130]), .Z(n2497) );
  NAND U2684 ( .A(n2490), .B(n2497), .Z(n5665) );
  ANDN U2685 ( .B(y[128]), .A(x[128]), .Z(n2488) );
  ANDN U2686 ( .B(y[129]), .A(x[129]), .Z(n2496) );
  NOR U2687 ( .A(n2488), .B(n2496), .Z(n5663) );
  NANDN U2688 ( .A(y[127]), .B(x[127]), .Z(n2006) );
  NANDN U2689 ( .A(y[128]), .B(x[128]), .Z(n2491) );
  NAND U2690 ( .A(n2006), .B(n2491), .Z(n5661) );
  ANDN U2691 ( .B(y[126]), .A(x[126]), .Z(n2480) );
  ANDN U2692 ( .B(y[127]), .A(x[127]), .Z(n2485) );
  NOR U2693 ( .A(n2480), .B(n2485), .Z(n5659) );
  NANDN U2694 ( .A(y[125]), .B(x[125]), .Z(n2476) );
  NANDN U2695 ( .A(y[126]), .B(x[126]), .Z(n2005) );
  NAND U2696 ( .A(n2476), .B(n2005), .Z(n5657) );
  ANDN U2697 ( .B(y[124]), .A(x[124]), .Z(n2471) );
  ANDN U2698 ( .B(y[125]), .A(x[125]), .Z(n2481) );
  NOR U2699 ( .A(n2471), .B(n2481), .Z(n5655) );
  NANDN U2700 ( .A(y[123]), .B(x[123]), .Z(n2468) );
  NANDN U2701 ( .A(y[124]), .B(x[124]), .Z(n2475) );
  NAND U2702 ( .A(n2468), .B(n2475), .Z(n5653) );
  ANDN U2703 ( .B(y[122]), .A(x[122]), .Z(n2466) );
  ANDN U2704 ( .B(y[123]), .A(x[123]), .Z(n2474) );
  NOR U2705 ( .A(n2466), .B(n2474), .Z(n5651) );
  NANDN U2706 ( .A(y[121]), .B(x[121]), .Z(n2008) );
  NANDN U2707 ( .A(y[122]), .B(x[122]), .Z(n2469) );
  NAND U2708 ( .A(n2008), .B(n2469), .Z(n5649) );
  ANDN U2709 ( .B(y[120]), .A(x[120]), .Z(n2458) );
  ANDN U2710 ( .B(y[121]), .A(x[121]), .Z(n2463) );
  NOR U2711 ( .A(n2458), .B(n2463), .Z(n5647) );
  NANDN U2712 ( .A(y[119]), .B(x[119]), .Z(n2454) );
  NANDN U2713 ( .A(y[120]), .B(x[120]), .Z(n2007) );
  NAND U2714 ( .A(n2454), .B(n2007), .Z(n5645) );
  ANDN U2715 ( .B(y[118]), .A(x[118]), .Z(n2449) );
  ANDN U2716 ( .B(y[119]), .A(x[119]), .Z(n2459) );
  NOR U2717 ( .A(n2449), .B(n2459), .Z(n5643) );
  NANDN U2718 ( .A(y[117]), .B(x[117]), .Z(n2446) );
  NANDN U2719 ( .A(y[118]), .B(x[118]), .Z(n2453) );
  NAND U2720 ( .A(n2446), .B(n2453), .Z(n5641) );
  ANDN U2721 ( .B(y[116]), .A(x[116]), .Z(n2444) );
  ANDN U2722 ( .B(y[117]), .A(x[117]), .Z(n2452) );
  NOR U2723 ( .A(n2444), .B(n2452), .Z(n5639) );
  NANDN U2724 ( .A(y[115]), .B(x[115]), .Z(n2009) );
  NANDN U2725 ( .A(y[116]), .B(x[116]), .Z(n2447) );
  NAND U2726 ( .A(n2009), .B(n2447), .Z(n5637) );
  NANDN U2727 ( .A(x[114]), .B(y[114]), .Z(n376) );
  ANDN U2728 ( .B(y[115]), .A(x[115]), .Z(n2441) );
  ANDN U2729 ( .B(n376), .A(n2441), .Z(n5635) );
  XOR U2730 ( .A(x[114]), .B(y[114]), .Z(n2436) );
  NANDN U2731 ( .A(y[113]), .B(x[113]), .Z(n2432) );
  NANDN U2732 ( .A(n2436), .B(n2432), .Z(n5633) );
  ANDN U2733 ( .B(y[112]), .A(x[112]), .Z(n2427) );
  ANDN U2734 ( .B(y[113]), .A(x[113]), .Z(n2437) );
  NOR U2735 ( .A(n2427), .B(n2437), .Z(n5631) );
  NANDN U2736 ( .A(y[111]), .B(x[111]), .Z(n2424) );
  NANDN U2737 ( .A(y[112]), .B(x[112]), .Z(n2434) );
  NAND U2738 ( .A(n2424), .B(n2434), .Z(n5629) );
  NANDN U2739 ( .A(x[110]), .B(y[110]), .Z(n377) );
  ANDN U2740 ( .B(y[111]), .A(x[111]), .Z(n2430) );
  ANDN U2741 ( .B(n377), .A(n2430), .Z(n5627) );
  XOR U2742 ( .A(x[110]), .B(y[110]), .Z(n2420) );
  NANDN U2743 ( .A(y[109]), .B(x[109]), .Z(n2012) );
  NANDN U2744 ( .A(n2420), .B(n2012), .Z(n5625) );
  ANDN U2745 ( .B(y[108]), .A(x[108]), .Z(n2414) );
  ANDN U2746 ( .B(y[109]), .A(x[109]), .Z(n2422) );
  NOR U2747 ( .A(n2414), .B(n2422), .Z(n5623) );
  NANDN U2748 ( .A(y[107]), .B(x[107]), .Z(n2410) );
  NANDN U2749 ( .A(y[108]), .B(x[108]), .Z(n2011) );
  NAND U2750 ( .A(n2410), .B(n2011), .Z(n5621) );
  NANDN U2751 ( .A(x[106]), .B(y[106]), .Z(n378) );
  ANDN U2752 ( .B(y[107]), .A(x[107]), .Z(n2415) );
  ANDN U2753 ( .B(n378), .A(n2415), .Z(n5619) );
  XOR U2754 ( .A(x[106]), .B(y[106]), .Z(n2408) );
  NANDN U2755 ( .A(y[105]), .B(x[105]), .Z(n2402) );
  NANDN U2756 ( .A(n2408), .B(n2402), .Z(n5617) );
  NANDN U2757 ( .A(x[104]), .B(y[104]), .Z(n379) );
  ANDN U2758 ( .B(y[105]), .A(x[105]), .Z(n2405) );
  ANDN U2759 ( .B(n379), .A(n2405), .Z(n5615) );
  XOR U2760 ( .A(x[104]), .B(y[104]), .Z(n2398) );
  NANDN U2761 ( .A(y[103]), .B(x[103]), .Z(n2014) );
  NANDN U2762 ( .A(n2398), .B(n2014), .Z(n5613) );
  ANDN U2763 ( .B(y[102]), .A(x[102]), .Z(n2392) );
  ANDN U2764 ( .B(y[103]), .A(x[103]), .Z(n2400) );
  NOR U2765 ( .A(n2392), .B(n2400), .Z(n5611) );
  NANDN U2766 ( .A(y[101]), .B(x[101]), .Z(n2388) );
  NANDN U2767 ( .A(y[102]), .B(x[102]), .Z(n2013) );
  NAND U2768 ( .A(n2388), .B(n2013), .Z(n5609) );
  NANDN U2769 ( .A(x[100]), .B(y[100]), .Z(n380) );
  ANDN U2770 ( .B(y[101]), .A(x[101]), .Z(n2393) );
  ANDN U2771 ( .B(n380), .A(n2393), .Z(n5607) );
  XOR U2772 ( .A(x[100]), .B(y[100]), .Z(n2386) );
  NANDN U2773 ( .A(y[99]), .B(x[99]), .Z(n2380) );
  NANDN U2774 ( .A(n2386), .B(n2380), .Z(n5605) );
  ANDN U2775 ( .B(y[98]), .A(x[98]), .Z(n2378) );
  ANDN U2776 ( .B(y[99]), .A(x[99]), .Z(n2383) );
  NOR U2777 ( .A(n2378), .B(n2383), .Z(n5603) );
  NANDN U2778 ( .A(y[97]), .B(x[97]), .Z(n2016) );
  NANDN U2779 ( .A(y[98]), .B(x[98]), .Z(n2381) );
  NAND U2780 ( .A(n2016), .B(n2381), .Z(n5601) );
  ANDN U2781 ( .B(y[96]), .A(x[96]), .Z(n2370) );
  ANDN U2782 ( .B(y[97]), .A(x[97]), .Z(n2375) );
  NOR U2783 ( .A(n2370), .B(n2375), .Z(n5599) );
  NANDN U2784 ( .A(y[95]), .B(x[95]), .Z(n2366) );
  NANDN U2785 ( .A(y[96]), .B(x[96]), .Z(n2015) );
  NAND U2786 ( .A(n2366), .B(n2015), .Z(n5597) );
  ANDN U2787 ( .B(y[94]), .A(x[94]), .Z(n2361) );
  ANDN U2788 ( .B(y[95]), .A(x[95]), .Z(n2371) );
  NOR U2789 ( .A(n2361), .B(n2371), .Z(n5595) );
  NANDN U2790 ( .A(y[93]), .B(x[93]), .Z(n2358) );
  NANDN U2791 ( .A(y[94]), .B(x[94]), .Z(n2365) );
  NAND U2792 ( .A(n2358), .B(n2365), .Z(n5593) );
  ANDN U2793 ( .B(y[92]), .A(x[92]), .Z(n2356) );
  ANDN U2794 ( .B(y[93]), .A(x[93]), .Z(n2364) );
  NOR U2795 ( .A(n2356), .B(n2364), .Z(n5591) );
  NANDN U2796 ( .A(y[91]), .B(x[91]), .Z(n2017) );
  NANDN U2797 ( .A(y[92]), .B(x[92]), .Z(n2359) );
  NAND U2798 ( .A(n2017), .B(n2359), .Z(n5589) );
  NANDN U2799 ( .A(x[90]), .B(y[90]), .Z(n381) );
  ANDN U2800 ( .B(y[91]), .A(x[91]), .Z(n2353) );
  ANDN U2801 ( .B(n381), .A(n2353), .Z(n5587) );
  XOR U2802 ( .A(x[90]), .B(y[90]), .Z(n2348) );
  NANDN U2803 ( .A(y[89]), .B(x[89]), .Z(n2344) );
  NANDN U2804 ( .A(n2348), .B(n2344), .Z(n5585) );
  ANDN U2805 ( .B(y[88]), .A(x[88]), .Z(n2339) );
  ANDN U2806 ( .B(y[89]), .A(x[89]), .Z(n2349) );
  NOR U2807 ( .A(n2339), .B(n2349), .Z(n5583) );
  NANDN U2808 ( .A(y[87]), .B(x[87]), .Z(n2336) );
  NANDN U2809 ( .A(y[88]), .B(x[88]), .Z(n2346) );
  NAND U2810 ( .A(n2336), .B(n2346), .Z(n5581) );
  NANDN U2811 ( .A(x[86]), .B(y[86]), .Z(n382) );
  ANDN U2812 ( .B(y[87]), .A(x[87]), .Z(n2342) );
  ANDN U2813 ( .B(n382), .A(n2342), .Z(n5579) );
  XOR U2814 ( .A(x[86]), .B(y[86]), .Z(n2332) );
  NANDN U2815 ( .A(y[85]), .B(x[85]), .Z(n2020) );
  NANDN U2816 ( .A(n2332), .B(n2020), .Z(n5577) );
  ANDN U2817 ( .B(y[84]), .A(x[84]), .Z(n2326) );
  ANDN U2818 ( .B(y[85]), .A(x[85]), .Z(n2334) );
  NOR U2819 ( .A(n2326), .B(n2334), .Z(n5575) );
  NANDN U2820 ( .A(y[83]), .B(x[83]), .Z(n2322) );
  NANDN U2821 ( .A(y[84]), .B(x[84]), .Z(n2019) );
  NAND U2822 ( .A(n2322), .B(n2019), .Z(n5573) );
  ANDN U2823 ( .B(y[82]), .A(x[82]), .Z(n2317) );
  ANDN U2824 ( .B(y[83]), .A(x[83]), .Z(n2327) );
  NOR U2825 ( .A(n2317), .B(n2327), .Z(n5571) );
  NANDN U2826 ( .A(y[81]), .B(x[81]), .Z(n2314) );
  NANDN U2827 ( .A(y[82]), .B(x[82]), .Z(n2321) );
  NAND U2828 ( .A(n2314), .B(n2321), .Z(n5569) );
  NANDN U2829 ( .A(x[80]), .B(y[80]), .Z(n383) );
  ANDN U2830 ( .B(y[81]), .A(x[81]), .Z(n2320) );
  ANDN U2831 ( .B(n383), .A(n2320), .Z(n5567) );
  XOR U2832 ( .A(x[80]), .B(y[80]), .Z(n2310) );
  NANDN U2833 ( .A(y[79]), .B(x[79]), .Z(n2022) );
  NANDN U2834 ( .A(n2310), .B(n2022), .Z(n5565) );
  ANDN U2835 ( .B(y[78]), .A(x[78]), .Z(n2304) );
  ANDN U2836 ( .B(y[79]), .A(x[79]), .Z(n2312) );
  NOR U2837 ( .A(n2304), .B(n2312), .Z(n5563) );
  NANDN U2838 ( .A(y[77]), .B(x[77]), .Z(n2300) );
  NANDN U2839 ( .A(y[78]), .B(x[78]), .Z(n2021) );
  NAND U2840 ( .A(n2300), .B(n2021), .Z(n5561) );
  ANDN U2841 ( .B(y[76]), .A(x[76]), .Z(n2295) );
  ANDN U2842 ( .B(y[77]), .A(x[77]), .Z(n2305) );
  NOR U2843 ( .A(n2295), .B(n2305), .Z(n5559) );
  NANDN U2844 ( .A(y[75]), .B(x[75]), .Z(n2292) );
  NANDN U2845 ( .A(y[76]), .B(x[76]), .Z(n2299) );
  NAND U2846 ( .A(n2292), .B(n2299), .Z(n5557) );
  ANDN U2847 ( .B(y[74]), .A(x[74]), .Z(n2290) );
  ANDN U2848 ( .B(y[75]), .A(x[75]), .Z(n2298) );
  NOR U2849 ( .A(n2290), .B(n2298), .Z(n5555) );
  NANDN U2850 ( .A(y[73]), .B(x[73]), .Z(n2024) );
  NANDN U2851 ( .A(y[74]), .B(x[74]), .Z(n2293) );
  NAND U2852 ( .A(n2024), .B(n2293), .Z(n5553) );
  ANDN U2853 ( .B(y[72]), .A(x[72]), .Z(n2282) );
  ANDN U2854 ( .B(y[73]), .A(x[73]), .Z(n2287) );
  NOR U2855 ( .A(n2282), .B(n2287), .Z(n5551) );
  NANDN U2856 ( .A(y[71]), .B(x[71]), .Z(n2278) );
  NANDN U2857 ( .A(y[72]), .B(x[72]), .Z(n2023) );
  NAND U2858 ( .A(n2278), .B(n2023), .Z(n5549) );
  ANDN U2859 ( .B(y[70]), .A(x[70]), .Z(n2273) );
  ANDN U2860 ( .B(y[71]), .A(x[71]), .Z(n2283) );
  NOR U2861 ( .A(n2273), .B(n2283), .Z(n5547) );
  NANDN U2862 ( .A(y[69]), .B(x[69]), .Z(n2270) );
  NANDN U2863 ( .A(y[70]), .B(x[70]), .Z(n2277) );
  NAND U2864 ( .A(n2270), .B(n2277), .Z(n5545) );
  ANDN U2865 ( .B(y[68]), .A(x[68]), .Z(n2268) );
  ANDN U2866 ( .B(y[69]), .A(x[69]), .Z(n2276) );
  NOR U2867 ( .A(n2268), .B(n2276), .Z(n5543) );
  NANDN U2868 ( .A(y[67]), .B(x[67]), .Z(n2026) );
  NANDN U2869 ( .A(y[68]), .B(x[68]), .Z(n2271) );
  NAND U2870 ( .A(n2026), .B(n2271), .Z(n5541) );
  ANDN U2871 ( .B(y[66]), .A(x[66]), .Z(n2260) );
  ANDN U2872 ( .B(y[67]), .A(x[67]), .Z(n2265) );
  NOR U2873 ( .A(n2260), .B(n2265), .Z(n5539) );
  NANDN U2874 ( .A(y[65]), .B(x[65]), .Z(n2256) );
  NANDN U2875 ( .A(y[66]), .B(x[66]), .Z(n2025) );
  NAND U2876 ( .A(n2256), .B(n2025), .Z(n5537) );
  ANDN U2877 ( .B(y[64]), .A(x[64]), .Z(n2251) );
  ANDN U2878 ( .B(y[65]), .A(x[65]), .Z(n2261) );
  NOR U2879 ( .A(n2251), .B(n2261), .Z(n5535) );
  NANDN U2880 ( .A(y[63]), .B(x[63]), .Z(n2248) );
  NANDN U2881 ( .A(y[64]), .B(x[64]), .Z(n2255) );
  NAND U2882 ( .A(n2248), .B(n2255), .Z(n5533) );
  ANDN U2883 ( .B(y[62]), .A(x[62]), .Z(n2246) );
  ANDN U2884 ( .B(y[63]), .A(x[63]), .Z(n2254) );
  NOR U2885 ( .A(n2246), .B(n2254), .Z(n5531) );
  NANDN U2886 ( .A(y[61]), .B(x[61]), .Z(n2028) );
  NANDN U2887 ( .A(y[62]), .B(x[62]), .Z(n2249) );
  NAND U2888 ( .A(n2028), .B(n2249), .Z(n5529) );
  ANDN U2889 ( .B(y[60]), .A(x[60]), .Z(n2238) );
  ANDN U2890 ( .B(y[61]), .A(x[61]), .Z(n2243) );
  NOR U2891 ( .A(n2238), .B(n2243), .Z(n5527) );
  NANDN U2892 ( .A(y[59]), .B(x[59]), .Z(n2234) );
  NANDN U2893 ( .A(y[60]), .B(x[60]), .Z(n2027) );
  NAND U2894 ( .A(n2234), .B(n2027), .Z(n5525) );
  ANDN U2895 ( .B(y[58]), .A(x[58]), .Z(n2229) );
  ANDN U2896 ( .B(y[59]), .A(x[59]), .Z(n2239) );
  NOR U2897 ( .A(n2229), .B(n2239), .Z(n5523) );
  NANDN U2898 ( .A(y[57]), .B(x[57]), .Z(n2226) );
  NANDN U2899 ( .A(y[58]), .B(x[58]), .Z(n2233) );
  NAND U2900 ( .A(n2226), .B(n2233), .Z(n5521) );
  ANDN U2901 ( .B(y[56]), .A(x[56]), .Z(n2224) );
  ANDN U2902 ( .B(y[57]), .A(x[57]), .Z(n2232) );
  NOR U2903 ( .A(n2224), .B(n2232), .Z(n5519) );
  NANDN U2904 ( .A(y[55]), .B(x[55]), .Z(n2030) );
  NANDN U2905 ( .A(y[56]), .B(x[56]), .Z(n2227) );
  NAND U2906 ( .A(n2030), .B(n2227), .Z(n5517) );
  ANDN U2907 ( .B(y[54]), .A(x[54]), .Z(n2216) );
  ANDN U2908 ( .B(y[55]), .A(x[55]), .Z(n2221) );
  NOR U2909 ( .A(n2216), .B(n2221), .Z(n5515) );
  NANDN U2910 ( .A(y[53]), .B(x[53]), .Z(n2212) );
  NANDN U2911 ( .A(y[54]), .B(x[54]), .Z(n2029) );
  NAND U2912 ( .A(n2212), .B(n2029), .Z(n5513) );
  ANDN U2913 ( .B(y[52]), .A(x[52]), .Z(n2207) );
  ANDN U2914 ( .B(y[53]), .A(x[53]), .Z(n2217) );
  NOR U2915 ( .A(n2207), .B(n2217), .Z(n5511) );
  NANDN U2916 ( .A(y[51]), .B(x[51]), .Z(n2204) );
  NANDN U2917 ( .A(y[52]), .B(x[52]), .Z(n2211) );
  NAND U2918 ( .A(n2204), .B(n2211), .Z(n5509) );
  ANDN U2919 ( .B(y[50]), .A(x[50]), .Z(n2202) );
  ANDN U2920 ( .B(y[51]), .A(x[51]), .Z(n2210) );
  NOR U2921 ( .A(n2202), .B(n2210), .Z(n5507) );
  NANDN U2922 ( .A(y[49]), .B(x[49]), .Z(n2032) );
  NANDN U2923 ( .A(y[50]), .B(x[50]), .Z(n2205) );
  NAND U2924 ( .A(n2032), .B(n2205), .Z(n5505) );
  ANDN U2925 ( .B(y[48]), .A(x[48]), .Z(n2194) );
  ANDN U2926 ( .B(y[49]), .A(x[49]), .Z(n2199) );
  NOR U2927 ( .A(n2194), .B(n2199), .Z(n5503) );
  NANDN U2928 ( .A(y[47]), .B(x[47]), .Z(n2190) );
  NANDN U2929 ( .A(y[48]), .B(x[48]), .Z(n2031) );
  NAND U2930 ( .A(n2190), .B(n2031), .Z(n5501) );
  ANDN U2931 ( .B(y[46]), .A(x[46]), .Z(n2185) );
  ANDN U2932 ( .B(y[47]), .A(x[47]), .Z(n2195) );
  NOR U2933 ( .A(n2185), .B(n2195), .Z(n5499) );
  NANDN U2934 ( .A(y[45]), .B(x[45]), .Z(n2182) );
  NANDN U2935 ( .A(y[46]), .B(x[46]), .Z(n2189) );
  NAND U2936 ( .A(n2182), .B(n2189), .Z(n5497) );
  ANDN U2937 ( .B(y[44]), .A(x[44]), .Z(n2180) );
  ANDN U2938 ( .B(y[45]), .A(x[45]), .Z(n2188) );
  NOR U2939 ( .A(n2180), .B(n2188), .Z(n5495) );
  NANDN U2940 ( .A(y[43]), .B(x[43]), .Z(n2034) );
  NANDN U2941 ( .A(y[44]), .B(x[44]), .Z(n2183) );
  NAND U2942 ( .A(n2034), .B(n2183), .Z(n5493) );
  ANDN U2943 ( .B(y[42]), .A(x[42]), .Z(n2172) );
  ANDN U2944 ( .B(y[43]), .A(x[43]), .Z(n2177) );
  NOR U2945 ( .A(n2172), .B(n2177), .Z(n5491) );
  NANDN U2946 ( .A(y[41]), .B(x[41]), .Z(n2168) );
  NANDN U2947 ( .A(y[42]), .B(x[42]), .Z(n2033) );
  NAND U2948 ( .A(n2168), .B(n2033), .Z(n5489) );
  ANDN U2949 ( .B(y[40]), .A(x[40]), .Z(n2163) );
  ANDN U2950 ( .B(y[41]), .A(x[41]), .Z(n2173) );
  NOR U2951 ( .A(n2163), .B(n2173), .Z(n5487) );
  NANDN U2952 ( .A(y[39]), .B(x[39]), .Z(n2160) );
  NANDN U2953 ( .A(y[40]), .B(x[40]), .Z(n2167) );
  NAND U2954 ( .A(n2160), .B(n2167), .Z(n5485) );
  ANDN U2955 ( .B(y[38]), .A(x[38]), .Z(n2158) );
  ANDN U2956 ( .B(y[39]), .A(x[39]), .Z(n2166) );
  NOR U2957 ( .A(n2158), .B(n2166), .Z(n5483) );
  NANDN U2958 ( .A(y[37]), .B(x[37]), .Z(n2036) );
  NANDN U2959 ( .A(y[38]), .B(x[38]), .Z(n2161) );
  NAND U2960 ( .A(n2036), .B(n2161), .Z(n5481) );
  ANDN U2961 ( .B(y[36]), .A(x[36]), .Z(n2150) );
  ANDN U2962 ( .B(y[37]), .A(x[37]), .Z(n2155) );
  NOR U2963 ( .A(n2150), .B(n2155), .Z(n5479) );
  NANDN U2964 ( .A(y[35]), .B(x[35]), .Z(n2146) );
  NANDN U2965 ( .A(y[36]), .B(x[36]), .Z(n2035) );
  NAND U2966 ( .A(n2146), .B(n2035), .Z(n5477) );
  ANDN U2967 ( .B(y[34]), .A(x[34]), .Z(n2141) );
  ANDN U2968 ( .B(y[35]), .A(x[35]), .Z(n2151) );
  NOR U2969 ( .A(n2141), .B(n2151), .Z(n5475) );
  NANDN U2970 ( .A(y[33]), .B(x[33]), .Z(n2138) );
  NANDN U2971 ( .A(y[34]), .B(x[34]), .Z(n2145) );
  NAND U2972 ( .A(n2138), .B(n2145), .Z(n5473) );
  ANDN U2973 ( .B(y[32]), .A(x[32]), .Z(n2136) );
  ANDN U2974 ( .B(y[33]), .A(x[33]), .Z(n2144) );
  NOR U2975 ( .A(n2136), .B(n2144), .Z(n5471) );
  NANDN U2976 ( .A(y[31]), .B(x[31]), .Z(n2038) );
  NANDN U2977 ( .A(y[32]), .B(x[32]), .Z(n2139) );
  NAND U2978 ( .A(n2038), .B(n2139), .Z(n5469) );
  ANDN U2979 ( .B(y[30]), .A(x[30]), .Z(n2128) );
  ANDN U2980 ( .B(y[31]), .A(x[31]), .Z(n2133) );
  NOR U2981 ( .A(n2128), .B(n2133), .Z(n5467) );
  NANDN U2982 ( .A(y[29]), .B(x[29]), .Z(n2124) );
  NANDN U2983 ( .A(y[30]), .B(x[30]), .Z(n2037) );
  NAND U2984 ( .A(n2124), .B(n2037), .Z(n5465) );
  ANDN U2985 ( .B(y[28]), .A(x[28]), .Z(n2119) );
  ANDN U2986 ( .B(y[29]), .A(x[29]), .Z(n2129) );
  NOR U2987 ( .A(n2119), .B(n2129), .Z(n5463) );
  NANDN U2988 ( .A(y[27]), .B(x[27]), .Z(n2116) );
  NANDN U2989 ( .A(y[28]), .B(x[28]), .Z(n2123) );
  NAND U2990 ( .A(n2116), .B(n2123), .Z(n5461) );
  ANDN U2991 ( .B(y[26]), .A(x[26]), .Z(n2114) );
  ANDN U2992 ( .B(y[27]), .A(x[27]), .Z(n2122) );
  NOR U2993 ( .A(n2114), .B(n2122), .Z(n5459) );
  NANDN U2994 ( .A(y[25]), .B(x[25]), .Z(n2040) );
  NANDN U2995 ( .A(y[26]), .B(x[26]), .Z(n2117) );
  NAND U2996 ( .A(n2040), .B(n2117), .Z(n5457) );
  ANDN U2997 ( .B(y[24]), .A(x[24]), .Z(n2106) );
  ANDN U2998 ( .B(y[25]), .A(x[25]), .Z(n2111) );
  NOR U2999 ( .A(n2106), .B(n2111), .Z(n5455) );
  NANDN U3000 ( .A(y[23]), .B(x[23]), .Z(n2102) );
  NANDN U3001 ( .A(y[24]), .B(x[24]), .Z(n2039) );
  NAND U3002 ( .A(n2102), .B(n2039), .Z(n5453) );
  ANDN U3003 ( .B(y[22]), .A(x[22]), .Z(n2097) );
  ANDN U3004 ( .B(y[23]), .A(x[23]), .Z(n2107) );
  NOR U3005 ( .A(n2097), .B(n2107), .Z(n5451) );
  NANDN U3006 ( .A(y[21]), .B(x[21]), .Z(n2094) );
  NANDN U3007 ( .A(y[22]), .B(x[22]), .Z(n2101) );
  NAND U3008 ( .A(n2094), .B(n2101), .Z(n5449) );
  ANDN U3009 ( .B(y[20]), .A(x[20]), .Z(n2092) );
  ANDN U3010 ( .B(y[21]), .A(x[21]), .Z(n2100) );
  NOR U3011 ( .A(n2092), .B(n2100), .Z(n5447) );
  NANDN U3012 ( .A(y[19]), .B(x[19]), .Z(n2042) );
  NANDN U3013 ( .A(y[20]), .B(x[20]), .Z(n2095) );
  NAND U3014 ( .A(n2042), .B(n2095), .Z(n5445) );
  ANDN U3015 ( .B(y[18]), .A(x[18]), .Z(n2084) );
  ANDN U3016 ( .B(y[19]), .A(x[19]), .Z(n2089) );
  NOR U3017 ( .A(n2084), .B(n2089), .Z(n5443) );
  NANDN U3018 ( .A(y[17]), .B(x[17]), .Z(n2080) );
  NANDN U3019 ( .A(y[18]), .B(x[18]), .Z(n2041) );
  NAND U3020 ( .A(n2080), .B(n2041), .Z(n5441) );
  ANDN U3021 ( .B(y[16]), .A(x[16]), .Z(n2075) );
  ANDN U3022 ( .B(y[17]), .A(x[17]), .Z(n2085) );
  NOR U3023 ( .A(n2075), .B(n2085), .Z(n5439) );
  NANDN U3024 ( .A(y[15]), .B(x[15]), .Z(n2072) );
  NANDN U3025 ( .A(y[16]), .B(x[16]), .Z(n2079) );
  NAND U3026 ( .A(n2072), .B(n2079), .Z(n5437) );
  ANDN U3027 ( .B(y[14]), .A(x[14]), .Z(n2070) );
  ANDN U3028 ( .B(y[15]), .A(x[15]), .Z(n2078) );
  NOR U3029 ( .A(n2070), .B(n2078), .Z(n5435) );
  NANDN U3030 ( .A(y[13]), .B(x[13]), .Z(n2044) );
  NANDN U3031 ( .A(y[14]), .B(x[14]), .Z(n2073) );
  NAND U3032 ( .A(n2044), .B(n2073), .Z(n5433) );
  ANDN U3033 ( .B(y[12]), .A(x[12]), .Z(n2062) );
  ANDN U3034 ( .B(y[13]), .A(x[13]), .Z(n2067) );
  NOR U3035 ( .A(n2062), .B(n2067), .Z(n5431) );
  NANDN U3036 ( .A(y[11]), .B(x[11]), .Z(n2060) );
  NANDN U3037 ( .A(y[12]), .B(x[12]), .Z(n2043) );
  NAND U3038 ( .A(n2060), .B(n2043), .Z(n5429) );
  ANDN U3039 ( .B(y[10]), .A(x[10]), .Z(n2058) );
  ANDN U3040 ( .B(y[11]), .A(x[11]), .Z(n2063) );
  NOR U3041 ( .A(n2058), .B(n2063), .Z(n5426) );
  NANDN U3042 ( .A(y[9]), .B(x[9]), .Z(n385) );
  NANDN U3043 ( .A(y[10]), .B(x[10]), .Z(n384) );
  NAND U3044 ( .A(n385), .B(n384), .Z(n2057) );
  NANDN U3045 ( .A(x[9]), .B(y[9]), .Z(n387) );
  NANDN U3046 ( .A(x[8]), .B(y[8]), .Z(n386) );
  AND U3047 ( .A(n387), .B(n386), .Z(n2045) );
  NANDN U3048 ( .A(y[7]), .B(x[7]), .Z(n389) );
  NANDN U3049 ( .A(y[8]), .B(x[8]), .Z(n388) );
  NAND U3050 ( .A(n389), .B(n388), .Z(n2046) );
  NANDN U3051 ( .A(x[7]), .B(y[7]), .Z(n391) );
  NANDN U3052 ( .A(x[6]), .B(y[6]), .Z(n390) );
  AND U3053 ( .A(n391), .B(n390), .Z(n2047) );
  NANDN U3054 ( .A(y[3]), .B(x[3]), .Z(n393) );
  NANDN U3055 ( .A(y[4]), .B(x[4]), .Z(n392) );
  NAND U3056 ( .A(n393), .B(n392), .Z(n2055) );
  NANDN U3057 ( .A(x[3]), .B(y[3]), .Z(n2049) );
  NANDN U3058 ( .A(x[2]), .B(y[2]), .Z(n2051) );
  NANDN U3059 ( .A(y[2]), .B(x[2]), .Z(n2054) );
  NANDN U3060 ( .A(y[1]), .B(x[1]), .Z(n2053) );
  NAND U3061 ( .A(n2054), .B(n2053), .Z(n396) );
  NANDN U3062 ( .A(x[0]), .B(y[0]), .Z(n394) );
  NANDN U3063 ( .A(x[1]), .B(y[1]), .Z(n2050) );
  NAND U3064 ( .A(n394), .B(n2050), .Z(n395) );
  NANDN U3065 ( .A(n396), .B(n395), .Z(n397) );
  AND U3066 ( .A(n2051), .B(n397), .Z(n398) );
  NAND U3067 ( .A(n2049), .B(n398), .Z(n399) );
  NANDN U3068 ( .A(n2055), .B(n399), .Z(n402) );
  NANDN U3069 ( .A(x[5]), .B(y[5]), .Z(n401) );
  NANDN U3070 ( .A(x[4]), .B(y[4]), .Z(n400) );
  AND U3071 ( .A(n401), .B(n400), .Z(n2056) );
  AND U3072 ( .A(n402), .B(n2056), .Z(n405) );
  NANDN U3073 ( .A(y[5]), .B(x[5]), .Z(n404) );
  NANDN U3074 ( .A(y[6]), .B(x[6]), .Z(n403) );
  NAND U3075 ( .A(n404), .B(n403), .Z(n2048) );
  OR U3076 ( .A(n405), .B(n2048), .Z(n406) );
  NAND U3077 ( .A(n2047), .B(n406), .Z(n407) );
  NANDN U3078 ( .A(n2046), .B(n407), .Z(n408) );
  NAND U3079 ( .A(n2045), .B(n408), .Z(n409) );
  NANDN U3080 ( .A(n2057), .B(n409), .Z(n410) );
  AND U3081 ( .A(n5426), .B(n410), .Z(n411) );
  OR U3082 ( .A(n5429), .B(n411), .Z(n412) );
  NAND U3083 ( .A(n5431), .B(n412), .Z(n413) );
  NANDN U3084 ( .A(n5433), .B(n413), .Z(n414) );
  NAND U3085 ( .A(n5435), .B(n414), .Z(n415) );
  NANDN U3086 ( .A(n5437), .B(n415), .Z(n416) );
  AND U3087 ( .A(n5439), .B(n416), .Z(n417) );
  OR U3088 ( .A(n5441), .B(n417), .Z(n418) );
  NAND U3089 ( .A(n5443), .B(n418), .Z(n419) );
  NANDN U3090 ( .A(n5445), .B(n419), .Z(n420) );
  NAND U3091 ( .A(n5447), .B(n420), .Z(n421) );
  NANDN U3092 ( .A(n5449), .B(n421), .Z(n422) );
  AND U3093 ( .A(n5451), .B(n422), .Z(n423) );
  OR U3094 ( .A(n5453), .B(n423), .Z(n424) );
  NAND U3095 ( .A(n5455), .B(n424), .Z(n425) );
  NANDN U3096 ( .A(n5457), .B(n425), .Z(n426) );
  NAND U3097 ( .A(n5459), .B(n426), .Z(n427) );
  NANDN U3098 ( .A(n5461), .B(n427), .Z(n428) );
  AND U3099 ( .A(n5463), .B(n428), .Z(n429) );
  OR U3100 ( .A(n5465), .B(n429), .Z(n430) );
  NAND U3101 ( .A(n5467), .B(n430), .Z(n431) );
  NANDN U3102 ( .A(n5469), .B(n431), .Z(n432) );
  NAND U3103 ( .A(n5471), .B(n432), .Z(n433) );
  NANDN U3104 ( .A(n5473), .B(n433), .Z(n434) );
  AND U3105 ( .A(n5475), .B(n434), .Z(n435) );
  OR U3106 ( .A(n5477), .B(n435), .Z(n436) );
  NAND U3107 ( .A(n5479), .B(n436), .Z(n437) );
  NANDN U3108 ( .A(n5481), .B(n437), .Z(n438) );
  NAND U3109 ( .A(n5483), .B(n438), .Z(n439) );
  NANDN U3110 ( .A(n5485), .B(n439), .Z(n440) );
  AND U3111 ( .A(n5487), .B(n440), .Z(n441) );
  OR U3112 ( .A(n5489), .B(n441), .Z(n442) );
  NAND U3113 ( .A(n5491), .B(n442), .Z(n443) );
  NANDN U3114 ( .A(n5493), .B(n443), .Z(n444) );
  NAND U3115 ( .A(n5495), .B(n444), .Z(n445) );
  NANDN U3116 ( .A(n5497), .B(n445), .Z(n446) );
  AND U3117 ( .A(n5499), .B(n446), .Z(n447) );
  OR U3118 ( .A(n5501), .B(n447), .Z(n448) );
  NAND U3119 ( .A(n5503), .B(n448), .Z(n449) );
  NANDN U3120 ( .A(n5505), .B(n449), .Z(n450) );
  NAND U3121 ( .A(n5507), .B(n450), .Z(n451) );
  NANDN U3122 ( .A(n5509), .B(n451), .Z(n452) );
  AND U3123 ( .A(n5511), .B(n452), .Z(n453) );
  OR U3124 ( .A(n5513), .B(n453), .Z(n454) );
  NAND U3125 ( .A(n5515), .B(n454), .Z(n455) );
  NANDN U3126 ( .A(n5517), .B(n455), .Z(n456) );
  NAND U3127 ( .A(n5519), .B(n456), .Z(n457) );
  NANDN U3128 ( .A(n5521), .B(n457), .Z(n458) );
  AND U3129 ( .A(n5523), .B(n458), .Z(n459) );
  OR U3130 ( .A(n5525), .B(n459), .Z(n460) );
  NAND U3131 ( .A(n5527), .B(n460), .Z(n461) );
  NANDN U3132 ( .A(n5529), .B(n461), .Z(n462) );
  NAND U3133 ( .A(n5531), .B(n462), .Z(n463) );
  NANDN U3134 ( .A(n5533), .B(n463), .Z(n464) );
  AND U3135 ( .A(n5535), .B(n464), .Z(n465) );
  OR U3136 ( .A(n5537), .B(n465), .Z(n466) );
  NAND U3137 ( .A(n5539), .B(n466), .Z(n467) );
  NANDN U3138 ( .A(n5541), .B(n467), .Z(n468) );
  NAND U3139 ( .A(n5543), .B(n468), .Z(n469) );
  NANDN U3140 ( .A(n5545), .B(n469), .Z(n470) );
  AND U3141 ( .A(n5547), .B(n470), .Z(n471) );
  OR U3142 ( .A(n5549), .B(n471), .Z(n472) );
  NAND U3143 ( .A(n5551), .B(n472), .Z(n473) );
  NANDN U3144 ( .A(n5553), .B(n473), .Z(n474) );
  NAND U3145 ( .A(n5555), .B(n474), .Z(n475) );
  NANDN U3146 ( .A(n5557), .B(n475), .Z(n476) );
  AND U3147 ( .A(n5559), .B(n476), .Z(n477) );
  OR U3148 ( .A(n5561), .B(n477), .Z(n478) );
  NAND U3149 ( .A(n5563), .B(n478), .Z(n479) );
  NANDN U3150 ( .A(n5565), .B(n479), .Z(n480) );
  NAND U3151 ( .A(n5567), .B(n480), .Z(n481) );
  NANDN U3152 ( .A(n5569), .B(n481), .Z(n482) );
  AND U3153 ( .A(n5571), .B(n482), .Z(n483) );
  OR U3154 ( .A(n5573), .B(n483), .Z(n484) );
  NAND U3155 ( .A(n5575), .B(n484), .Z(n485) );
  NANDN U3156 ( .A(n5577), .B(n485), .Z(n486) );
  NAND U3157 ( .A(n5579), .B(n486), .Z(n487) );
  NANDN U3158 ( .A(n5581), .B(n487), .Z(n488) );
  AND U3159 ( .A(n5583), .B(n488), .Z(n489) );
  OR U3160 ( .A(n5585), .B(n489), .Z(n490) );
  NAND U3161 ( .A(n5587), .B(n490), .Z(n491) );
  NANDN U3162 ( .A(n5589), .B(n491), .Z(n492) );
  NAND U3163 ( .A(n5591), .B(n492), .Z(n493) );
  NANDN U3164 ( .A(n5593), .B(n493), .Z(n494) );
  AND U3165 ( .A(n5595), .B(n494), .Z(n495) );
  OR U3166 ( .A(n5597), .B(n495), .Z(n496) );
  NAND U3167 ( .A(n5599), .B(n496), .Z(n497) );
  NANDN U3168 ( .A(n5601), .B(n497), .Z(n498) );
  NAND U3169 ( .A(n5603), .B(n498), .Z(n499) );
  NANDN U3170 ( .A(n5605), .B(n499), .Z(n500) );
  AND U3171 ( .A(n5607), .B(n500), .Z(n501) );
  OR U3172 ( .A(n5609), .B(n501), .Z(n502) );
  NAND U3173 ( .A(n5611), .B(n502), .Z(n503) );
  NANDN U3174 ( .A(n5613), .B(n503), .Z(n504) );
  NAND U3175 ( .A(n5615), .B(n504), .Z(n505) );
  NANDN U3176 ( .A(n5617), .B(n505), .Z(n506) );
  AND U3177 ( .A(n5619), .B(n506), .Z(n507) );
  OR U3178 ( .A(n5621), .B(n507), .Z(n508) );
  NAND U3179 ( .A(n5623), .B(n508), .Z(n509) );
  NANDN U3180 ( .A(n5625), .B(n509), .Z(n510) );
  NAND U3181 ( .A(n5627), .B(n510), .Z(n511) );
  NANDN U3182 ( .A(n5629), .B(n511), .Z(n512) );
  AND U3183 ( .A(n5631), .B(n512), .Z(n513) );
  OR U3184 ( .A(n5633), .B(n513), .Z(n514) );
  NAND U3185 ( .A(n5635), .B(n514), .Z(n515) );
  NANDN U3186 ( .A(n5637), .B(n515), .Z(n516) );
  NAND U3187 ( .A(n5639), .B(n516), .Z(n517) );
  NANDN U3188 ( .A(n5641), .B(n517), .Z(n518) );
  AND U3189 ( .A(n5643), .B(n518), .Z(n519) );
  OR U3190 ( .A(n5645), .B(n519), .Z(n520) );
  NAND U3191 ( .A(n5647), .B(n520), .Z(n521) );
  NANDN U3192 ( .A(n5649), .B(n521), .Z(n522) );
  NAND U3193 ( .A(n5651), .B(n522), .Z(n523) );
  NANDN U3194 ( .A(n5653), .B(n523), .Z(n524) );
  AND U3195 ( .A(n5655), .B(n524), .Z(n525) );
  OR U3196 ( .A(n5657), .B(n525), .Z(n526) );
  NAND U3197 ( .A(n5659), .B(n526), .Z(n527) );
  NANDN U3198 ( .A(n5661), .B(n527), .Z(n528) );
  NAND U3199 ( .A(n5663), .B(n528), .Z(n529) );
  NANDN U3200 ( .A(n5665), .B(n529), .Z(n530) );
  AND U3201 ( .A(n5667), .B(n530), .Z(n531) );
  OR U3202 ( .A(n5669), .B(n531), .Z(n532) );
  NAND U3203 ( .A(n5671), .B(n532), .Z(n533) );
  NANDN U3204 ( .A(n5673), .B(n533), .Z(n534) );
  NAND U3205 ( .A(n5675), .B(n534), .Z(n535) );
  NANDN U3206 ( .A(n5677), .B(n535), .Z(n536) );
  AND U3207 ( .A(n5679), .B(n536), .Z(n537) );
  OR U3208 ( .A(n5681), .B(n537), .Z(n538) );
  NAND U3209 ( .A(n5683), .B(n538), .Z(n539) );
  NANDN U3210 ( .A(n5685), .B(n539), .Z(n540) );
  NAND U3211 ( .A(n5687), .B(n540), .Z(n541) );
  NANDN U3212 ( .A(n5689), .B(n541), .Z(n542) );
  AND U3213 ( .A(n5691), .B(n542), .Z(n543) );
  OR U3214 ( .A(n5693), .B(n543), .Z(n544) );
  NAND U3215 ( .A(n5695), .B(n544), .Z(n545) );
  NANDN U3216 ( .A(n5697), .B(n545), .Z(n546) );
  NAND U3217 ( .A(n5699), .B(n546), .Z(n547) );
  NANDN U3218 ( .A(n5701), .B(n547), .Z(n548) );
  AND U3219 ( .A(n5703), .B(n548), .Z(n549) );
  OR U3220 ( .A(n5705), .B(n549), .Z(n550) );
  NAND U3221 ( .A(n5707), .B(n550), .Z(n551) );
  NANDN U3222 ( .A(n5709), .B(n551), .Z(n552) );
  NAND U3223 ( .A(n5711), .B(n552), .Z(n553) );
  NANDN U3224 ( .A(n5713), .B(n553), .Z(n554) );
  AND U3225 ( .A(n5715), .B(n554), .Z(n555) );
  OR U3226 ( .A(n5717), .B(n555), .Z(n556) );
  NAND U3227 ( .A(n5719), .B(n556), .Z(n557) );
  NANDN U3228 ( .A(n5721), .B(n557), .Z(n558) );
  NAND U3229 ( .A(n5723), .B(n558), .Z(n559) );
  NANDN U3230 ( .A(n5725), .B(n559), .Z(n560) );
  AND U3231 ( .A(n5727), .B(n560), .Z(n561) );
  OR U3232 ( .A(n5729), .B(n561), .Z(n562) );
  NAND U3233 ( .A(n5731), .B(n562), .Z(n563) );
  NANDN U3234 ( .A(n5733), .B(n563), .Z(n564) );
  NAND U3235 ( .A(n5735), .B(n564), .Z(n565) );
  NANDN U3236 ( .A(n5737), .B(n565), .Z(n566) );
  AND U3237 ( .A(n5739), .B(n566), .Z(n567) );
  OR U3238 ( .A(n5741), .B(n567), .Z(n568) );
  NAND U3239 ( .A(n5743), .B(n568), .Z(n569) );
  NANDN U3240 ( .A(n5745), .B(n569), .Z(n570) );
  NAND U3241 ( .A(n5747), .B(n570), .Z(n571) );
  NANDN U3242 ( .A(n5749), .B(n571), .Z(n572) );
  AND U3243 ( .A(n5751), .B(n572), .Z(n573) );
  OR U3244 ( .A(n5753), .B(n573), .Z(n574) );
  NAND U3245 ( .A(n5755), .B(n574), .Z(n575) );
  NANDN U3246 ( .A(n5757), .B(n575), .Z(n576) );
  NAND U3247 ( .A(n5759), .B(n576), .Z(n577) );
  NANDN U3248 ( .A(n5761), .B(n577), .Z(n578) );
  AND U3249 ( .A(n5763), .B(n578), .Z(n579) );
  OR U3250 ( .A(n5765), .B(n579), .Z(n580) );
  NAND U3251 ( .A(n5767), .B(n580), .Z(n581) );
  NANDN U3252 ( .A(n5769), .B(n581), .Z(n582) );
  NAND U3253 ( .A(n5771), .B(n582), .Z(n583) );
  NANDN U3254 ( .A(n5773), .B(n583), .Z(n584) );
  AND U3255 ( .A(n5775), .B(n584), .Z(n585) );
  OR U3256 ( .A(n5777), .B(n585), .Z(n586) );
  NAND U3257 ( .A(n5779), .B(n586), .Z(n587) );
  NANDN U3258 ( .A(n5781), .B(n587), .Z(n588) );
  NAND U3259 ( .A(n5783), .B(n588), .Z(n589) );
  NANDN U3260 ( .A(n5785), .B(n589), .Z(n590) );
  AND U3261 ( .A(n5787), .B(n590), .Z(n591) );
  OR U3262 ( .A(n5789), .B(n591), .Z(n592) );
  NAND U3263 ( .A(n5791), .B(n592), .Z(n593) );
  NANDN U3264 ( .A(n5793), .B(n593), .Z(n594) );
  NAND U3265 ( .A(n5795), .B(n594), .Z(n595) );
  NANDN U3266 ( .A(n5797), .B(n595), .Z(n596) );
  AND U3267 ( .A(n5799), .B(n596), .Z(n597) );
  OR U3268 ( .A(n5801), .B(n597), .Z(n598) );
  NAND U3269 ( .A(n5803), .B(n598), .Z(n599) );
  NANDN U3270 ( .A(n5805), .B(n599), .Z(n600) );
  NAND U3271 ( .A(n5807), .B(n600), .Z(n601) );
  NANDN U3272 ( .A(n5809), .B(n601), .Z(n602) );
  AND U3273 ( .A(n5811), .B(n602), .Z(n603) );
  OR U3274 ( .A(n5813), .B(n603), .Z(n604) );
  NAND U3275 ( .A(n5815), .B(n604), .Z(n605) );
  NANDN U3276 ( .A(n5817), .B(n605), .Z(n606) );
  NAND U3277 ( .A(n5819), .B(n606), .Z(n607) );
  NANDN U3278 ( .A(n5821), .B(n607), .Z(n608) );
  AND U3279 ( .A(n5823), .B(n608), .Z(n609) );
  OR U3280 ( .A(n5825), .B(n609), .Z(n610) );
  NAND U3281 ( .A(n5827), .B(n610), .Z(n611) );
  NANDN U3282 ( .A(n5829), .B(n611), .Z(n612) );
  NAND U3283 ( .A(n5831), .B(n612), .Z(n613) );
  NANDN U3284 ( .A(n5833), .B(n613), .Z(n614) );
  AND U3285 ( .A(n5835), .B(n614), .Z(n615) );
  OR U3286 ( .A(n5837), .B(n615), .Z(n616) );
  NAND U3287 ( .A(n5839), .B(n616), .Z(n617) );
  NANDN U3288 ( .A(n5841), .B(n617), .Z(n618) );
  NAND U3289 ( .A(n5843), .B(n618), .Z(n619) );
  NANDN U3290 ( .A(n5845), .B(n619), .Z(n620) );
  AND U3291 ( .A(n5847), .B(n620), .Z(n621) );
  OR U3292 ( .A(n5849), .B(n621), .Z(n622) );
  NAND U3293 ( .A(n5851), .B(n622), .Z(n623) );
  NANDN U3294 ( .A(n5853), .B(n623), .Z(n624) );
  NAND U3295 ( .A(n5855), .B(n624), .Z(n625) );
  NANDN U3296 ( .A(n5857), .B(n625), .Z(n626) );
  AND U3297 ( .A(n5859), .B(n626), .Z(n627) );
  OR U3298 ( .A(n5861), .B(n627), .Z(n628) );
  NAND U3299 ( .A(n5863), .B(n628), .Z(n629) );
  NANDN U3300 ( .A(n5865), .B(n629), .Z(n630) );
  NAND U3301 ( .A(n5867), .B(n630), .Z(n631) );
  NANDN U3302 ( .A(n5869), .B(n631), .Z(n632) );
  AND U3303 ( .A(n5871), .B(n632), .Z(n633) );
  OR U3304 ( .A(n5873), .B(n633), .Z(n634) );
  NAND U3305 ( .A(n5875), .B(n634), .Z(n635) );
  NANDN U3306 ( .A(n5877), .B(n635), .Z(n636) );
  NAND U3307 ( .A(n5879), .B(n636), .Z(n637) );
  NANDN U3308 ( .A(n5881), .B(n637), .Z(n638) );
  AND U3309 ( .A(n5883), .B(n638), .Z(n639) );
  OR U3310 ( .A(n5885), .B(n639), .Z(n640) );
  NAND U3311 ( .A(n5887), .B(n640), .Z(n641) );
  NANDN U3312 ( .A(n5889), .B(n641), .Z(n642) );
  NAND U3313 ( .A(n5891), .B(n642), .Z(n643) );
  NANDN U3314 ( .A(n5893), .B(n643), .Z(n644) );
  AND U3315 ( .A(n5895), .B(n644), .Z(n645) );
  OR U3316 ( .A(n5897), .B(n645), .Z(n646) );
  NAND U3317 ( .A(n5899), .B(n646), .Z(n647) );
  NANDN U3318 ( .A(n5901), .B(n647), .Z(n648) );
  NAND U3319 ( .A(n5903), .B(n648), .Z(n649) );
  NANDN U3320 ( .A(n5905), .B(n649), .Z(n650) );
  AND U3321 ( .A(n5907), .B(n650), .Z(n651) );
  OR U3322 ( .A(n5909), .B(n651), .Z(n652) );
  NAND U3323 ( .A(n5911), .B(n652), .Z(n653) );
  NANDN U3324 ( .A(n5913), .B(n653), .Z(n654) );
  NAND U3325 ( .A(n5915), .B(n654), .Z(n655) );
  NANDN U3326 ( .A(n5917), .B(n655), .Z(n656) );
  AND U3327 ( .A(n5919), .B(n656), .Z(n657) );
  OR U3328 ( .A(n5921), .B(n657), .Z(n658) );
  NAND U3329 ( .A(n5923), .B(n658), .Z(n659) );
  NANDN U3330 ( .A(n5925), .B(n659), .Z(n660) );
  NAND U3331 ( .A(n5927), .B(n660), .Z(n661) );
  NANDN U3332 ( .A(n5929), .B(n661), .Z(n662) );
  AND U3333 ( .A(n5931), .B(n662), .Z(n663) );
  OR U3334 ( .A(n5933), .B(n663), .Z(n664) );
  NAND U3335 ( .A(n5935), .B(n664), .Z(n665) );
  NANDN U3336 ( .A(n5937), .B(n665), .Z(n666) );
  NAND U3337 ( .A(n5939), .B(n666), .Z(n667) );
  NANDN U3338 ( .A(n5941), .B(n667), .Z(n668) );
  AND U3339 ( .A(n5943), .B(n668), .Z(n669) );
  OR U3340 ( .A(n5945), .B(n669), .Z(n670) );
  NAND U3341 ( .A(n5947), .B(n670), .Z(n671) );
  NANDN U3342 ( .A(n5949), .B(n671), .Z(n672) );
  NAND U3343 ( .A(n5951), .B(n672), .Z(n673) );
  NANDN U3344 ( .A(n5953), .B(n673), .Z(n674) );
  AND U3345 ( .A(n5955), .B(n674), .Z(n675) );
  OR U3346 ( .A(n5957), .B(n675), .Z(n676) );
  NAND U3347 ( .A(n5959), .B(n676), .Z(n677) );
  NANDN U3348 ( .A(n5961), .B(n677), .Z(n678) );
  NAND U3349 ( .A(n5963), .B(n678), .Z(n679) );
  NANDN U3350 ( .A(n5965), .B(n679), .Z(n680) );
  AND U3351 ( .A(n5967), .B(n680), .Z(n681) );
  OR U3352 ( .A(n5969), .B(n681), .Z(n682) );
  NAND U3353 ( .A(n5971), .B(n682), .Z(n683) );
  NANDN U3354 ( .A(n5973), .B(n683), .Z(n684) );
  NAND U3355 ( .A(n5975), .B(n684), .Z(n685) );
  NANDN U3356 ( .A(n5977), .B(n685), .Z(n686) );
  AND U3357 ( .A(n5979), .B(n686), .Z(n687) );
  OR U3358 ( .A(n5981), .B(n687), .Z(n688) );
  NAND U3359 ( .A(n5983), .B(n688), .Z(n689) );
  NANDN U3360 ( .A(n5985), .B(n689), .Z(n690) );
  NAND U3361 ( .A(n5987), .B(n690), .Z(n691) );
  NANDN U3362 ( .A(n5989), .B(n691), .Z(n692) );
  AND U3363 ( .A(n5991), .B(n692), .Z(n693) );
  OR U3364 ( .A(n5993), .B(n693), .Z(n694) );
  NAND U3365 ( .A(n5995), .B(n694), .Z(n695) );
  NANDN U3366 ( .A(n5997), .B(n695), .Z(n696) );
  NAND U3367 ( .A(n5999), .B(n696), .Z(n697) );
  NANDN U3368 ( .A(n6001), .B(n697), .Z(n698) );
  AND U3369 ( .A(n6003), .B(n698), .Z(n701) );
  NANDN U3370 ( .A(y[299]), .B(x[299]), .Z(n700) );
  NANDN U3371 ( .A(y[300]), .B(x[300]), .Z(n699) );
  AND U3372 ( .A(n700), .B(n699), .Z(n6005) );
  NANDN U3373 ( .A(n701), .B(n6005), .Z(n702) );
  NAND U3374 ( .A(n6007), .B(n702), .Z(n703) );
  NANDN U3375 ( .A(n6009), .B(n703), .Z(n704) );
  NAND U3376 ( .A(n6011), .B(n704), .Z(n705) );
  NANDN U3377 ( .A(n6013), .B(n705), .Z(n706) );
  AND U3378 ( .A(n6015), .B(n706), .Z(n707) );
  OR U3379 ( .A(n6017), .B(n707), .Z(n708) );
  NAND U3380 ( .A(n6019), .B(n708), .Z(n709) );
  NANDN U3381 ( .A(n6021), .B(n709), .Z(n710) );
  NAND U3382 ( .A(n6023), .B(n710), .Z(n711) );
  NANDN U3383 ( .A(n6025), .B(n711), .Z(n712) );
  AND U3384 ( .A(n6027), .B(n712), .Z(n713) );
  OR U3385 ( .A(n6029), .B(n713), .Z(n714) );
  NAND U3386 ( .A(n6031), .B(n714), .Z(n715) );
  NANDN U3387 ( .A(n6033), .B(n715), .Z(n716) );
  NAND U3388 ( .A(n6035), .B(n716), .Z(n717) );
  NANDN U3389 ( .A(n6037), .B(n717), .Z(n718) );
  AND U3390 ( .A(n6039), .B(n718), .Z(n719) );
  OR U3391 ( .A(n6041), .B(n719), .Z(n720) );
  NAND U3392 ( .A(n6043), .B(n720), .Z(n721) );
  NANDN U3393 ( .A(n6045), .B(n721), .Z(n722) );
  NAND U3394 ( .A(n6047), .B(n722), .Z(n723) );
  NANDN U3395 ( .A(n6049), .B(n723), .Z(n724) );
  AND U3396 ( .A(n6051), .B(n724), .Z(n725) );
  OR U3397 ( .A(n6053), .B(n725), .Z(n726) );
  NAND U3398 ( .A(n6055), .B(n726), .Z(n727) );
  NANDN U3399 ( .A(n6057), .B(n727), .Z(n728) );
  NAND U3400 ( .A(n6059), .B(n728), .Z(n729) );
  NANDN U3401 ( .A(n6061), .B(n729), .Z(n730) );
  AND U3402 ( .A(n6063), .B(n730), .Z(n731) );
  OR U3403 ( .A(n6065), .B(n731), .Z(n732) );
  NAND U3404 ( .A(n6067), .B(n732), .Z(n733) );
  NANDN U3405 ( .A(n6069), .B(n733), .Z(n734) );
  NAND U3406 ( .A(n6071), .B(n734), .Z(n735) );
  NANDN U3407 ( .A(n6073), .B(n735), .Z(n736) );
  AND U3408 ( .A(n6075), .B(n736), .Z(n737) );
  OR U3409 ( .A(n6077), .B(n737), .Z(n738) );
  NAND U3410 ( .A(n6079), .B(n738), .Z(n739) );
  NANDN U3411 ( .A(n6081), .B(n739), .Z(n740) );
  NAND U3412 ( .A(n6083), .B(n740), .Z(n741) );
  NANDN U3413 ( .A(n6085), .B(n741), .Z(n742) );
  AND U3414 ( .A(n6087), .B(n742), .Z(n743) );
  OR U3415 ( .A(n6089), .B(n743), .Z(n744) );
  NAND U3416 ( .A(n6091), .B(n744), .Z(n745) );
  NANDN U3417 ( .A(n6093), .B(n745), .Z(n746) );
  NAND U3418 ( .A(n6095), .B(n746), .Z(n747) );
  NANDN U3419 ( .A(n6097), .B(n747), .Z(n748) );
  AND U3420 ( .A(n6099), .B(n748), .Z(n749) );
  OR U3421 ( .A(n6101), .B(n749), .Z(n750) );
  NAND U3422 ( .A(n6103), .B(n750), .Z(n751) );
  NANDN U3423 ( .A(n6105), .B(n751), .Z(n752) );
  NAND U3424 ( .A(n6107), .B(n752), .Z(n753) );
  NANDN U3425 ( .A(n6109), .B(n753), .Z(n754) );
  AND U3426 ( .A(n6111), .B(n754), .Z(n755) );
  OR U3427 ( .A(n6113), .B(n755), .Z(n756) );
  NAND U3428 ( .A(n6115), .B(n756), .Z(n757) );
  NANDN U3429 ( .A(n6117), .B(n757), .Z(n758) );
  NAND U3430 ( .A(n6119), .B(n758), .Z(n759) );
  NANDN U3431 ( .A(n6121), .B(n759), .Z(n760) );
  AND U3432 ( .A(n6123), .B(n760), .Z(n761) );
  OR U3433 ( .A(n6125), .B(n761), .Z(n762) );
  NAND U3434 ( .A(n6127), .B(n762), .Z(n763) );
  NANDN U3435 ( .A(n6129), .B(n763), .Z(n764) );
  NAND U3436 ( .A(n6131), .B(n764), .Z(n765) );
  NANDN U3437 ( .A(n6133), .B(n765), .Z(n766) );
  AND U3438 ( .A(n6135), .B(n766), .Z(n767) );
  OR U3439 ( .A(n6137), .B(n767), .Z(n768) );
  NAND U3440 ( .A(n6139), .B(n768), .Z(n769) );
  NANDN U3441 ( .A(n6141), .B(n769), .Z(n770) );
  NAND U3442 ( .A(n6143), .B(n770), .Z(n771) );
  NANDN U3443 ( .A(n6145), .B(n771), .Z(n772) );
  AND U3444 ( .A(n6147), .B(n772), .Z(n773) );
  OR U3445 ( .A(n6149), .B(n773), .Z(n774) );
  NAND U3446 ( .A(n6151), .B(n774), .Z(n775) );
  NANDN U3447 ( .A(n6153), .B(n775), .Z(n776) );
  NAND U3448 ( .A(n6155), .B(n776), .Z(n777) );
  NANDN U3449 ( .A(n6157), .B(n777), .Z(n778) );
  AND U3450 ( .A(n6159), .B(n778), .Z(n779) );
  OR U3451 ( .A(n6161), .B(n779), .Z(n780) );
  NAND U3452 ( .A(n6163), .B(n780), .Z(n781) );
  NANDN U3453 ( .A(n6165), .B(n781), .Z(n782) );
  NAND U3454 ( .A(n6167), .B(n782), .Z(n783) );
  NANDN U3455 ( .A(n6169), .B(n783), .Z(n784) );
  AND U3456 ( .A(n6171), .B(n784), .Z(n785) );
  OR U3457 ( .A(n6173), .B(n785), .Z(n786) );
  NAND U3458 ( .A(n6175), .B(n786), .Z(n787) );
  NANDN U3459 ( .A(n6177), .B(n787), .Z(n788) );
  NAND U3460 ( .A(n6179), .B(n788), .Z(n789) );
  NANDN U3461 ( .A(n6181), .B(n789), .Z(n790) );
  AND U3462 ( .A(n6183), .B(n790), .Z(n791) );
  OR U3463 ( .A(n6185), .B(n791), .Z(n792) );
  NAND U3464 ( .A(n6187), .B(n792), .Z(n793) );
  NANDN U3465 ( .A(n6189), .B(n793), .Z(n794) );
  NAND U3466 ( .A(n6191), .B(n794), .Z(n795) );
  NANDN U3467 ( .A(n6193), .B(n795), .Z(n796) );
  AND U3468 ( .A(n6195), .B(n796), .Z(n797) );
  OR U3469 ( .A(n6197), .B(n797), .Z(n798) );
  NAND U3470 ( .A(n6199), .B(n798), .Z(n799) );
  NANDN U3471 ( .A(n6201), .B(n799), .Z(n800) );
  NAND U3472 ( .A(n6203), .B(n800), .Z(n801) );
  NANDN U3473 ( .A(n6205), .B(n801), .Z(n802) );
  AND U3474 ( .A(n6207), .B(n802), .Z(n803) );
  OR U3475 ( .A(n6209), .B(n803), .Z(n804) );
  NAND U3476 ( .A(n6211), .B(n804), .Z(n805) );
  NANDN U3477 ( .A(n6213), .B(n805), .Z(n806) );
  NAND U3478 ( .A(n6215), .B(n806), .Z(n807) );
  NANDN U3479 ( .A(n6217), .B(n807), .Z(n808) );
  AND U3480 ( .A(n6219), .B(n808), .Z(n809) );
  OR U3481 ( .A(n6221), .B(n809), .Z(n810) );
  NAND U3482 ( .A(n6223), .B(n810), .Z(n811) );
  NANDN U3483 ( .A(n6225), .B(n811), .Z(n812) );
  NAND U3484 ( .A(n6227), .B(n812), .Z(n813) );
  NANDN U3485 ( .A(n6229), .B(n813), .Z(n814) );
  AND U3486 ( .A(n6231), .B(n814), .Z(n815) );
  OR U3487 ( .A(n6233), .B(n815), .Z(n816) );
  NAND U3488 ( .A(n6235), .B(n816), .Z(n817) );
  NANDN U3489 ( .A(n6237), .B(n817), .Z(n818) );
  NAND U3490 ( .A(n6239), .B(n818), .Z(n819) );
  NANDN U3491 ( .A(n6241), .B(n819), .Z(n820) );
  AND U3492 ( .A(n6243), .B(n820), .Z(n821) );
  OR U3493 ( .A(n6245), .B(n821), .Z(n822) );
  NAND U3494 ( .A(n6247), .B(n822), .Z(n823) );
  NANDN U3495 ( .A(n6249), .B(n823), .Z(n824) );
  NAND U3496 ( .A(n6251), .B(n824), .Z(n825) );
  NANDN U3497 ( .A(n6253), .B(n825), .Z(n826) );
  AND U3498 ( .A(n6255), .B(n826), .Z(n827) );
  OR U3499 ( .A(n6257), .B(n827), .Z(n828) );
  NAND U3500 ( .A(n6259), .B(n828), .Z(n829) );
  NANDN U3501 ( .A(n6261), .B(n829), .Z(n830) );
  NAND U3502 ( .A(n6263), .B(n830), .Z(n831) );
  NANDN U3503 ( .A(n6265), .B(n831), .Z(n832) );
  AND U3504 ( .A(n6267), .B(n832), .Z(n833) );
  OR U3505 ( .A(n6269), .B(n833), .Z(n834) );
  NAND U3506 ( .A(n6271), .B(n834), .Z(n835) );
  NANDN U3507 ( .A(n6273), .B(n835), .Z(n836) );
  NAND U3508 ( .A(n6275), .B(n836), .Z(n837) );
  NANDN U3509 ( .A(n6277), .B(n837), .Z(n838) );
  AND U3510 ( .A(n6279), .B(n838), .Z(n839) );
  OR U3511 ( .A(n6281), .B(n839), .Z(n840) );
  NAND U3512 ( .A(n6283), .B(n840), .Z(n841) );
  NANDN U3513 ( .A(n6285), .B(n841), .Z(n842) );
  NAND U3514 ( .A(n6287), .B(n842), .Z(n843) );
  NANDN U3515 ( .A(n6289), .B(n843), .Z(n844) );
  AND U3516 ( .A(n6291), .B(n844), .Z(n845) );
  OR U3517 ( .A(n6293), .B(n845), .Z(n846) );
  NAND U3518 ( .A(n6295), .B(n846), .Z(n847) );
  NANDN U3519 ( .A(n6297), .B(n847), .Z(n848) );
  NAND U3520 ( .A(n6299), .B(n848), .Z(n849) );
  NANDN U3521 ( .A(n6301), .B(n849), .Z(n850) );
  AND U3522 ( .A(n6303), .B(n850), .Z(n851) );
  OR U3523 ( .A(n6305), .B(n851), .Z(n852) );
  NAND U3524 ( .A(n6307), .B(n852), .Z(n853) );
  NANDN U3525 ( .A(n6309), .B(n853), .Z(n854) );
  NAND U3526 ( .A(n6311), .B(n854), .Z(n855) );
  NANDN U3527 ( .A(n6313), .B(n855), .Z(n856) );
  AND U3528 ( .A(n6315), .B(n856), .Z(n857) );
  OR U3529 ( .A(n6317), .B(n857), .Z(n858) );
  NAND U3530 ( .A(n6319), .B(n858), .Z(n859) );
  NANDN U3531 ( .A(n6321), .B(n859), .Z(n860) );
  NAND U3532 ( .A(n6323), .B(n860), .Z(n861) );
  NANDN U3533 ( .A(n6325), .B(n861), .Z(n862) );
  AND U3534 ( .A(n6327), .B(n862), .Z(n863) );
  OR U3535 ( .A(n6329), .B(n863), .Z(n864) );
  NAND U3536 ( .A(n6331), .B(n864), .Z(n865) );
  NANDN U3537 ( .A(n6333), .B(n865), .Z(n866) );
  NAND U3538 ( .A(n6335), .B(n866), .Z(n867) );
  NANDN U3539 ( .A(n6337), .B(n867), .Z(n868) );
  AND U3540 ( .A(n6339), .B(n868), .Z(n869) );
  OR U3541 ( .A(n6341), .B(n869), .Z(n870) );
  NAND U3542 ( .A(n6343), .B(n870), .Z(n871) );
  NANDN U3543 ( .A(n6345), .B(n871), .Z(n872) );
  NAND U3544 ( .A(n6347), .B(n872), .Z(n873) );
  NANDN U3545 ( .A(n6349), .B(n873), .Z(n874) );
  AND U3546 ( .A(n6351), .B(n874), .Z(n875) );
  OR U3547 ( .A(n6353), .B(n875), .Z(n876) );
  NAND U3548 ( .A(n6355), .B(n876), .Z(n877) );
  NANDN U3549 ( .A(n6357), .B(n877), .Z(n878) );
  NAND U3550 ( .A(n6359), .B(n878), .Z(n879) );
  NANDN U3551 ( .A(n6361), .B(n879), .Z(n880) );
  AND U3552 ( .A(n6363), .B(n880), .Z(n881) );
  OR U3553 ( .A(n6365), .B(n881), .Z(n882) );
  NAND U3554 ( .A(n6367), .B(n882), .Z(n883) );
  NANDN U3555 ( .A(n6369), .B(n883), .Z(n884) );
  NAND U3556 ( .A(n6371), .B(n884), .Z(n885) );
  NANDN U3557 ( .A(n6373), .B(n885), .Z(n886) );
  AND U3558 ( .A(n6375), .B(n886), .Z(n887) );
  OR U3559 ( .A(n6377), .B(n887), .Z(n888) );
  NAND U3560 ( .A(n6379), .B(n888), .Z(n889) );
  NANDN U3561 ( .A(n6381), .B(n889), .Z(n890) );
  NAND U3562 ( .A(n6383), .B(n890), .Z(n891) );
  NANDN U3563 ( .A(n6385), .B(n891), .Z(n892) );
  AND U3564 ( .A(n6387), .B(n892), .Z(n893) );
  OR U3565 ( .A(n6389), .B(n893), .Z(n894) );
  NAND U3566 ( .A(n6391), .B(n894), .Z(n895) );
  NANDN U3567 ( .A(n6393), .B(n895), .Z(n896) );
  NAND U3568 ( .A(n6395), .B(n896), .Z(n897) );
  NANDN U3569 ( .A(n6397), .B(n897), .Z(n898) );
  AND U3570 ( .A(n6399), .B(n898), .Z(n899) );
  OR U3571 ( .A(n6401), .B(n899), .Z(n900) );
  NAND U3572 ( .A(n6403), .B(n900), .Z(n901) );
  NANDN U3573 ( .A(n6405), .B(n901), .Z(n902) );
  NAND U3574 ( .A(n6407), .B(n902), .Z(n903) );
  NANDN U3575 ( .A(n6409), .B(n903), .Z(n904) );
  AND U3576 ( .A(n6411), .B(n904), .Z(n905) );
  OR U3577 ( .A(n6413), .B(n905), .Z(n906) );
  NAND U3578 ( .A(n6415), .B(n906), .Z(n907) );
  NANDN U3579 ( .A(n6417), .B(n907), .Z(n908) );
  NAND U3580 ( .A(n6419), .B(n908), .Z(n909) );
  NANDN U3581 ( .A(n6421), .B(n909), .Z(n910) );
  AND U3582 ( .A(n6423), .B(n910), .Z(n911) );
  OR U3583 ( .A(n6425), .B(n911), .Z(n912) );
  NAND U3584 ( .A(n6427), .B(n912), .Z(n913) );
  NANDN U3585 ( .A(n6429), .B(n913), .Z(n914) );
  NAND U3586 ( .A(n6431), .B(n914), .Z(n915) );
  NANDN U3587 ( .A(n6433), .B(n915), .Z(n916) );
  AND U3588 ( .A(n6435), .B(n916), .Z(n917) );
  OR U3589 ( .A(n6437), .B(n917), .Z(n918) );
  NAND U3590 ( .A(n6439), .B(n918), .Z(n919) );
  NANDN U3591 ( .A(n6441), .B(n919), .Z(n920) );
  NAND U3592 ( .A(n6443), .B(n920), .Z(n921) );
  NANDN U3593 ( .A(n6445), .B(n921), .Z(n922) );
  AND U3594 ( .A(n6447), .B(n922), .Z(n923) );
  OR U3595 ( .A(n6449), .B(n923), .Z(n924) );
  NAND U3596 ( .A(n6451), .B(n924), .Z(n925) );
  NANDN U3597 ( .A(n6453), .B(n925), .Z(n926) );
  NAND U3598 ( .A(n6455), .B(n926), .Z(n927) );
  NANDN U3599 ( .A(n6457), .B(n927), .Z(n928) );
  AND U3600 ( .A(n6459), .B(n928), .Z(n929) );
  OR U3601 ( .A(n6461), .B(n929), .Z(n930) );
  NAND U3602 ( .A(n6463), .B(n930), .Z(n931) );
  NANDN U3603 ( .A(n6465), .B(n931), .Z(n932) );
  NAND U3604 ( .A(n6467), .B(n932), .Z(n933) );
  NANDN U3605 ( .A(n6469), .B(n933), .Z(n934) );
  AND U3606 ( .A(n6471), .B(n934), .Z(n935) );
  OR U3607 ( .A(n6473), .B(n935), .Z(n936) );
  NAND U3608 ( .A(n6475), .B(n936), .Z(n937) );
  NANDN U3609 ( .A(n6477), .B(n937), .Z(n938) );
  NAND U3610 ( .A(n6479), .B(n938), .Z(n939) );
  NANDN U3611 ( .A(n6481), .B(n939), .Z(n940) );
  AND U3612 ( .A(n6483), .B(n940), .Z(n941) );
  OR U3613 ( .A(n6485), .B(n941), .Z(n942) );
  NAND U3614 ( .A(n6487), .B(n942), .Z(n943) );
  NANDN U3615 ( .A(n6489), .B(n943), .Z(n944) );
  NAND U3616 ( .A(n6491), .B(n944), .Z(n945) );
  NANDN U3617 ( .A(n6493), .B(n945), .Z(n946) );
  AND U3618 ( .A(n6495), .B(n946), .Z(n947) );
  OR U3619 ( .A(n6497), .B(n947), .Z(n948) );
  NAND U3620 ( .A(n6499), .B(n948), .Z(n949) );
  NANDN U3621 ( .A(n6501), .B(n949), .Z(n950) );
  NAND U3622 ( .A(n6503), .B(n950), .Z(n951) );
  NANDN U3623 ( .A(n6505), .B(n951), .Z(n952) );
  AND U3624 ( .A(n6507), .B(n952), .Z(n953) );
  OR U3625 ( .A(n6509), .B(n953), .Z(n954) );
  NAND U3626 ( .A(n6511), .B(n954), .Z(n955) );
  NANDN U3627 ( .A(n6513), .B(n955), .Z(n956) );
  NAND U3628 ( .A(n6515), .B(n956), .Z(n957) );
  NANDN U3629 ( .A(n6517), .B(n957), .Z(n958) );
  AND U3630 ( .A(n6519), .B(n958), .Z(n959) );
  OR U3631 ( .A(n6521), .B(n959), .Z(n960) );
  NAND U3632 ( .A(n6523), .B(n960), .Z(n961) );
  NANDN U3633 ( .A(n6525), .B(n961), .Z(n962) );
  NAND U3634 ( .A(n6527), .B(n962), .Z(n963) );
  NANDN U3635 ( .A(n6529), .B(n963), .Z(n964) );
  AND U3636 ( .A(n6531), .B(n964), .Z(n965) );
  OR U3637 ( .A(n6533), .B(n965), .Z(n966) );
  NAND U3638 ( .A(n6535), .B(n966), .Z(n967) );
  NANDN U3639 ( .A(n6537), .B(n967), .Z(n968) );
  NAND U3640 ( .A(n6539), .B(n968), .Z(n969) );
  NANDN U3641 ( .A(n6541), .B(n969), .Z(n970) );
  AND U3642 ( .A(n6543), .B(n970), .Z(n971) );
  OR U3643 ( .A(n6545), .B(n971), .Z(n972) );
  NAND U3644 ( .A(n6547), .B(n972), .Z(n973) );
  NANDN U3645 ( .A(n6549), .B(n973), .Z(n974) );
  NAND U3646 ( .A(n6551), .B(n974), .Z(n975) );
  NANDN U3647 ( .A(n6553), .B(n975), .Z(n976) );
  AND U3648 ( .A(n6555), .B(n976), .Z(n979) );
  NANDN U3649 ( .A(y[575]), .B(x[575]), .Z(n978) );
  NANDN U3650 ( .A(y[576]), .B(x[576]), .Z(n977) );
  AND U3651 ( .A(n978), .B(n977), .Z(n6557) );
  NANDN U3652 ( .A(n979), .B(n6557), .Z(n980) );
  NANDN U3653 ( .A(n6558), .B(n980), .Z(n981) );
  NANDN U3654 ( .A(n6561), .B(n981), .Z(n982) );
  NAND U3655 ( .A(n6563), .B(n982), .Z(n983) );
  NANDN U3656 ( .A(n6565), .B(n983), .Z(n984) );
  AND U3657 ( .A(n6567), .B(n984), .Z(n985) );
  OR U3658 ( .A(n6569), .B(n985), .Z(n986) );
  NAND U3659 ( .A(n6571), .B(n986), .Z(n987) );
  NANDN U3660 ( .A(n6573), .B(n987), .Z(n988) );
  NAND U3661 ( .A(n6575), .B(n988), .Z(n989) );
  NANDN U3662 ( .A(n6577), .B(n989), .Z(n990) );
  AND U3663 ( .A(n6579), .B(n990), .Z(n991) );
  OR U3664 ( .A(n6581), .B(n991), .Z(n992) );
  NAND U3665 ( .A(n6583), .B(n992), .Z(n993) );
  NANDN U3666 ( .A(n6585), .B(n993), .Z(n994) );
  NAND U3667 ( .A(n6587), .B(n994), .Z(n995) );
  NANDN U3668 ( .A(n6589), .B(n995), .Z(n996) );
  AND U3669 ( .A(n6591), .B(n996), .Z(n997) );
  OR U3670 ( .A(n6593), .B(n997), .Z(n998) );
  NAND U3671 ( .A(n6595), .B(n998), .Z(n999) );
  NANDN U3672 ( .A(n6597), .B(n999), .Z(n1000) );
  NAND U3673 ( .A(n6599), .B(n1000), .Z(n1001) );
  NANDN U3674 ( .A(n6601), .B(n1001), .Z(n1002) );
  AND U3675 ( .A(n6603), .B(n1002), .Z(n1003) );
  OR U3676 ( .A(n6605), .B(n1003), .Z(n1004) );
  NAND U3677 ( .A(n6607), .B(n1004), .Z(n1005) );
  NANDN U3678 ( .A(n6609), .B(n1005), .Z(n1006) );
  NAND U3679 ( .A(n6611), .B(n1006), .Z(n1007) );
  NANDN U3680 ( .A(n6613), .B(n1007), .Z(n1008) );
  AND U3681 ( .A(n6615), .B(n1008), .Z(n1009) );
  OR U3682 ( .A(n6617), .B(n1009), .Z(n1010) );
  NAND U3683 ( .A(n6619), .B(n1010), .Z(n1011) );
  NANDN U3684 ( .A(n6621), .B(n1011), .Z(n1012) );
  NAND U3685 ( .A(n6623), .B(n1012), .Z(n1013) );
  NANDN U3686 ( .A(n6625), .B(n1013), .Z(n1014) );
  AND U3687 ( .A(n6627), .B(n1014), .Z(n1015) );
  OR U3688 ( .A(n6629), .B(n1015), .Z(n1016) );
  NAND U3689 ( .A(n6631), .B(n1016), .Z(n1017) );
  NANDN U3690 ( .A(n6633), .B(n1017), .Z(n1018) );
  NAND U3691 ( .A(n6635), .B(n1018), .Z(n1019) );
  NANDN U3692 ( .A(n6637), .B(n1019), .Z(n1020) );
  AND U3693 ( .A(n6639), .B(n1020), .Z(n1021) );
  OR U3694 ( .A(n6641), .B(n1021), .Z(n1022) );
  NAND U3695 ( .A(n6643), .B(n1022), .Z(n1023) );
  NANDN U3696 ( .A(n6645), .B(n1023), .Z(n1024) );
  NAND U3697 ( .A(n6647), .B(n1024), .Z(n1025) );
  NANDN U3698 ( .A(n6649), .B(n1025), .Z(n1026) );
  AND U3699 ( .A(n6651), .B(n1026), .Z(n1027) );
  OR U3700 ( .A(n6653), .B(n1027), .Z(n1028) );
  NAND U3701 ( .A(n6655), .B(n1028), .Z(n1029) );
  NANDN U3702 ( .A(n6657), .B(n1029), .Z(n1030) );
  NAND U3703 ( .A(n6659), .B(n1030), .Z(n1031) );
  NANDN U3704 ( .A(n6661), .B(n1031), .Z(n1032) );
  AND U3705 ( .A(n6663), .B(n1032), .Z(n1033) );
  OR U3706 ( .A(n6665), .B(n1033), .Z(n1034) );
  NAND U3707 ( .A(n6667), .B(n1034), .Z(n1035) );
  NANDN U3708 ( .A(n6669), .B(n1035), .Z(n1036) );
  NAND U3709 ( .A(n6671), .B(n1036), .Z(n1037) );
  NANDN U3710 ( .A(n6673), .B(n1037), .Z(n1038) );
  AND U3711 ( .A(n6675), .B(n1038), .Z(n1039) );
  OR U3712 ( .A(n6677), .B(n1039), .Z(n1040) );
  NAND U3713 ( .A(n6679), .B(n1040), .Z(n1041) );
  NANDN U3714 ( .A(n6681), .B(n1041), .Z(n1042) );
  NAND U3715 ( .A(n6683), .B(n1042), .Z(n1043) );
  NANDN U3716 ( .A(n6685), .B(n1043), .Z(n1044) );
  AND U3717 ( .A(n6687), .B(n1044), .Z(n1045) );
  OR U3718 ( .A(n6689), .B(n1045), .Z(n1046) );
  NAND U3719 ( .A(n6691), .B(n1046), .Z(n1047) );
  NANDN U3720 ( .A(n6693), .B(n1047), .Z(n1048) );
  NAND U3721 ( .A(n6695), .B(n1048), .Z(n1049) );
  NANDN U3722 ( .A(n6697), .B(n1049), .Z(n1050) );
  AND U3723 ( .A(n6698), .B(n1050), .Z(n1051) );
  OR U3724 ( .A(n6699), .B(n1051), .Z(n1052) );
  NAND U3725 ( .A(n6700), .B(n1052), .Z(n1053) );
  NANDN U3726 ( .A(n6701), .B(n1053), .Z(n1054) );
  NAND U3727 ( .A(n6702), .B(n1054), .Z(n1055) );
  NANDN U3728 ( .A(n6703), .B(n1055), .Z(n1056) );
  AND U3729 ( .A(n6704), .B(n1056), .Z(n1057) );
  OR U3730 ( .A(n6705), .B(n1057), .Z(n1058) );
  AND U3731 ( .A(n1059), .B(n1058), .Z(n1061) );
  NANDN U3732 ( .A(y[655]), .B(x[655]), .Z(n6707) );
  NANDN U3733 ( .A(y[656]), .B(x[656]), .Z(n1837) );
  AND U3734 ( .A(n6707), .B(n1837), .Z(n1060) );
  NANDN U3735 ( .A(n1061), .B(n1060), .Z(n1062) );
  ANDN U3736 ( .B(y[657]), .A(x[657]), .Z(n6709) );
  ANDN U3737 ( .B(n1062), .A(n6709), .Z(n1063) );
  NANDN U3738 ( .A(x[656]), .B(y[656]), .Z(n4419) );
  NAND U3739 ( .A(n1063), .B(n4419), .Z(n1064) );
  ANDN U3740 ( .B(x[657]), .A(y[657]), .Z(n1836) );
  ANDN U3741 ( .B(n1064), .A(n1836), .Z(n1065) );
  NAND U3742 ( .A(n6710), .B(n1065), .Z(n1066) );
  NAND U3743 ( .A(n6711), .B(n1066), .Z(n1067) );
  NANDN U3744 ( .A(n6712), .B(n1067), .Z(n1068) );
  AND U3745 ( .A(n6713), .B(n1068), .Z(n1069) );
  OR U3746 ( .A(n6714), .B(n1069), .Z(n1070) );
  NAND U3747 ( .A(n6716), .B(n1070), .Z(n1071) );
  NANDN U3748 ( .A(n6718), .B(n1071), .Z(n1072) );
  NAND U3749 ( .A(n6720), .B(n1072), .Z(n1073) );
  NANDN U3750 ( .A(n6722), .B(n1073), .Z(n1074) );
  AND U3751 ( .A(n6724), .B(n1074), .Z(n1075) );
  OR U3752 ( .A(n6726), .B(n1075), .Z(n1076) );
  NAND U3753 ( .A(n6728), .B(n1076), .Z(n1077) );
  NANDN U3754 ( .A(n6730), .B(n1077), .Z(n1078) );
  NAND U3755 ( .A(n6732), .B(n1078), .Z(n1079) );
  NANDN U3756 ( .A(n6734), .B(n1079), .Z(n1080) );
  AND U3757 ( .A(n6736), .B(n1080), .Z(n1081) );
  OR U3758 ( .A(n6738), .B(n1081), .Z(n1082) );
  NAND U3759 ( .A(n6740), .B(n1082), .Z(n1083) );
  NANDN U3760 ( .A(n6742), .B(n1083), .Z(n1084) );
  NAND U3761 ( .A(n6744), .B(n1084), .Z(n1085) );
  NANDN U3762 ( .A(n6746), .B(n1085), .Z(n1086) );
  AND U3763 ( .A(n6748), .B(n1086), .Z(n1087) );
  OR U3764 ( .A(n6750), .B(n1087), .Z(n1088) );
  NAND U3765 ( .A(n6752), .B(n1088), .Z(n1089) );
  NANDN U3766 ( .A(n6754), .B(n1089), .Z(n1090) );
  NAND U3767 ( .A(n6756), .B(n1090), .Z(n1091) );
  NANDN U3768 ( .A(n6758), .B(n1091), .Z(n1092) );
  AND U3769 ( .A(n6760), .B(n1092), .Z(n1093) );
  OR U3770 ( .A(n6762), .B(n1093), .Z(n1094) );
  NAND U3771 ( .A(n6764), .B(n1094), .Z(n1095) );
  NANDN U3772 ( .A(n6766), .B(n1095), .Z(n1096) );
  NAND U3773 ( .A(n6768), .B(n1096), .Z(n1097) );
  NANDN U3774 ( .A(n6770), .B(n1097), .Z(n1098) );
  AND U3775 ( .A(n6772), .B(n1098), .Z(n1099) );
  OR U3776 ( .A(n6774), .B(n1099), .Z(n1100) );
  NAND U3777 ( .A(n6776), .B(n1100), .Z(n1101) );
  NANDN U3778 ( .A(n6778), .B(n1101), .Z(n1102) );
  NAND U3779 ( .A(n6780), .B(n1102), .Z(n1103) );
  NANDN U3780 ( .A(n6782), .B(n1103), .Z(n1104) );
  AND U3781 ( .A(n6784), .B(n1104), .Z(n1105) );
  OR U3782 ( .A(n6786), .B(n1105), .Z(n1106) );
  NAND U3783 ( .A(n6788), .B(n1106), .Z(n1107) );
  NANDN U3784 ( .A(n6790), .B(n1107), .Z(n1108) );
  NAND U3785 ( .A(n6792), .B(n1108), .Z(n1109) );
  NANDN U3786 ( .A(n6794), .B(n1109), .Z(n1110) );
  AND U3787 ( .A(n6796), .B(n1110), .Z(n1111) );
  OR U3788 ( .A(n6798), .B(n1111), .Z(n1112) );
  NAND U3789 ( .A(n6800), .B(n1112), .Z(n1113) );
  NANDN U3790 ( .A(n6802), .B(n1113), .Z(n1114) );
  NAND U3791 ( .A(n6804), .B(n1114), .Z(n1115) );
  NANDN U3792 ( .A(n6806), .B(n1115), .Z(n1116) );
  AND U3793 ( .A(n6808), .B(n1116), .Z(n1117) );
  OR U3794 ( .A(n6810), .B(n1117), .Z(n1118) );
  NAND U3795 ( .A(n6812), .B(n1118), .Z(n1119) );
  NANDN U3796 ( .A(n6814), .B(n1119), .Z(n1120) );
  NAND U3797 ( .A(n6816), .B(n1120), .Z(n1121) );
  NANDN U3798 ( .A(n6818), .B(n1121), .Z(n1122) );
  AND U3799 ( .A(n6820), .B(n1122), .Z(n1123) );
  OR U3800 ( .A(n6822), .B(n1123), .Z(n1124) );
  NAND U3801 ( .A(n6824), .B(n1124), .Z(n1125) );
  NANDN U3802 ( .A(n6826), .B(n1125), .Z(n1126) );
  NAND U3803 ( .A(n6828), .B(n1126), .Z(n1127) );
  NANDN U3804 ( .A(n6830), .B(n1127), .Z(n1128) );
  AND U3805 ( .A(n6832), .B(n1128), .Z(n1129) );
  OR U3806 ( .A(n6834), .B(n1129), .Z(n1130) );
  NAND U3807 ( .A(n6836), .B(n1130), .Z(n1131) );
  NANDN U3808 ( .A(n6838), .B(n1131), .Z(n1132) );
  NANDN U3809 ( .A(n6839), .B(n1132), .Z(n1133) );
  NANDN U3810 ( .A(n6842), .B(n1133), .Z(n1134) );
  AND U3811 ( .A(n6844), .B(n1134), .Z(n1135) );
  OR U3812 ( .A(n6846), .B(n1135), .Z(n1136) );
  NAND U3813 ( .A(n6848), .B(n1136), .Z(n1137) );
  NANDN U3814 ( .A(n6850), .B(n1137), .Z(n1138) );
  NAND U3815 ( .A(n6852), .B(n1138), .Z(n1139) );
  NANDN U3816 ( .A(n6854), .B(n1139), .Z(n1140) );
  AND U3817 ( .A(n6856), .B(n1140), .Z(n1141) );
  OR U3818 ( .A(n6858), .B(n1141), .Z(n1142) );
  NAND U3819 ( .A(n6860), .B(n1142), .Z(n1143) );
  NANDN U3820 ( .A(n6862), .B(n1143), .Z(n1144) );
  NAND U3821 ( .A(n6864), .B(n1144), .Z(n1145) );
  NANDN U3822 ( .A(n6866), .B(n1145), .Z(n1146) );
  AND U3823 ( .A(n6868), .B(n1146), .Z(n1147) );
  OR U3824 ( .A(n6870), .B(n1147), .Z(n1148) );
  NAND U3825 ( .A(n6872), .B(n1148), .Z(n1149) );
  NANDN U3826 ( .A(n6874), .B(n1149), .Z(n1150) );
  NAND U3827 ( .A(n6876), .B(n1150), .Z(n1151) );
  NANDN U3828 ( .A(n6878), .B(n1151), .Z(n1152) );
  AND U3829 ( .A(n6880), .B(n1152), .Z(n1153) );
  OR U3830 ( .A(n6882), .B(n1153), .Z(n1154) );
  NAND U3831 ( .A(n6884), .B(n1154), .Z(n1155) );
  NANDN U3832 ( .A(n6886), .B(n1155), .Z(n1156) );
  NAND U3833 ( .A(n6888), .B(n1156), .Z(n1157) );
  NANDN U3834 ( .A(n6890), .B(n1157), .Z(n1158) );
  AND U3835 ( .A(n6892), .B(n1158), .Z(n1159) );
  OR U3836 ( .A(n6894), .B(n1159), .Z(n1160) );
  NAND U3837 ( .A(n6896), .B(n1160), .Z(n1161) );
  NANDN U3838 ( .A(n6898), .B(n1161), .Z(n1162) );
  NAND U3839 ( .A(n6900), .B(n1162), .Z(n1163) );
  NANDN U3840 ( .A(n6902), .B(n1163), .Z(n1164) );
  AND U3841 ( .A(n6904), .B(n1164), .Z(n1165) );
  OR U3842 ( .A(n6906), .B(n1165), .Z(n1166) );
  NAND U3843 ( .A(n6908), .B(n1166), .Z(n1167) );
  NANDN U3844 ( .A(n6910), .B(n1167), .Z(n1168) );
  NAND U3845 ( .A(n6912), .B(n1168), .Z(n1169) );
  NANDN U3846 ( .A(n6914), .B(n1169), .Z(n1170) );
  AND U3847 ( .A(n6916), .B(n1170), .Z(n1171) );
  OR U3848 ( .A(n6918), .B(n1171), .Z(n1172) );
  NAND U3849 ( .A(n6920), .B(n1172), .Z(n1173) );
  NANDN U3850 ( .A(n6922), .B(n1173), .Z(n1174) );
  NAND U3851 ( .A(n6924), .B(n1174), .Z(n1175) );
  NANDN U3852 ( .A(n6926), .B(n1175), .Z(n1176) );
  AND U3853 ( .A(n6928), .B(n1176), .Z(n1177) );
  OR U3854 ( .A(n6930), .B(n1177), .Z(n1178) );
  NAND U3855 ( .A(n6932), .B(n1178), .Z(n1179) );
  NANDN U3856 ( .A(n6934), .B(n1179), .Z(n1180) );
  NAND U3857 ( .A(n6936), .B(n1180), .Z(n1181) );
  NANDN U3858 ( .A(n6938), .B(n1181), .Z(n1182) );
  AND U3859 ( .A(n6940), .B(n1182), .Z(n1183) );
  OR U3860 ( .A(n6942), .B(n1183), .Z(n1184) );
  NAND U3861 ( .A(n6944), .B(n1184), .Z(n1185) );
  NANDN U3862 ( .A(n6946), .B(n1185), .Z(n1186) );
  NAND U3863 ( .A(n6948), .B(n1186), .Z(n1187) );
  NANDN U3864 ( .A(n6950), .B(n1187), .Z(n1188) );
  AND U3865 ( .A(n6952), .B(n1188), .Z(n1189) );
  OR U3866 ( .A(n6954), .B(n1189), .Z(n1190) );
  NAND U3867 ( .A(n6956), .B(n1190), .Z(n1191) );
  NANDN U3868 ( .A(n6958), .B(n1191), .Z(n1192) );
  NAND U3869 ( .A(n6960), .B(n1192), .Z(n1193) );
  NANDN U3870 ( .A(n6962), .B(n1193), .Z(n1194) );
  AND U3871 ( .A(n6964), .B(n1194), .Z(n1195) );
  OR U3872 ( .A(n6966), .B(n1195), .Z(n1196) );
  NAND U3873 ( .A(n6968), .B(n1196), .Z(n1197) );
  NANDN U3874 ( .A(n6970), .B(n1197), .Z(n1198) );
  NAND U3875 ( .A(n6972), .B(n1198), .Z(n1199) );
  NANDN U3876 ( .A(n6974), .B(n1199), .Z(n1200) );
  AND U3877 ( .A(n6976), .B(n1200), .Z(n1201) );
  OR U3878 ( .A(n6978), .B(n1201), .Z(n1202) );
  NAND U3879 ( .A(n6980), .B(n1202), .Z(n1203) );
  NANDN U3880 ( .A(n6982), .B(n1203), .Z(n1204) );
  NAND U3881 ( .A(n6984), .B(n1204), .Z(n1205) );
  NANDN U3882 ( .A(n6986), .B(n1205), .Z(n1206) );
  AND U3883 ( .A(n6988), .B(n1206), .Z(n1207) );
  OR U3884 ( .A(n6990), .B(n1207), .Z(n1208) );
  NAND U3885 ( .A(n6992), .B(n1208), .Z(n1209) );
  NANDN U3886 ( .A(n6994), .B(n1209), .Z(n1210) );
  NAND U3887 ( .A(n6996), .B(n1210), .Z(n1211) );
  NANDN U3888 ( .A(n6998), .B(n1211), .Z(n1212) );
  AND U3889 ( .A(n7000), .B(n1212), .Z(n1213) );
  OR U3890 ( .A(n7002), .B(n1213), .Z(n1214) );
  NAND U3891 ( .A(n7004), .B(n1214), .Z(n1215) );
  NANDN U3892 ( .A(n7006), .B(n1215), .Z(n1216) );
  NAND U3893 ( .A(n7008), .B(n1216), .Z(n1217) );
  NANDN U3894 ( .A(n7010), .B(n1217), .Z(n1218) );
  AND U3895 ( .A(n7012), .B(n1218), .Z(n1219) );
  OR U3896 ( .A(n7014), .B(n1219), .Z(n1220) );
  NAND U3897 ( .A(n7016), .B(n1220), .Z(n1221) );
  NANDN U3898 ( .A(n7018), .B(n1221), .Z(n1222) );
  NAND U3899 ( .A(n7020), .B(n1222), .Z(n1223) );
  NANDN U3900 ( .A(n7022), .B(n1223), .Z(n1224) );
  AND U3901 ( .A(n7024), .B(n1224), .Z(n1225) );
  OR U3902 ( .A(n7026), .B(n1225), .Z(n1226) );
  NAND U3903 ( .A(n7028), .B(n1226), .Z(n1227) );
  NANDN U3904 ( .A(n7030), .B(n1227), .Z(n1228) );
  NAND U3905 ( .A(n7032), .B(n1228), .Z(n1229) );
  NANDN U3906 ( .A(n7034), .B(n1229), .Z(n1230) );
  AND U3907 ( .A(n7036), .B(n1230), .Z(n1232) );
  NANDN U3908 ( .A(y[823]), .B(x[823]), .Z(n7037) );
  ANDN U3909 ( .B(x[824]), .A(y[824]), .Z(n1765) );
  ANDN U3910 ( .B(n7037), .A(n1765), .Z(n1231) );
  NANDN U3911 ( .A(n1232), .B(n1231), .Z(n1233) );
  ANDN U3912 ( .B(y[824]), .A(x[824]), .Z(n7038) );
  ANDN U3913 ( .B(n1233), .A(n7038), .Z(n1234) );
  NANDN U3914 ( .A(x[825]), .B(y[825]), .Z(n1764) );
  NAND U3915 ( .A(n1234), .B(n1764), .Z(n1235) );
  NANDN U3916 ( .A(y[826]), .B(x[826]), .Z(n1762) );
  AND U3917 ( .A(n1235), .B(n1762), .Z(n1236) );
  NAND U3918 ( .A(n1767), .B(n1236), .Z(n1237) );
  NANDN U3919 ( .A(x[826]), .B(y[826]), .Z(n1763) );
  AND U3920 ( .A(n1237), .B(n1763), .Z(n1238) );
  NANDN U3921 ( .A(n5423), .B(n1238), .Z(n1239) );
  NANDN U3922 ( .A(n5023), .B(n1239), .Z(n1240) );
  ANDN U3923 ( .B(x[827]), .A(y[827]), .Z(n1761) );
  OR U3924 ( .A(n1240), .B(n1761), .Z(n1241) );
  AND U3925 ( .A(n5424), .B(n1241), .Z(n1242) );
  NANDN U3926 ( .A(x[829]), .B(y[829]), .Z(n1756) );
  NAND U3927 ( .A(n1242), .B(n1756), .Z(n1243) );
  ANDN U3928 ( .B(x[830]), .A(y[830]), .Z(n1751) );
  ANDN U3929 ( .B(n1243), .A(n1751), .Z(n1244) );
  NANDN U3930 ( .A(n1758), .B(n1244), .Z(n1245) );
  NAND U3931 ( .A(n1757), .B(n1245), .Z(n1246) );
  NANDN U3932 ( .A(y[832]), .B(x[832]), .Z(n1749) );
  AND U3933 ( .A(n1246), .B(n1749), .Z(n1247) );
  NANDN U3934 ( .A(n1753), .B(n1247), .Z(n1248) );
  ANDN U3935 ( .B(y[832]), .A(x[832]), .Z(n7044) );
  ANDN U3936 ( .B(n1248), .A(n7044), .Z(n1249) );
  NAND U3937 ( .A(n7046), .B(n1249), .Z(n1250) );
  NAND U3938 ( .A(n5029), .B(n1250), .Z(n1251) );
  ANDN U3939 ( .B(x[833]), .A(y[833]), .Z(n1748) );
  OR U3940 ( .A(n1251), .B(n1748), .Z(n1252) );
  NAND U3941 ( .A(n1253), .B(n1252), .Z(n1254) );
  NANDN U3942 ( .A(n7050), .B(n1254), .Z(n1255) );
  ANDN U3943 ( .B(x[835]), .A(y[835]), .Z(n1747) );
  OR U3944 ( .A(n1255), .B(n1747), .Z(n1256) );
  NAND U3945 ( .A(n7052), .B(n1256), .Z(n1257) );
  NANDN U3946 ( .A(n7053), .B(n1257), .Z(n1258) );
  NAND U3947 ( .A(n7054), .B(n1258), .Z(n1259) );
  ANDN U3948 ( .B(x[840]), .A(y[840]), .Z(n1745) );
  ANDN U3949 ( .B(n1259), .A(n1745), .Z(n1260) );
  NANDN U3950 ( .A(n7055), .B(n1260), .Z(n1261) );
  NANDN U3951 ( .A(x[840]), .B(y[840]), .Z(n7056) );
  AND U3952 ( .A(n1261), .B(n7056), .Z(n1262) );
  NAND U3953 ( .A(n1743), .B(n1262), .Z(n1263) );
  NAND U3954 ( .A(n1746), .B(n1263), .Z(n1264) );
  ANDN U3955 ( .B(x[842]), .A(y[842]), .Z(n1741) );
  OR U3956 ( .A(n1264), .B(n1741), .Z(n1265) );
  NAND U3957 ( .A(n1744), .B(n1265), .Z(n1266) );
  NANDN U3958 ( .A(n1742), .B(n1266), .Z(n1267) );
  NANDN U3959 ( .A(y[844]), .B(x[844]), .Z(n1739) );
  NANDN U3960 ( .A(n1267), .B(n1739), .Z(n1268) );
  AND U3961 ( .A(n1269), .B(n1268), .Z(n1271) );
  NANDN U3962 ( .A(y[846]), .B(x[846]), .Z(n1735) );
  ANDN U3963 ( .B(x[845]), .A(y[845]), .Z(n1738) );
  ANDN U3964 ( .B(n1735), .A(n1738), .Z(n1270) );
  NANDN U3965 ( .A(n1271), .B(n1270), .Z(n1272) );
  AND U3966 ( .A(n1736), .B(n1272), .Z(n1273) );
  NANDN U3967 ( .A(x[847]), .B(y[847]), .Z(n1732) );
  NAND U3968 ( .A(n1273), .B(n1732), .Z(n1274) );
  ANDN U3969 ( .B(x[848]), .A(y[848]), .Z(n1730) );
  ANDN U3970 ( .B(n1274), .A(n1730), .Z(n1275) );
  NAND U3971 ( .A(n1734), .B(n1275), .Z(n1276) );
  NAND U3972 ( .A(n1733), .B(n1276), .Z(n1277) );
  NANDN U3973 ( .A(n7064), .B(n1277), .Z(n1278) );
  AND U3974 ( .A(n7066), .B(n1278), .Z(n1279) );
  OR U3975 ( .A(n7067), .B(n1279), .Z(n1280) );
  NAND U3976 ( .A(n7068), .B(n1280), .Z(n1281) );
  NAND U3977 ( .A(n7069), .B(n1281), .Z(n1282) );
  ANDN U3978 ( .B(x[856]), .A(y[856]), .Z(n1727) );
  OR U3979 ( .A(n1282), .B(n1727), .Z(n1283) );
  NAND U3980 ( .A(n1284), .B(n1283), .Z(n1285) );
  NANDN U3981 ( .A(y[857]), .B(x[857]), .Z(n1728) );
  AND U3982 ( .A(n1285), .B(n1728), .Z(n1286) );
  NAND U3983 ( .A(n1725), .B(n1286), .Z(n1287) );
  NANDN U3984 ( .A(n5076), .B(n1287), .Z(n1288) );
  ANDN U3985 ( .B(y[859]), .A(x[859]), .Z(n1723) );
  OR U3986 ( .A(n1288), .B(n1723), .Z(n1289) );
  AND U3987 ( .A(n1290), .B(n1289), .Z(n1292) );
  NANDN U3988 ( .A(x[861]), .B(y[861]), .Z(n1719) );
  ANDN U3989 ( .B(y[860]), .A(x[860]), .Z(n1724) );
  ANDN U3990 ( .B(n1719), .A(n1724), .Z(n1291) );
  NANDN U3991 ( .A(n1292), .B(n1291), .Z(n1293) );
  AND U3992 ( .A(n1722), .B(n1293), .Z(n1294) );
  NAND U3993 ( .A(n5083), .B(n1294), .Z(n1295) );
  NAND U3994 ( .A(n1720), .B(n1295), .Z(n1296) );
  AND U3995 ( .A(n5085), .B(n1296), .Z(n1297) );
  NANDN U3996 ( .A(y[864]), .B(x[864]), .Z(n1717) );
  NAND U3997 ( .A(n1297), .B(n1717), .Z(n1298) );
  NANDN U3998 ( .A(x[865]), .B(y[865]), .Z(n5419) );
  AND U3999 ( .A(n1298), .B(n5419), .Z(n1299) );
  NANDN U4000 ( .A(n1718), .B(n1299), .Z(n1300) );
  NANDN U4001 ( .A(y[866]), .B(x[866]), .Z(n1715) );
  AND U4002 ( .A(n1300), .B(n1715), .Z(n1301) );
  NAND U4003 ( .A(n1716), .B(n1301), .Z(n1302) );
  NANDN U4004 ( .A(n5417), .B(n1302), .Z(n1303) );
  NANDN U4005 ( .A(y[867]), .B(x[867]), .Z(n1714) );
  AND U4006 ( .A(n1303), .B(n1714), .Z(n1304) );
  NAND U4007 ( .A(n5098), .B(n1304), .Z(n1305) );
  NANDN U4008 ( .A(n5414), .B(n1305), .Z(n1306) );
  NAND U4009 ( .A(n7101), .B(n1306), .Z(n1307) );
  NANDN U4010 ( .A(n7102), .B(n1307), .Z(n1308) );
  NANDN U4011 ( .A(y[871]), .B(x[871]), .Z(n5104) );
  AND U4012 ( .A(n1308), .B(n5104), .Z(n1309) );
  NANDN U4013 ( .A(y[872]), .B(x[872]), .Z(n1708) );
  NAND U4014 ( .A(n1309), .B(n1708), .Z(n1310) );
  NANDN U4015 ( .A(x[873]), .B(y[873]), .Z(n1707) );
  AND U4016 ( .A(n1310), .B(n1707), .Z(n1311) );
  NANDN U4017 ( .A(n1710), .B(n1311), .Z(n1312) );
  NANDN U4018 ( .A(y[873]), .B(x[873]), .Z(n1709) );
  AND U4019 ( .A(n1312), .B(n1709), .Z(n1313) );
  NAND U4020 ( .A(n1704), .B(n1313), .Z(n1314) );
  NANDN U4021 ( .A(n1706), .B(n1314), .Z(n1315) );
  ANDN U4022 ( .B(y[875]), .A(x[875]), .Z(n1701) );
  OR U4023 ( .A(n1315), .B(n1701), .Z(n1316) );
  NAND U4024 ( .A(n1317), .B(n1316), .Z(n1318) );
  NANDN U4025 ( .A(x[876]), .B(y[876]), .Z(n1702) );
  AND U4026 ( .A(n1318), .B(n1702), .Z(n1319) );
  NAND U4027 ( .A(n1698), .B(n1319), .Z(n1320) );
  NANDN U4028 ( .A(n1699), .B(n1320), .Z(n1321) );
  ANDN U4029 ( .B(x[878]), .A(y[878]), .Z(n1695) );
  OR U4030 ( .A(n1321), .B(n1695), .Z(n1322) );
  AND U4031 ( .A(n7126), .B(n1322), .Z(n1323) );
  NANDN U4032 ( .A(n1697), .B(n1323), .Z(n1324) );
  AND U4033 ( .A(n1325), .B(n1324), .Z(n1327) );
  NANDN U4034 ( .A(x[880]), .B(y[880]), .Z(n1326) );
  NANDN U4035 ( .A(x[881]), .B(y[881]), .Z(n5413) );
  NAND U4036 ( .A(n1326), .B(n5413), .Z(n7123) );
  OR U4037 ( .A(n1327), .B(n7123), .Z(n1328) );
  AND U4038 ( .A(n1692), .B(n1328), .Z(n1329) );
  NAND U4039 ( .A(n1691), .B(n1329), .Z(n1330) );
  NANDN U4040 ( .A(n5411), .B(n1330), .Z(n1331) );
  AND U4041 ( .A(n7135), .B(n1331), .Z(n1332) );
  ANDN U4042 ( .B(y[885]), .A(x[885]), .Z(n5130) );
  NANDN U4043 ( .A(x[884]), .B(y[884]), .Z(n5125) );
  NANDN U4044 ( .A(n5130), .B(n5125), .Z(n5410) );
  OR U4045 ( .A(n1332), .B(n5410), .Z(n1333) );
  NAND U4046 ( .A(n5409), .B(n1333), .Z(n1334) );
  NANDN U4047 ( .A(n7140), .B(n1334), .Z(n1335) );
  NANDN U4048 ( .A(y[887]), .B(x[887]), .Z(n1688) );
  AND U4049 ( .A(n1335), .B(n1688), .Z(n1336) );
  NAND U4050 ( .A(n1685), .B(n1336), .Z(n1337) );
  NANDN U4051 ( .A(n1686), .B(n1337), .Z(n1338) );
  ANDN U4052 ( .B(y[889]), .A(x[889]), .Z(n1682) );
  OR U4053 ( .A(n1338), .B(n1682), .Z(n1339) );
  NAND U4054 ( .A(n1340), .B(n1339), .Z(n1341) );
  NANDN U4055 ( .A(x[890]), .B(y[890]), .Z(n1683) );
  AND U4056 ( .A(n1341), .B(n1683), .Z(n1342) );
  NAND U4057 ( .A(n1679), .B(n1342), .Z(n1343) );
  NANDN U4058 ( .A(n1680), .B(n1343), .Z(n1344) );
  ANDN U4059 ( .B(x[892]), .A(y[892]), .Z(n1676) );
  OR U4060 ( .A(n1344), .B(n1676), .Z(n1345) );
  AND U4061 ( .A(n1678), .B(n1345), .Z(n1346) );
  NANDN U4062 ( .A(x[893]), .B(y[893]), .Z(n1674) );
  NAND U4063 ( .A(n1346), .B(n1674), .Z(n1347) );
  NAND U4064 ( .A(n1677), .B(n1347), .Z(n1348) );
  ANDN U4065 ( .B(x[894]), .A(y[894]), .Z(n5146) );
  OR U4066 ( .A(n1348), .B(n5146), .Z(n1349) );
  NAND U4067 ( .A(n1675), .B(n1349), .Z(n1350) );
  NANDN U4068 ( .A(n5147), .B(n1350), .Z(n1351) );
  NANDN U4069 ( .A(y[896]), .B(x[896]), .Z(n1672) );
  NANDN U4070 ( .A(n1351), .B(n1672), .Z(n1352) );
  AND U4071 ( .A(n1353), .B(n1352), .Z(n1355) );
  NANDN U4072 ( .A(y[897]), .B(x[897]), .Z(n1673) );
  ANDN U4073 ( .B(x[898]), .A(y[898]), .Z(n1669) );
  ANDN U4074 ( .B(n1673), .A(n1669), .Z(n1354) );
  NANDN U4075 ( .A(n1355), .B(n1354), .Z(n1356) );
  NANDN U4076 ( .A(n7166), .B(n1356), .Z(n1357) );
  NANDN U4077 ( .A(y[899]), .B(x[899]), .Z(n1670) );
  AND U4078 ( .A(n1357), .B(n1670), .Z(n1358) );
  NAND U4079 ( .A(n5160), .B(n1358), .Z(n1359) );
  NANDN U4080 ( .A(n7175), .B(n1359), .Z(n1360) );
  NANDN U4081 ( .A(n7178), .B(n1360), .Z(n1361) );
  AND U4082 ( .A(n7181), .B(n1361), .Z(n1363) );
  NANDN U4083 ( .A(y[903]), .B(x[903]), .Z(n7182) );
  ANDN U4084 ( .B(x[904]), .A(y[904]), .Z(n1664) );
  ANDN U4085 ( .B(n7182), .A(n1664), .Z(n1362) );
  NANDN U4086 ( .A(n1363), .B(n1362), .Z(n1364) );
  ANDN U4087 ( .B(y[904]), .A(x[904]), .Z(n7185) );
  ANDN U4088 ( .B(n1364), .A(n7185), .Z(n1365) );
  NANDN U4089 ( .A(x[905]), .B(y[905]), .Z(n1663) );
  NAND U4090 ( .A(n1365), .B(n1663), .Z(n1366) );
  AND U4091 ( .A(n1666), .B(n1366), .Z(n1367) );
  NANDN U4092 ( .A(y[906]), .B(x[906]), .Z(n1661) );
  NAND U4093 ( .A(n1367), .B(n1661), .Z(n1368) );
  ANDN U4094 ( .B(y[907]), .A(x[907]), .Z(n1658) );
  ANDN U4095 ( .B(n1368), .A(n1658), .Z(n1369) );
  NANDN U4096 ( .A(n1662), .B(n1369), .Z(n1370) );
  NANDN U4097 ( .A(y[908]), .B(x[908]), .Z(n1656) );
  AND U4098 ( .A(n1370), .B(n1656), .Z(n1371) );
  NAND U4099 ( .A(n1660), .B(n1371), .Z(n1372) );
  NAND U4100 ( .A(n1659), .B(n1372), .Z(n1373) );
  NANDN U4101 ( .A(y[910]), .B(x[910]), .Z(n1653) );
  AND U4102 ( .A(n1373), .B(n1653), .Z(n1374) );
  NAND U4103 ( .A(n1657), .B(n1374), .Z(n1375) );
  NAND U4104 ( .A(n7197), .B(n1375), .Z(n1376) );
  NANDN U4105 ( .A(y[912]), .B(x[912]), .Z(n1651) );
  AND U4106 ( .A(n1376), .B(n1651), .Z(n1377) );
  NAND U4107 ( .A(n1654), .B(n1377), .Z(n1378) );
  NANDN U4108 ( .A(n1379), .B(n1378), .Z(n1381) );
  NANDN U4109 ( .A(y[913]), .B(x[913]), .Z(n1650) );
  NANDN U4110 ( .A(y[914]), .B(x[914]), .Z(n7206) );
  AND U4111 ( .A(n1650), .B(n7206), .Z(n1380) );
  NAND U4112 ( .A(n1381), .B(n1380), .Z(n1382) );
  AND U4113 ( .A(n7208), .B(n1382), .Z(n1383) );
  OR U4114 ( .A(n7209), .B(n1383), .Z(n1384) );
  NAND U4115 ( .A(n7210), .B(n1384), .Z(n1385) );
  NANDN U4116 ( .A(n7211), .B(n1385), .Z(n1386) );
  NAND U4117 ( .A(n7212), .B(n1386), .Z(n1387) );
  NANDN U4118 ( .A(y[920]), .B(x[920]), .Z(n1649) );
  AND U4119 ( .A(n1387), .B(n1649), .Z(n1388) );
  NAND U4120 ( .A(n7213), .B(n1388), .Z(n1389) );
  ANDN U4121 ( .B(y[920]), .A(x[920]), .Z(n7214) );
  ANDN U4122 ( .B(n1389), .A(n7214), .Z(n1390) );
  NAND U4123 ( .A(n1645), .B(n1390), .Z(n1391) );
  NANDN U4124 ( .A(n1647), .B(n1391), .Z(n1392) );
  ANDN U4125 ( .B(x[922]), .A(y[922]), .Z(n1640) );
  OR U4126 ( .A(n1392), .B(n1640), .Z(n1393) );
  NAND U4127 ( .A(n1646), .B(n1393), .Z(n1394) );
  NANDN U4128 ( .A(n1642), .B(n1394), .Z(n1395) );
  NANDN U4129 ( .A(y[924]), .B(x[924]), .Z(n1638) );
  NANDN U4130 ( .A(n1395), .B(n1638), .Z(n1396) );
  AND U4131 ( .A(n1636), .B(n1396), .Z(n1397) );
  NANDN U4132 ( .A(x[924]), .B(y[924]), .Z(n7218) );
  NAND U4133 ( .A(n1397), .B(n7218), .Z(n1398) );
  ANDN U4134 ( .B(x[926]), .A(y[926]), .Z(n1632) );
  ANDN U4135 ( .B(n1398), .A(n1632), .Z(n1399) );
  NANDN U4136 ( .A(n1637), .B(n1399), .Z(n1400) );
  NANDN U4137 ( .A(x[926]), .B(y[926]), .Z(n1635) );
  AND U4138 ( .A(n1400), .B(n1635), .Z(n1401) );
  NAND U4139 ( .A(n1631), .B(n1401), .Z(n1402) );
  NANDN U4140 ( .A(n1633), .B(n1402), .Z(n1403) );
  ANDN U4141 ( .B(x[928]), .A(y[928]), .Z(n5211) );
  OR U4142 ( .A(n1403), .B(n5211), .Z(n1404) );
  NAND U4143 ( .A(n1405), .B(n1404), .Z(n1406) );
  NANDN U4144 ( .A(y[929]), .B(x[929]), .Z(n5212) );
  AND U4145 ( .A(n1406), .B(n5212), .Z(n1407) );
  NAND U4146 ( .A(n1627), .B(n1407), .Z(n1408) );
  NANDN U4147 ( .A(n7227), .B(n1408), .Z(n1409) );
  ANDN U4148 ( .B(y[930]), .A(x[930]), .Z(n1628) );
  OR U4149 ( .A(n1409), .B(n1628), .Z(n1410) );
  AND U4150 ( .A(n1626), .B(n1410), .Z(n1411) );
  NAND U4151 ( .A(n7228), .B(n1411), .Z(n1412) );
  NANDN U4152 ( .A(n7229), .B(n1412), .Z(n1413) );
  AND U4153 ( .A(n7230), .B(n1413), .Z(n1415) );
  ANDN U4154 ( .B(y[935]), .A(x[935]), .Z(n5230) );
  NANDN U4155 ( .A(x[934]), .B(y[934]), .Z(n1414) );
  NANDN U4156 ( .A(n5230), .B(n1414), .Z(n7231) );
  OR U4157 ( .A(n1415), .B(n7231), .Z(n1416) );
  AND U4158 ( .A(n7232), .B(n1416), .Z(n1417) );
  NANDN U4159 ( .A(y[936]), .B(x[936]), .Z(n1624) );
  NAND U4160 ( .A(n1417), .B(n1624), .Z(n1418) );
  NANDN U4161 ( .A(x[937]), .B(y[937]), .Z(n5236) );
  AND U4162 ( .A(n1418), .B(n5236), .Z(n1419) );
  NANDN U4163 ( .A(n7233), .B(n1419), .Z(n1420) );
  NANDN U4164 ( .A(y[937]), .B(x[937]), .Z(n1625) );
  AND U4165 ( .A(n1420), .B(n1625), .Z(n1421) );
  NAND U4166 ( .A(n5239), .B(n1421), .Z(n1422) );
  NANDN U4167 ( .A(n5235), .B(n1422), .Z(n1423) );
  NANDN U4168 ( .A(x[939]), .B(y[939]), .Z(n5234) );
  NANDN U4169 ( .A(n1423), .B(n5234), .Z(n1424) );
  AND U4170 ( .A(n1425), .B(n1424), .Z(n1427) );
  NANDN U4171 ( .A(x[941]), .B(y[941]), .Z(n1623) );
  ANDN U4172 ( .B(y[940]), .A(x[940]), .Z(n5233) );
  ANDN U4173 ( .B(n1623), .A(n5233), .Z(n1426) );
  NANDN U4174 ( .A(n1427), .B(n1426), .Z(n1428) );
  AND U4175 ( .A(n5243), .B(n1428), .Z(n1429) );
  NAND U4176 ( .A(n5248), .B(n1429), .Z(n1430) );
  NANDN U4177 ( .A(n1622), .B(n1430), .Z(n1431) );
  AND U4178 ( .A(n5250), .B(n1431), .Z(n1432) );
  NANDN U4179 ( .A(y[944]), .B(x[944]), .Z(n1620) );
  NAND U4180 ( .A(n1432), .B(n1620), .Z(n1433) );
  ANDN U4181 ( .B(y[945]), .A(x[945]), .Z(n1617) );
  ANDN U4182 ( .B(n1433), .A(n1617), .Z(n1434) );
  NANDN U4183 ( .A(n1621), .B(n1434), .Z(n1435) );
  AND U4184 ( .A(n1618), .B(n1435), .Z(n1436) );
  NAND U4185 ( .A(n1619), .B(n1436), .Z(n1437) );
  NANDN U4186 ( .A(n7240), .B(n1437), .Z(n1438) );
  NANDN U4187 ( .A(y[947]), .B(x[947]), .Z(n5256) );
  AND U4188 ( .A(n1438), .B(n5256), .Z(n1439) );
  NAND U4189 ( .A(n1616), .B(n1439), .Z(n1440) );
  NANDN U4190 ( .A(n5401), .B(n1440), .Z(n1441) );
  NANDN U4191 ( .A(n7252), .B(n1441), .Z(n1442) );
  AND U4192 ( .A(n7254), .B(n1442), .Z(n1444) );
  ANDN U4193 ( .B(x[952]), .A(y[952]), .Z(n1612) );
  ANDN U4194 ( .B(x[951]), .A(y[951]), .Z(n7256) );
  NOR U4195 ( .A(n1612), .B(n7256), .Z(n1443) );
  NANDN U4196 ( .A(n1444), .B(n1443), .Z(n1445) );
  NANDN U4197 ( .A(n5399), .B(n1445), .Z(n1446) );
  ANDN U4198 ( .B(y[952]), .A(x[952]), .Z(n5400) );
  OR U4199 ( .A(n1446), .B(n5400), .Z(n1447) );
  AND U4200 ( .A(n1614), .B(n1447), .Z(n1448) );
  NAND U4201 ( .A(n1613), .B(n1448), .Z(n1449) );
  NAND U4202 ( .A(n1450), .B(n1449), .Z(n1451) );
  NANDN U4203 ( .A(y[955]), .B(x[955]), .Z(n1615) );
  AND U4204 ( .A(n1451), .B(n1615), .Z(n1452) );
  NAND U4205 ( .A(n1610), .B(n1452), .Z(n1453) );
  NANDN U4206 ( .A(n5277), .B(n1453), .Z(n1454) );
  ANDN U4207 ( .B(y[957]), .A(x[957]), .Z(n1607) );
  OR U4208 ( .A(n1454), .B(n1607), .Z(n1455) );
  AND U4209 ( .A(n1611), .B(n1455), .Z(n1456) );
  NANDN U4210 ( .A(n1604), .B(n1456), .Z(n1457) );
  NAND U4211 ( .A(n1458), .B(n1457), .Z(n1459) );
  NANDN U4212 ( .A(y[959]), .B(x[959]), .Z(n1606) );
  AND U4213 ( .A(n1459), .B(n1606), .Z(n1460) );
  NAND U4214 ( .A(n1600), .B(n1460), .Z(n1461) );
  NANDN U4215 ( .A(n1601), .B(n1461), .Z(n1462) );
  ANDN U4216 ( .B(y[961]), .A(x[961]), .Z(n1596) );
  OR U4217 ( .A(n1462), .B(n1596), .Z(n1463) );
  NANDN U4218 ( .A(y[962]), .B(x[962]), .Z(n1592) );
  AND U4219 ( .A(n1463), .B(n1592), .Z(n1464) );
  NANDN U4220 ( .A(n1598), .B(n1464), .Z(n1465) );
  AND U4221 ( .A(n1597), .B(n1465), .Z(n1466) );
  NANDN U4222 ( .A(y[963]), .B(x[963]), .Z(n1593) );
  NANDN U4223 ( .A(n1466), .B(n1593), .Z(n1467) );
  ANDN U4224 ( .B(x[964]), .A(y[964]), .Z(n1595) );
  OR U4225 ( .A(n1467), .B(n1595), .Z(n1468) );
  NAND U4226 ( .A(n5396), .B(n1468), .Z(n1469) );
  NANDN U4227 ( .A(n7277), .B(n1469), .Z(n1470) );
  NAND U4228 ( .A(n7278), .B(n1470), .Z(n1471) );
  ANDN U4229 ( .B(x[967]), .A(y[967]), .Z(n7279) );
  ANDN U4230 ( .B(n1471), .A(n7279), .Z(n1472) );
  NANDN U4231 ( .A(n1588), .B(n1472), .Z(n1473) );
  AND U4232 ( .A(n7283), .B(n1473), .Z(n1474) );
  NANDN U4233 ( .A(n7280), .B(n1474), .Z(n1475) );
  NANDN U4234 ( .A(n1590), .B(n1475), .Z(n1476) );
  NANDN U4235 ( .A(y[969]), .B(x[969]), .Z(n1589) );
  NANDN U4236 ( .A(n1476), .B(n1589), .Z(n1477) );
  AND U4237 ( .A(n7282), .B(n1477), .Z(n1478) );
  NANDN U4238 ( .A(x[971]), .B(y[971]), .Z(n5302) );
  NAND U4239 ( .A(n1478), .B(n5302), .Z(n1479) );
  NANDN U4240 ( .A(y[972]), .B(x[972]), .Z(n1587) );
  AND U4241 ( .A(n1479), .B(n1587), .Z(n1480) );
  NAND U4242 ( .A(n1591), .B(n1480), .Z(n1481) );
  NANDN U4243 ( .A(x[972]), .B(y[972]), .Z(n5301) );
  AND U4244 ( .A(n1481), .B(n5301), .Z(n1482) );
  NAND U4245 ( .A(n1583), .B(n1482), .Z(n1483) );
  NANDN U4246 ( .A(n5311), .B(n1483), .Z(n1484) );
  ANDN U4247 ( .B(x[973]), .A(y[973]), .Z(n1585) );
  OR U4248 ( .A(n1484), .B(n1585), .Z(n1485) );
  NAND U4249 ( .A(n1584), .B(n1485), .Z(n1486) );
  AND U4250 ( .A(n5306), .B(n1486), .Z(n1487) );
  NANDN U4251 ( .A(y[975]), .B(x[975]), .Z(n5312) );
  NAND U4252 ( .A(n1487), .B(n5312), .Z(n1488) );
  NANDN U4253 ( .A(n1489), .B(n1488), .Z(n1490) );
  AND U4254 ( .A(n7298), .B(n1490), .Z(n1491) );
  OR U4255 ( .A(n7300), .B(n1491), .Z(n1492) );
  NAND U4256 ( .A(n7302), .B(n1492), .Z(n1493) );
  NANDN U4257 ( .A(n7303), .B(n1493), .Z(n1494) );
  NANDN U4258 ( .A(n7306), .B(n1494), .Z(n1495) );
  AND U4259 ( .A(n7315), .B(n1495), .Z(n1496) );
  NANDN U4260 ( .A(n7309), .B(n1496), .Z(n1497) );
  ANDN U4261 ( .B(x[985]), .A(y[985]), .Z(n1580) );
  ANDN U4262 ( .B(n1497), .A(n1580), .Z(n1498) );
  NAND U4263 ( .A(n5337), .B(n1498), .Z(n1499) );
  NANDN U4264 ( .A(x[986]), .B(y[986]), .Z(n7312) );
  AND U4265 ( .A(n1499), .B(n7312), .Z(n1500) );
  NAND U4266 ( .A(n5342), .B(n1500), .Z(n1501) );
  NANDN U4267 ( .A(n1579), .B(n1501), .Z(n1502) );
  ANDN U4268 ( .B(x[988]), .A(y[988]), .Z(n1576) );
  OR U4269 ( .A(n1502), .B(n1576), .Z(n1503) );
  NAND U4270 ( .A(n1504), .B(n1503), .Z(n1505) );
  NANDN U4271 ( .A(n1563), .B(n1505), .Z(n1506) );
  NANDN U4272 ( .A(x[990]), .B(y[990]), .Z(n1572) );
  AND U4273 ( .A(n1506), .B(n1572), .Z(n1507) );
  NAND U4274 ( .A(n1566), .B(n1507), .Z(n1508) );
  NANDN U4275 ( .A(n1560), .B(n1508), .Z(n1509) );
  NANDN U4276 ( .A(x[992]), .B(y[992]), .Z(n1567) );
  AND U4277 ( .A(n1509), .B(n1567), .Z(n1510) );
  NAND U4278 ( .A(n1555), .B(n1510), .Z(n1511) );
  NAND U4279 ( .A(n1562), .B(n1511), .Z(n1512) );
  ANDN U4280 ( .B(x[994]), .A(y[994]), .Z(n5348) );
  OR U4281 ( .A(n1512), .B(n5348), .Z(n1513) );
  AND U4282 ( .A(n1556), .B(n1513), .Z(n1514) );
  NANDN U4283 ( .A(n1558), .B(n1514), .Z(n1515) );
  NAND U4284 ( .A(n1516), .B(n1515), .Z(n1517) );
  NANDN U4285 ( .A(n1557), .B(n1517), .Z(n1518) );
  ANDN U4286 ( .B(y[997]), .A(x[997]), .Z(n5360) );
  OR U4287 ( .A(n1518), .B(n5360), .Z(n1519) );
  NAND U4288 ( .A(n1549), .B(n1519), .Z(n1520) );
  NANDN U4289 ( .A(n5363), .B(n1520), .Z(n1521) );
  ANDN U4290 ( .B(y[999]), .A(x[999]), .Z(n1551) );
  OR U4291 ( .A(n1521), .B(n1551), .Z(n1522) );
  AND U4292 ( .A(n1553), .B(n1522), .Z(n1523) );
  NANDN U4293 ( .A(n1550), .B(n1523), .Z(n1524) );
  NAND U4294 ( .A(n1525), .B(n1524), .Z(n1526) );
  NAND U4295 ( .A(n1554), .B(n1526), .Z(n1527) );
  ANDN U4296 ( .B(x[1001]), .A(y[1001]), .Z(n1548) );
  OR U4297 ( .A(n1527), .B(n1548), .Z(n1528) );
  AND U4298 ( .A(n1547), .B(n1528), .Z(n1529) );
  ANDN U4299 ( .B(x[1004]), .A(y[1004]), .Z(n5367) );
  OR U4300 ( .A(n1529), .B(n5367), .Z(n1530) );
  AND U4301 ( .A(n1531), .B(n1530), .Z(n1533) );
  NANDN U4302 ( .A(y[1005]), .B(x[1005]), .Z(n5369) );
  ANDN U4303 ( .B(x[1006]), .A(y[1006]), .Z(n5370) );
  ANDN U4304 ( .B(n5369), .A(n5370), .Z(n1532) );
  NANDN U4305 ( .A(n1533), .B(n1532), .Z(n1534) );
  AND U4306 ( .A(n7329), .B(n1534), .Z(n1536) );
  OR U4307 ( .A(n1536), .B(n1535), .Z(n1539) );
  NANDN U4308 ( .A(x[1008]), .B(y[1008]), .Z(n1537) );
  NANDN U4309 ( .A(n1538), .B(n1537), .Z(n5375) );
  IV U4310 ( .A(n5375), .Z(n7331) );
  AND U4311 ( .A(n1539), .B(n7331), .Z(n1543) );
  ANDN U4312 ( .B(n1541), .A(n1540), .Z(n1542) );
  NANDN U4313 ( .A(n1543), .B(n1542), .Z(n1544) );
  AND U4314 ( .A(n1545), .B(n1544), .Z(n5377) );
  NAND U4315 ( .A(n1547), .B(n1546), .Z(n5358) );
  AND U4316 ( .A(n1556), .B(n1555), .Z(n1559) );
  AND U4317 ( .A(n1559), .B(n5352), .Z(n7323) );
  IV U4318 ( .A(n1560), .Z(n1561) );
  AND U4319 ( .A(n1562), .B(n1561), .Z(n1571) );
  NANDN U4320 ( .A(y[991]), .B(x[991]), .Z(n1565) );
  IV U4321 ( .A(n1563), .Z(n1564) );
  AND U4322 ( .A(n1565), .B(n1564), .Z(n1569) );
  AND U4323 ( .A(n1567), .B(n1566), .Z(n1575) );
  IV U4324 ( .A(n1575), .Z(n1568) );
  OR U4325 ( .A(n1569), .B(n1568), .Z(n1570) );
  AND U4326 ( .A(n1571), .B(n1570), .Z(n5391) );
  AND U4327 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U4328 ( .A(n1575), .B(n1574), .Z(n7322) );
  NANDN U4329 ( .A(y[989]), .B(x[989]), .Z(n1578) );
  IV U4330 ( .A(n1576), .Z(n1577) );
  AND U4331 ( .A(n1578), .B(n1577), .Z(n7321) );
  ANDN U4332 ( .B(x[982]), .A(y[982]), .Z(n5332) );
  NOR U4333 ( .A(n1582), .B(n1581), .Z(n5325) );
  NAND U4334 ( .A(n1584), .B(n1583), .Z(n7288) );
  IV U4335 ( .A(n1585), .Z(n1586) );
  AND U4336 ( .A(n1587), .B(n1586), .Z(n7286) );
  AND U4337 ( .A(n7281), .B(n7284), .Z(n5300) );
  IV U4338 ( .A(n1598), .Z(n1599) );
  AND U4339 ( .A(n1600), .B(n1599), .Z(n7275) );
  IV U4340 ( .A(n1601), .Z(n1602) );
  AND U4341 ( .A(n1603), .B(n1602), .Z(n7274) );
  IV U4342 ( .A(n1604), .Z(n1605) );
  AND U4343 ( .A(n1606), .B(n1605), .Z(n7273) );
  IV U4344 ( .A(n1607), .Z(n1608) );
  AND U4345 ( .A(n1609), .B(n1608), .Z(n7272) );
  AND U4346 ( .A(n1611), .B(n1610), .Z(n7269) );
  AND U4347 ( .A(n1615), .B(n1614), .Z(n5398) );
  AND U4348 ( .A(n7260), .B(n5398), .Z(n5276) );
  IV U4349 ( .A(n1616), .Z(n7247) );
  IV U4350 ( .A(n1617), .Z(n7244) );
  AND U4351 ( .A(n1618), .B(n7244), .Z(n5255) );
  NAND U4352 ( .A(n1620), .B(n1619), .Z(n7239) );
  IV U4353 ( .A(n1621), .Z(n7237) );
  NAND U4354 ( .A(n1625), .B(n1624), .Z(n7234) );
  NANDN U4355 ( .A(y[934]), .B(x[934]), .Z(n5228) );
  NAND U4356 ( .A(n1627), .B(n1626), .Z(n7225) );
  IV U4357 ( .A(n1632), .Z(n1634) );
  ANDN U4358 ( .B(n1634), .A(n1633), .Z(n7221) );
  AND U4359 ( .A(n1636), .B(n1635), .Z(n7220) );
  IV U4360 ( .A(n1637), .Z(n1639) );
  NAND U4361 ( .A(n1639), .B(n1638), .Z(n7219) );
  NANDN U4362 ( .A(n1641), .B(n1640), .Z(n1644) );
  IV U4363 ( .A(n1642), .Z(n1643) );
  AND U4364 ( .A(n1644), .B(n1643), .Z(n7217) );
  NAND U4365 ( .A(n1646), .B(n1645), .Z(n7216) );
  IV U4366 ( .A(n1647), .Z(n1648) );
  AND U4367 ( .A(n1649), .B(n1648), .Z(n7215) );
  AND U4368 ( .A(n1651), .B(n1650), .Z(n5406) );
  AND U4369 ( .A(n1661), .B(n1660), .Z(n7191) );
  IV U4370 ( .A(n1664), .Z(n1665) );
  AND U4371 ( .A(n1666), .B(n1665), .Z(n7187) );
  NANDN U4372 ( .A(y[902]), .B(x[902]), .Z(n5166) );
  AND U4373 ( .A(n1668), .B(n1667), .Z(n5163) );
  IV U4374 ( .A(n1669), .Z(n1671) );
  NAND U4375 ( .A(n1671), .B(n1670), .Z(n5407) );
  NAND U4376 ( .A(n1673), .B(n1672), .Z(n7165) );
  AND U4377 ( .A(n1675), .B(n1674), .Z(n7159) );
  NAND U4378 ( .A(n1679), .B(n1678), .Z(n7153) );
  IV U4379 ( .A(n1686), .Z(n7146) );
  AND U4380 ( .A(n1687), .B(n7146), .Z(n5138) );
  IV U4381 ( .A(n1688), .Z(n7143) );
  NANDN U4382 ( .A(y[886]), .B(x[886]), .Z(n5135) );
  AND U4383 ( .A(n1690), .B(n1689), .Z(n5129) );
  IV U4384 ( .A(n1691), .Z(n7130) );
  NANDN U4385 ( .A(y[880]), .B(x[880]), .Z(n1693) );
  NAND U4386 ( .A(n1693), .B(n1692), .Z(n5412) );
  AND U4387 ( .A(n1694), .B(n7126), .Z(n5116) );
  IV U4388 ( .A(n1703), .Z(n1705) );
  NAND U4389 ( .A(n1705), .B(n1704), .Z(n7114) );
  NAND U4390 ( .A(n1709), .B(n1708), .Z(n7110) );
  IV U4391 ( .A(n1710), .Z(n7108) );
  AND U4392 ( .A(n1711), .B(n7108), .Z(n5107) );
  AND U4393 ( .A(n1713), .B(n1712), .Z(n5101) );
  NAND U4394 ( .A(n1715), .B(n1714), .Z(n5415) );
  NAND U4395 ( .A(n1717), .B(n1716), .Z(n7091) );
  IV U4396 ( .A(n1718), .Z(n7088) );
  AND U4397 ( .A(n1720), .B(n1719), .Z(n7084) );
  NAND U4398 ( .A(n1722), .B(n1721), .Z(n7082) );
  AND U4399 ( .A(n1726), .B(n1725), .Z(n5420) );
  AND U4400 ( .A(n1729), .B(n7069), .Z(n5071) );
  AND U4401 ( .A(n1731), .B(n1730), .Z(n7065) );
  NAND U4402 ( .A(n1733), .B(n1732), .Z(n5421) );
  NAND U4403 ( .A(n1735), .B(n1734), .Z(n7063) );
  AND U4404 ( .A(n1737), .B(n1736), .Z(n7062) );
  AND U4405 ( .A(n1744), .B(n1743), .Z(n7058) );
  IV U4406 ( .A(n1750), .Z(n1752) );
  NANDN U4407 ( .A(n1752), .B(n1751), .Z(n1755) );
  IV U4408 ( .A(n1753), .Z(n1754) );
  AND U4409 ( .A(n1755), .B(n1754), .Z(n7043) );
  NAND U4410 ( .A(n1757), .B(n1756), .Z(n5422) );
  NANDN U4411 ( .A(y[828]), .B(x[828]), .Z(n1760) );
  IV U4412 ( .A(n1758), .Z(n1759) );
  AND U4413 ( .A(n1760), .B(n1759), .Z(n7042) );
  NAND U4414 ( .A(n1764), .B(n1763), .Z(n7040) );
  IV U4415 ( .A(n1765), .Z(n1766) );
  AND U4416 ( .A(n1767), .B(n1766), .Z(n7039) );
  NOR U4417 ( .A(n1769), .B(n1768), .Z(n5011) );
  ANDN U4418 ( .B(x[818]), .A(y[818]), .Z(n5001) );
  ANDN U4419 ( .B(x[816]), .A(y[816]), .Z(n4993) );
  ANDN U4420 ( .B(x[814]), .A(y[814]), .Z(n1771) );
  NOR U4421 ( .A(n1771), .B(n1770), .Z(n4985) );
  NANDN U4422 ( .A(y[810]), .B(x[810]), .Z(n1773) );
  AND U4423 ( .A(n1773), .B(n1772), .Z(n4971) );
  NOR U4424 ( .A(n1775), .B(n1774), .Z(n4945) );
  ANDN U4425 ( .B(x[802]), .A(y[802]), .Z(n4941) );
  NANDN U4426 ( .A(y[796]), .B(x[796]), .Z(n4919) );
  NOR U4427 ( .A(n1777), .B(n1776), .Z(n4915) );
  NANDN U4428 ( .A(y[788]), .B(x[788]), .Z(n4889) );
  NOR U4429 ( .A(n1779), .B(n1778), .Z(n4885) );
  NANDN U4430 ( .A(y[780]), .B(x[780]), .Z(n4859) );
  NOR U4431 ( .A(n1781), .B(n1780), .Z(n4855) );
  ANDN U4432 ( .B(x[778]), .A(y[778]), .Z(n4851) );
  ANDN U4433 ( .B(x[774]), .A(y[774]), .Z(n4837) );
  ANDN U4434 ( .B(x[772]), .A(y[772]), .Z(n1783) );
  NOR U4435 ( .A(n1783), .B(n1782), .Z(n4829) );
  AND U4436 ( .A(n1785), .B(n1784), .Z(n4815) );
  ANDN U4437 ( .B(x[764]), .A(y[764]), .Z(n1786) );
  NOR U4438 ( .A(n1787), .B(n1786), .Z(n4801) );
  NANDN U4439 ( .A(y[762]), .B(x[762]), .Z(n4795) );
  NAND U4440 ( .A(n1789), .B(n1788), .Z(n4783) );
  AND U4441 ( .A(n1791), .B(n1790), .Z(n4769) );
  ANDN U4442 ( .B(x[754]), .A(y[754]), .Z(n4767) );
  NANDN U4443 ( .A(y[752]), .B(x[752]), .Z(n4759) );
  AND U4444 ( .A(n1793), .B(n1792), .Z(n4755) );
  ANDN U4445 ( .B(x[750]), .A(y[750]), .Z(n4753) );
  NOR U4446 ( .A(n1795), .B(n1794), .Z(n4741) );
  ANDN U4447 ( .B(x[744]), .A(y[744]), .Z(n4731) );
  NAND U4448 ( .A(n1797), .B(n1796), .Z(n4715) );
  AND U4449 ( .A(n1799), .B(n1798), .Z(n4713) );
  NAND U4450 ( .A(n1801), .B(n1800), .Z(n4703) );
  AND U4451 ( .A(n1803), .B(n1802), .Z(n4701) );
  AND U4452 ( .A(n1805), .B(n1804), .Z(n4691) );
  NANDN U4453 ( .A(y[730]), .B(x[730]), .Z(n4685) );
  AND U4454 ( .A(n1807), .B(n1806), .Z(n4669) );
  NANDN U4455 ( .A(y[722]), .B(x[722]), .Z(n4656) );
  NAND U4456 ( .A(n1809), .B(n1808), .Z(n4628) );
  ANDN U4457 ( .B(x[712]), .A(y[712]), .Z(n4618) );
  NOR U4458 ( .A(n1811), .B(n1810), .Z(n4610) );
  AND U4459 ( .A(n1813), .B(n1812), .Z(n4584) );
  ANDN U4460 ( .B(x[702]), .A(y[702]), .Z(n4582) );
  NAND U4461 ( .A(n1815), .B(n1814), .Z(n4570) );
  AND U4462 ( .A(n1817), .B(n1816), .Z(n4568) );
  NAND U4463 ( .A(n1819), .B(n1818), .Z(n4558) );
  AND U4464 ( .A(n1821), .B(n1820), .Z(n4556) );
  XNOR U4465 ( .A(x[690]), .B(y[690]), .Z(n4538) );
  AND U4466 ( .A(n1823), .B(n1822), .Z(n4530) );
  ANDN U4467 ( .B(x[682]), .A(y[682]), .Z(n4512) );
  NANDN U4468 ( .A(y[680]), .B(x[680]), .Z(n1825) );
  AND U4469 ( .A(n1825), .B(n1824), .Z(n4504) );
  ANDN U4470 ( .B(x[676]), .A(y[676]), .Z(n4490) );
  NANDN U4471 ( .A(y[674]), .B(x[674]), .Z(n1827) );
  AND U4472 ( .A(n1827), .B(n1826), .Z(n4482) );
  ANDN U4473 ( .B(x[672]), .A(y[672]), .Z(n4476) );
  NAND U4474 ( .A(n1829), .B(n1828), .Z(n4468) );
  AND U4475 ( .A(n1831), .B(n1830), .Z(n4466) );
  ANDN U4476 ( .B(x[666]), .A(y[666]), .Z(n1833) );
  NOR U4477 ( .A(n1833), .B(n1832), .Z(n4456) );
  AND U4478 ( .A(n1835), .B(n1834), .Z(n4442) );
  AND U4479 ( .A(n1838), .B(n6707), .Z(n4418) );
  AND U4480 ( .A(n1840), .B(n1839), .Z(n4381) );
  AND U4481 ( .A(n1842), .B(n1841), .Z(n4359) );
  AND U4482 ( .A(n1844), .B(n1843), .Z(n4337) );
  NANDN U4483 ( .A(y[630]), .B(x[630]), .Z(n4331) );
  NANDN U4484 ( .A(y[626]), .B(x[626]), .Z(n1846) );
  AND U4485 ( .A(n1846), .B(n1845), .Z(n4315) );
  AND U4486 ( .A(n1848), .B(n1847), .Z(n4293) );
  AND U4487 ( .A(n1850), .B(n1849), .Z(n4271) );
  NANDN U4488 ( .A(y[608]), .B(x[608]), .Z(n1852) );
  AND U4489 ( .A(n1852), .B(n1851), .Z(n4249) );
  AND U4490 ( .A(n1854), .B(n1853), .Z(n4227) );
  AND U4491 ( .A(n1856), .B(n1855), .Z(n4205) );
  AND U4492 ( .A(n1858), .B(n1857), .Z(n4183) );
  NANDN U4493 ( .A(y[584]), .B(x[584]), .Z(n1860) );
  AND U4494 ( .A(n1860), .B(n1859), .Z(n4161) );
  AND U4495 ( .A(n1862), .B(n1861), .Z(n4139) );
  AND U4496 ( .A(n1864), .B(n1863), .Z(n4091) );
  NANDN U4497 ( .A(y[562]), .B(x[562]), .Z(n4085) );
  AND U4498 ( .A(n1866), .B(n1865), .Z(n4069) );
  AND U4499 ( .A(n1868), .B(n1867), .Z(n4047) );
  NANDN U4500 ( .A(y[550]), .B(x[550]), .Z(n4041) );
  AND U4501 ( .A(n1870), .B(n1869), .Z(n4025) );
  AND U4502 ( .A(n1872), .B(n1871), .Z(n4003) );
  NANDN U4503 ( .A(y[538]), .B(x[538]), .Z(n3997) );
  AND U4504 ( .A(n1874), .B(n1873), .Z(n3981) );
  NANDN U4505 ( .A(y[532]), .B(x[532]), .Z(n3975) );
  NANDN U4506 ( .A(y[528]), .B(x[528]), .Z(n1876) );
  AND U4507 ( .A(n1876), .B(n1875), .Z(n3959) );
  AND U4508 ( .A(n1878), .B(n1877), .Z(n3937) );
  AND U4509 ( .A(n1880), .B(n1879), .Z(n3915) );
  NANDN U4510 ( .A(y[514]), .B(x[514]), .Z(n3909) );
  AND U4511 ( .A(n1882), .B(n1881), .Z(n3893) );
  NANDN U4512 ( .A(y[508]), .B(x[508]), .Z(n3887) );
  AND U4513 ( .A(n1884), .B(n1883), .Z(n3871) );
  AND U4514 ( .A(n1886), .B(n1885), .Z(n3849) );
  NANDN U4515 ( .A(y[496]), .B(x[496]), .Z(n3843) );
  AND U4516 ( .A(n1888), .B(n1887), .Z(n3827) );
  NANDN U4517 ( .A(y[490]), .B(x[490]), .Z(n3821) );
  NANDN U4518 ( .A(y[486]), .B(x[486]), .Z(n1890) );
  AND U4519 ( .A(n1890), .B(n1889), .Z(n3805) );
  NANDN U4520 ( .A(y[480]), .B(x[480]), .Z(n1892) );
  AND U4521 ( .A(n1892), .B(n1891), .Z(n3783) );
  NANDN U4522 ( .A(y[474]), .B(x[474]), .Z(n1894) );
  AND U4523 ( .A(n1894), .B(n1893), .Z(n3761) );
  NANDN U4524 ( .A(y[468]), .B(x[468]), .Z(n1896) );
  AND U4525 ( .A(n1896), .B(n1895), .Z(n3739) );
  NANDN U4526 ( .A(y[462]), .B(x[462]), .Z(n1898) );
  AND U4527 ( .A(n1898), .B(n1897), .Z(n3717) );
  AND U4528 ( .A(n1900), .B(n1899), .Z(n3695) );
  AND U4529 ( .A(n1902), .B(n1901), .Z(n3673) );
  AND U4530 ( .A(n1904), .B(n1903), .Z(n3651) );
  NANDN U4531 ( .A(y[442]), .B(x[442]), .Z(n3645) );
  AND U4532 ( .A(n1906), .B(n1905), .Z(n3629) );
  NANDN U4533 ( .A(y[436]), .B(x[436]), .Z(n3623) );
  AND U4534 ( .A(n1908), .B(n1907), .Z(n3607) );
  AND U4535 ( .A(n1910), .B(n1909), .Z(n3585) );
  AND U4536 ( .A(n1912), .B(n1911), .Z(n3563) );
  NANDN U4537 ( .A(y[418]), .B(x[418]), .Z(n3557) );
  AND U4538 ( .A(n1914), .B(n1913), .Z(n3541) );
  AND U4539 ( .A(n1916), .B(n1915), .Z(n3519) );
  NANDN U4540 ( .A(y[406]), .B(x[406]), .Z(n3513) );
  NANDN U4541 ( .A(y[402]), .B(x[402]), .Z(n1918) );
  AND U4542 ( .A(n1918), .B(n1917), .Z(n3497) );
  AND U4543 ( .A(n1920), .B(n1919), .Z(n3475) );
  NANDN U4544 ( .A(y[394]), .B(x[394]), .Z(n3469) );
  AND U4545 ( .A(n1922), .B(n1921), .Z(n3453) );
  AND U4546 ( .A(n1924), .B(n1923), .Z(n3431) );
  NANDN U4547 ( .A(y[382]), .B(x[382]), .Z(n3425) );
  NANDN U4548 ( .A(y[378]), .B(x[378]), .Z(n1926) );
  AND U4549 ( .A(n1926), .B(n1925), .Z(n3409) );
  NANDN U4550 ( .A(y[372]), .B(x[372]), .Z(n1928) );
  AND U4551 ( .A(n1928), .B(n1927), .Z(n3387) );
  AND U4552 ( .A(n1930), .B(n1929), .Z(n3365) );
  NANDN U4553 ( .A(y[364]), .B(x[364]), .Z(n3359) );
  AND U4554 ( .A(n1932), .B(n1931), .Z(n3343) );
  NANDN U4555 ( .A(y[358]), .B(x[358]), .Z(n3337) );
  NANDN U4556 ( .A(y[354]), .B(x[354]), .Z(n1934) );
  AND U4557 ( .A(n1934), .B(n1933), .Z(n3321) );
  NANDN U4558 ( .A(y[348]), .B(x[348]), .Z(n1936) );
  AND U4559 ( .A(n1936), .B(n1935), .Z(n3299) );
  AND U4560 ( .A(n1938), .B(n1937), .Z(n3277) );
  AND U4561 ( .A(n1940), .B(n1939), .Z(n3255) );
  NANDN U4562 ( .A(y[330]), .B(x[330]), .Z(n1942) );
  AND U4563 ( .A(n1942), .B(n1941), .Z(n3233) );
  AND U4564 ( .A(n1944), .B(n1943), .Z(n3211) );
  AND U4565 ( .A(n1946), .B(n1945), .Z(n3189) );
  NANDN U4566 ( .A(y[312]), .B(x[312]), .Z(n1948) );
  AND U4567 ( .A(n1948), .B(n1947), .Z(n3167) );
  AND U4568 ( .A(n1950), .B(n1949), .Z(n3145) );
  NANDN U4569 ( .A(y[288]), .B(x[288]), .Z(n1952) );
  AND U4570 ( .A(n1952), .B(n1951), .Z(n3078) );
  AND U4571 ( .A(n1954), .B(n1953), .Z(n3056) );
  AND U4572 ( .A(n1956), .B(n1955), .Z(n3034) );
  AND U4573 ( .A(n1958), .B(n1957), .Z(n3012) );
  AND U4574 ( .A(n1960), .B(n1959), .Z(n2990) );
  AND U4575 ( .A(n1962), .B(n1961), .Z(n2968) );
  AND U4576 ( .A(n1964), .B(n1963), .Z(n2946) );
  NANDN U4577 ( .A(y[250]), .B(x[250]), .Z(n2940) );
  AND U4578 ( .A(n1966), .B(n1965), .Z(n2924) );
  AND U4579 ( .A(n1968), .B(n1967), .Z(n2902) );
  AND U4580 ( .A(n1970), .B(n1969), .Z(n2880) );
  NANDN U4581 ( .A(y[228]), .B(x[228]), .Z(n1972) );
  AND U4582 ( .A(n1972), .B(n1971), .Z(n2858) );
  AND U4583 ( .A(n1974), .B(n1973), .Z(n2836) );
  NANDN U4584 ( .A(y[220]), .B(x[220]), .Z(n2830) );
  AND U4585 ( .A(n1976), .B(n1975), .Z(n2814) );
  AND U4586 ( .A(n1978), .B(n1977), .Z(n2792) );
  NANDN U4587 ( .A(y[208]), .B(x[208]), .Z(n2786) );
  AND U4588 ( .A(n1980), .B(n1979), .Z(n2770) );
  AND U4589 ( .A(n1982), .B(n1981), .Z(n2748) );
  AND U4590 ( .A(n1984), .B(n1983), .Z(n2726) );
  AND U4591 ( .A(n1986), .B(n1985), .Z(n2704) );
  NANDN U4592 ( .A(y[184]), .B(x[184]), .Z(n2698) );
  AND U4593 ( .A(n1988), .B(n1987), .Z(n2682) );
  AND U4594 ( .A(n1990), .B(n1989), .Z(n2660) );
  NANDN U4595 ( .A(y[168]), .B(x[168]), .Z(n1992) );
  AND U4596 ( .A(n1992), .B(n1991), .Z(n2638) );
  NANDN U4597 ( .A(y[162]), .B(x[162]), .Z(n1994) );
  AND U4598 ( .A(n1994), .B(n1993), .Z(n2616) );
  AND U4599 ( .A(n1996), .B(n1995), .Z(n2594) );
  AND U4600 ( .A(n1998), .B(n1997), .Z(n2572) );
  AND U4601 ( .A(n2000), .B(n1999), .Z(n2550) );
  AND U4602 ( .A(n2002), .B(n2001), .Z(n2528) );
  AND U4603 ( .A(n2004), .B(n2003), .Z(n2506) );
  AND U4604 ( .A(n2006), .B(n2005), .Z(n2484) );
  AND U4605 ( .A(n2008), .B(n2007), .Z(n2462) );
  NANDN U4606 ( .A(y[114]), .B(x[114]), .Z(n2010) );
  AND U4607 ( .A(n2010), .B(n2009), .Z(n2440) );
  AND U4608 ( .A(n2012), .B(n2011), .Z(n2418) );
  NANDN U4609 ( .A(y[106]), .B(x[106]), .Z(n2412) );
  AND U4610 ( .A(n2014), .B(n2013), .Z(n2396) );
  NANDN U4611 ( .A(y[100]), .B(x[100]), .Z(n2390) );
  AND U4612 ( .A(n2016), .B(n2015), .Z(n2374) );
  NANDN U4613 ( .A(y[90]), .B(x[90]), .Z(n2018) );
  AND U4614 ( .A(n2018), .B(n2017), .Z(n2352) );
  AND U4615 ( .A(n2020), .B(n2019), .Z(n2330) );
  AND U4616 ( .A(n2022), .B(n2021), .Z(n2308) );
  AND U4617 ( .A(n2024), .B(n2023), .Z(n2286) );
  AND U4618 ( .A(n2026), .B(n2025), .Z(n2264) );
  AND U4619 ( .A(n2028), .B(n2027), .Z(n2242) );
  AND U4620 ( .A(n2030), .B(n2029), .Z(n2220) );
  AND U4621 ( .A(n2032), .B(n2031), .Z(n2198) );
  AND U4622 ( .A(n2034), .B(n2033), .Z(n2176) );
  AND U4623 ( .A(n2036), .B(n2035), .Z(n2154) );
  AND U4624 ( .A(n2038), .B(n2037), .Z(n2132) );
  AND U4625 ( .A(n2040), .B(n2039), .Z(n2110) );
  AND U4626 ( .A(n2042), .B(n2041), .Z(n2088) );
  AND U4627 ( .A(n2044), .B(n2043), .Z(n2066) );
  NANDN U4628 ( .A(y[0]), .B(x[0]), .Z(n2052) );
  OR U4629 ( .A(n5427), .B(n2058), .Z(n2059) );
  NAND U4630 ( .A(n2060), .B(n2059), .Z(n2061) );
  NANDN U4631 ( .A(n2062), .B(n2061), .Z(n2064) );
  OR U4632 ( .A(n2064), .B(n2063), .Z(n2065) );
  AND U4633 ( .A(n2066), .B(n2065), .Z(n2068) );
  NOR U4634 ( .A(n2068), .B(n2067), .Z(n2069) );
  NANDN U4635 ( .A(n2070), .B(n2069), .Z(n2071) );
  AND U4636 ( .A(n2072), .B(n2071), .Z(n2074) );
  NAND U4637 ( .A(n2074), .B(n2073), .Z(n2076) );
  ANDN U4638 ( .B(n2076), .A(n2075), .Z(n2077) );
  NANDN U4639 ( .A(n2078), .B(n2077), .Z(n2082) );
  AND U4640 ( .A(n2080), .B(n2079), .Z(n2081) );
  NAND U4641 ( .A(n2082), .B(n2081), .Z(n2083) );
  NANDN U4642 ( .A(n2084), .B(n2083), .Z(n2086) );
  OR U4643 ( .A(n2086), .B(n2085), .Z(n2087) );
  AND U4644 ( .A(n2088), .B(n2087), .Z(n2090) );
  NOR U4645 ( .A(n2090), .B(n2089), .Z(n2091) );
  NANDN U4646 ( .A(n2092), .B(n2091), .Z(n2093) );
  AND U4647 ( .A(n2094), .B(n2093), .Z(n2096) );
  NAND U4648 ( .A(n2096), .B(n2095), .Z(n2098) );
  ANDN U4649 ( .B(n2098), .A(n2097), .Z(n2099) );
  NANDN U4650 ( .A(n2100), .B(n2099), .Z(n2104) );
  AND U4651 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U4652 ( .A(n2104), .B(n2103), .Z(n2105) );
  NANDN U4653 ( .A(n2106), .B(n2105), .Z(n2108) );
  OR U4654 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U4655 ( .A(n2110), .B(n2109), .Z(n2112) );
  NOR U4656 ( .A(n2112), .B(n2111), .Z(n2113) );
  NANDN U4657 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U4658 ( .A(n2116), .B(n2115), .Z(n2118) );
  NAND U4659 ( .A(n2118), .B(n2117), .Z(n2120) );
  ANDN U4660 ( .B(n2120), .A(n2119), .Z(n2121) );
  NANDN U4661 ( .A(n2122), .B(n2121), .Z(n2126) );
  AND U4662 ( .A(n2124), .B(n2123), .Z(n2125) );
  NAND U4663 ( .A(n2126), .B(n2125), .Z(n2127) );
  NANDN U4664 ( .A(n2128), .B(n2127), .Z(n2130) );
  OR U4665 ( .A(n2130), .B(n2129), .Z(n2131) );
  AND U4666 ( .A(n2132), .B(n2131), .Z(n2134) );
  NOR U4667 ( .A(n2134), .B(n2133), .Z(n2135) );
  NANDN U4668 ( .A(n2136), .B(n2135), .Z(n2137) );
  AND U4669 ( .A(n2138), .B(n2137), .Z(n2140) );
  NAND U4670 ( .A(n2140), .B(n2139), .Z(n2142) );
  ANDN U4671 ( .B(n2142), .A(n2141), .Z(n2143) );
  NANDN U4672 ( .A(n2144), .B(n2143), .Z(n2148) );
  AND U4673 ( .A(n2146), .B(n2145), .Z(n2147) );
  NAND U4674 ( .A(n2148), .B(n2147), .Z(n2149) );
  NANDN U4675 ( .A(n2150), .B(n2149), .Z(n2152) );
  OR U4676 ( .A(n2152), .B(n2151), .Z(n2153) );
  AND U4677 ( .A(n2154), .B(n2153), .Z(n2156) );
  NOR U4678 ( .A(n2156), .B(n2155), .Z(n2157) );
  NANDN U4679 ( .A(n2158), .B(n2157), .Z(n2159) );
  AND U4680 ( .A(n2160), .B(n2159), .Z(n2162) );
  NAND U4681 ( .A(n2162), .B(n2161), .Z(n2164) );
  ANDN U4682 ( .B(n2164), .A(n2163), .Z(n2165) );
  NANDN U4683 ( .A(n2166), .B(n2165), .Z(n2170) );
  AND U4684 ( .A(n2168), .B(n2167), .Z(n2169) );
  NAND U4685 ( .A(n2170), .B(n2169), .Z(n2171) );
  NANDN U4686 ( .A(n2172), .B(n2171), .Z(n2174) );
  OR U4687 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U4688 ( .A(n2176), .B(n2175), .Z(n2178) );
  NOR U4689 ( .A(n2178), .B(n2177), .Z(n2179) );
  NANDN U4690 ( .A(n2180), .B(n2179), .Z(n2181) );
  AND U4691 ( .A(n2182), .B(n2181), .Z(n2184) );
  NAND U4692 ( .A(n2184), .B(n2183), .Z(n2186) );
  ANDN U4693 ( .B(n2186), .A(n2185), .Z(n2187) );
  NANDN U4694 ( .A(n2188), .B(n2187), .Z(n2192) );
  AND U4695 ( .A(n2190), .B(n2189), .Z(n2191) );
  NAND U4696 ( .A(n2192), .B(n2191), .Z(n2193) );
  NANDN U4697 ( .A(n2194), .B(n2193), .Z(n2196) );
  OR U4698 ( .A(n2196), .B(n2195), .Z(n2197) );
  AND U4699 ( .A(n2198), .B(n2197), .Z(n2200) );
  NOR U4700 ( .A(n2200), .B(n2199), .Z(n2201) );
  NANDN U4701 ( .A(n2202), .B(n2201), .Z(n2203) );
  AND U4702 ( .A(n2204), .B(n2203), .Z(n2206) );
  NAND U4703 ( .A(n2206), .B(n2205), .Z(n2208) );
  ANDN U4704 ( .B(n2208), .A(n2207), .Z(n2209) );
  NANDN U4705 ( .A(n2210), .B(n2209), .Z(n2214) );
  AND U4706 ( .A(n2212), .B(n2211), .Z(n2213) );
  NAND U4707 ( .A(n2214), .B(n2213), .Z(n2215) );
  NANDN U4708 ( .A(n2216), .B(n2215), .Z(n2218) );
  OR U4709 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U4710 ( .A(n2220), .B(n2219), .Z(n2222) );
  NOR U4711 ( .A(n2222), .B(n2221), .Z(n2223) );
  NANDN U4712 ( .A(n2224), .B(n2223), .Z(n2225) );
  AND U4713 ( .A(n2226), .B(n2225), .Z(n2228) );
  NAND U4714 ( .A(n2228), .B(n2227), .Z(n2230) );
  ANDN U4715 ( .B(n2230), .A(n2229), .Z(n2231) );
  NANDN U4716 ( .A(n2232), .B(n2231), .Z(n2236) );
  AND U4717 ( .A(n2234), .B(n2233), .Z(n2235) );
  NAND U4718 ( .A(n2236), .B(n2235), .Z(n2237) );
  NANDN U4719 ( .A(n2238), .B(n2237), .Z(n2240) );
  OR U4720 ( .A(n2240), .B(n2239), .Z(n2241) );
  AND U4721 ( .A(n2242), .B(n2241), .Z(n2244) );
  NOR U4722 ( .A(n2244), .B(n2243), .Z(n2245) );
  NANDN U4723 ( .A(n2246), .B(n2245), .Z(n2247) );
  AND U4724 ( .A(n2248), .B(n2247), .Z(n2250) );
  NAND U4725 ( .A(n2250), .B(n2249), .Z(n2252) );
  ANDN U4726 ( .B(n2252), .A(n2251), .Z(n2253) );
  NANDN U4727 ( .A(n2254), .B(n2253), .Z(n2258) );
  AND U4728 ( .A(n2256), .B(n2255), .Z(n2257) );
  NAND U4729 ( .A(n2258), .B(n2257), .Z(n2259) );
  NANDN U4730 ( .A(n2260), .B(n2259), .Z(n2262) );
  OR U4731 ( .A(n2262), .B(n2261), .Z(n2263) );
  AND U4732 ( .A(n2264), .B(n2263), .Z(n2266) );
  NOR U4733 ( .A(n2266), .B(n2265), .Z(n2267) );
  NANDN U4734 ( .A(n2268), .B(n2267), .Z(n2269) );
  AND U4735 ( .A(n2270), .B(n2269), .Z(n2272) );
  NAND U4736 ( .A(n2272), .B(n2271), .Z(n2274) );
  ANDN U4737 ( .B(n2274), .A(n2273), .Z(n2275) );
  NANDN U4738 ( .A(n2276), .B(n2275), .Z(n2280) );
  AND U4739 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U4740 ( .A(n2280), .B(n2279), .Z(n2281) );
  NANDN U4741 ( .A(n2282), .B(n2281), .Z(n2284) );
  OR U4742 ( .A(n2284), .B(n2283), .Z(n2285) );
  AND U4743 ( .A(n2286), .B(n2285), .Z(n2288) );
  NOR U4744 ( .A(n2288), .B(n2287), .Z(n2289) );
  NANDN U4745 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U4746 ( .A(n2292), .B(n2291), .Z(n2294) );
  NAND U4747 ( .A(n2294), .B(n2293), .Z(n2296) );
  ANDN U4748 ( .B(n2296), .A(n2295), .Z(n2297) );
  NANDN U4749 ( .A(n2298), .B(n2297), .Z(n2302) );
  AND U4750 ( .A(n2300), .B(n2299), .Z(n2301) );
  NAND U4751 ( .A(n2302), .B(n2301), .Z(n2303) );
  NANDN U4752 ( .A(n2304), .B(n2303), .Z(n2306) );
  OR U4753 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U4754 ( .A(n2308), .B(n2307), .Z(n2309) );
  NOR U4755 ( .A(n2310), .B(n2309), .Z(n2311) );
  NANDN U4756 ( .A(n2312), .B(n2311), .Z(n2313) );
  AND U4757 ( .A(n2314), .B(n2313), .Z(n2316) );
  NANDN U4758 ( .A(y[80]), .B(x[80]), .Z(n2315) );
  NAND U4759 ( .A(n2316), .B(n2315), .Z(n2318) );
  ANDN U4760 ( .B(n2318), .A(n2317), .Z(n2319) );
  NANDN U4761 ( .A(n2320), .B(n2319), .Z(n2324) );
  AND U4762 ( .A(n2322), .B(n2321), .Z(n2323) );
  NAND U4763 ( .A(n2324), .B(n2323), .Z(n2325) );
  NANDN U4764 ( .A(n2326), .B(n2325), .Z(n2328) );
  OR U4765 ( .A(n2328), .B(n2327), .Z(n2329) );
  AND U4766 ( .A(n2330), .B(n2329), .Z(n2331) );
  NOR U4767 ( .A(n2332), .B(n2331), .Z(n2333) );
  NANDN U4768 ( .A(n2334), .B(n2333), .Z(n2335) );
  AND U4769 ( .A(n2336), .B(n2335), .Z(n2338) );
  NANDN U4770 ( .A(y[86]), .B(x[86]), .Z(n2337) );
  NAND U4771 ( .A(n2338), .B(n2337), .Z(n2340) );
  ANDN U4772 ( .B(n2340), .A(n2339), .Z(n2341) );
  NANDN U4773 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U4774 ( .A(n2344), .B(n2343), .Z(n2345) );
  NAND U4775 ( .A(n2346), .B(n2345), .Z(n2347) );
  NANDN U4776 ( .A(n2348), .B(n2347), .Z(n2350) );
  OR U4777 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U4778 ( .A(n2352), .B(n2351), .Z(n2354) );
  NOR U4779 ( .A(n2354), .B(n2353), .Z(n2355) );
  NANDN U4780 ( .A(n2356), .B(n2355), .Z(n2357) );
  AND U4781 ( .A(n2358), .B(n2357), .Z(n2360) );
  NAND U4782 ( .A(n2360), .B(n2359), .Z(n2362) );
  ANDN U4783 ( .B(n2362), .A(n2361), .Z(n2363) );
  NANDN U4784 ( .A(n2364), .B(n2363), .Z(n2368) );
  AND U4785 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U4786 ( .A(n2368), .B(n2367), .Z(n2369) );
  NANDN U4787 ( .A(n2370), .B(n2369), .Z(n2372) );
  OR U4788 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U4789 ( .A(n2374), .B(n2373), .Z(n2376) );
  NOR U4790 ( .A(n2376), .B(n2375), .Z(n2377) );
  NANDN U4791 ( .A(n2378), .B(n2377), .Z(n2379) );
  AND U4792 ( .A(n2380), .B(n2379), .Z(n2382) );
  NAND U4793 ( .A(n2382), .B(n2381), .Z(n2384) );
  ANDN U4794 ( .B(n2384), .A(n2383), .Z(n2385) );
  NANDN U4795 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U4796 ( .A(n2388), .B(n2387), .Z(n2389) );
  NAND U4797 ( .A(n2390), .B(n2389), .Z(n2391) );
  NANDN U4798 ( .A(n2392), .B(n2391), .Z(n2394) );
  OR U4799 ( .A(n2394), .B(n2393), .Z(n2395) );
  AND U4800 ( .A(n2396), .B(n2395), .Z(n2397) );
  NOR U4801 ( .A(n2398), .B(n2397), .Z(n2399) );
  NANDN U4802 ( .A(n2400), .B(n2399), .Z(n2401) );
  AND U4803 ( .A(n2402), .B(n2401), .Z(n2404) );
  NANDN U4804 ( .A(y[104]), .B(x[104]), .Z(n2403) );
  NAND U4805 ( .A(n2404), .B(n2403), .Z(n2406) );
  ANDN U4806 ( .B(n2406), .A(n2405), .Z(n2407) );
  NANDN U4807 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U4808 ( .A(n2410), .B(n2409), .Z(n2411) );
  NAND U4809 ( .A(n2412), .B(n2411), .Z(n2413) );
  NANDN U4810 ( .A(n2414), .B(n2413), .Z(n2416) );
  OR U4811 ( .A(n2416), .B(n2415), .Z(n2417) );
  AND U4812 ( .A(n2418), .B(n2417), .Z(n2419) );
  NOR U4813 ( .A(n2420), .B(n2419), .Z(n2421) );
  NANDN U4814 ( .A(n2422), .B(n2421), .Z(n2423) );
  AND U4815 ( .A(n2424), .B(n2423), .Z(n2426) );
  NANDN U4816 ( .A(y[110]), .B(x[110]), .Z(n2425) );
  NAND U4817 ( .A(n2426), .B(n2425), .Z(n2428) );
  ANDN U4818 ( .B(n2428), .A(n2427), .Z(n2429) );
  NANDN U4819 ( .A(n2430), .B(n2429), .Z(n2431) );
  AND U4820 ( .A(n2432), .B(n2431), .Z(n2433) );
  NAND U4821 ( .A(n2434), .B(n2433), .Z(n2435) );
  NANDN U4822 ( .A(n2436), .B(n2435), .Z(n2438) );
  OR U4823 ( .A(n2438), .B(n2437), .Z(n2439) );
  AND U4824 ( .A(n2440), .B(n2439), .Z(n2442) );
  NOR U4825 ( .A(n2442), .B(n2441), .Z(n2443) );
  NANDN U4826 ( .A(n2444), .B(n2443), .Z(n2445) );
  AND U4827 ( .A(n2446), .B(n2445), .Z(n2448) );
  NAND U4828 ( .A(n2448), .B(n2447), .Z(n2450) );
  ANDN U4829 ( .B(n2450), .A(n2449), .Z(n2451) );
  NANDN U4830 ( .A(n2452), .B(n2451), .Z(n2456) );
  AND U4831 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U4832 ( .A(n2456), .B(n2455), .Z(n2457) );
  NANDN U4833 ( .A(n2458), .B(n2457), .Z(n2460) );
  OR U4834 ( .A(n2460), .B(n2459), .Z(n2461) );
  AND U4835 ( .A(n2462), .B(n2461), .Z(n2464) );
  NOR U4836 ( .A(n2464), .B(n2463), .Z(n2465) );
  NANDN U4837 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U4838 ( .A(n2468), .B(n2467), .Z(n2470) );
  NAND U4839 ( .A(n2470), .B(n2469), .Z(n2472) );
  ANDN U4840 ( .B(n2472), .A(n2471), .Z(n2473) );
  NANDN U4841 ( .A(n2474), .B(n2473), .Z(n2478) );
  AND U4842 ( .A(n2476), .B(n2475), .Z(n2477) );
  NAND U4843 ( .A(n2478), .B(n2477), .Z(n2479) );
  NANDN U4844 ( .A(n2480), .B(n2479), .Z(n2482) );
  OR U4845 ( .A(n2482), .B(n2481), .Z(n2483) );
  AND U4846 ( .A(n2484), .B(n2483), .Z(n2486) );
  NOR U4847 ( .A(n2486), .B(n2485), .Z(n2487) );
  NANDN U4848 ( .A(n2488), .B(n2487), .Z(n2489) );
  AND U4849 ( .A(n2490), .B(n2489), .Z(n2492) );
  NAND U4850 ( .A(n2492), .B(n2491), .Z(n2494) );
  ANDN U4851 ( .B(n2494), .A(n2493), .Z(n2495) );
  NANDN U4852 ( .A(n2496), .B(n2495), .Z(n2500) );
  AND U4853 ( .A(n2498), .B(n2497), .Z(n2499) );
  NAND U4854 ( .A(n2500), .B(n2499), .Z(n2501) );
  NANDN U4855 ( .A(n2502), .B(n2501), .Z(n2504) );
  OR U4856 ( .A(n2504), .B(n2503), .Z(n2505) );
  AND U4857 ( .A(n2506), .B(n2505), .Z(n2508) );
  NOR U4858 ( .A(n2508), .B(n2507), .Z(n2509) );
  NANDN U4859 ( .A(n2510), .B(n2509), .Z(n2511) );
  AND U4860 ( .A(n2512), .B(n2511), .Z(n2514) );
  NAND U4861 ( .A(n2514), .B(n2513), .Z(n2516) );
  ANDN U4862 ( .B(n2516), .A(n2515), .Z(n2517) );
  NANDN U4863 ( .A(n2518), .B(n2517), .Z(n2522) );
  AND U4864 ( .A(n2520), .B(n2519), .Z(n2521) );
  NAND U4865 ( .A(n2522), .B(n2521), .Z(n2523) );
  NANDN U4866 ( .A(n2524), .B(n2523), .Z(n2526) );
  OR U4867 ( .A(n2526), .B(n2525), .Z(n2527) );
  AND U4868 ( .A(n2528), .B(n2527), .Z(n2530) );
  NOR U4869 ( .A(n2530), .B(n2529), .Z(n2531) );
  NANDN U4870 ( .A(n2532), .B(n2531), .Z(n2533) );
  AND U4871 ( .A(n2534), .B(n2533), .Z(n2536) );
  NAND U4872 ( .A(n2536), .B(n2535), .Z(n2538) );
  ANDN U4873 ( .B(n2538), .A(n2537), .Z(n2539) );
  NANDN U4874 ( .A(n2540), .B(n2539), .Z(n2544) );
  AND U4875 ( .A(n2542), .B(n2541), .Z(n2543) );
  NAND U4876 ( .A(n2544), .B(n2543), .Z(n2545) );
  NANDN U4877 ( .A(n2546), .B(n2545), .Z(n2548) );
  OR U4878 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U4879 ( .A(n2550), .B(n2549), .Z(n2551) );
  NOR U4880 ( .A(n2552), .B(n2551), .Z(n2553) );
  NANDN U4881 ( .A(n2554), .B(n2553), .Z(n2555) );
  AND U4882 ( .A(n2556), .B(n2555), .Z(n2558) );
  NANDN U4883 ( .A(y[146]), .B(x[146]), .Z(n2557) );
  NAND U4884 ( .A(n2558), .B(n2557), .Z(n2560) );
  ANDN U4885 ( .B(n2560), .A(n2559), .Z(n2561) );
  NANDN U4886 ( .A(n2562), .B(n2561), .Z(n2566) );
  AND U4887 ( .A(n2564), .B(n2563), .Z(n2565) );
  NAND U4888 ( .A(n2566), .B(n2565), .Z(n2567) );
  NANDN U4889 ( .A(n2568), .B(n2567), .Z(n2570) );
  OR U4890 ( .A(n2570), .B(n2569), .Z(n2571) );
  AND U4891 ( .A(n2572), .B(n2571), .Z(n2574) );
  NOR U4892 ( .A(n2574), .B(n2573), .Z(n2575) );
  NANDN U4893 ( .A(n2576), .B(n2575), .Z(n2577) );
  AND U4894 ( .A(n2578), .B(n2577), .Z(n2580) );
  NAND U4895 ( .A(n2580), .B(n2579), .Z(n2582) );
  ANDN U4896 ( .B(n2582), .A(n2581), .Z(n2583) );
  NANDN U4897 ( .A(n2584), .B(n2583), .Z(n2588) );
  AND U4898 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U4899 ( .A(n2588), .B(n2587), .Z(n2589) );
  NANDN U4900 ( .A(n2590), .B(n2589), .Z(n2592) );
  OR U4901 ( .A(n2592), .B(n2591), .Z(n2593) );
  AND U4902 ( .A(n2594), .B(n2593), .Z(n2596) );
  NOR U4903 ( .A(n2596), .B(n2595), .Z(n2597) );
  NANDN U4904 ( .A(n2598), .B(n2597), .Z(n2599) );
  AND U4905 ( .A(n2600), .B(n2599), .Z(n2602) );
  NAND U4906 ( .A(n2602), .B(n2601), .Z(n2604) );
  ANDN U4907 ( .B(n2604), .A(n2603), .Z(n2605) );
  NANDN U4908 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U4909 ( .A(n2608), .B(n2607), .Z(n2609) );
  NAND U4910 ( .A(n2610), .B(n2609), .Z(n2611) );
  NANDN U4911 ( .A(n2612), .B(n2611), .Z(n2614) );
  OR U4912 ( .A(n2614), .B(n2613), .Z(n2615) );
  AND U4913 ( .A(n2616), .B(n2615), .Z(n2618) );
  NOR U4914 ( .A(n2618), .B(n2617), .Z(n2619) );
  NANDN U4915 ( .A(n2620), .B(n2619), .Z(n2621) );
  AND U4916 ( .A(n2622), .B(n2621), .Z(n2624) );
  NAND U4917 ( .A(n2624), .B(n2623), .Z(n2626) );
  ANDN U4918 ( .B(n2626), .A(n2625), .Z(n2627) );
  NANDN U4919 ( .A(n2628), .B(n2627), .Z(n2632) );
  NANDN U4920 ( .A(y[166]), .B(x[166]), .Z(n2629) );
  AND U4921 ( .A(n2630), .B(n2629), .Z(n2631) );
  NAND U4922 ( .A(n2632), .B(n2631), .Z(n2633) );
  NANDN U4923 ( .A(n2634), .B(n2633), .Z(n2636) );
  OR U4924 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U4925 ( .A(n2638), .B(n2637), .Z(n2639) );
  NOR U4926 ( .A(n2640), .B(n2639), .Z(n2641) );
  NANDN U4927 ( .A(n2642), .B(n2641), .Z(n2643) );
  AND U4928 ( .A(n2644), .B(n2643), .Z(n2646) );
  NANDN U4929 ( .A(y[170]), .B(x[170]), .Z(n2645) );
  NAND U4930 ( .A(n2646), .B(n2645), .Z(n2648) );
  ANDN U4931 ( .B(n2648), .A(n2647), .Z(n2649) );
  NANDN U4932 ( .A(n2650), .B(n2649), .Z(n2654) );
  AND U4933 ( .A(n2652), .B(n2651), .Z(n2653) );
  NAND U4934 ( .A(n2654), .B(n2653), .Z(n2655) );
  NANDN U4935 ( .A(n2656), .B(n2655), .Z(n2658) );
  OR U4936 ( .A(n2658), .B(n2657), .Z(n2659) );
  AND U4937 ( .A(n2660), .B(n2659), .Z(n2661) );
  NOR U4938 ( .A(n2662), .B(n2661), .Z(n2663) );
  NANDN U4939 ( .A(n2664), .B(n2663), .Z(n2665) );
  AND U4940 ( .A(n2666), .B(n2665), .Z(n2668) );
  NANDN U4941 ( .A(y[176]), .B(x[176]), .Z(n2667) );
  NAND U4942 ( .A(n2668), .B(n2667), .Z(n2670) );
  ANDN U4943 ( .B(n2670), .A(n2669), .Z(n2671) );
  NANDN U4944 ( .A(n2672), .B(n2671), .Z(n2676) );
  AND U4945 ( .A(n2674), .B(n2673), .Z(n2675) );
  NAND U4946 ( .A(n2676), .B(n2675), .Z(n2677) );
  NANDN U4947 ( .A(n2678), .B(n2677), .Z(n2680) );
  OR U4948 ( .A(n2680), .B(n2679), .Z(n2681) );
  AND U4949 ( .A(n2682), .B(n2681), .Z(n2684) );
  NOR U4950 ( .A(n2684), .B(n2683), .Z(n2685) );
  NANDN U4951 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U4952 ( .A(n2688), .B(n2687), .Z(n2690) );
  NAND U4953 ( .A(n2690), .B(n2689), .Z(n2692) );
  ANDN U4954 ( .B(n2692), .A(n2691), .Z(n2693) );
  NANDN U4955 ( .A(n2694), .B(n2693), .Z(n2695) );
  AND U4956 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U4957 ( .A(n2698), .B(n2697), .Z(n2699) );
  NANDN U4958 ( .A(n2700), .B(n2699), .Z(n2702) );
  OR U4959 ( .A(n2702), .B(n2701), .Z(n2703) );
  AND U4960 ( .A(n2704), .B(n2703), .Z(n2706) );
  NOR U4961 ( .A(n2706), .B(n2705), .Z(n2707) );
  NANDN U4962 ( .A(n2708), .B(n2707), .Z(n2709) );
  AND U4963 ( .A(n2710), .B(n2709), .Z(n2712) );
  NAND U4964 ( .A(n2712), .B(n2711), .Z(n2714) );
  ANDN U4965 ( .B(n2714), .A(n2713), .Z(n2715) );
  NANDN U4966 ( .A(n2716), .B(n2715), .Z(n2720) );
  AND U4967 ( .A(n2718), .B(n2717), .Z(n2719) );
  NAND U4968 ( .A(n2720), .B(n2719), .Z(n2721) );
  NANDN U4969 ( .A(n2722), .B(n2721), .Z(n2724) );
  OR U4970 ( .A(n2724), .B(n2723), .Z(n2725) );
  AND U4971 ( .A(n2726), .B(n2725), .Z(n2728) );
  NOR U4972 ( .A(n2728), .B(n2727), .Z(n2729) );
  NANDN U4973 ( .A(n2730), .B(n2729), .Z(n2731) );
  AND U4974 ( .A(n2732), .B(n2731), .Z(n2734) );
  NAND U4975 ( .A(n2734), .B(n2733), .Z(n2736) );
  ANDN U4976 ( .B(n2736), .A(n2735), .Z(n2737) );
  NANDN U4977 ( .A(n2738), .B(n2737), .Z(n2742) );
  AND U4978 ( .A(n2740), .B(n2739), .Z(n2741) );
  NAND U4979 ( .A(n2742), .B(n2741), .Z(n2743) );
  NANDN U4980 ( .A(n2744), .B(n2743), .Z(n2746) );
  OR U4981 ( .A(n2746), .B(n2745), .Z(n2747) );
  AND U4982 ( .A(n2748), .B(n2747), .Z(n2750) );
  NOR U4983 ( .A(n2750), .B(n2749), .Z(n2751) );
  NANDN U4984 ( .A(n2752), .B(n2751), .Z(n2753) );
  AND U4985 ( .A(n2754), .B(n2753), .Z(n2756) );
  NAND U4986 ( .A(n2756), .B(n2755), .Z(n2758) );
  ANDN U4987 ( .B(n2758), .A(n2757), .Z(n2759) );
  NANDN U4988 ( .A(n2760), .B(n2759), .Z(n2764) );
  AND U4989 ( .A(n2762), .B(n2761), .Z(n2763) );
  NAND U4990 ( .A(n2764), .B(n2763), .Z(n2765) );
  NANDN U4991 ( .A(n2766), .B(n2765), .Z(n2768) );
  OR U4992 ( .A(n2768), .B(n2767), .Z(n2769) );
  AND U4993 ( .A(n2770), .B(n2769), .Z(n2772) );
  NOR U4994 ( .A(n2772), .B(n2771), .Z(n2773) );
  NANDN U4995 ( .A(n2774), .B(n2773), .Z(n2775) );
  AND U4996 ( .A(n2776), .B(n2775), .Z(n2778) );
  NAND U4997 ( .A(n2778), .B(n2777), .Z(n2780) );
  ANDN U4998 ( .B(n2780), .A(n2779), .Z(n2781) );
  NANDN U4999 ( .A(n2782), .B(n2781), .Z(n2783) );
  AND U5000 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U5001 ( .A(n2786), .B(n2785), .Z(n2787) );
  NANDN U5002 ( .A(n2788), .B(n2787), .Z(n2790) );
  OR U5003 ( .A(n2790), .B(n2789), .Z(n2791) );
  AND U5004 ( .A(n2792), .B(n2791), .Z(n2794) );
  NOR U5005 ( .A(n2794), .B(n2793), .Z(n2795) );
  NANDN U5006 ( .A(n2796), .B(n2795), .Z(n2797) );
  AND U5007 ( .A(n2798), .B(n2797), .Z(n2800) );
  NAND U5008 ( .A(n2800), .B(n2799), .Z(n2802) );
  ANDN U5009 ( .B(n2802), .A(n2801), .Z(n2803) );
  NANDN U5010 ( .A(n2804), .B(n2803), .Z(n2808) );
  AND U5011 ( .A(n2806), .B(n2805), .Z(n2807) );
  NAND U5012 ( .A(n2808), .B(n2807), .Z(n2809) );
  NANDN U5013 ( .A(n2810), .B(n2809), .Z(n2812) );
  OR U5014 ( .A(n2812), .B(n2811), .Z(n2813) );
  AND U5015 ( .A(n2814), .B(n2813), .Z(n2815) );
  NOR U5016 ( .A(n2816), .B(n2815), .Z(n2817) );
  NANDN U5017 ( .A(n2818), .B(n2817), .Z(n2819) );
  AND U5018 ( .A(n2820), .B(n2819), .Z(n2822) );
  NANDN U5019 ( .A(y[218]), .B(x[218]), .Z(n2821) );
  NAND U5020 ( .A(n2822), .B(n2821), .Z(n2824) );
  ANDN U5021 ( .B(n2824), .A(n2823), .Z(n2825) );
  NANDN U5022 ( .A(n2826), .B(n2825), .Z(n2827) );
  AND U5023 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U5024 ( .A(n2830), .B(n2829), .Z(n2831) );
  NANDN U5025 ( .A(n2832), .B(n2831), .Z(n2834) );
  OR U5026 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U5027 ( .A(n2836), .B(n2835), .Z(n2837) );
  NOR U5028 ( .A(n2838), .B(n2837), .Z(n2839) );
  NANDN U5029 ( .A(n2840), .B(n2839), .Z(n2841) );
  AND U5030 ( .A(n2842), .B(n2841), .Z(n2844) );
  NANDN U5031 ( .A(y[224]), .B(x[224]), .Z(n2843) );
  NAND U5032 ( .A(n2844), .B(n2843), .Z(n2846) );
  ANDN U5033 ( .B(n2846), .A(n2845), .Z(n2847) );
  NANDN U5034 ( .A(n2848), .B(n2847), .Z(n2849) );
  AND U5035 ( .A(n2850), .B(n2849), .Z(n2851) );
  NAND U5036 ( .A(n2852), .B(n2851), .Z(n2853) );
  NANDN U5037 ( .A(n2854), .B(n2853), .Z(n2856) );
  OR U5038 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U5039 ( .A(n2858), .B(n2857), .Z(n2860) );
  NOR U5040 ( .A(n2860), .B(n2859), .Z(n2861) );
  NANDN U5041 ( .A(n2862), .B(n2861), .Z(n2863) );
  AND U5042 ( .A(n2864), .B(n2863), .Z(n2866) );
  NAND U5043 ( .A(n2866), .B(n2865), .Z(n2868) );
  ANDN U5044 ( .B(n2868), .A(n2867), .Z(n2869) );
  NANDN U5045 ( .A(n2870), .B(n2869), .Z(n2874) );
  AND U5046 ( .A(n2872), .B(n2871), .Z(n2873) );
  NAND U5047 ( .A(n2874), .B(n2873), .Z(n2875) );
  NANDN U5048 ( .A(n2876), .B(n2875), .Z(n2878) );
  OR U5049 ( .A(n2878), .B(n2877), .Z(n2879) );
  AND U5050 ( .A(n2880), .B(n2879), .Z(n2882) );
  NOR U5051 ( .A(n2882), .B(n2881), .Z(n2883) );
  NANDN U5052 ( .A(n2884), .B(n2883), .Z(n2885) );
  AND U5053 ( .A(n2886), .B(n2885), .Z(n2888) );
  NAND U5054 ( .A(n2888), .B(n2887), .Z(n2890) );
  ANDN U5055 ( .B(n2890), .A(n2889), .Z(n2891) );
  NANDN U5056 ( .A(n2892), .B(n2891), .Z(n2896) );
  AND U5057 ( .A(n2894), .B(n2893), .Z(n2895) );
  NAND U5058 ( .A(n2896), .B(n2895), .Z(n2897) );
  NANDN U5059 ( .A(n2898), .B(n2897), .Z(n2900) );
  OR U5060 ( .A(n2900), .B(n2899), .Z(n2901) );
  AND U5061 ( .A(n2902), .B(n2901), .Z(n2904) );
  NOR U5062 ( .A(n2904), .B(n2903), .Z(n2905) );
  NANDN U5063 ( .A(n2906), .B(n2905), .Z(n2907) );
  AND U5064 ( .A(n2908), .B(n2907), .Z(n2910) );
  NAND U5065 ( .A(n2910), .B(n2909), .Z(n2912) );
  ANDN U5066 ( .B(n2912), .A(n2911), .Z(n2913) );
  NANDN U5067 ( .A(n2914), .B(n2913), .Z(n2918) );
  AND U5068 ( .A(n2916), .B(n2915), .Z(n2917) );
  NAND U5069 ( .A(n2918), .B(n2917), .Z(n2919) );
  NANDN U5070 ( .A(n2920), .B(n2919), .Z(n2922) );
  OR U5071 ( .A(n2922), .B(n2921), .Z(n2923) );
  AND U5072 ( .A(n2924), .B(n2923), .Z(n2926) );
  NOR U5073 ( .A(n2926), .B(n2925), .Z(n2927) );
  NANDN U5074 ( .A(n2928), .B(n2927), .Z(n2929) );
  AND U5075 ( .A(n2930), .B(n2929), .Z(n2932) );
  NAND U5076 ( .A(n2932), .B(n2931), .Z(n2934) );
  ANDN U5077 ( .B(n2934), .A(n2933), .Z(n2935) );
  NANDN U5078 ( .A(n2936), .B(n2935), .Z(n2937) );
  AND U5079 ( .A(n2938), .B(n2937), .Z(n2939) );
  NAND U5080 ( .A(n2940), .B(n2939), .Z(n2941) );
  NANDN U5081 ( .A(n2942), .B(n2941), .Z(n2944) );
  OR U5082 ( .A(n2944), .B(n2943), .Z(n2945) );
  AND U5083 ( .A(n2946), .B(n2945), .Z(n2947) );
  NOR U5084 ( .A(n2948), .B(n2947), .Z(n2949) );
  NANDN U5085 ( .A(n2950), .B(n2949), .Z(n2951) );
  AND U5086 ( .A(n2952), .B(n2951), .Z(n2954) );
  NANDN U5087 ( .A(y[254]), .B(x[254]), .Z(n2953) );
  NAND U5088 ( .A(n2954), .B(n2953), .Z(n2956) );
  ANDN U5089 ( .B(n2956), .A(n2955), .Z(n2957) );
  NANDN U5090 ( .A(n2958), .B(n2957), .Z(n2962) );
  AND U5091 ( .A(n2960), .B(n2959), .Z(n2961) );
  NAND U5092 ( .A(n2962), .B(n2961), .Z(n2963) );
  NANDN U5093 ( .A(n2964), .B(n2963), .Z(n2966) );
  OR U5094 ( .A(n2966), .B(n2965), .Z(n2967) );
  AND U5095 ( .A(n2968), .B(n2967), .Z(n2970) );
  NOR U5096 ( .A(n2970), .B(n2969), .Z(n2971) );
  NANDN U5097 ( .A(n2972), .B(n2971), .Z(n2973) );
  AND U5098 ( .A(n2974), .B(n2973), .Z(n2976) );
  NAND U5099 ( .A(n2976), .B(n2975), .Z(n2978) );
  ANDN U5100 ( .B(n2978), .A(n2977), .Z(n2979) );
  NANDN U5101 ( .A(n2980), .B(n2979), .Z(n2984) );
  AND U5102 ( .A(n2982), .B(n2981), .Z(n2983) );
  NAND U5103 ( .A(n2984), .B(n2983), .Z(n2985) );
  NANDN U5104 ( .A(n2986), .B(n2985), .Z(n2988) );
  OR U5105 ( .A(n2988), .B(n2987), .Z(n2989) );
  AND U5106 ( .A(n2990), .B(n2989), .Z(n2991) );
  NOR U5107 ( .A(n2992), .B(n2991), .Z(n2993) );
  NANDN U5108 ( .A(n2994), .B(n2993), .Z(n2995) );
  AND U5109 ( .A(n2996), .B(n2995), .Z(n2998) );
  NANDN U5110 ( .A(y[266]), .B(x[266]), .Z(n2997) );
  NAND U5111 ( .A(n2998), .B(n2997), .Z(n3000) );
  ANDN U5112 ( .B(n3000), .A(n2999), .Z(n3001) );
  NANDN U5113 ( .A(n3002), .B(n3001), .Z(n3006) );
  AND U5114 ( .A(n3004), .B(n3003), .Z(n3005) );
  NAND U5115 ( .A(n3006), .B(n3005), .Z(n3007) );
  NANDN U5116 ( .A(n3008), .B(n3007), .Z(n3010) );
  OR U5117 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U5118 ( .A(n3012), .B(n3011), .Z(n3013) );
  NOR U5119 ( .A(n3014), .B(n3013), .Z(n3015) );
  NANDN U5120 ( .A(n3016), .B(n3015), .Z(n3017) );
  AND U5121 ( .A(n3018), .B(n3017), .Z(n3020) );
  NANDN U5122 ( .A(y[272]), .B(x[272]), .Z(n3019) );
  NAND U5123 ( .A(n3020), .B(n3019), .Z(n3022) );
  ANDN U5124 ( .B(n3022), .A(n3021), .Z(n3023) );
  NANDN U5125 ( .A(n3024), .B(n3023), .Z(n3028) );
  AND U5126 ( .A(n3026), .B(n3025), .Z(n3027) );
  NAND U5127 ( .A(n3028), .B(n3027), .Z(n3029) );
  NANDN U5128 ( .A(n3030), .B(n3029), .Z(n3032) );
  OR U5129 ( .A(n3032), .B(n3031), .Z(n3033) );
  AND U5130 ( .A(n3034), .B(n3033), .Z(n3035) );
  NOR U5131 ( .A(n3036), .B(n3035), .Z(n3037) );
  NANDN U5132 ( .A(n3038), .B(n3037), .Z(n3039) );
  AND U5133 ( .A(n3040), .B(n3039), .Z(n3042) );
  NANDN U5134 ( .A(y[278]), .B(x[278]), .Z(n3041) );
  NAND U5135 ( .A(n3042), .B(n3041), .Z(n3044) );
  ANDN U5136 ( .B(n3044), .A(n3043), .Z(n3045) );
  NANDN U5137 ( .A(n3046), .B(n3045), .Z(n3050) );
  AND U5138 ( .A(n3048), .B(n3047), .Z(n3049) );
  NAND U5139 ( .A(n3050), .B(n3049), .Z(n3051) );
  NANDN U5140 ( .A(n3052), .B(n3051), .Z(n3054) );
  OR U5141 ( .A(n3054), .B(n3053), .Z(n3055) );
  AND U5142 ( .A(n3056), .B(n3055), .Z(n3058) );
  NOR U5143 ( .A(n3058), .B(n3057), .Z(n3059) );
  NANDN U5144 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U5145 ( .A(n3062), .B(n3061), .Z(n3064) );
  NAND U5146 ( .A(n3064), .B(n3063), .Z(n3066) );
  ANDN U5147 ( .B(n3066), .A(n3065), .Z(n3067) );
  NANDN U5148 ( .A(n3068), .B(n3067), .Z(n3069) );
  AND U5149 ( .A(n3070), .B(n3069), .Z(n3071) );
  NAND U5150 ( .A(n3072), .B(n3071), .Z(n3073) );
  NANDN U5151 ( .A(n3074), .B(n3073), .Z(n3076) );
  OR U5152 ( .A(n3076), .B(n3075), .Z(n3077) );
  AND U5153 ( .A(n3078), .B(n3077), .Z(n3080) );
  NOR U5154 ( .A(n3080), .B(n3079), .Z(n3081) );
  NANDN U5155 ( .A(n3082), .B(n3081), .Z(n3083) );
  AND U5156 ( .A(n3084), .B(n3083), .Z(n3086) );
  NAND U5157 ( .A(n3086), .B(n3085), .Z(n3088) );
  ANDN U5158 ( .B(n3088), .A(n3087), .Z(n3089) );
  NANDN U5159 ( .A(n3090), .B(n3089), .Z(n3094) );
  AND U5160 ( .A(n3092), .B(n3091), .Z(n3093) );
  NAND U5161 ( .A(n3094), .B(n3093), .Z(n3095) );
  NANDN U5162 ( .A(n3096), .B(n3095), .Z(n3097) );
  OR U5163 ( .A(n3098), .B(n3097), .Z(n3099) );
  AND U5164 ( .A(n3100), .B(n3099), .Z(n3102) );
  NAND U5165 ( .A(n3102), .B(n3101), .Z(n3104) );
  ANDN U5166 ( .B(n3104), .A(n3103), .Z(n3105) );
  NANDN U5167 ( .A(n3106), .B(n3105), .Z(n3110) );
  AND U5168 ( .A(n3108), .B(n3107), .Z(n3109) );
  NAND U5169 ( .A(n3110), .B(n3109), .Z(n3111) );
  NANDN U5170 ( .A(n3112), .B(n3111), .Z(n3115) );
  NANDN U5171 ( .A(x[298]), .B(n3115), .Z(n3114) );
  ANDN U5172 ( .B(n3114), .A(n3113), .Z(n3118) );
  XNOR U5173 ( .A(n3115), .B(x[298]), .Z(n3116) );
  NAND U5174 ( .A(n3116), .B(y[298]), .Z(n3117) );
  NAND U5175 ( .A(n3118), .B(n3117), .Z(n3119) );
  NAND U5176 ( .A(n6005), .B(n3119), .Z(n3120) );
  NANDN U5177 ( .A(n3121), .B(n3120), .Z(n3122) );
  AND U5178 ( .A(n3123), .B(n3122), .Z(n3125) );
  NOR U5179 ( .A(n3125), .B(n3124), .Z(n3126) );
  NANDN U5180 ( .A(n3127), .B(n3126), .Z(n3128) );
  AND U5181 ( .A(n3129), .B(n3128), .Z(n3131) );
  NAND U5182 ( .A(n3131), .B(n3130), .Z(n3133) );
  ANDN U5183 ( .B(n3133), .A(n3132), .Z(n3134) );
  NANDN U5184 ( .A(n3135), .B(n3134), .Z(n3139) );
  AND U5185 ( .A(n3137), .B(n3136), .Z(n3138) );
  NAND U5186 ( .A(n3139), .B(n3138), .Z(n3140) );
  NANDN U5187 ( .A(n3141), .B(n3140), .Z(n3143) );
  OR U5188 ( .A(n3143), .B(n3142), .Z(n3144) );
  AND U5189 ( .A(n3145), .B(n3144), .Z(n3147) );
  NOR U5190 ( .A(n3147), .B(n3146), .Z(n3148) );
  NANDN U5191 ( .A(n3149), .B(n3148), .Z(n3150) );
  AND U5192 ( .A(n3151), .B(n3150), .Z(n3153) );
  NAND U5193 ( .A(n3153), .B(n3152), .Z(n3155) );
  ANDN U5194 ( .B(n3155), .A(n3154), .Z(n3156) );
  NANDN U5195 ( .A(n3157), .B(n3156), .Z(n3158) );
  AND U5196 ( .A(n3159), .B(n3158), .Z(n3160) );
  NAND U5197 ( .A(n3161), .B(n3160), .Z(n3162) );
  NANDN U5198 ( .A(n3163), .B(n3162), .Z(n3165) );
  OR U5199 ( .A(n3165), .B(n3164), .Z(n3166) );
  AND U5200 ( .A(n3167), .B(n3166), .Z(n3168) );
  NOR U5201 ( .A(n3169), .B(n3168), .Z(n3170) );
  NANDN U5202 ( .A(n3171), .B(n3170), .Z(n3172) );
  AND U5203 ( .A(n3173), .B(n3172), .Z(n3175) );
  NANDN U5204 ( .A(y[314]), .B(x[314]), .Z(n3174) );
  NAND U5205 ( .A(n3175), .B(n3174), .Z(n3177) );
  ANDN U5206 ( .B(n3177), .A(n3176), .Z(n3178) );
  NANDN U5207 ( .A(n3179), .B(n3178), .Z(n3183) );
  AND U5208 ( .A(n3181), .B(n3180), .Z(n3182) );
  NAND U5209 ( .A(n3183), .B(n3182), .Z(n3184) );
  NANDN U5210 ( .A(n3185), .B(n3184), .Z(n3187) );
  OR U5211 ( .A(n3187), .B(n3186), .Z(n3188) );
  AND U5212 ( .A(n3189), .B(n3188), .Z(n3191) );
  NOR U5213 ( .A(n3191), .B(n3190), .Z(n3192) );
  NANDN U5214 ( .A(n3193), .B(n3192), .Z(n3194) );
  AND U5215 ( .A(n3195), .B(n3194), .Z(n3197) );
  NAND U5216 ( .A(n3197), .B(n3196), .Z(n3199) );
  ANDN U5217 ( .B(n3199), .A(n3198), .Z(n3200) );
  NANDN U5218 ( .A(n3201), .B(n3200), .Z(n3205) );
  AND U5219 ( .A(n3203), .B(n3202), .Z(n3204) );
  NAND U5220 ( .A(n3205), .B(n3204), .Z(n3206) );
  NANDN U5221 ( .A(n3207), .B(n3206), .Z(n3209) );
  OR U5222 ( .A(n3209), .B(n3208), .Z(n3210) );
  AND U5223 ( .A(n3211), .B(n3210), .Z(n3213) );
  NOR U5224 ( .A(n3213), .B(n3212), .Z(n3214) );
  NANDN U5225 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U5226 ( .A(n3217), .B(n3216), .Z(n3219) );
  NAND U5227 ( .A(n3219), .B(n3218), .Z(n3221) );
  ANDN U5228 ( .B(n3221), .A(n3220), .Z(n3222) );
  NANDN U5229 ( .A(n3223), .B(n3222), .Z(n3224) );
  AND U5230 ( .A(n3225), .B(n3224), .Z(n3226) );
  NAND U5231 ( .A(n3227), .B(n3226), .Z(n3228) );
  NANDN U5232 ( .A(n3229), .B(n3228), .Z(n3231) );
  OR U5233 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U5234 ( .A(n3233), .B(n3232), .Z(n3235) );
  NOR U5235 ( .A(n3235), .B(n3234), .Z(n3236) );
  NANDN U5236 ( .A(n3237), .B(n3236), .Z(n3238) );
  AND U5237 ( .A(n3239), .B(n3238), .Z(n3241) );
  NAND U5238 ( .A(n3241), .B(n3240), .Z(n3243) );
  ANDN U5239 ( .B(n3243), .A(n3242), .Z(n3244) );
  NANDN U5240 ( .A(n3245), .B(n3244), .Z(n3249) );
  AND U5241 ( .A(n3247), .B(n3246), .Z(n3248) );
  NAND U5242 ( .A(n3249), .B(n3248), .Z(n3250) );
  NANDN U5243 ( .A(n3251), .B(n3250), .Z(n3253) );
  OR U5244 ( .A(n3253), .B(n3252), .Z(n3254) );
  AND U5245 ( .A(n3255), .B(n3254), .Z(n3256) );
  NOR U5246 ( .A(n3257), .B(n3256), .Z(n3258) );
  NANDN U5247 ( .A(n3259), .B(n3258), .Z(n3260) );
  AND U5248 ( .A(n3261), .B(n3260), .Z(n3263) );
  NANDN U5249 ( .A(y[338]), .B(x[338]), .Z(n3262) );
  NAND U5250 ( .A(n3263), .B(n3262), .Z(n3265) );
  ANDN U5251 ( .B(n3265), .A(n3264), .Z(n3266) );
  NANDN U5252 ( .A(n3267), .B(n3266), .Z(n3271) );
  AND U5253 ( .A(n3269), .B(n3268), .Z(n3270) );
  NAND U5254 ( .A(n3271), .B(n3270), .Z(n3272) );
  NANDN U5255 ( .A(n3273), .B(n3272), .Z(n3275) );
  OR U5256 ( .A(n3275), .B(n3274), .Z(n3276) );
  AND U5257 ( .A(n3277), .B(n3276), .Z(n3278) );
  NOR U5258 ( .A(n3279), .B(n3278), .Z(n3280) );
  NANDN U5259 ( .A(n3281), .B(n3280), .Z(n3282) );
  AND U5260 ( .A(n3283), .B(n3282), .Z(n3285) );
  NANDN U5261 ( .A(y[344]), .B(x[344]), .Z(n3284) );
  NAND U5262 ( .A(n3285), .B(n3284), .Z(n3287) );
  ANDN U5263 ( .B(n3287), .A(n3286), .Z(n3288) );
  NANDN U5264 ( .A(n3289), .B(n3288), .Z(n3290) );
  AND U5265 ( .A(n3291), .B(n3290), .Z(n3292) );
  NAND U5266 ( .A(n3293), .B(n3292), .Z(n3294) );
  NANDN U5267 ( .A(n3295), .B(n3294), .Z(n3297) );
  OR U5268 ( .A(n3297), .B(n3296), .Z(n3298) );
  AND U5269 ( .A(n3299), .B(n3298), .Z(n3301) );
  NOR U5270 ( .A(n3301), .B(n3300), .Z(n3302) );
  NANDN U5271 ( .A(n3303), .B(n3302), .Z(n3304) );
  AND U5272 ( .A(n3305), .B(n3304), .Z(n3307) );
  NAND U5273 ( .A(n3307), .B(n3306), .Z(n3309) );
  ANDN U5274 ( .B(n3309), .A(n3308), .Z(n3310) );
  NANDN U5275 ( .A(n3311), .B(n3310), .Z(n3315) );
  NANDN U5276 ( .A(y[352]), .B(x[352]), .Z(n3312) );
  AND U5277 ( .A(n3313), .B(n3312), .Z(n3314) );
  NAND U5278 ( .A(n3315), .B(n3314), .Z(n3316) );
  NANDN U5279 ( .A(n3317), .B(n3316), .Z(n3319) );
  OR U5280 ( .A(n3319), .B(n3318), .Z(n3320) );
  AND U5281 ( .A(n3321), .B(n3320), .Z(n3322) );
  NOR U5282 ( .A(n3323), .B(n3322), .Z(n3324) );
  NANDN U5283 ( .A(n3325), .B(n3324), .Z(n3326) );
  AND U5284 ( .A(n3327), .B(n3326), .Z(n3329) );
  NANDN U5285 ( .A(y[356]), .B(x[356]), .Z(n3328) );
  NAND U5286 ( .A(n3329), .B(n3328), .Z(n3331) );
  ANDN U5287 ( .B(n3331), .A(n3330), .Z(n3332) );
  NANDN U5288 ( .A(n3333), .B(n3332), .Z(n3334) );
  AND U5289 ( .A(n3335), .B(n3334), .Z(n3336) );
  NAND U5290 ( .A(n3337), .B(n3336), .Z(n3338) );
  NANDN U5291 ( .A(n3339), .B(n3338), .Z(n3341) );
  OR U5292 ( .A(n3341), .B(n3340), .Z(n3342) );
  AND U5293 ( .A(n3343), .B(n3342), .Z(n3344) );
  NOR U5294 ( .A(n3345), .B(n3344), .Z(n3346) );
  NANDN U5295 ( .A(n3347), .B(n3346), .Z(n3348) );
  AND U5296 ( .A(n3349), .B(n3348), .Z(n3351) );
  NANDN U5297 ( .A(y[362]), .B(x[362]), .Z(n3350) );
  NAND U5298 ( .A(n3351), .B(n3350), .Z(n3353) );
  ANDN U5299 ( .B(n3353), .A(n3352), .Z(n3354) );
  NANDN U5300 ( .A(n3355), .B(n3354), .Z(n3356) );
  AND U5301 ( .A(n3357), .B(n3356), .Z(n3358) );
  NAND U5302 ( .A(n3359), .B(n3358), .Z(n3360) );
  NANDN U5303 ( .A(n3361), .B(n3360), .Z(n3363) );
  OR U5304 ( .A(n3363), .B(n3362), .Z(n3364) );
  AND U5305 ( .A(n3365), .B(n3364), .Z(n3367) );
  NOR U5306 ( .A(n3367), .B(n3366), .Z(n3368) );
  NANDN U5307 ( .A(n3369), .B(n3368), .Z(n3370) );
  AND U5308 ( .A(n3371), .B(n3370), .Z(n3373) );
  NAND U5309 ( .A(n3373), .B(n3372), .Z(n3375) );
  ANDN U5310 ( .B(n3375), .A(n3374), .Z(n3376) );
  NANDN U5311 ( .A(n3377), .B(n3376), .Z(n3381) );
  NANDN U5312 ( .A(y[370]), .B(x[370]), .Z(n3378) );
  AND U5313 ( .A(n3379), .B(n3378), .Z(n3380) );
  NAND U5314 ( .A(n3381), .B(n3380), .Z(n3382) );
  NANDN U5315 ( .A(n3383), .B(n3382), .Z(n3385) );
  OR U5316 ( .A(n3385), .B(n3384), .Z(n3386) );
  AND U5317 ( .A(n3387), .B(n3386), .Z(n3389) );
  NOR U5318 ( .A(n3389), .B(n3388), .Z(n3390) );
  NANDN U5319 ( .A(n3391), .B(n3390), .Z(n3392) );
  AND U5320 ( .A(n3393), .B(n3392), .Z(n3395) );
  NAND U5321 ( .A(n3395), .B(n3394), .Z(n3397) );
  ANDN U5322 ( .B(n3397), .A(n3396), .Z(n3398) );
  NANDN U5323 ( .A(n3399), .B(n3398), .Z(n3403) );
  NANDN U5324 ( .A(y[376]), .B(x[376]), .Z(n3400) );
  AND U5325 ( .A(n3401), .B(n3400), .Z(n3402) );
  NAND U5326 ( .A(n3403), .B(n3402), .Z(n3404) );
  NANDN U5327 ( .A(n3405), .B(n3404), .Z(n3407) );
  OR U5328 ( .A(n3407), .B(n3406), .Z(n3408) );
  AND U5329 ( .A(n3409), .B(n3408), .Z(n3411) );
  NOR U5330 ( .A(n3411), .B(n3410), .Z(n3412) );
  NANDN U5331 ( .A(n3413), .B(n3412), .Z(n3414) );
  AND U5332 ( .A(n3415), .B(n3414), .Z(n3417) );
  NAND U5333 ( .A(n3417), .B(n3416), .Z(n3419) );
  ANDN U5334 ( .B(n3419), .A(n3418), .Z(n3420) );
  NANDN U5335 ( .A(n3421), .B(n3420), .Z(n3422) );
  AND U5336 ( .A(n3423), .B(n3422), .Z(n3424) );
  NAND U5337 ( .A(n3425), .B(n3424), .Z(n3426) );
  NANDN U5338 ( .A(n3427), .B(n3426), .Z(n3429) );
  OR U5339 ( .A(n3429), .B(n3428), .Z(n3430) );
  AND U5340 ( .A(n3431), .B(n3430), .Z(n3433) );
  NOR U5341 ( .A(n3433), .B(n3432), .Z(n3434) );
  NANDN U5342 ( .A(n3435), .B(n3434), .Z(n3436) );
  AND U5343 ( .A(n3437), .B(n3436), .Z(n3439) );
  NAND U5344 ( .A(n3439), .B(n3438), .Z(n3441) );
  ANDN U5345 ( .B(n3441), .A(n3440), .Z(n3442) );
  NANDN U5346 ( .A(n3443), .B(n3442), .Z(n3447) );
  AND U5347 ( .A(n3445), .B(n3444), .Z(n3446) );
  NAND U5348 ( .A(n3447), .B(n3446), .Z(n3448) );
  NANDN U5349 ( .A(n3449), .B(n3448), .Z(n3451) );
  OR U5350 ( .A(n3451), .B(n3450), .Z(n3452) );
  AND U5351 ( .A(n3453), .B(n3452), .Z(n3454) );
  NOR U5352 ( .A(n3455), .B(n3454), .Z(n3456) );
  NANDN U5353 ( .A(n3457), .B(n3456), .Z(n3458) );
  AND U5354 ( .A(n3459), .B(n3458), .Z(n3461) );
  NANDN U5355 ( .A(y[392]), .B(x[392]), .Z(n3460) );
  NAND U5356 ( .A(n3461), .B(n3460), .Z(n3463) );
  ANDN U5357 ( .B(n3463), .A(n3462), .Z(n3464) );
  NANDN U5358 ( .A(n3465), .B(n3464), .Z(n3466) );
  AND U5359 ( .A(n3467), .B(n3466), .Z(n3468) );
  NAND U5360 ( .A(n3469), .B(n3468), .Z(n3470) );
  NANDN U5361 ( .A(n3471), .B(n3470), .Z(n3473) );
  OR U5362 ( .A(n3473), .B(n3472), .Z(n3474) );
  AND U5363 ( .A(n3475), .B(n3474), .Z(n3476) );
  NOR U5364 ( .A(n3477), .B(n3476), .Z(n3478) );
  NANDN U5365 ( .A(n3479), .B(n3478), .Z(n3480) );
  AND U5366 ( .A(n3481), .B(n3480), .Z(n3483) );
  NANDN U5367 ( .A(y[398]), .B(x[398]), .Z(n3482) );
  NAND U5368 ( .A(n3483), .B(n3482), .Z(n3485) );
  ANDN U5369 ( .B(n3485), .A(n3484), .Z(n3486) );
  NANDN U5370 ( .A(n3487), .B(n3486), .Z(n3491) );
  NANDN U5371 ( .A(y[400]), .B(x[400]), .Z(n3488) );
  AND U5372 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND U5373 ( .A(n3491), .B(n3490), .Z(n3492) );
  NANDN U5374 ( .A(n3493), .B(n3492), .Z(n3495) );
  OR U5375 ( .A(n3495), .B(n3494), .Z(n3496) );
  AND U5376 ( .A(n3497), .B(n3496), .Z(n3499) );
  NOR U5377 ( .A(n3499), .B(n3498), .Z(n3500) );
  NANDN U5378 ( .A(n3501), .B(n3500), .Z(n3502) );
  AND U5379 ( .A(n3503), .B(n3502), .Z(n3505) );
  NAND U5380 ( .A(n3505), .B(n3504), .Z(n3507) );
  ANDN U5381 ( .B(n3507), .A(n3506), .Z(n3508) );
  NANDN U5382 ( .A(n3509), .B(n3508), .Z(n3510) );
  AND U5383 ( .A(n3511), .B(n3510), .Z(n3512) );
  NAND U5384 ( .A(n3513), .B(n3512), .Z(n3514) );
  NANDN U5385 ( .A(n3515), .B(n3514), .Z(n3517) );
  OR U5386 ( .A(n3517), .B(n3516), .Z(n3518) );
  AND U5387 ( .A(n3519), .B(n3518), .Z(n3521) );
  NOR U5388 ( .A(n3521), .B(n3520), .Z(n3522) );
  NANDN U5389 ( .A(n3523), .B(n3522), .Z(n3524) );
  AND U5390 ( .A(n3525), .B(n3524), .Z(n3527) );
  NAND U5391 ( .A(n3527), .B(n3526), .Z(n3529) );
  ANDN U5392 ( .B(n3529), .A(n3528), .Z(n3530) );
  NANDN U5393 ( .A(n3531), .B(n3530), .Z(n3535) );
  AND U5394 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U5395 ( .A(n3535), .B(n3534), .Z(n3536) );
  NANDN U5396 ( .A(n3537), .B(n3536), .Z(n3539) );
  OR U5397 ( .A(n3539), .B(n3538), .Z(n3540) );
  AND U5398 ( .A(n3541), .B(n3540), .Z(n3543) );
  NOR U5399 ( .A(n3543), .B(n3542), .Z(n3544) );
  NANDN U5400 ( .A(n3545), .B(n3544), .Z(n3546) );
  AND U5401 ( .A(n3547), .B(n3546), .Z(n3549) );
  NAND U5402 ( .A(n3549), .B(n3548), .Z(n3551) );
  ANDN U5403 ( .B(n3551), .A(n3550), .Z(n3552) );
  NANDN U5404 ( .A(n3553), .B(n3552), .Z(n3554) );
  AND U5405 ( .A(n3555), .B(n3554), .Z(n3556) );
  NAND U5406 ( .A(n3557), .B(n3556), .Z(n3558) );
  NANDN U5407 ( .A(n3559), .B(n3558), .Z(n3561) );
  OR U5408 ( .A(n3561), .B(n3560), .Z(n3562) );
  AND U5409 ( .A(n3563), .B(n3562), .Z(n3565) );
  NOR U5410 ( .A(n3565), .B(n3564), .Z(n3566) );
  NANDN U5411 ( .A(n3567), .B(n3566), .Z(n3568) );
  AND U5412 ( .A(n3569), .B(n3568), .Z(n3571) );
  NAND U5413 ( .A(n3571), .B(n3570), .Z(n3573) );
  ANDN U5414 ( .B(n3573), .A(n3572), .Z(n3574) );
  NANDN U5415 ( .A(n3575), .B(n3574), .Z(n3579) );
  AND U5416 ( .A(n3577), .B(n3576), .Z(n3578) );
  NAND U5417 ( .A(n3579), .B(n3578), .Z(n3580) );
  NANDN U5418 ( .A(n3581), .B(n3580), .Z(n3583) );
  OR U5419 ( .A(n3583), .B(n3582), .Z(n3584) );
  AND U5420 ( .A(n3585), .B(n3584), .Z(n3587) );
  NOR U5421 ( .A(n3587), .B(n3586), .Z(n3588) );
  NANDN U5422 ( .A(n3589), .B(n3588), .Z(n3590) );
  AND U5423 ( .A(n3591), .B(n3590), .Z(n3593) );
  NAND U5424 ( .A(n3593), .B(n3592), .Z(n3595) );
  ANDN U5425 ( .B(n3595), .A(n3594), .Z(n3596) );
  NANDN U5426 ( .A(n3597), .B(n3596), .Z(n3601) );
  AND U5427 ( .A(n3599), .B(n3598), .Z(n3600) );
  NAND U5428 ( .A(n3601), .B(n3600), .Z(n3602) );
  NANDN U5429 ( .A(n3603), .B(n3602), .Z(n3605) );
  OR U5430 ( .A(n3605), .B(n3604), .Z(n3606) );
  AND U5431 ( .A(n3607), .B(n3606), .Z(n3608) );
  NOR U5432 ( .A(n3609), .B(n3608), .Z(n3610) );
  NANDN U5433 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U5434 ( .A(n3613), .B(n3612), .Z(n3615) );
  NANDN U5435 ( .A(y[434]), .B(x[434]), .Z(n3614) );
  NAND U5436 ( .A(n3615), .B(n3614), .Z(n3617) );
  ANDN U5437 ( .B(n3617), .A(n3616), .Z(n3618) );
  NANDN U5438 ( .A(n3619), .B(n3618), .Z(n3620) );
  AND U5439 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U5440 ( .A(n3623), .B(n3622), .Z(n3624) );
  NANDN U5441 ( .A(n3625), .B(n3624), .Z(n3627) );
  OR U5442 ( .A(n3627), .B(n3626), .Z(n3628) );
  AND U5443 ( .A(n3629), .B(n3628), .Z(n3631) );
  NOR U5444 ( .A(n3631), .B(n3630), .Z(n3632) );
  NANDN U5445 ( .A(n3633), .B(n3632), .Z(n3634) );
  AND U5446 ( .A(n3635), .B(n3634), .Z(n3637) );
  NAND U5447 ( .A(n3637), .B(n3636), .Z(n3639) );
  ANDN U5448 ( .B(n3639), .A(n3638), .Z(n3640) );
  NANDN U5449 ( .A(n3641), .B(n3640), .Z(n3642) );
  AND U5450 ( .A(n3643), .B(n3642), .Z(n3644) );
  NAND U5451 ( .A(n3645), .B(n3644), .Z(n3646) );
  NANDN U5452 ( .A(n3647), .B(n3646), .Z(n3649) );
  OR U5453 ( .A(n3649), .B(n3648), .Z(n3650) );
  AND U5454 ( .A(n3651), .B(n3650), .Z(n3653) );
  NOR U5455 ( .A(n3653), .B(n3652), .Z(n3654) );
  NANDN U5456 ( .A(n3655), .B(n3654), .Z(n3656) );
  AND U5457 ( .A(n3657), .B(n3656), .Z(n3659) );
  NAND U5458 ( .A(n3659), .B(n3658), .Z(n3661) );
  ANDN U5459 ( .B(n3661), .A(n3660), .Z(n3662) );
  NANDN U5460 ( .A(n3663), .B(n3662), .Z(n3667) );
  AND U5461 ( .A(n3665), .B(n3664), .Z(n3666) );
  NAND U5462 ( .A(n3667), .B(n3666), .Z(n3668) );
  NANDN U5463 ( .A(n3669), .B(n3668), .Z(n3671) );
  OR U5464 ( .A(n3671), .B(n3670), .Z(n3672) );
  AND U5465 ( .A(n3673), .B(n3672), .Z(n3675) );
  NOR U5466 ( .A(n3675), .B(n3674), .Z(n3676) );
  NANDN U5467 ( .A(n3677), .B(n3676), .Z(n3678) );
  AND U5468 ( .A(n3679), .B(n3678), .Z(n3681) );
  NAND U5469 ( .A(n3681), .B(n3680), .Z(n3683) );
  ANDN U5470 ( .B(n3683), .A(n3682), .Z(n3684) );
  NANDN U5471 ( .A(n3685), .B(n3684), .Z(n3689) );
  AND U5472 ( .A(n3687), .B(n3686), .Z(n3688) );
  NAND U5473 ( .A(n3689), .B(n3688), .Z(n3690) );
  NANDN U5474 ( .A(n3691), .B(n3690), .Z(n3693) );
  OR U5475 ( .A(n3693), .B(n3692), .Z(n3694) );
  AND U5476 ( .A(n3695), .B(n3694), .Z(n3697) );
  NOR U5477 ( .A(n3697), .B(n3696), .Z(n3698) );
  NANDN U5478 ( .A(n3699), .B(n3698), .Z(n3700) );
  AND U5479 ( .A(n3701), .B(n3700), .Z(n3703) );
  NAND U5480 ( .A(n3703), .B(n3702), .Z(n3705) );
  ANDN U5481 ( .B(n3705), .A(n3704), .Z(n3706) );
  NANDN U5482 ( .A(n3707), .B(n3706), .Z(n3708) );
  AND U5483 ( .A(n3709), .B(n3708), .Z(n3710) );
  NAND U5484 ( .A(n3711), .B(n3710), .Z(n3712) );
  NANDN U5485 ( .A(n3713), .B(n3712), .Z(n3715) );
  OR U5486 ( .A(n3715), .B(n3714), .Z(n3716) );
  AND U5487 ( .A(n3717), .B(n3716), .Z(n3718) );
  NOR U5488 ( .A(n3719), .B(n3718), .Z(n3720) );
  NANDN U5489 ( .A(n3721), .B(n3720), .Z(n3722) );
  AND U5490 ( .A(n3723), .B(n3722), .Z(n3725) );
  NANDN U5491 ( .A(y[464]), .B(x[464]), .Z(n3724) );
  NAND U5492 ( .A(n3725), .B(n3724), .Z(n3727) );
  ANDN U5493 ( .B(n3727), .A(n3726), .Z(n3728) );
  NANDN U5494 ( .A(n3729), .B(n3728), .Z(n3733) );
  NANDN U5495 ( .A(y[466]), .B(x[466]), .Z(n3730) );
  AND U5496 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U5497 ( .A(n3733), .B(n3732), .Z(n3734) );
  NANDN U5498 ( .A(n3735), .B(n3734), .Z(n3737) );
  OR U5499 ( .A(n3737), .B(n3736), .Z(n3738) );
  AND U5500 ( .A(n3739), .B(n3738), .Z(n3741) );
  NOR U5501 ( .A(n3741), .B(n3740), .Z(n3742) );
  NANDN U5502 ( .A(n3743), .B(n3742), .Z(n3744) );
  AND U5503 ( .A(n3745), .B(n3744), .Z(n3747) );
  NAND U5504 ( .A(n3747), .B(n3746), .Z(n3749) );
  ANDN U5505 ( .B(n3749), .A(n3748), .Z(n3750) );
  NANDN U5506 ( .A(n3751), .B(n3750), .Z(n3755) );
  NANDN U5507 ( .A(y[472]), .B(x[472]), .Z(n3752) );
  AND U5508 ( .A(n3753), .B(n3752), .Z(n3754) );
  NAND U5509 ( .A(n3755), .B(n3754), .Z(n3756) );
  NANDN U5510 ( .A(n3757), .B(n3756), .Z(n3759) );
  OR U5511 ( .A(n3759), .B(n3758), .Z(n3760) );
  AND U5512 ( .A(n3761), .B(n3760), .Z(n3763) );
  NOR U5513 ( .A(n3763), .B(n3762), .Z(n3764) );
  NANDN U5514 ( .A(n3765), .B(n3764), .Z(n3766) );
  AND U5515 ( .A(n3767), .B(n3766), .Z(n3769) );
  NAND U5516 ( .A(n3769), .B(n3768), .Z(n3771) );
  ANDN U5517 ( .B(n3771), .A(n3770), .Z(n3772) );
  NANDN U5518 ( .A(n3773), .B(n3772), .Z(n3774) );
  AND U5519 ( .A(n3775), .B(n3774), .Z(n3776) );
  NAND U5520 ( .A(n3777), .B(n3776), .Z(n3778) );
  NANDN U5521 ( .A(n3779), .B(n3778), .Z(n3781) );
  OR U5522 ( .A(n3781), .B(n3780), .Z(n3782) );
  AND U5523 ( .A(n3783), .B(n3782), .Z(n3785) );
  NOR U5524 ( .A(n3785), .B(n3784), .Z(n3786) );
  NANDN U5525 ( .A(n3787), .B(n3786), .Z(n3788) );
  AND U5526 ( .A(n3789), .B(n3788), .Z(n3791) );
  NAND U5527 ( .A(n3791), .B(n3790), .Z(n3793) );
  ANDN U5528 ( .B(n3793), .A(n3792), .Z(n3794) );
  NANDN U5529 ( .A(n3795), .B(n3794), .Z(n3799) );
  NANDN U5530 ( .A(y[484]), .B(x[484]), .Z(n3796) );
  AND U5531 ( .A(n3797), .B(n3796), .Z(n3798) );
  NAND U5532 ( .A(n3799), .B(n3798), .Z(n3800) );
  NANDN U5533 ( .A(n3801), .B(n3800), .Z(n3803) );
  OR U5534 ( .A(n3803), .B(n3802), .Z(n3804) );
  AND U5535 ( .A(n3805), .B(n3804), .Z(n3806) );
  NOR U5536 ( .A(n3807), .B(n3806), .Z(n3808) );
  NANDN U5537 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U5538 ( .A(n3811), .B(n3810), .Z(n3813) );
  NANDN U5539 ( .A(y[488]), .B(x[488]), .Z(n3812) );
  NAND U5540 ( .A(n3813), .B(n3812), .Z(n3815) );
  ANDN U5541 ( .B(n3815), .A(n3814), .Z(n3816) );
  NANDN U5542 ( .A(n3817), .B(n3816), .Z(n3818) );
  AND U5543 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U5544 ( .A(n3821), .B(n3820), .Z(n3822) );
  NANDN U5545 ( .A(n3823), .B(n3822), .Z(n3825) );
  OR U5546 ( .A(n3825), .B(n3824), .Z(n3826) );
  AND U5547 ( .A(n3827), .B(n3826), .Z(n3829) );
  NOR U5548 ( .A(n3829), .B(n3828), .Z(n3830) );
  NANDN U5549 ( .A(n3831), .B(n3830), .Z(n3832) );
  AND U5550 ( .A(n3833), .B(n3832), .Z(n3835) );
  NAND U5551 ( .A(n3835), .B(n3834), .Z(n3837) );
  ANDN U5552 ( .B(n3837), .A(n3836), .Z(n3838) );
  NANDN U5553 ( .A(n3839), .B(n3838), .Z(n3840) );
  AND U5554 ( .A(n3841), .B(n3840), .Z(n3842) );
  NAND U5555 ( .A(n3843), .B(n3842), .Z(n3844) );
  NANDN U5556 ( .A(n3845), .B(n3844), .Z(n3847) );
  OR U5557 ( .A(n3847), .B(n3846), .Z(n3848) );
  AND U5558 ( .A(n3849), .B(n3848), .Z(n3851) );
  NOR U5559 ( .A(n3851), .B(n3850), .Z(n3852) );
  NANDN U5560 ( .A(n3853), .B(n3852), .Z(n3854) );
  AND U5561 ( .A(n3855), .B(n3854), .Z(n3857) );
  NAND U5562 ( .A(n3857), .B(n3856), .Z(n3859) );
  ANDN U5563 ( .B(n3859), .A(n3858), .Z(n3860) );
  NANDN U5564 ( .A(n3861), .B(n3860), .Z(n3865) );
  AND U5565 ( .A(n3863), .B(n3862), .Z(n3864) );
  NAND U5566 ( .A(n3865), .B(n3864), .Z(n3866) );
  NANDN U5567 ( .A(n3867), .B(n3866), .Z(n3869) );
  OR U5568 ( .A(n3869), .B(n3868), .Z(n3870) );
  AND U5569 ( .A(n3871), .B(n3870), .Z(n3873) );
  NOR U5570 ( .A(n3873), .B(n3872), .Z(n3874) );
  NANDN U5571 ( .A(n3875), .B(n3874), .Z(n3876) );
  AND U5572 ( .A(n3877), .B(n3876), .Z(n3879) );
  NAND U5573 ( .A(n3879), .B(n3878), .Z(n3881) );
  ANDN U5574 ( .B(n3881), .A(n3880), .Z(n3882) );
  NANDN U5575 ( .A(n3883), .B(n3882), .Z(n3884) );
  AND U5576 ( .A(n3885), .B(n3884), .Z(n3886) );
  NAND U5577 ( .A(n3887), .B(n3886), .Z(n3888) );
  NANDN U5578 ( .A(n3889), .B(n3888), .Z(n3891) );
  OR U5579 ( .A(n3891), .B(n3890), .Z(n3892) );
  AND U5580 ( .A(n3893), .B(n3892), .Z(n3895) );
  NOR U5581 ( .A(n3895), .B(n3894), .Z(n3896) );
  NANDN U5582 ( .A(n3897), .B(n3896), .Z(n3898) );
  AND U5583 ( .A(n3899), .B(n3898), .Z(n3901) );
  NAND U5584 ( .A(n3901), .B(n3900), .Z(n3903) );
  ANDN U5585 ( .B(n3903), .A(n3902), .Z(n3904) );
  NANDN U5586 ( .A(n3905), .B(n3904), .Z(n3906) );
  AND U5587 ( .A(n3907), .B(n3906), .Z(n3908) );
  NAND U5588 ( .A(n3909), .B(n3908), .Z(n3910) );
  NANDN U5589 ( .A(n3911), .B(n3910), .Z(n3913) );
  OR U5590 ( .A(n3913), .B(n3912), .Z(n3914) );
  AND U5591 ( .A(n3915), .B(n3914), .Z(n3917) );
  NOR U5592 ( .A(n3917), .B(n3916), .Z(n3918) );
  NANDN U5593 ( .A(n3919), .B(n3918), .Z(n3920) );
  AND U5594 ( .A(n3921), .B(n3920), .Z(n3923) );
  NAND U5595 ( .A(n3923), .B(n3922), .Z(n3925) );
  ANDN U5596 ( .B(n3925), .A(n3924), .Z(n3926) );
  NANDN U5597 ( .A(n3927), .B(n3926), .Z(n3931) );
  AND U5598 ( .A(n3929), .B(n3928), .Z(n3930) );
  NAND U5599 ( .A(n3931), .B(n3930), .Z(n3932) );
  NANDN U5600 ( .A(n3933), .B(n3932), .Z(n3935) );
  OR U5601 ( .A(n3935), .B(n3934), .Z(n3936) );
  AND U5602 ( .A(n3937), .B(n3936), .Z(n3939) );
  NOR U5603 ( .A(n3939), .B(n3938), .Z(n3940) );
  NANDN U5604 ( .A(n3941), .B(n3940), .Z(n3942) );
  AND U5605 ( .A(n3943), .B(n3942), .Z(n3945) );
  NAND U5606 ( .A(n3945), .B(n3944), .Z(n3947) );
  ANDN U5607 ( .B(n3947), .A(n3946), .Z(n3948) );
  NANDN U5608 ( .A(n3949), .B(n3948), .Z(n3953) );
  NANDN U5609 ( .A(y[526]), .B(x[526]), .Z(n3950) );
  AND U5610 ( .A(n3951), .B(n3950), .Z(n3952) );
  NAND U5611 ( .A(n3953), .B(n3952), .Z(n3954) );
  NANDN U5612 ( .A(n3955), .B(n3954), .Z(n3957) );
  OR U5613 ( .A(n3957), .B(n3956), .Z(n3958) );
  AND U5614 ( .A(n3959), .B(n3958), .Z(n3960) );
  NOR U5615 ( .A(n3961), .B(n3960), .Z(n3962) );
  NANDN U5616 ( .A(n3963), .B(n3962), .Z(n3964) );
  AND U5617 ( .A(n3965), .B(n3964), .Z(n3967) );
  NANDN U5618 ( .A(y[530]), .B(x[530]), .Z(n3966) );
  NAND U5619 ( .A(n3967), .B(n3966), .Z(n3969) );
  ANDN U5620 ( .B(n3969), .A(n3968), .Z(n3970) );
  NANDN U5621 ( .A(n3971), .B(n3970), .Z(n3972) );
  AND U5622 ( .A(n3973), .B(n3972), .Z(n3974) );
  NAND U5623 ( .A(n3975), .B(n3974), .Z(n3976) );
  NANDN U5624 ( .A(n3977), .B(n3976), .Z(n3979) );
  OR U5625 ( .A(n3979), .B(n3978), .Z(n3980) );
  AND U5626 ( .A(n3981), .B(n3980), .Z(n3983) );
  NOR U5627 ( .A(n3983), .B(n3982), .Z(n3984) );
  NANDN U5628 ( .A(n3985), .B(n3984), .Z(n3986) );
  AND U5629 ( .A(n3987), .B(n3986), .Z(n3989) );
  NAND U5630 ( .A(n3989), .B(n3988), .Z(n3991) );
  ANDN U5631 ( .B(n3991), .A(n3990), .Z(n3992) );
  NANDN U5632 ( .A(n3993), .B(n3992), .Z(n3994) );
  AND U5633 ( .A(n3995), .B(n3994), .Z(n3996) );
  NAND U5634 ( .A(n3997), .B(n3996), .Z(n3998) );
  NANDN U5635 ( .A(n3999), .B(n3998), .Z(n4001) );
  OR U5636 ( .A(n4001), .B(n4000), .Z(n4002) );
  AND U5637 ( .A(n4003), .B(n4002), .Z(n4005) );
  NOR U5638 ( .A(n4005), .B(n4004), .Z(n4006) );
  NANDN U5639 ( .A(n4007), .B(n4006), .Z(n4008) );
  AND U5640 ( .A(n4009), .B(n4008), .Z(n4011) );
  NAND U5641 ( .A(n4011), .B(n4010), .Z(n4013) );
  ANDN U5642 ( .B(n4013), .A(n4012), .Z(n4014) );
  NANDN U5643 ( .A(n4015), .B(n4014), .Z(n4019) );
  AND U5644 ( .A(n4017), .B(n4016), .Z(n4018) );
  NAND U5645 ( .A(n4019), .B(n4018), .Z(n4020) );
  NANDN U5646 ( .A(n4021), .B(n4020), .Z(n4023) );
  OR U5647 ( .A(n4023), .B(n4022), .Z(n4024) );
  AND U5648 ( .A(n4025), .B(n4024), .Z(n4027) );
  NOR U5649 ( .A(n4027), .B(n4026), .Z(n4028) );
  NANDN U5650 ( .A(n4029), .B(n4028), .Z(n4030) );
  AND U5651 ( .A(n4031), .B(n4030), .Z(n4033) );
  NAND U5652 ( .A(n4033), .B(n4032), .Z(n4035) );
  ANDN U5653 ( .B(n4035), .A(n4034), .Z(n4036) );
  NANDN U5654 ( .A(n4037), .B(n4036), .Z(n4038) );
  AND U5655 ( .A(n4039), .B(n4038), .Z(n4040) );
  NAND U5656 ( .A(n4041), .B(n4040), .Z(n4042) );
  NANDN U5657 ( .A(n4043), .B(n4042), .Z(n4045) );
  OR U5658 ( .A(n4045), .B(n4044), .Z(n4046) );
  AND U5659 ( .A(n4047), .B(n4046), .Z(n4049) );
  NOR U5660 ( .A(n4049), .B(n4048), .Z(n4050) );
  NANDN U5661 ( .A(n4051), .B(n4050), .Z(n4052) );
  AND U5662 ( .A(n4053), .B(n4052), .Z(n4055) );
  NAND U5663 ( .A(n4055), .B(n4054), .Z(n4057) );
  ANDN U5664 ( .B(n4057), .A(n4056), .Z(n4058) );
  NANDN U5665 ( .A(n4059), .B(n4058), .Z(n4063) );
  AND U5666 ( .A(n4061), .B(n4060), .Z(n4062) );
  NAND U5667 ( .A(n4063), .B(n4062), .Z(n4064) );
  NANDN U5668 ( .A(n4065), .B(n4064), .Z(n4067) );
  OR U5669 ( .A(n4067), .B(n4066), .Z(n4068) );
  AND U5670 ( .A(n4069), .B(n4068), .Z(n4070) );
  NOR U5671 ( .A(n4071), .B(n4070), .Z(n4072) );
  NANDN U5672 ( .A(n4073), .B(n4072), .Z(n4074) );
  AND U5673 ( .A(n4075), .B(n4074), .Z(n4077) );
  NANDN U5674 ( .A(y[560]), .B(x[560]), .Z(n4076) );
  NAND U5675 ( .A(n4077), .B(n4076), .Z(n4079) );
  ANDN U5676 ( .B(n4079), .A(n4078), .Z(n4080) );
  NANDN U5677 ( .A(n4081), .B(n4080), .Z(n4082) );
  AND U5678 ( .A(n4083), .B(n4082), .Z(n4084) );
  NAND U5679 ( .A(n4085), .B(n4084), .Z(n4086) );
  NANDN U5680 ( .A(n4087), .B(n4086), .Z(n4089) );
  OR U5681 ( .A(n4089), .B(n4088), .Z(n4090) );
  AND U5682 ( .A(n4091), .B(n4090), .Z(n4093) );
  NOR U5683 ( .A(n4093), .B(n4092), .Z(n4094) );
  NANDN U5684 ( .A(n4095), .B(n4094), .Z(n4096) );
  AND U5685 ( .A(n4097), .B(n4096), .Z(n4099) );
  NAND U5686 ( .A(n4099), .B(n4098), .Z(n4101) );
  ANDN U5687 ( .B(n4101), .A(n4100), .Z(n4102) );
  NANDN U5688 ( .A(n4103), .B(n4102), .Z(n4107) );
  AND U5689 ( .A(n4105), .B(n4104), .Z(n4106) );
  NAND U5690 ( .A(n4107), .B(n4106), .Z(n4108) );
  NANDN U5691 ( .A(n4109), .B(n4108), .Z(n4110) );
  OR U5692 ( .A(n4111), .B(n4110), .Z(n4112) );
  AND U5693 ( .A(n4113), .B(n4112), .Z(n4115) );
  NAND U5694 ( .A(n4115), .B(n4114), .Z(n4117) );
  ANDN U5695 ( .B(n4117), .A(n4116), .Z(n4118) );
  NANDN U5696 ( .A(n4119), .B(n4118), .Z(n4123) );
  AND U5697 ( .A(n4121), .B(n4120), .Z(n4122) );
  NAND U5698 ( .A(n4123), .B(n4122), .Z(n4124) );
  NANDN U5699 ( .A(n4125), .B(n4124), .Z(n4128) );
  NANDN U5700 ( .A(x[574]), .B(n4128), .Z(n4127) );
  ANDN U5701 ( .B(n4127), .A(n4126), .Z(n4131) );
  XNOR U5702 ( .A(n4128), .B(x[574]), .Z(n4129) );
  NAND U5703 ( .A(n4129), .B(y[574]), .Z(n4130) );
  NAND U5704 ( .A(n4131), .B(n4130), .Z(n4132) );
  NAND U5705 ( .A(n6557), .B(n4132), .Z(n4133) );
  NANDN U5706 ( .A(n6558), .B(n4133), .Z(n4134) );
  AND U5707 ( .A(n4135), .B(n4134), .Z(n4136) );
  OR U5708 ( .A(n4137), .B(n4136), .Z(n4138) );
  AND U5709 ( .A(n4139), .B(n4138), .Z(n4140) );
  NOR U5710 ( .A(n4141), .B(n4140), .Z(n4142) );
  NANDN U5711 ( .A(n4143), .B(n4142), .Z(n4144) );
  AND U5712 ( .A(n4145), .B(n4144), .Z(n4147) );
  NANDN U5713 ( .A(y[580]), .B(x[580]), .Z(n4146) );
  NAND U5714 ( .A(n4147), .B(n4146), .Z(n4149) );
  ANDN U5715 ( .B(n4149), .A(n4148), .Z(n4150) );
  NANDN U5716 ( .A(n4151), .B(n4150), .Z(n4155) );
  NANDN U5717 ( .A(y[582]), .B(x[582]), .Z(n4152) );
  AND U5718 ( .A(n4153), .B(n4152), .Z(n4154) );
  NAND U5719 ( .A(n4155), .B(n4154), .Z(n4156) );
  NANDN U5720 ( .A(n4157), .B(n4156), .Z(n4159) );
  OR U5721 ( .A(n4159), .B(n4158), .Z(n4160) );
  AND U5722 ( .A(n4161), .B(n4160), .Z(n4162) );
  NOR U5723 ( .A(n4163), .B(n4162), .Z(n4164) );
  NANDN U5724 ( .A(n4165), .B(n4164), .Z(n4166) );
  AND U5725 ( .A(n4167), .B(n4166), .Z(n4169) );
  NANDN U5726 ( .A(y[586]), .B(x[586]), .Z(n4168) );
  NAND U5727 ( .A(n4169), .B(n4168), .Z(n4171) );
  ANDN U5728 ( .B(n4171), .A(n4170), .Z(n4172) );
  NANDN U5729 ( .A(n4173), .B(n4172), .Z(n4177) );
  AND U5730 ( .A(n4175), .B(n4174), .Z(n4176) );
  NAND U5731 ( .A(n4177), .B(n4176), .Z(n4178) );
  NANDN U5732 ( .A(n4179), .B(n4178), .Z(n4181) );
  OR U5733 ( .A(n4181), .B(n4180), .Z(n4182) );
  AND U5734 ( .A(n4183), .B(n4182), .Z(n4185) );
  NOR U5735 ( .A(n4185), .B(n4184), .Z(n4186) );
  NANDN U5736 ( .A(n4187), .B(n4186), .Z(n4188) );
  AND U5737 ( .A(n4189), .B(n4188), .Z(n4191) );
  NAND U5738 ( .A(n4191), .B(n4190), .Z(n4193) );
  ANDN U5739 ( .B(n4193), .A(n4192), .Z(n4194) );
  NANDN U5740 ( .A(n4195), .B(n4194), .Z(n4199) );
  AND U5741 ( .A(n4197), .B(n4196), .Z(n4198) );
  NAND U5742 ( .A(n4199), .B(n4198), .Z(n4200) );
  NANDN U5743 ( .A(n4201), .B(n4200), .Z(n4203) );
  OR U5744 ( .A(n4203), .B(n4202), .Z(n4204) );
  AND U5745 ( .A(n4205), .B(n4204), .Z(n4207) );
  NOR U5746 ( .A(n4207), .B(n4206), .Z(n4208) );
  NANDN U5747 ( .A(n4209), .B(n4208), .Z(n4210) );
  AND U5748 ( .A(n4211), .B(n4210), .Z(n4213) );
  NAND U5749 ( .A(n4213), .B(n4212), .Z(n4215) );
  ANDN U5750 ( .B(n4215), .A(n4214), .Z(n4216) );
  NANDN U5751 ( .A(n4217), .B(n4216), .Z(n4221) );
  AND U5752 ( .A(n4219), .B(n4218), .Z(n4220) );
  NAND U5753 ( .A(n4221), .B(n4220), .Z(n4222) );
  NANDN U5754 ( .A(n4223), .B(n4222), .Z(n4225) );
  OR U5755 ( .A(n4225), .B(n4224), .Z(n4226) );
  AND U5756 ( .A(n4227), .B(n4226), .Z(n4229) );
  NOR U5757 ( .A(n4229), .B(n4228), .Z(n4230) );
  NANDN U5758 ( .A(n4231), .B(n4230), .Z(n4232) );
  AND U5759 ( .A(n4233), .B(n4232), .Z(n4235) );
  NAND U5760 ( .A(n4235), .B(n4234), .Z(n4237) );
  ANDN U5761 ( .B(n4237), .A(n4236), .Z(n4238) );
  NANDN U5762 ( .A(n4239), .B(n4238), .Z(n4240) );
  AND U5763 ( .A(n4241), .B(n4240), .Z(n4242) );
  NAND U5764 ( .A(n4243), .B(n4242), .Z(n4244) );
  NANDN U5765 ( .A(n4245), .B(n4244), .Z(n4247) );
  OR U5766 ( .A(n4247), .B(n4246), .Z(n4248) );
  AND U5767 ( .A(n4249), .B(n4248), .Z(n4250) );
  NOR U5768 ( .A(n4251), .B(n4250), .Z(n4252) );
  NANDN U5769 ( .A(n4253), .B(n4252), .Z(n4254) );
  AND U5770 ( .A(n4255), .B(n4254), .Z(n4257) );
  NANDN U5771 ( .A(y[610]), .B(x[610]), .Z(n4256) );
  NAND U5772 ( .A(n4257), .B(n4256), .Z(n4259) );
  ANDN U5773 ( .B(n4259), .A(n4258), .Z(n4260) );
  NANDN U5774 ( .A(n4261), .B(n4260), .Z(n4265) );
  AND U5775 ( .A(n4263), .B(n4262), .Z(n4264) );
  NAND U5776 ( .A(n4265), .B(n4264), .Z(n4266) );
  NANDN U5777 ( .A(n4267), .B(n4266), .Z(n4269) );
  OR U5778 ( .A(n4269), .B(n4268), .Z(n4270) );
  AND U5779 ( .A(n4271), .B(n4270), .Z(n4272) );
  NOR U5780 ( .A(n4273), .B(n4272), .Z(n4274) );
  NANDN U5781 ( .A(n4275), .B(n4274), .Z(n4276) );
  AND U5782 ( .A(n4277), .B(n4276), .Z(n4279) );
  NANDN U5783 ( .A(y[616]), .B(x[616]), .Z(n4278) );
  NAND U5784 ( .A(n4279), .B(n4278), .Z(n4281) );
  ANDN U5785 ( .B(n4281), .A(n4280), .Z(n4282) );
  NANDN U5786 ( .A(n4283), .B(n4282), .Z(n4287) );
  AND U5787 ( .A(n4285), .B(n4284), .Z(n4286) );
  NAND U5788 ( .A(n4287), .B(n4286), .Z(n4288) );
  NANDN U5789 ( .A(n4289), .B(n4288), .Z(n4291) );
  OR U5790 ( .A(n4291), .B(n4290), .Z(n4292) );
  AND U5791 ( .A(n4293), .B(n4292), .Z(n4295) );
  NOR U5792 ( .A(n4295), .B(n4294), .Z(n4296) );
  NANDN U5793 ( .A(n4297), .B(n4296), .Z(n4298) );
  AND U5794 ( .A(n4299), .B(n4298), .Z(n4301) );
  NAND U5795 ( .A(n4301), .B(n4300), .Z(n4303) );
  ANDN U5796 ( .B(n4303), .A(n4302), .Z(n4304) );
  NANDN U5797 ( .A(n4305), .B(n4304), .Z(n4306) );
  AND U5798 ( .A(n4307), .B(n4306), .Z(n4308) );
  NAND U5799 ( .A(n4309), .B(n4308), .Z(n4310) );
  NANDN U5800 ( .A(n4311), .B(n4310), .Z(n4313) );
  OR U5801 ( .A(n4313), .B(n4312), .Z(n4314) );
  AND U5802 ( .A(n4315), .B(n4314), .Z(n4317) );
  NOR U5803 ( .A(n4317), .B(n4316), .Z(n4318) );
  NANDN U5804 ( .A(n4319), .B(n4318), .Z(n4320) );
  AND U5805 ( .A(n4321), .B(n4320), .Z(n4323) );
  NAND U5806 ( .A(n4323), .B(n4322), .Z(n4325) );
  ANDN U5807 ( .B(n4325), .A(n4324), .Z(n4326) );
  NANDN U5808 ( .A(n4327), .B(n4326), .Z(n4328) );
  AND U5809 ( .A(n4329), .B(n4328), .Z(n4330) );
  NAND U5810 ( .A(n4331), .B(n4330), .Z(n4332) );
  NANDN U5811 ( .A(n4333), .B(n4332), .Z(n4335) );
  OR U5812 ( .A(n4335), .B(n4334), .Z(n4336) );
  AND U5813 ( .A(n4337), .B(n4336), .Z(n4339) );
  NOR U5814 ( .A(n4339), .B(n4338), .Z(n4340) );
  NANDN U5815 ( .A(n4341), .B(n4340), .Z(n4342) );
  AND U5816 ( .A(n4343), .B(n4342), .Z(n4345) );
  NAND U5817 ( .A(n4345), .B(n4344), .Z(n4347) );
  ANDN U5818 ( .B(n4347), .A(n4346), .Z(n4348) );
  NANDN U5819 ( .A(n4349), .B(n4348), .Z(n4353) );
  AND U5820 ( .A(n4351), .B(n4350), .Z(n4352) );
  NAND U5821 ( .A(n4353), .B(n4352), .Z(n4354) );
  NANDN U5822 ( .A(n4355), .B(n4354), .Z(n4357) );
  OR U5823 ( .A(n4357), .B(n4356), .Z(n4358) );
  AND U5824 ( .A(n4359), .B(n4358), .Z(n4361) );
  NOR U5825 ( .A(n4361), .B(n4360), .Z(n4362) );
  NANDN U5826 ( .A(n4363), .B(n4362), .Z(n4364) );
  AND U5827 ( .A(n4365), .B(n4364), .Z(n4367) );
  NAND U5828 ( .A(n4367), .B(n4366), .Z(n4369) );
  ANDN U5829 ( .B(n4369), .A(n4368), .Z(n4370) );
  NANDN U5830 ( .A(n4371), .B(n4370), .Z(n4375) );
  AND U5831 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U5832 ( .A(n4375), .B(n4374), .Z(n4376) );
  NANDN U5833 ( .A(n4377), .B(n4376), .Z(n4379) );
  OR U5834 ( .A(n4379), .B(n4378), .Z(n4380) );
  AND U5835 ( .A(n4381), .B(n4380), .Z(n4382) );
  NOR U5836 ( .A(n4383), .B(n4382), .Z(n4384) );
  NANDN U5837 ( .A(n4385), .B(n4384), .Z(n4386) );
  AND U5838 ( .A(n4387), .B(n4386), .Z(n4389) );
  NANDN U5839 ( .A(y[646]), .B(x[646]), .Z(n4388) );
  NAND U5840 ( .A(n4389), .B(n4388), .Z(n4391) );
  ANDN U5841 ( .B(n4391), .A(n4390), .Z(n4392) );
  NANDN U5842 ( .A(n4393), .B(n4392), .Z(n4397) );
  NANDN U5843 ( .A(y[648]), .B(x[648]), .Z(n4394) );
  AND U5844 ( .A(n4395), .B(n4394), .Z(n4396) );
  NAND U5845 ( .A(n4397), .B(n4396), .Z(n4398) );
  NANDN U5846 ( .A(n4399), .B(n4398), .Z(n4400) );
  OR U5847 ( .A(n4401), .B(n4400), .Z(n4402) );
  AND U5848 ( .A(n4403), .B(n4402), .Z(n4405) );
  NANDN U5849 ( .A(y[650]), .B(x[650]), .Z(n4404) );
  NAND U5850 ( .A(n4405), .B(n4404), .Z(n4407) );
  ANDN U5851 ( .B(n4407), .A(n4406), .Z(n4408) );
  NANDN U5852 ( .A(n4409), .B(n4408), .Z(n4413) );
  AND U5853 ( .A(n4411), .B(n4410), .Z(n4412) );
  NAND U5854 ( .A(n4413), .B(n4412), .Z(n4414) );
  NANDN U5855 ( .A(n4415), .B(n4414), .Z(n4416) );
  OR U5856 ( .A(n4416), .B(n6706), .Z(n4417) );
  AND U5857 ( .A(n4418), .B(n4417), .Z(n4421) );
  NAND U5858 ( .A(n4420), .B(n4419), .Z(n5425) );
  OR U5859 ( .A(n4421), .B(n5425), .Z(n4422) );
  NAND U5860 ( .A(n6708), .B(n4422), .Z(n4423) );
  NANDN U5861 ( .A(n4424), .B(n4423), .Z(n4425) );
  OR U5862 ( .A(n6709), .B(n4425), .Z(n4426) );
  AND U5863 ( .A(n4427), .B(n4426), .Z(n4428) );
  NAND U5864 ( .A(n4428), .B(n6710), .Z(n4430) );
  ANDN U5865 ( .B(n4430), .A(n4429), .Z(n4431) );
  NANDN U5866 ( .A(n4432), .B(n4431), .Z(n4436) );
  AND U5867 ( .A(n4434), .B(n4433), .Z(n4435) );
  NAND U5868 ( .A(n4436), .B(n4435), .Z(n4437) );
  NANDN U5869 ( .A(n4438), .B(n4437), .Z(n4440) );
  OR U5870 ( .A(n4440), .B(n4439), .Z(n4441) );
  AND U5871 ( .A(n4442), .B(n4441), .Z(n4444) );
  NOR U5872 ( .A(n4444), .B(n4443), .Z(n4445) );
  NANDN U5873 ( .A(n4446), .B(n4445), .Z(n4447) );
  AND U5874 ( .A(n4448), .B(n4447), .Z(n4450) );
  AND U5875 ( .A(n4450), .B(n4449), .Z(n4454) );
  AND U5876 ( .A(n4452), .B(n4451), .Z(n4453) );
  NANDN U5877 ( .A(n4454), .B(n4453), .Z(n4455) );
  NAND U5878 ( .A(n4456), .B(n4455), .Z(n4460) );
  AND U5879 ( .A(n4458), .B(n4457), .Z(n4459) );
  NAND U5880 ( .A(n4460), .B(n4459), .Z(n4461) );
  NANDN U5881 ( .A(n4462), .B(n4461), .Z(n4464) );
  OR U5882 ( .A(n4464), .B(n4463), .Z(n4465) );
  NAND U5883 ( .A(n4466), .B(n4465), .Z(n4467) );
  NANDN U5884 ( .A(n4468), .B(n4467), .Z(n4472) );
  AND U5885 ( .A(n4470), .B(n4469), .Z(n4471) );
  NAND U5886 ( .A(n4472), .B(n4471), .Z(n4473) );
  NANDN U5887 ( .A(n4474), .B(n4473), .Z(n4475) );
  OR U5888 ( .A(n4476), .B(n4475), .Z(n4477) );
  AND U5889 ( .A(n4478), .B(n4477), .Z(n4479) );
  NANDN U5890 ( .A(n4480), .B(n4479), .Z(n4481) );
  NAND U5891 ( .A(n4482), .B(n4481), .Z(n4486) );
  AND U5892 ( .A(n4484), .B(n4483), .Z(n4485) );
  NAND U5893 ( .A(n4486), .B(n4485), .Z(n4487) );
  NANDN U5894 ( .A(n4488), .B(n4487), .Z(n4489) );
  OR U5895 ( .A(n4490), .B(n4489), .Z(n4491) );
  AND U5896 ( .A(n4492), .B(n4491), .Z(n4494) );
  NAND U5897 ( .A(n4494), .B(n4493), .Z(n4496) );
  AND U5898 ( .A(n4496), .B(n4495), .Z(n4498) );
  NANDN U5899 ( .A(y[678]), .B(x[678]), .Z(n4497) );
  NAND U5900 ( .A(n4498), .B(n4497), .Z(n4499) );
  NAND U5901 ( .A(n4500), .B(n4499), .Z(n4502) );
  OR U5902 ( .A(n4502), .B(n4501), .Z(n4503) );
  AND U5903 ( .A(n4504), .B(n4503), .Z(n4508) );
  NAND U5904 ( .A(n4506), .B(n4505), .Z(n4507) );
  OR U5905 ( .A(n4508), .B(n4507), .Z(n4509) );
  AND U5906 ( .A(n4510), .B(n4509), .Z(n4511) );
  NANDN U5907 ( .A(n4512), .B(n4511), .Z(n4513) );
  AND U5908 ( .A(n4514), .B(n4513), .Z(n4516) );
  NAND U5909 ( .A(n4516), .B(n4515), .Z(n4518) );
  ANDN U5910 ( .B(x[684]), .A(y[684]), .Z(n4517) );
  ANDN U5911 ( .B(n4518), .A(n4517), .Z(n4519) );
  NANDN U5912 ( .A(n4520), .B(n4519), .Z(n4524) );
  AND U5913 ( .A(n4522), .B(n4521), .Z(n4523) );
  NAND U5914 ( .A(n4524), .B(n4523), .Z(n4525) );
  NANDN U5915 ( .A(n4526), .B(n4525), .Z(n4528) );
  OR U5916 ( .A(n4528), .B(n4527), .Z(n4529) );
  AND U5917 ( .A(n4530), .B(n4529), .Z(n4532) );
  ANDN U5918 ( .B(x[688]), .A(y[688]), .Z(n4531) );
  NOR U5919 ( .A(n4532), .B(n4531), .Z(n4533) );
  NANDN U5920 ( .A(n4534), .B(n4533), .Z(n4535) );
  AND U5921 ( .A(n4536), .B(n4535), .Z(n4537) );
  NAND U5922 ( .A(n4538), .B(n4537), .Z(n4539) );
  NAND U5923 ( .A(n4540), .B(n4539), .Z(n4541) );
  AND U5924 ( .A(n4542), .B(n4541), .Z(n4543) );
  OR U5925 ( .A(n4544), .B(n4543), .Z(n4545) );
  AND U5926 ( .A(n4546), .B(n4545), .Z(n4547) );
  ANDN U5927 ( .B(n4548), .A(n4547), .Z(n4549) );
  NAND U5928 ( .A(n4550), .B(n4549), .Z(n4551) );
  NANDN U5929 ( .A(n4552), .B(n4551), .Z(n4554) );
  OR U5930 ( .A(n4554), .B(n4553), .Z(n4555) );
  NAND U5931 ( .A(n4556), .B(n4555), .Z(n4557) );
  NANDN U5932 ( .A(n4558), .B(n4557), .Z(n4562) );
  AND U5933 ( .A(n4560), .B(n4559), .Z(n4561) );
  NAND U5934 ( .A(n4562), .B(n4561), .Z(n4563) );
  NANDN U5935 ( .A(n4564), .B(n4563), .Z(n4566) );
  OR U5936 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U5937 ( .A(n4568), .B(n4567), .Z(n4569) );
  NANDN U5938 ( .A(n4570), .B(n4569), .Z(n4571) );
  AND U5939 ( .A(n4572), .B(n4571), .Z(n4573) );
  NAND U5940 ( .A(n4574), .B(n4573), .Z(n4575) );
  NANDN U5941 ( .A(n4576), .B(n4575), .Z(n4577) );
  OR U5942 ( .A(n4578), .B(n4577), .Z(n4579) );
  AND U5943 ( .A(n4580), .B(n4579), .Z(n4581) );
  NANDN U5944 ( .A(n4582), .B(n4581), .Z(n4583) );
  AND U5945 ( .A(n4584), .B(n4583), .Z(n4585) );
  ANDN U5946 ( .B(n4586), .A(n4585), .Z(n4587) );
  NAND U5947 ( .A(n4588), .B(n4587), .Z(n4589) );
  NANDN U5948 ( .A(n4590), .B(n4589), .Z(n4591) );
  OR U5949 ( .A(n4592), .B(n4591), .Z(n4593) );
  AND U5950 ( .A(n4594), .B(n4593), .Z(n4596) );
  NANDN U5951 ( .A(y[706]), .B(x[706]), .Z(n4595) );
  NAND U5952 ( .A(n4596), .B(n4595), .Z(n4598) );
  ANDN U5953 ( .B(n4598), .A(n4597), .Z(n4599) );
  NANDN U5954 ( .A(n4600), .B(n4599), .Z(n4604) );
  NANDN U5955 ( .A(y[708]), .B(x[708]), .Z(n4601) );
  AND U5956 ( .A(n4602), .B(n4601), .Z(n4603) );
  NAND U5957 ( .A(n4604), .B(n4603), .Z(n4605) );
  NANDN U5958 ( .A(n4606), .B(n4605), .Z(n4608) );
  OR U5959 ( .A(n4608), .B(n4607), .Z(n4609) );
  NAND U5960 ( .A(n4610), .B(n4609), .Z(n4614) );
  AND U5961 ( .A(n4612), .B(n4611), .Z(n4613) );
  NAND U5962 ( .A(n4614), .B(n4613), .Z(n4615) );
  NANDN U5963 ( .A(n4616), .B(n4615), .Z(n4617) );
  OR U5964 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U5965 ( .A(n4620), .B(n4619), .Z(n4622) );
  NAND U5966 ( .A(n4622), .B(n4621), .Z(n4624) );
  AND U5967 ( .A(n4624), .B(n4623), .Z(n4626) );
  NANDN U5968 ( .A(y[714]), .B(x[714]), .Z(n4625) );
  NAND U5969 ( .A(n4626), .B(n4625), .Z(n4627) );
  NANDN U5970 ( .A(n4628), .B(n4627), .Z(n4629) );
  AND U5971 ( .A(n4630), .B(n4629), .Z(n4632) );
  NAND U5972 ( .A(n4632), .B(n4631), .Z(n4634) );
  ANDN U5973 ( .B(n4634), .A(n4633), .Z(n4635) );
  NANDN U5974 ( .A(n4636), .B(n4635), .Z(n4640) );
  NANDN U5975 ( .A(y[718]), .B(x[718]), .Z(n4637) );
  AND U5976 ( .A(n4638), .B(n4637), .Z(n4639) );
  NAND U5977 ( .A(n4640), .B(n4639), .Z(n4641) );
  NANDN U5978 ( .A(n4642), .B(n4641), .Z(n4645) );
  NAND U5979 ( .A(n4645), .B(y[720]), .Z(n4643) );
  AND U5980 ( .A(n4644), .B(n4643), .Z(n4648) );
  XOR U5981 ( .A(n4645), .B(y[720]), .Z(n4646) );
  NANDN U5982 ( .A(x[720]), .B(n4646), .Z(n4647) );
  AND U5983 ( .A(n4648), .B(n4647), .Z(n4649) );
  OR U5984 ( .A(n4650), .B(n4649), .Z(n4651) );
  AND U5985 ( .A(n4652), .B(n4651), .Z(n4653) );
  ANDN U5986 ( .B(n4654), .A(n4653), .Z(n4655) );
  NAND U5987 ( .A(n4656), .B(n4655), .Z(n4657) );
  NANDN U5988 ( .A(n4658), .B(n4657), .Z(n4659) );
  OR U5989 ( .A(n4659), .B(n6839), .Z(n4665) );
  OR U5990 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U5991 ( .A(n4663), .B(n4662), .Z(n4664) );
  ANDN U5992 ( .B(n4665), .A(n4664), .Z(n4666) );
  OR U5993 ( .A(n4667), .B(n4666), .Z(n4668) );
  AND U5994 ( .A(n4669), .B(n4668), .Z(n4670) );
  NOR U5995 ( .A(n4671), .B(n4670), .Z(n4672) );
  NANDN U5996 ( .A(n4673), .B(n4672), .Z(n4674) );
  AND U5997 ( .A(n4675), .B(n4674), .Z(n4677) );
  NANDN U5998 ( .A(y[728]), .B(x[728]), .Z(n4676) );
  NAND U5999 ( .A(n4677), .B(n4676), .Z(n4679) );
  ANDN U6000 ( .B(n4679), .A(n4678), .Z(n4680) );
  NANDN U6001 ( .A(n4681), .B(n4680), .Z(n4682) );
  AND U6002 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U6003 ( .A(n4685), .B(n4684), .Z(n4686) );
  NANDN U6004 ( .A(n4687), .B(n4686), .Z(n4689) );
  OR U6005 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U6006 ( .A(n4691), .B(n4690), .Z(n4695) );
  AND U6007 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U6008 ( .A(n4695), .B(n4694), .Z(n4696) );
  NANDN U6009 ( .A(n4697), .B(n4696), .Z(n4699) );
  OR U6010 ( .A(n4699), .B(n4698), .Z(n4700) );
  NAND U6011 ( .A(n4701), .B(n4700), .Z(n4702) );
  NANDN U6012 ( .A(n4703), .B(n4702), .Z(n4707) );
  AND U6013 ( .A(n4705), .B(n4704), .Z(n4706) );
  NAND U6014 ( .A(n4707), .B(n4706), .Z(n4708) );
  NANDN U6015 ( .A(n4709), .B(n4708), .Z(n4711) );
  OR U6016 ( .A(n4711), .B(n4710), .Z(n4712) );
  NAND U6017 ( .A(n4713), .B(n4712), .Z(n4714) );
  NANDN U6018 ( .A(n4715), .B(n4714), .Z(n4719) );
  AND U6019 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U6020 ( .A(n4719), .B(n4718), .Z(n4720) );
  NANDN U6021 ( .A(n4721), .B(n4720), .Z(n4722) );
  OR U6022 ( .A(n4723), .B(n4722), .Z(n4724) );
  AND U6023 ( .A(n4725), .B(n4724), .Z(n4727) );
  NAND U6024 ( .A(n4727), .B(n4726), .Z(n4729) );
  ANDN U6025 ( .B(n4729), .A(n4728), .Z(n4730) );
  NANDN U6026 ( .A(n4731), .B(n4730), .Z(n4735) );
  AND U6027 ( .A(n4733), .B(n4732), .Z(n4734) );
  NAND U6028 ( .A(n4735), .B(n4734), .Z(n4736) );
  NANDN U6029 ( .A(n4737), .B(n4736), .Z(n4739) );
  ANDN U6030 ( .B(x[746]), .A(y[746]), .Z(n4738) );
  OR U6031 ( .A(n4739), .B(n4738), .Z(n4740) );
  NAND U6032 ( .A(n4741), .B(n4740), .Z(n4745) );
  NANDN U6033 ( .A(y[748]), .B(x[748]), .Z(n4742) );
  AND U6034 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U6035 ( .A(n4745), .B(n4744), .Z(n4746) );
  NANDN U6036 ( .A(n4747), .B(n4746), .Z(n4748) );
  OR U6037 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U6038 ( .A(n4751), .B(n4750), .Z(n4752) );
  NANDN U6039 ( .A(n4753), .B(n4752), .Z(n4754) );
  AND U6040 ( .A(n4755), .B(n4754), .Z(n4756) );
  ANDN U6041 ( .B(n4757), .A(n4756), .Z(n4758) );
  NAND U6042 ( .A(n4759), .B(n4758), .Z(n4760) );
  NANDN U6043 ( .A(n4761), .B(n4760), .Z(n4762) );
  OR U6044 ( .A(n4763), .B(n4762), .Z(n4764) );
  AND U6045 ( .A(n4765), .B(n4764), .Z(n4766) );
  NANDN U6046 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U6047 ( .A(n4769), .B(n4768), .Z(n4771) );
  NOR U6048 ( .A(n4771), .B(n4770), .Z(n4772) );
  NANDN U6049 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U6050 ( .A(n4775), .B(n4774), .Z(n4777) );
  AND U6051 ( .A(n4777), .B(n4776), .Z(n4781) );
  AND U6052 ( .A(n4779), .B(n4778), .Z(n4780) );
  NANDN U6053 ( .A(n4781), .B(n4780), .Z(n4782) );
  NANDN U6054 ( .A(n4783), .B(n4782), .Z(n4784) );
  AND U6055 ( .A(n4785), .B(n4784), .Z(n4787) );
  NANDN U6056 ( .A(y[760]), .B(x[760]), .Z(n4786) );
  NAND U6057 ( .A(n4787), .B(n4786), .Z(n4789) );
  ANDN U6058 ( .B(n4789), .A(n4788), .Z(n4790) );
  NANDN U6059 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U6060 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U6061 ( .A(n4795), .B(n4794), .Z(n4796) );
  NANDN U6062 ( .A(n4797), .B(n4796), .Z(n4799) );
  OR U6063 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U6064 ( .A(n4801), .B(n4800), .Z(n4805) );
  AND U6065 ( .A(n4803), .B(n4802), .Z(n4804) );
  NAND U6066 ( .A(n4805), .B(n4804), .Z(n4806) );
  NANDN U6067 ( .A(n4807), .B(n4806), .Z(n4808) );
  OR U6068 ( .A(n4809), .B(n4808), .Z(n4810) );
  AND U6069 ( .A(n4811), .B(n4810), .Z(n4812) );
  NANDN U6070 ( .A(n4813), .B(n4812), .Z(n4814) );
  AND U6071 ( .A(n4815), .B(n4814), .Z(n4817) );
  NOR U6072 ( .A(n4817), .B(n4816), .Z(n4818) );
  NANDN U6073 ( .A(n4819), .B(n4818), .Z(n4820) );
  AND U6074 ( .A(n4821), .B(n4820), .Z(n4823) );
  AND U6075 ( .A(n4823), .B(n4822), .Z(n4827) );
  AND U6076 ( .A(n4825), .B(n4824), .Z(n4826) );
  NANDN U6077 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U6078 ( .A(n4829), .B(n4828), .Z(n4833) );
  AND U6079 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U6080 ( .A(n4833), .B(n4832), .Z(n4834) );
  NANDN U6081 ( .A(n4835), .B(n4834), .Z(n4836) );
  OR U6082 ( .A(n4837), .B(n4836), .Z(n4838) );
  AND U6083 ( .A(n4839), .B(n4838), .Z(n4841) );
  NAND U6084 ( .A(n4841), .B(n4840), .Z(n4843) );
  ANDN U6085 ( .B(n4843), .A(n4842), .Z(n4844) );
  NANDN U6086 ( .A(n4845), .B(n4844), .Z(n4849) );
  AND U6087 ( .A(n4847), .B(n4846), .Z(n4848) );
  NAND U6088 ( .A(n4849), .B(n4848), .Z(n4850) );
  NANDN U6089 ( .A(n4851), .B(n4850), .Z(n4853) );
  OR U6090 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U6091 ( .A(n4855), .B(n4854), .Z(n4856) );
  AND U6092 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U6093 ( .A(n4859), .B(n4858), .Z(n4860) );
  NANDN U6094 ( .A(n4861), .B(n4860), .Z(n4862) );
  OR U6095 ( .A(n4863), .B(n4862), .Z(n4864) );
  AND U6096 ( .A(n4865), .B(n4864), .Z(n4866) );
  NANDN U6097 ( .A(n4867), .B(n4866), .Z(n4868) );
  AND U6098 ( .A(n4869), .B(n4868), .Z(n4871) );
  NAND U6099 ( .A(n4871), .B(n4870), .Z(n4873) );
  ANDN U6100 ( .B(n4873), .A(n4872), .Z(n4874) );
  NANDN U6101 ( .A(n4875), .B(n4874), .Z(n4879) );
  AND U6102 ( .A(n4877), .B(n4876), .Z(n4878) );
  NAND U6103 ( .A(n4879), .B(n4878), .Z(n4880) );
  NANDN U6104 ( .A(n4881), .B(n4880), .Z(n4883) );
  OR U6105 ( .A(n4883), .B(n4882), .Z(n4884) );
  NAND U6106 ( .A(n4885), .B(n4884), .Z(n4886) );
  AND U6107 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U6108 ( .A(n4889), .B(n4888), .Z(n4890) );
  NANDN U6109 ( .A(n4891), .B(n4890), .Z(n4892) );
  OR U6110 ( .A(n4893), .B(n4892), .Z(n4894) );
  AND U6111 ( .A(n4895), .B(n4894), .Z(n4896) );
  NANDN U6112 ( .A(n4897), .B(n4896), .Z(n4898) );
  AND U6113 ( .A(n4899), .B(n4898), .Z(n4901) );
  NAND U6114 ( .A(n4901), .B(n4900), .Z(n4903) );
  ANDN U6115 ( .B(n4903), .A(n4902), .Z(n4904) );
  NANDN U6116 ( .A(n4905), .B(n4904), .Z(n4909) );
  AND U6117 ( .A(n4907), .B(n4906), .Z(n4908) );
  NAND U6118 ( .A(n4909), .B(n4908), .Z(n4910) );
  NANDN U6119 ( .A(n4911), .B(n4910), .Z(n4913) );
  OR U6120 ( .A(n4913), .B(n4912), .Z(n4914) );
  NAND U6121 ( .A(n4915), .B(n4914), .Z(n4916) );
  AND U6122 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U6123 ( .A(n4919), .B(n4918), .Z(n4920) );
  NANDN U6124 ( .A(n4921), .B(n4920), .Z(n4922) );
  OR U6125 ( .A(n4923), .B(n4922), .Z(n4924) );
  AND U6126 ( .A(n4925), .B(n4924), .Z(n4926) );
  NANDN U6127 ( .A(n4927), .B(n4926), .Z(n4928) );
  AND U6128 ( .A(n4929), .B(n4928), .Z(n4931) );
  NAND U6129 ( .A(n4931), .B(n4930), .Z(n4933) );
  ANDN U6130 ( .B(x[800]), .A(y[800]), .Z(n4932) );
  ANDN U6131 ( .B(n4933), .A(n4932), .Z(n4934) );
  NANDN U6132 ( .A(n4935), .B(n4934), .Z(n4939) );
  AND U6133 ( .A(n4937), .B(n4936), .Z(n4938) );
  NAND U6134 ( .A(n4939), .B(n4938), .Z(n4940) );
  NANDN U6135 ( .A(n4941), .B(n4940), .Z(n4943) );
  OR U6136 ( .A(n4943), .B(n4942), .Z(n4944) );
  NAND U6137 ( .A(n4945), .B(n4944), .Z(n4949) );
  NANDN U6138 ( .A(y[804]), .B(x[804]), .Z(n4946) );
  AND U6139 ( .A(n4947), .B(n4946), .Z(n4948) );
  NAND U6140 ( .A(n4949), .B(n4948), .Z(n4950) );
  NANDN U6141 ( .A(n4951), .B(n4950), .Z(n4952) );
  OR U6142 ( .A(n4953), .B(n4952), .Z(n4954) );
  AND U6143 ( .A(n4955), .B(n4954), .Z(n4957) );
  NANDN U6144 ( .A(y[806]), .B(x[806]), .Z(n4956) );
  NAND U6145 ( .A(n4957), .B(n4956), .Z(n4959) );
  ANDN U6146 ( .B(n4959), .A(n4958), .Z(n4960) );
  NANDN U6147 ( .A(n4961), .B(n4960), .Z(n4965) );
  NANDN U6148 ( .A(y[808]), .B(x[808]), .Z(n4962) );
  AND U6149 ( .A(n4963), .B(n4962), .Z(n4964) );
  NAND U6150 ( .A(n4965), .B(n4964), .Z(n4966) );
  NANDN U6151 ( .A(n4967), .B(n4966), .Z(n4969) );
  OR U6152 ( .A(n4969), .B(n4968), .Z(n4970) );
  AND U6153 ( .A(n4971), .B(n4970), .Z(n4973) );
  NOR U6154 ( .A(n4973), .B(n4972), .Z(n4974) );
  NANDN U6155 ( .A(n4975), .B(n4974), .Z(n4976) );
  AND U6156 ( .A(n4977), .B(n4976), .Z(n4979) );
  AND U6157 ( .A(n4979), .B(n4978), .Z(n4983) );
  AND U6158 ( .A(n4981), .B(n4980), .Z(n4982) );
  NANDN U6159 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U6160 ( .A(n4985), .B(n4984), .Z(n4989) );
  AND U6161 ( .A(n4987), .B(n4986), .Z(n4988) );
  NAND U6162 ( .A(n4989), .B(n4988), .Z(n4990) );
  NANDN U6163 ( .A(n4991), .B(n4990), .Z(n4992) );
  OR U6164 ( .A(n4993), .B(n4992), .Z(n4994) );
  AND U6165 ( .A(n4995), .B(n4994), .Z(n4997) );
  NAND U6166 ( .A(n4997), .B(n4996), .Z(n4999) );
  ANDN U6167 ( .B(n4999), .A(n4998), .Z(n5000) );
  NANDN U6168 ( .A(n5001), .B(n5000), .Z(n5005) );
  AND U6169 ( .A(n5003), .B(n5002), .Z(n5004) );
  NAND U6170 ( .A(n5005), .B(n5004), .Z(n5006) );
  NANDN U6171 ( .A(n5007), .B(n5006), .Z(n5009) );
  OR U6172 ( .A(n5009), .B(n5008), .Z(n5010) );
  NAND U6173 ( .A(n5011), .B(n5010), .Z(n5014) );
  AND U6174 ( .A(n5012), .B(n7037), .Z(n5013) );
  NAND U6175 ( .A(n5014), .B(n5013), .Z(n5015) );
  NANDN U6176 ( .A(n5016), .B(n5015), .Z(n5017) );
  OR U6177 ( .A(n5017), .B(n7038), .Z(n5018) );
  NAND U6178 ( .A(n7039), .B(n5018), .Z(n5019) );
  NANDN U6179 ( .A(n7040), .B(n5019), .Z(n5020) );
  NAND U6180 ( .A(n7041), .B(n5020), .Z(n5021) );
  ANDN U6181 ( .B(n5021), .A(n5423), .Z(n5022) );
  NANDN U6182 ( .A(n5023), .B(n5022), .Z(n5024) );
  NAND U6183 ( .A(n7042), .B(n5024), .Z(n5025) );
  NANDN U6184 ( .A(n5422), .B(n5025), .Z(n5026) );
  AND U6185 ( .A(n7043), .B(n5026), .Z(n5027) );
  OR U6186 ( .A(n7044), .B(n5027), .Z(n5028) );
  AND U6187 ( .A(n7045), .B(n5028), .Z(n5031) );
  NAND U6188 ( .A(n5029), .B(n7046), .Z(n5030) );
  OR U6189 ( .A(n5031), .B(n5030), .Z(n5032) );
  AND U6190 ( .A(n7048), .B(n5032), .Z(n5033) );
  ANDN U6191 ( .B(n5034), .A(n5033), .Z(n5035) );
  NAND U6192 ( .A(n7049), .B(n5035), .Z(n5036) );
  NANDN U6193 ( .A(n5037), .B(n5036), .Z(n5038) );
  OR U6194 ( .A(n7050), .B(n5038), .Z(n5039) );
  AND U6195 ( .A(n5040), .B(n5039), .Z(n5042) );
  NAND U6196 ( .A(n5042), .B(n5041), .Z(n5044) );
  ANDN U6197 ( .B(x[838]), .A(y[838]), .Z(n5043) );
  ANDN U6198 ( .B(n5044), .A(n5043), .Z(n5045) );
  NANDN U6199 ( .A(n7055), .B(n5045), .Z(n5048) );
  AND U6200 ( .A(n5046), .B(n7056), .Z(n5047) );
  NAND U6201 ( .A(n5048), .B(n5047), .Z(n5049) );
  NANDN U6202 ( .A(n7057), .B(n5049), .Z(n5050) );
  NAND U6203 ( .A(n7058), .B(n5050), .Z(n5051) );
  NAND U6204 ( .A(n7059), .B(n5051), .Z(n5052) );
  AND U6205 ( .A(n7060), .B(n5052), .Z(n5053) );
  OR U6206 ( .A(n7061), .B(n5053), .Z(n5054) );
  NAND U6207 ( .A(n7062), .B(n5054), .Z(n5055) );
  NANDN U6208 ( .A(n7063), .B(n5055), .Z(n5056) );
  NANDN U6209 ( .A(n5421), .B(n5056), .Z(n5057) );
  AND U6210 ( .A(n5058), .B(n5057), .Z(n5059) );
  NANDN U6211 ( .A(n7065), .B(n5059), .Z(n5060) );
  NAND U6212 ( .A(n5061), .B(n5060), .Z(n5062) );
  NANDN U6213 ( .A(n5063), .B(n5062), .Z(n5064) );
  OR U6214 ( .A(n5065), .B(n5064), .Z(n5066) );
  AND U6215 ( .A(n5067), .B(n5066), .Z(n5068) );
  NANDN U6216 ( .A(n5069), .B(n5068), .Z(n5070) );
  AND U6217 ( .A(n5071), .B(n5070), .Z(n5072) );
  NOR U6218 ( .A(n7070), .B(n5072), .Z(n5073) );
  NANDN U6219 ( .A(n5074), .B(n5073), .Z(n5075) );
  AND U6220 ( .A(n7073), .B(n5075), .Z(n5078) );
  ANDN U6221 ( .B(n5077), .A(n5076), .Z(n7076) );
  NANDN U6222 ( .A(n5078), .B(n7076), .Z(n5079) );
  NAND U6223 ( .A(n5420), .B(n5079), .Z(n5080) );
  NAND U6224 ( .A(n7080), .B(n5080), .Z(n5081) );
  NANDN U6225 ( .A(n7082), .B(n5081), .Z(n5082) );
  AND U6226 ( .A(n7084), .B(n5082), .Z(n5086) );
  OR U6227 ( .A(n5086), .B(n7085), .Z(n5087) );
  NAND U6228 ( .A(n7088), .B(n5087), .Z(n5088) );
  NANDN U6229 ( .A(n7091), .B(n5088), .Z(n5091) );
  AND U6230 ( .A(n5089), .B(n5419), .Z(n5090) );
  NAND U6231 ( .A(n5091), .B(n5090), .Z(n5092) );
  NANDN U6232 ( .A(n5415), .B(n5092), .Z(n5095) );
  AND U6233 ( .A(n5093), .B(n5416), .Z(n5094) );
  NAND U6234 ( .A(n5095), .B(n5094), .Z(n5096) );
  NANDN U6235 ( .A(n5097), .B(n5096), .Z(n5099) );
  IV U6236 ( .A(n5098), .Z(n7097) );
  OR U6237 ( .A(n5099), .B(n7097), .Z(n5100) );
  NAND U6238 ( .A(n5101), .B(n5100), .Z(n5102) );
  NANDN U6239 ( .A(n5103), .B(n5102), .Z(n5105) );
  IV U6240 ( .A(n5104), .Z(n7105) );
  OR U6241 ( .A(n5105), .B(n7105), .Z(n5106) );
  AND U6242 ( .A(n5107), .B(n5106), .Z(n5108) );
  OR U6243 ( .A(n7110), .B(n5108), .Z(n5109) );
  NAND U6244 ( .A(n7112), .B(n5109), .Z(n5110) );
  NANDN U6245 ( .A(n7114), .B(n5110), .Z(n5111) );
  NAND U6246 ( .A(n7116), .B(n5111), .Z(n5112) );
  NANDN U6247 ( .A(n7118), .B(n5112), .Z(n5113) );
  AND U6248 ( .A(n7120), .B(n5113), .Z(n5114) );
  OR U6249 ( .A(n7122), .B(n5114), .Z(n5115) );
  NAND U6250 ( .A(n5116), .B(n5115), .Z(n5117) );
  NANDN U6251 ( .A(n5412), .B(n5117), .Z(n5120) );
  AND U6252 ( .A(n5118), .B(n5413), .Z(n5119) );
  NAND U6253 ( .A(n5120), .B(n5119), .Z(n5121) );
  NANDN U6254 ( .A(n7130), .B(n5121), .Z(n5122) );
  OR U6255 ( .A(n5123), .B(n5122), .Z(n5124) );
  AND U6256 ( .A(n5125), .B(n5124), .Z(n5126) );
  NANDN U6257 ( .A(n5127), .B(n5126), .Z(n5128) );
  AND U6258 ( .A(n5129), .B(n5128), .Z(n5131) );
  NOR U6259 ( .A(n5131), .B(n5130), .Z(n5132) );
  NANDN U6260 ( .A(n5133), .B(n5132), .Z(n5134) );
  AND U6261 ( .A(n5135), .B(n5134), .Z(n5136) );
  NANDN U6262 ( .A(n7143), .B(n5136), .Z(n5137) );
  AND U6263 ( .A(n5138), .B(n5137), .Z(n5139) );
  OR U6264 ( .A(n7148), .B(n5139), .Z(n5140) );
  NAND U6265 ( .A(n7150), .B(n5140), .Z(n5141) );
  NANDN U6266 ( .A(n7152), .B(n5141), .Z(n5142) );
  NANDN U6267 ( .A(n7153), .B(n5142), .Z(n5143) );
  AND U6268 ( .A(n7156), .B(n5143), .Z(n5144) );
  ANDN U6269 ( .B(n7159), .A(n5144), .Z(n5148) );
  NANDN U6270 ( .A(n5148), .B(n7161), .Z(n5149) );
  NAND U6271 ( .A(n7162), .B(n5149), .Z(n5150) );
  NANDN U6272 ( .A(n7165), .B(n5150), .Z(n5153) );
  AND U6273 ( .A(n5151), .B(n7169), .Z(n5152) );
  NAND U6274 ( .A(n5153), .B(n5152), .Z(n5154) );
  NANDN U6275 ( .A(n5407), .B(n5154), .Z(n5157) );
  AND U6276 ( .A(n5155), .B(n5408), .Z(n5156) );
  NAND U6277 ( .A(n5157), .B(n5156), .Z(n5158) );
  NANDN U6278 ( .A(n5159), .B(n5158), .Z(n5161) );
  IV U6279 ( .A(n5160), .Z(n7173) );
  OR U6280 ( .A(n5161), .B(n7173), .Z(n5162) );
  NAND U6281 ( .A(n5163), .B(n5162), .Z(n5164) );
  AND U6282 ( .A(n7182), .B(n5164), .Z(n5165) );
  NAND U6283 ( .A(n5166), .B(n5165), .Z(n5167) );
  NANDN U6284 ( .A(n5168), .B(n5167), .Z(n5169) );
  OR U6285 ( .A(n5169), .B(n7185), .Z(n5170) );
  NAND U6286 ( .A(n7187), .B(n5170), .Z(n5171) );
  NANDN U6287 ( .A(n7189), .B(n5171), .Z(n5172) );
  NAND U6288 ( .A(n7191), .B(n5172), .Z(n5173) );
  NANDN U6289 ( .A(n7193), .B(n5173), .Z(n5174) );
  AND U6290 ( .A(n7195), .B(n5174), .Z(n5175) );
  NANDN U6291 ( .A(n5175), .B(n7197), .Z(n5176) );
  NAND U6292 ( .A(n7199), .B(n5176), .Z(n5177) );
  NANDN U6293 ( .A(n7201), .B(n5177), .Z(n5178) );
  NAND U6294 ( .A(n5406), .B(n5178), .Z(n5179) );
  ANDN U6295 ( .B(n5179), .A(n7204), .Z(n5180) );
  NANDN U6296 ( .A(n5181), .B(n5180), .Z(n5184) );
  AND U6297 ( .A(n5182), .B(n7206), .Z(n5183) );
  NAND U6298 ( .A(n5184), .B(n5183), .Z(n5185) );
  NANDN U6299 ( .A(n5186), .B(n5185), .Z(n5187) );
  OR U6300 ( .A(n5188), .B(n5187), .Z(n5189) );
  AND U6301 ( .A(n5190), .B(n5189), .Z(n5192) );
  NAND U6302 ( .A(n5192), .B(n5191), .Z(n5194) );
  ANDN U6303 ( .B(n5194), .A(n5193), .Z(n5195) );
  NANDN U6304 ( .A(n5196), .B(n5195), .Z(n5199) );
  NANDN U6305 ( .A(y[918]), .B(x[918]), .Z(n5197) );
  AND U6306 ( .A(n5197), .B(n7213), .Z(n5198) );
  NAND U6307 ( .A(n5199), .B(n5198), .Z(n5200) );
  NANDN U6308 ( .A(n5201), .B(n5200), .Z(n5202) );
  OR U6309 ( .A(n5202), .B(n7214), .Z(n5203) );
  NAND U6310 ( .A(n7215), .B(n5203), .Z(n5204) );
  NANDN U6311 ( .A(n7216), .B(n5204), .Z(n5205) );
  NAND U6312 ( .A(n7217), .B(n5205), .Z(n5206) );
  NAND U6313 ( .A(n7218), .B(n5206), .Z(n5207) );
  NANDN U6314 ( .A(n7219), .B(n5207), .Z(n5208) );
  NAND U6315 ( .A(n7220), .B(n5208), .Z(n5209) );
  NAND U6316 ( .A(n7221), .B(n5209), .Z(n5210) );
  AND U6317 ( .A(n7222), .B(n5210), .Z(n5213) );
  NANDN U6318 ( .A(n5213), .B(n7223), .Z(n5214) );
  NAND U6319 ( .A(n7224), .B(n5214), .Z(n5215) );
  NANDN U6320 ( .A(n7225), .B(n5215), .Z(n5218) );
  NOR U6321 ( .A(n7227), .B(n5216), .Z(n5217) );
  NAND U6322 ( .A(n5218), .B(n5217), .Z(n5219) );
  AND U6323 ( .A(n5220), .B(n5219), .Z(n5221) );
  NAND U6324 ( .A(n7228), .B(n5221), .Z(n5223) );
  ANDN U6325 ( .B(n5223), .A(n5222), .Z(n5224) );
  NANDN U6326 ( .A(n5225), .B(n5224), .Z(n5226) );
  AND U6327 ( .A(n7232), .B(n5226), .Z(n5227) );
  NAND U6328 ( .A(n5228), .B(n5227), .Z(n5229) );
  NANDN U6329 ( .A(n5230), .B(n5229), .Z(n5231) );
  OR U6330 ( .A(n5231), .B(n7233), .Z(n5232) );
  NANDN U6331 ( .A(n7234), .B(n5232), .Z(n5237) );
  AND U6332 ( .A(n5237), .B(n7235), .Z(n5246) );
  NAND U6333 ( .A(n5239), .B(n5238), .Z(n5240) );
  NAND U6334 ( .A(n5241), .B(n5240), .Z(n5242) );
  AND U6335 ( .A(n5243), .B(n5242), .Z(n5245) );
  NAND U6336 ( .A(n5245), .B(n5244), .Z(n5405) );
  OR U6337 ( .A(n5246), .B(n5405), .Z(n5247) );
  AND U6338 ( .A(n7236), .B(n5247), .Z(n5251) );
  OR U6339 ( .A(n5251), .B(n5404), .Z(n5252) );
  NAND U6340 ( .A(n7237), .B(n5252), .Z(n5253) );
  NANDN U6341 ( .A(n7239), .B(n5253), .Z(n5254) );
  AND U6342 ( .A(n5255), .B(n5254), .Z(n5258) );
  NANDN U6343 ( .A(y[946]), .B(x[946]), .Z(n5257) );
  NAND U6344 ( .A(n5257), .B(n5256), .Z(n5402) );
  OR U6345 ( .A(n5258), .B(n5402), .Z(n5259) );
  AND U6346 ( .A(n5260), .B(n5259), .Z(n5261) );
  NAND U6347 ( .A(n5261), .B(n5403), .Z(n5263) );
  ANDN U6348 ( .B(n5263), .A(n5262), .Z(n5264) );
  NANDN U6349 ( .A(n7247), .B(n5264), .Z(n5268) );
  AND U6350 ( .A(n5266), .B(n5265), .Z(n5267) );
  NAND U6351 ( .A(n5268), .B(n5267), .Z(n5269) );
  NANDN U6352 ( .A(n5270), .B(n5269), .Z(n5271) );
  OR U6353 ( .A(n7256), .B(n5271), .Z(n5272) );
  AND U6354 ( .A(n5273), .B(n5272), .Z(n5274) );
  NANDN U6355 ( .A(n5400), .B(n5274), .Z(n5275) );
  AND U6356 ( .A(n5276), .B(n5275), .Z(n5279) );
  NANDN U6357 ( .A(n5279), .B(n7267), .Z(n5280) );
  NAND U6358 ( .A(n7269), .B(n5280), .Z(n5281) );
  NAND U6359 ( .A(n7272), .B(n5281), .Z(n5282) );
  NAND U6360 ( .A(n7273), .B(n5282), .Z(n5283) );
  NAND U6361 ( .A(n7274), .B(n5283), .Z(n5284) );
  NAND U6362 ( .A(n7275), .B(n5284), .Z(n5285) );
  NAND U6363 ( .A(n7276), .B(n5285), .Z(n5287) );
  ANDN U6364 ( .B(n5287), .A(n5286), .Z(n5288) );
  NANDN U6365 ( .A(n5397), .B(n5288), .Z(n5292) );
  AND U6366 ( .A(n5290), .B(n5289), .Z(n5291) );
  NAND U6367 ( .A(n5292), .B(n5291), .Z(n5293) );
  NANDN U6368 ( .A(n5294), .B(n5293), .Z(n5295) );
  OR U6369 ( .A(n7279), .B(n5295), .Z(n5296) );
  AND U6370 ( .A(n5297), .B(n5296), .Z(n5298) );
  NANDN U6371 ( .A(n7280), .B(n5298), .Z(n5299) );
  AND U6372 ( .A(n5300), .B(n5299), .Z(n5303) );
  NAND U6373 ( .A(n5302), .B(n5301), .Z(n5395) );
  OR U6374 ( .A(n5303), .B(n5395), .Z(n5304) );
  NAND U6375 ( .A(n7286), .B(n5304), .Z(n5305) );
  NANDN U6376 ( .A(n7288), .B(n5305), .Z(n5314) );
  XNOR U6377 ( .A(x[977]), .B(y[977]), .Z(n5307) );
  NAND U6378 ( .A(n5307), .B(n5306), .Z(n5308) );
  NAND U6379 ( .A(n5309), .B(n5308), .Z(n5393) );
  AND U6380 ( .A(n5393), .B(n7290), .Z(n5313) );
  NAND U6381 ( .A(n5314), .B(n5313), .Z(n5315) );
  NANDN U6382 ( .A(n5316), .B(n5315), .Z(n5319) );
  NANDN U6383 ( .A(y[978]), .B(x[978]), .Z(n5394) );
  AND U6384 ( .A(n5317), .B(n5394), .Z(n5318) );
  NAND U6385 ( .A(n5319), .B(n5318), .Z(n5320) );
  NANDN U6386 ( .A(n5321), .B(n5320), .Z(n5323) );
  OR U6387 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U6388 ( .A(n5325), .B(n5324), .Z(n5329) );
  AND U6389 ( .A(n5327), .B(n5326), .Z(n5328) );
  NAND U6390 ( .A(n5329), .B(n5328), .Z(n5330) );
  NANDN U6391 ( .A(n7306), .B(n5330), .Z(n5331) );
  OR U6392 ( .A(n5332), .B(n5331), .Z(n5333) );
  AND U6393 ( .A(n5334), .B(n5333), .Z(n5335) );
  NANDN U6394 ( .A(n7309), .B(n5335), .Z(n5336) );
  AND U6395 ( .A(n7311), .B(n5336), .Z(n5339) );
  NAND U6396 ( .A(n5337), .B(n7315), .Z(n5338) );
  OR U6397 ( .A(n5339), .B(n5338), .Z(n5340) );
  AND U6398 ( .A(n7317), .B(n5340), .Z(n5343) );
  NAND U6399 ( .A(n5342), .B(n5341), .Z(n5392) );
  OR U6400 ( .A(n5343), .B(n5392), .Z(n5344) );
  NAND U6401 ( .A(n7321), .B(n5344), .Z(n5345) );
  NANDN U6402 ( .A(n7322), .B(n5345), .Z(n5346) );
  NAND U6403 ( .A(n5391), .B(n5346), .Z(n5347) );
  NAND U6404 ( .A(n7323), .B(n5347), .Z(n5357) );
  IV U6405 ( .A(n5348), .Z(n5350) );
  NAND U6406 ( .A(n5350), .B(n5349), .Z(n5351) );
  NAND U6407 ( .A(n5352), .B(n5351), .Z(n5353) );
  AND U6408 ( .A(n5354), .B(n5353), .Z(n5356) );
  NANDN U6409 ( .A(y[997]), .B(x[997]), .Z(n5355) );
  AND U6410 ( .A(n5356), .B(n5355), .Z(n7324) );
  AND U6411 ( .A(n5357), .B(n7324), .Z(n5364) );
  ANDN U6412 ( .B(n5359), .A(n5358), .Z(n5361) );
  ANDN U6413 ( .B(n5361), .A(n5360), .Z(n5362) );
  NANDN U6414 ( .A(n5363), .B(n5362), .Z(n7325) );
  OR U6415 ( .A(n5364), .B(n7325), .Z(n5365) );
  NAND U6416 ( .A(n7326), .B(n5365), .Z(n5366) );
  NANDN U6417 ( .A(n7327), .B(n5366), .Z(n5373) );
  IV U6418 ( .A(n5367), .Z(n5368) );
  AND U6419 ( .A(n5369), .B(n5368), .Z(n7328) );
  AND U6420 ( .A(n7328), .B(n5390), .Z(n5372) );
  NAND U6421 ( .A(n5373), .B(n5372), .Z(n5374) );
  NANDN U6422 ( .A(n5375), .B(n5374), .Z(n5376) );
  NAND U6423 ( .A(n5377), .B(n5376), .Z(n7341) );
  NANDN U6424 ( .A(n7341), .B(e), .Z(n5) );
  NANDN U6425 ( .A(n5386), .B(n5385), .Z(n5387) );
  IV U6426 ( .A(n5389), .Z(n7335) );
  IV U6427 ( .A(n5392), .Z(n7319) );
  AND U6428 ( .A(n5394), .B(n5393), .Z(n7294) );
  IV U6429 ( .A(n5398), .Z(n7266) );
  IV U6430 ( .A(n5399), .Z(n7264) );
  IV U6431 ( .A(n5400), .Z(n7258) );
  IV U6432 ( .A(n5401), .Z(n7250) );
  NAND U6433 ( .A(n5403), .B(n5402), .Z(n7246) );
  IV U6434 ( .A(n5406), .Z(n7203) );
  NAND U6435 ( .A(n5408), .B(n5407), .Z(n7172) );
  IV U6436 ( .A(n5409), .Z(n7139) );
  IV U6437 ( .A(n5410), .Z(n7137) );
  IV U6438 ( .A(n5411), .Z(n7133) );
  NAND U6439 ( .A(n5413), .B(n5412), .Z(n7129) );
  IV U6440 ( .A(n5414), .Z(n7099) );
  NAND U6441 ( .A(n5416), .B(n5415), .Z(n7095) );
  IV U6442 ( .A(n5417), .Z(n5418) );
  AND U6443 ( .A(n5419), .B(n5418), .Z(n7093) );
  IV U6444 ( .A(n5420), .Z(n7078) );
  NANDN U6445 ( .A(n5427), .B(n5426), .Z(n5428) );
  NANDN U6446 ( .A(n5429), .B(n5428), .Z(n5430) );
  AND U6447 ( .A(n5431), .B(n5430), .Z(n5432) );
  OR U6448 ( .A(n5433), .B(n5432), .Z(n5434) );
  NAND U6449 ( .A(n5435), .B(n5434), .Z(n5436) );
  NANDN U6450 ( .A(n5437), .B(n5436), .Z(n5438) );
  NAND U6451 ( .A(n5439), .B(n5438), .Z(n5440) );
  NANDN U6452 ( .A(n5441), .B(n5440), .Z(n5442) );
  AND U6453 ( .A(n5443), .B(n5442), .Z(n5444) );
  OR U6454 ( .A(n5445), .B(n5444), .Z(n5446) );
  NAND U6455 ( .A(n5447), .B(n5446), .Z(n5448) );
  NANDN U6456 ( .A(n5449), .B(n5448), .Z(n5450) );
  NAND U6457 ( .A(n5451), .B(n5450), .Z(n5452) );
  NANDN U6458 ( .A(n5453), .B(n5452), .Z(n5454) );
  AND U6459 ( .A(n5455), .B(n5454), .Z(n5456) );
  OR U6460 ( .A(n5457), .B(n5456), .Z(n5458) );
  NAND U6461 ( .A(n5459), .B(n5458), .Z(n5460) );
  NANDN U6462 ( .A(n5461), .B(n5460), .Z(n5462) );
  NAND U6463 ( .A(n5463), .B(n5462), .Z(n5464) );
  NANDN U6464 ( .A(n5465), .B(n5464), .Z(n5466) );
  AND U6465 ( .A(n5467), .B(n5466), .Z(n5468) );
  OR U6466 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U6467 ( .A(n5471), .B(n5470), .Z(n5472) );
  NANDN U6468 ( .A(n5473), .B(n5472), .Z(n5474) );
  NAND U6469 ( .A(n5475), .B(n5474), .Z(n5476) );
  NANDN U6470 ( .A(n5477), .B(n5476), .Z(n5478) );
  AND U6471 ( .A(n5479), .B(n5478), .Z(n5480) );
  OR U6472 ( .A(n5481), .B(n5480), .Z(n5482) );
  NAND U6473 ( .A(n5483), .B(n5482), .Z(n5484) );
  NANDN U6474 ( .A(n5485), .B(n5484), .Z(n5486) );
  NAND U6475 ( .A(n5487), .B(n5486), .Z(n5488) );
  NANDN U6476 ( .A(n5489), .B(n5488), .Z(n5490) );
  AND U6477 ( .A(n5491), .B(n5490), .Z(n5492) );
  OR U6478 ( .A(n5493), .B(n5492), .Z(n5494) );
  NAND U6479 ( .A(n5495), .B(n5494), .Z(n5496) );
  NANDN U6480 ( .A(n5497), .B(n5496), .Z(n5498) );
  NAND U6481 ( .A(n5499), .B(n5498), .Z(n5500) );
  NANDN U6482 ( .A(n5501), .B(n5500), .Z(n5502) );
  AND U6483 ( .A(n5503), .B(n5502), .Z(n5504) );
  OR U6484 ( .A(n5505), .B(n5504), .Z(n5506) );
  NAND U6485 ( .A(n5507), .B(n5506), .Z(n5508) );
  NANDN U6486 ( .A(n5509), .B(n5508), .Z(n5510) );
  NAND U6487 ( .A(n5511), .B(n5510), .Z(n5512) );
  NANDN U6488 ( .A(n5513), .B(n5512), .Z(n5514) );
  AND U6489 ( .A(n5515), .B(n5514), .Z(n5516) );
  OR U6490 ( .A(n5517), .B(n5516), .Z(n5518) );
  NAND U6491 ( .A(n5519), .B(n5518), .Z(n5520) );
  NANDN U6492 ( .A(n5521), .B(n5520), .Z(n5522) );
  NAND U6493 ( .A(n5523), .B(n5522), .Z(n5524) );
  NANDN U6494 ( .A(n5525), .B(n5524), .Z(n5526) );
  AND U6495 ( .A(n5527), .B(n5526), .Z(n5528) );
  OR U6496 ( .A(n5529), .B(n5528), .Z(n5530) );
  NAND U6497 ( .A(n5531), .B(n5530), .Z(n5532) );
  NANDN U6498 ( .A(n5533), .B(n5532), .Z(n5534) );
  NAND U6499 ( .A(n5535), .B(n5534), .Z(n5536) );
  NANDN U6500 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U6501 ( .A(n5539), .B(n5538), .Z(n5540) );
  OR U6502 ( .A(n5541), .B(n5540), .Z(n5542) );
  NAND U6503 ( .A(n5543), .B(n5542), .Z(n5544) );
  NANDN U6504 ( .A(n5545), .B(n5544), .Z(n5546) );
  NAND U6505 ( .A(n5547), .B(n5546), .Z(n5548) );
  NANDN U6506 ( .A(n5549), .B(n5548), .Z(n5550) );
  AND U6507 ( .A(n5551), .B(n5550), .Z(n5552) );
  OR U6508 ( .A(n5553), .B(n5552), .Z(n5554) );
  NAND U6509 ( .A(n5555), .B(n5554), .Z(n5556) );
  NANDN U6510 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U6511 ( .A(n5559), .B(n5558), .Z(n5560) );
  NANDN U6512 ( .A(n5561), .B(n5560), .Z(n5562) );
  AND U6513 ( .A(n5563), .B(n5562), .Z(n5564) );
  OR U6514 ( .A(n5565), .B(n5564), .Z(n5566) );
  NAND U6515 ( .A(n5567), .B(n5566), .Z(n5568) );
  NANDN U6516 ( .A(n5569), .B(n5568), .Z(n5570) );
  NAND U6517 ( .A(n5571), .B(n5570), .Z(n5572) );
  NANDN U6518 ( .A(n5573), .B(n5572), .Z(n5574) );
  AND U6519 ( .A(n5575), .B(n5574), .Z(n5576) );
  OR U6520 ( .A(n5577), .B(n5576), .Z(n5578) );
  NAND U6521 ( .A(n5579), .B(n5578), .Z(n5580) );
  NANDN U6522 ( .A(n5581), .B(n5580), .Z(n5582) );
  NAND U6523 ( .A(n5583), .B(n5582), .Z(n5584) );
  NANDN U6524 ( .A(n5585), .B(n5584), .Z(n5586) );
  AND U6525 ( .A(n5587), .B(n5586), .Z(n5588) );
  OR U6526 ( .A(n5589), .B(n5588), .Z(n5590) );
  NAND U6527 ( .A(n5591), .B(n5590), .Z(n5592) );
  NANDN U6528 ( .A(n5593), .B(n5592), .Z(n5594) );
  NAND U6529 ( .A(n5595), .B(n5594), .Z(n5596) );
  NANDN U6530 ( .A(n5597), .B(n5596), .Z(n5598) );
  AND U6531 ( .A(n5599), .B(n5598), .Z(n5600) );
  OR U6532 ( .A(n5601), .B(n5600), .Z(n5602) );
  NAND U6533 ( .A(n5603), .B(n5602), .Z(n5604) );
  NANDN U6534 ( .A(n5605), .B(n5604), .Z(n5606) );
  NAND U6535 ( .A(n5607), .B(n5606), .Z(n5608) );
  NANDN U6536 ( .A(n5609), .B(n5608), .Z(n5610) );
  AND U6537 ( .A(n5611), .B(n5610), .Z(n5612) );
  OR U6538 ( .A(n5613), .B(n5612), .Z(n5614) );
  NAND U6539 ( .A(n5615), .B(n5614), .Z(n5616) );
  NANDN U6540 ( .A(n5617), .B(n5616), .Z(n5618) );
  NAND U6541 ( .A(n5619), .B(n5618), .Z(n5620) );
  NANDN U6542 ( .A(n5621), .B(n5620), .Z(n5622) );
  AND U6543 ( .A(n5623), .B(n5622), .Z(n5624) );
  OR U6544 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U6545 ( .A(n5627), .B(n5626), .Z(n5628) );
  NANDN U6546 ( .A(n5629), .B(n5628), .Z(n5630) );
  NAND U6547 ( .A(n5631), .B(n5630), .Z(n5632) );
  NANDN U6548 ( .A(n5633), .B(n5632), .Z(n5634) );
  AND U6549 ( .A(n5635), .B(n5634), .Z(n5636) );
  OR U6550 ( .A(n5637), .B(n5636), .Z(n5638) );
  NAND U6551 ( .A(n5639), .B(n5638), .Z(n5640) );
  NANDN U6552 ( .A(n5641), .B(n5640), .Z(n5642) );
  NAND U6553 ( .A(n5643), .B(n5642), .Z(n5644) );
  NANDN U6554 ( .A(n5645), .B(n5644), .Z(n5646) );
  AND U6555 ( .A(n5647), .B(n5646), .Z(n5648) );
  OR U6556 ( .A(n5649), .B(n5648), .Z(n5650) );
  NAND U6557 ( .A(n5651), .B(n5650), .Z(n5652) );
  NANDN U6558 ( .A(n5653), .B(n5652), .Z(n5654) );
  NAND U6559 ( .A(n5655), .B(n5654), .Z(n5656) );
  NANDN U6560 ( .A(n5657), .B(n5656), .Z(n5658) );
  AND U6561 ( .A(n5659), .B(n5658), .Z(n5660) );
  OR U6562 ( .A(n5661), .B(n5660), .Z(n5662) );
  NAND U6563 ( .A(n5663), .B(n5662), .Z(n5664) );
  NANDN U6564 ( .A(n5665), .B(n5664), .Z(n5666) );
  NAND U6565 ( .A(n5667), .B(n5666), .Z(n5668) );
  NANDN U6566 ( .A(n5669), .B(n5668), .Z(n5670) );
  AND U6567 ( .A(n5671), .B(n5670), .Z(n5672) );
  OR U6568 ( .A(n5673), .B(n5672), .Z(n5674) );
  NAND U6569 ( .A(n5675), .B(n5674), .Z(n5676) );
  NANDN U6570 ( .A(n5677), .B(n5676), .Z(n5678) );
  NAND U6571 ( .A(n5679), .B(n5678), .Z(n5680) );
  NANDN U6572 ( .A(n5681), .B(n5680), .Z(n5682) );
  AND U6573 ( .A(n5683), .B(n5682), .Z(n5684) );
  OR U6574 ( .A(n5685), .B(n5684), .Z(n5686) );
  NAND U6575 ( .A(n5687), .B(n5686), .Z(n5688) );
  NANDN U6576 ( .A(n5689), .B(n5688), .Z(n5690) );
  NAND U6577 ( .A(n5691), .B(n5690), .Z(n5692) );
  NANDN U6578 ( .A(n5693), .B(n5692), .Z(n5694) );
  AND U6579 ( .A(n5695), .B(n5694), .Z(n5696) );
  OR U6580 ( .A(n5697), .B(n5696), .Z(n5698) );
  NAND U6581 ( .A(n5699), .B(n5698), .Z(n5700) );
  NANDN U6582 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U6583 ( .A(n5703), .B(n5702), .Z(n5704) );
  NANDN U6584 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U6585 ( .A(n5707), .B(n5706), .Z(n5708) );
  OR U6586 ( .A(n5709), .B(n5708), .Z(n5710) );
  NAND U6587 ( .A(n5711), .B(n5710), .Z(n5712) );
  NANDN U6588 ( .A(n5713), .B(n5712), .Z(n5714) );
  NAND U6589 ( .A(n5715), .B(n5714), .Z(n5716) );
  NANDN U6590 ( .A(n5717), .B(n5716), .Z(n5718) );
  AND U6591 ( .A(n5719), .B(n5718), .Z(n5720) );
  OR U6592 ( .A(n5721), .B(n5720), .Z(n5722) );
  NAND U6593 ( .A(n5723), .B(n5722), .Z(n5724) );
  NANDN U6594 ( .A(n5725), .B(n5724), .Z(n5726) );
  NAND U6595 ( .A(n5727), .B(n5726), .Z(n5728) );
  NANDN U6596 ( .A(n5729), .B(n5728), .Z(n5730) );
  AND U6597 ( .A(n5731), .B(n5730), .Z(n5732) );
  OR U6598 ( .A(n5733), .B(n5732), .Z(n5734) );
  NAND U6599 ( .A(n5735), .B(n5734), .Z(n5736) );
  NANDN U6600 ( .A(n5737), .B(n5736), .Z(n5738) );
  NAND U6601 ( .A(n5739), .B(n5738), .Z(n5740) );
  NANDN U6602 ( .A(n5741), .B(n5740), .Z(n5742) );
  AND U6603 ( .A(n5743), .B(n5742), .Z(n5744) );
  OR U6604 ( .A(n5745), .B(n5744), .Z(n5746) );
  NAND U6605 ( .A(n5747), .B(n5746), .Z(n5748) );
  NANDN U6606 ( .A(n5749), .B(n5748), .Z(n5750) );
  NAND U6607 ( .A(n5751), .B(n5750), .Z(n5752) );
  NANDN U6608 ( .A(n5753), .B(n5752), .Z(n5754) );
  AND U6609 ( .A(n5755), .B(n5754), .Z(n5756) );
  OR U6610 ( .A(n5757), .B(n5756), .Z(n5758) );
  NAND U6611 ( .A(n5759), .B(n5758), .Z(n5760) );
  NANDN U6612 ( .A(n5761), .B(n5760), .Z(n5762) );
  NAND U6613 ( .A(n5763), .B(n5762), .Z(n5764) );
  NANDN U6614 ( .A(n5765), .B(n5764), .Z(n5766) );
  AND U6615 ( .A(n5767), .B(n5766), .Z(n5768) );
  OR U6616 ( .A(n5769), .B(n5768), .Z(n5770) );
  NAND U6617 ( .A(n5771), .B(n5770), .Z(n5772) );
  NANDN U6618 ( .A(n5773), .B(n5772), .Z(n5774) );
  NAND U6619 ( .A(n5775), .B(n5774), .Z(n5776) );
  NANDN U6620 ( .A(n5777), .B(n5776), .Z(n5778) );
  AND U6621 ( .A(n5779), .B(n5778), .Z(n5780) );
  OR U6622 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U6623 ( .A(n5783), .B(n5782), .Z(n5784) );
  NANDN U6624 ( .A(n5785), .B(n5784), .Z(n5786) );
  NAND U6625 ( .A(n5787), .B(n5786), .Z(n5788) );
  NANDN U6626 ( .A(n5789), .B(n5788), .Z(n5790) );
  AND U6627 ( .A(n5791), .B(n5790), .Z(n5792) );
  OR U6628 ( .A(n5793), .B(n5792), .Z(n5794) );
  NAND U6629 ( .A(n5795), .B(n5794), .Z(n5796) );
  NANDN U6630 ( .A(n5797), .B(n5796), .Z(n5798) );
  NAND U6631 ( .A(n5799), .B(n5798), .Z(n5800) );
  NANDN U6632 ( .A(n5801), .B(n5800), .Z(n5802) );
  AND U6633 ( .A(n5803), .B(n5802), .Z(n5804) );
  OR U6634 ( .A(n5805), .B(n5804), .Z(n5806) );
  NAND U6635 ( .A(n5807), .B(n5806), .Z(n5808) );
  NANDN U6636 ( .A(n5809), .B(n5808), .Z(n5810) );
  NAND U6637 ( .A(n5811), .B(n5810), .Z(n5812) );
  NANDN U6638 ( .A(n5813), .B(n5812), .Z(n5814) );
  AND U6639 ( .A(n5815), .B(n5814), .Z(n5816) );
  OR U6640 ( .A(n5817), .B(n5816), .Z(n5818) );
  NAND U6641 ( .A(n5819), .B(n5818), .Z(n5820) );
  NANDN U6642 ( .A(n5821), .B(n5820), .Z(n5822) );
  NAND U6643 ( .A(n5823), .B(n5822), .Z(n5824) );
  NANDN U6644 ( .A(n5825), .B(n5824), .Z(n5826) );
  AND U6645 ( .A(n5827), .B(n5826), .Z(n5828) );
  OR U6646 ( .A(n5829), .B(n5828), .Z(n5830) );
  NAND U6647 ( .A(n5831), .B(n5830), .Z(n5832) );
  NANDN U6648 ( .A(n5833), .B(n5832), .Z(n5834) );
  NAND U6649 ( .A(n5835), .B(n5834), .Z(n5836) );
  NANDN U6650 ( .A(n5837), .B(n5836), .Z(n5838) );
  AND U6651 ( .A(n5839), .B(n5838), .Z(n5840) );
  OR U6652 ( .A(n5841), .B(n5840), .Z(n5842) );
  NAND U6653 ( .A(n5843), .B(n5842), .Z(n5844) );
  NANDN U6654 ( .A(n5845), .B(n5844), .Z(n5846) );
  NAND U6655 ( .A(n5847), .B(n5846), .Z(n5848) );
  NANDN U6656 ( .A(n5849), .B(n5848), .Z(n5850) );
  AND U6657 ( .A(n5851), .B(n5850), .Z(n5852) );
  OR U6658 ( .A(n5853), .B(n5852), .Z(n5854) );
  NAND U6659 ( .A(n5855), .B(n5854), .Z(n5856) );
  NANDN U6660 ( .A(n5857), .B(n5856), .Z(n5858) );
  NAND U6661 ( .A(n5859), .B(n5858), .Z(n5860) );
  NANDN U6662 ( .A(n5861), .B(n5860), .Z(n5862) );
  AND U6663 ( .A(n5863), .B(n5862), .Z(n5864) );
  OR U6664 ( .A(n5865), .B(n5864), .Z(n5866) );
  NAND U6665 ( .A(n5867), .B(n5866), .Z(n5868) );
  NANDN U6666 ( .A(n5869), .B(n5868), .Z(n5870) );
  NAND U6667 ( .A(n5871), .B(n5870), .Z(n5872) );
  NANDN U6668 ( .A(n5873), .B(n5872), .Z(n5874) );
  AND U6669 ( .A(n5875), .B(n5874), .Z(n5876) );
  OR U6670 ( .A(n5877), .B(n5876), .Z(n5878) );
  NAND U6671 ( .A(n5879), .B(n5878), .Z(n5880) );
  NANDN U6672 ( .A(n5881), .B(n5880), .Z(n5882) );
  NAND U6673 ( .A(n5883), .B(n5882), .Z(n5884) );
  NANDN U6674 ( .A(n5885), .B(n5884), .Z(n5886) );
  AND U6675 ( .A(n5887), .B(n5886), .Z(n5888) );
  OR U6676 ( .A(n5889), .B(n5888), .Z(n5890) );
  NAND U6677 ( .A(n5891), .B(n5890), .Z(n5892) );
  NANDN U6678 ( .A(n5893), .B(n5892), .Z(n5894) );
  NAND U6679 ( .A(n5895), .B(n5894), .Z(n5896) );
  NANDN U6680 ( .A(n5897), .B(n5896), .Z(n5898) );
  AND U6681 ( .A(n5899), .B(n5898), .Z(n5900) );
  OR U6682 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U6683 ( .A(n5903), .B(n5902), .Z(n5904) );
  NANDN U6684 ( .A(n5905), .B(n5904), .Z(n5906) );
  NAND U6685 ( .A(n5907), .B(n5906), .Z(n5908) );
  NANDN U6686 ( .A(n5909), .B(n5908), .Z(n5910) );
  AND U6687 ( .A(n5911), .B(n5910), .Z(n5912) );
  OR U6688 ( .A(n5913), .B(n5912), .Z(n5914) );
  NAND U6689 ( .A(n5915), .B(n5914), .Z(n5916) );
  NANDN U6690 ( .A(n5917), .B(n5916), .Z(n5918) );
  NAND U6691 ( .A(n5919), .B(n5918), .Z(n5920) );
  NANDN U6692 ( .A(n5921), .B(n5920), .Z(n5922) );
  AND U6693 ( .A(n5923), .B(n5922), .Z(n5924) );
  OR U6694 ( .A(n5925), .B(n5924), .Z(n5926) );
  NAND U6695 ( .A(n5927), .B(n5926), .Z(n5928) );
  NANDN U6696 ( .A(n5929), .B(n5928), .Z(n5930) );
  NAND U6697 ( .A(n5931), .B(n5930), .Z(n5932) );
  NANDN U6698 ( .A(n5933), .B(n5932), .Z(n5934) );
  AND U6699 ( .A(n5935), .B(n5934), .Z(n5936) );
  OR U6700 ( .A(n5937), .B(n5936), .Z(n5938) );
  NAND U6701 ( .A(n5939), .B(n5938), .Z(n5940) );
  NANDN U6702 ( .A(n5941), .B(n5940), .Z(n5942) );
  NAND U6703 ( .A(n5943), .B(n5942), .Z(n5944) );
  NANDN U6704 ( .A(n5945), .B(n5944), .Z(n5946) );
  AND U6705 ( .A(n5947), .B(n5946), .Z(n5948) );
  OR U6706 ( .A(n5949), .B(n5948), .Z(n5950) );
  NAND U6707 ( .A(n5951), .B(n5950), .Z(n5952) );
  NANDN U6708 ( .A(n5953), .B(n5952), .Z(n5954) );
  NAND U6709 ( .A(n5955), .B(n5954), .Z(n5956) );
  NANDN U6710 ( .A(n5957), .B(n5956), .Z(n5958) );
  AND U6711 ( .A(n5959), .B(n5958), .Z(n5960) );
  OR U6712 ( .A(n5961), .B(n5960), .Z(n5962) );
  NAND U6713 ( .A(n5963), .B(n5962), .Z(n5964) );
  NANDN U6714 ( .A(n5965), .B(n5964), .Z(n5966) );
  NAND U6715 ( .A(n5967), .B(n5966), .Z(n5968) );
  NANDN U6716 ( .A(n5969), .B(n5968), .Z(n5970) );
  AND U6717 ( .A(n5971), .B(n5970), .Z(n5972) );
  OR U6718 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U6719 ( .A(n5975), .B(n5974), .Z(n5976) );
  NANDN U6720 ( .A(n5977), .B(n5976), .Z(n5978) );
  NAND U6721 ( .A(n5979), .B(n5978), .Z(n5980) );
  NANDN U6722 ( .A(n5981), .B(n5980), .Z(n5982) );
  AND U6723 ( .A(n5983), .B(n5982), .Z(n5984) );
  OR U6724 ( .A(n5985), .B(n5984), .Z(n5986) );
  NAND U6725 ( .A(n5987), .B(n5986), .Z(n5988) );
  NANDN U6726 ( .A(n5989), .B(n5988), .Z(n5990) );
  NAND U6727 ( .A(n5991), .B(n5990), .Z(n5992) );
  NANDN U6728 ( .A(n5993), .B(n5992), .Z(n5994) );
  AND U6729 ( .A(n5995), .B(n5994), .Z(n5996) );
  OR U6730 ( .A(n5997), .B(n5996), .Z(n5998) );
  NAND U6731 ( .A(n5999), .B(n5998), .Z(n6000) );
  NANDN U6732 ( .A(n6001), .B(n6000), .Z(n6002) );
  NAND U6733 ( .A(n6003), .B(n6002), .Z(n6004) );
  NAND U6734 ( .A(n6005), .B(n6004), .Z(n6006) );
  AND U6735 ( .A(n6007), .B(n6006), .Z(n6008) );
  OR U6736 ( .A(n6009), .B(n6008), .Z(n6010) );
  NAND U6737 ( .A(n6011), .B(n6010), .Z(n6012) );
  NANDN U6738 ( .A(n6013), .B(n6012), .Z(n6014) );
  NAND U6739 ( .A(n6015), .B(n6014), .Z(n6016) );
  NANDN U6740 ( .A(n6017), .B(n6016), .Z(n6018) );
  AND U6741 ( .A(n6019), .B(n6018), .Z(n6020) );
  OR U6742 ( .A(n6021), .B(n6020), .Z(n6022) );
  NAND U6743 ( .A(n6023), .B(n6022), .Z(n6024) );
  NANDN U6744 ( .A(n6025), .B(n6024), .Z(n6026) );
  NAND U6745 ( .A(n6027), .B(n6026), .Z(n6028) );
  NANDN U6746 ( .A(n6029), .B(n6028), .Z(n6030) );
  AND U6747 ( .A(n6031), .B(n6030), .Z(n6032) );
  OR U6748 ( .A(n6033), .B(n6032), .Z(n6034) );
  NAND U6749 ( .A(n6035), .B(n6034), .Z(n6036) );
  NANDN U6750 ( .A(n6037), .B(n6036), .Z(n6038) );
  NAND U6751 ( .A(n6039), .B(n6038), .Z(n6040) );
  NANDN U6752 ( .A(n6041), .B(n6040), .Z(n6042) );
  AND U6753 ( .A(n6043), .B(n6042), .Z(n6044) );
  OR U6754 ( .A(n6045), .B(n6044), .Z(n6046) );
  NAND U6755 ( .A(n6047), .B(n6046), .Z(n6048) );
  NANDN U6756 ( .A(n6049), .B(n6048), .Z(n6050) );
  NAND U6757 ( .A(n6051), .B(n6050), .Z(n6052) );
  NANDN U6758 ( .A(n6053), .B(n6052), .Z(n6054) );
  AND U6759 ( .A(n6055), .B(n6054), .Z(n6056) );
  OR U6760 ( .A(n6057), .B(n6056), .Z(n6058) );
  NAND U6761 ( .A(n6059), .B(n6058), .Z(n6060) );
  NANDN U6762 ( .A(n6061), .B(n6060), .Z(n6062) );
  NAND U6763 ( .A(n6063), .B(n6062), .Z(n6064) );
  NANDN U6764 ( .A(n6065), .B(n6064), .Z(n6066) );
  AND U6765 ( .A(n6067), .B(n6066), .Z(n6068) );
  OR U6766 ( .A(n6069), .B(n6068), .Z(n6070) );
  NAND U6767 ( .A(n6071), .B(n6070), .Z(n6072) );
  NANDN U6768 ( .A(n6073), .B(n6072), .Z(n6074) );
  NAND U6769 ( .A(n6075), .B(n6074), .Z(n6076) );
  NANDN U6770 ( .A(n6077), .B(n6076), .Z(n6078) );
  AND U6771 ( .A(n6079), .B(n6078), .Z(n6080) );
  OR U6772 ( .A(n6081), .B(n6080), .Z(n6082) );
  NAND U6773 ( .A(n6083), .B(n6082), .Z(n6084) );
  NANDN U6774 ( .A(n6085), .B(n6084), .Z(n6086) );
  NAND U6775 ( .A(n6087), .B(n6086), .Z(n6088) );
  NANDN U6776 ( .A(n6089), .B(n6088), .Z(n6090) );
  AND U6777 ( .A(n6091), .B(n6090), .Z(n6092) );
  OR U6778 ( .A(n6093), .B(n6092), .Z(n6094) );
  NAND U6779 ( .A(n6095), .B(n6094), .Z(n6096) );
  NANDN U6780 ( .A(n6097), .B(n6096), .Z(n6098) );
  NAND U6781 ( .A(n6099), .B(n6098), .Z(n6100) );
  NANDN U6782 ( .A(n6101), .B(n6100), .Z(n6102) );
  AND U6783 ( .A(n6103), .B(n6102), .Z(n6104) );
  OR U6784 ( .A(n6105), .B(n6104), .Z(n6106) );
  NAND U6785 ( .A(n6107), .B(n6106), .Z(n6108) );
  NANDN U6786 ( .A(n6109), .B(n6108), .Z(n6110) );
  NAND U6787 ( .A(n6111), .B(n6110), .Z(n6112) );
  NANDN U6788 ( .A(n6113), .B(n6112), .Z(n6114) );
  AND U6789 ( .A(n6115), .B(n6114), .Z(n6116) );
  OR U6790 ( .A(n6117), .B(n6116), .Z(n6118) );
  NAND U6791 ( .A(n6119), .B(n6118), .Z(n6120) );
  NANDN U6792 ( .A(n6121), .B(n6120), .Z(n6122) );
  NAND U6793 ( .A(n6123), .B(n6122), .Z(n6124) );
  NANDN U6794 ( .A(n6125), .B(n6124), .Z(n6126) );
  AND U6795 ( .A(n6127), .B(n6126), .Z(n6128) );
  OR U6796 ( .A(n6129), .B(n6128), .Z(n6130) );
  NAND U6797 ( .A(n6131), .B(n6130), .Z(n6132) );
  NANDN U6798 ( .A(n6133), .B(n6132), .Z(n6134) );
  NAND U6799 ( .A(n6135), .B(n6134), .Z(n6136) );
  NANDN U6800 ( .A(n6137), .B(n6136), .Z(n6138) );
  AND U6801 ( .A(n6139), .B(n6138), .Z(n6140) );
  OR U6802 ( .A(n6141), .B(n6140), .Z(n6142) );
  NAND U6803 ( .A(n6143), .B(n6142), .Z(n6144) );
  NANDN U6804 ( .A(n6145), .B(n6144), .Z(n6146) );
  NAND U6805 ( .A(n6147), .B(n6146), .Z(n6148) );
  NANDN U6806 ( .A(n6149), .B(n6148), .Z(n6150) );
  AND U6807 ( .A(n6151), .B(n6150), .Z(n6152) );
  OR U6808 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U6809 ( .A(n6155), .B(n6154), .Z(n6156) );
  NANDN U6810 ( .A(n6157), .B(n6156), .Z(n6158) );
  NAND U6811 ( .A(n6159), .B(n6158), .Z(n6160) );
  NANDN U6812 ( .A(n6161), .B(n6160), .Z(n6162) );
  AND U6813 ( .A(n6163), .B(n6162), .Z(n6164) );
  OR U6814 ( .A(n6165), .B(n6164), .Z(n6166) );
  NAND U6815 ( .A(n6167), .B(n6166), .Z(n6168) );
  NANDN U6816 ( .A(n6169), .B(n6168), .Z(n6170) );
  NAND U6817 ( .A(n6171), .B(n6170), .Z(n6172) );
  NANDN U6818 ( .A(n6173), .B(n6172), .Z(n6174) );
  AND U6819 ( .A(n6175), .B(n6174), .Z(n6176) );
  OR U6820 ( .A(n6177), .B(n6176), .Z(n6178) );
  NAND U6821 ( .A(n6179), .B(n6178), .Z(n6180) );
  NANDN U6822 ( .A(n6181), .B(n6180), .Z(n6182) );
  NAND U6823 ( .A(n6183), .B(n6182), .Z(n6184) );
  NANDN U6824 ( .A(n6185), .B(n6184), .Z(n6186) );
  AND U6825 ( .A(n6187), .B(n6186), .Z(n6188) );
  OR U6826 ( .A(n6189), .B(n6188), .Z(n6190) );
  NAND U6827 ( .A(n6191), .B(n6190), .Z(n6192) );
  NANDN U6828 ( .A(n6193), .B(n6192), .Z(n6194) );
  NAND U6829 ( .A(n6195), .B(n6194), .Z(n6196) );
  NANDN U6830 ( .A(n6197), .B(n6196), .Z(n6198) );
  AND U6831 ( .A(n6199), .B(n6198), .Z(n6200) );
  OR U6832 ( .A(n6201), .B(n6200), .Z(n6202) );
  NAND U6833 ( .A(n6203), .B(n6202), .Z(n6204) );
  NANDN U6834 ( .A(n6205), .B(n6204), .Z(n6206) );
  NAND U6835 ( .A(n6207), .B(n6206), .Z(n6208) );
  NANDN U6836 ( .A(n6209), .B(n6208), .Z(n6210) );
  AND U6837 ( .A(n6211), .B(n6210), .Z(n6212) );
  OR U6838 ( .A(n6213), .B(n6212), .Z(n6214) );
  NAND U6839 ( .A(n6215), .B(n6214), .Z(n6216) );
  NANDN U6840 ( .A(n6217), .B(n6216), .Z(n6218) );
  NAND U6841 ( .A(n6219), .B(n6218), .Z(n6220) );
  NANDN U6842 ( .A(n6221), .B(n6220), .Z(n6222) );
  AND U6843 ( .A(n6223), .B(n6222), .Z(n6224) );
  OR U6844 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U6845 ( .A(n6227), .B(n6226), .Z(n6228) );
  NANDN U6846 ( .A(n6229), .B(n6228), .Z(n6230) );
  NAND U6847 ( .A(n6231), .B(n6230), .Z(n6232) );
  NANDN U6848 ( .A(n6233), .B(n6232), .Z(n6234) );
  AND U6849 ( .A(n6235), .B(n6234), .Z(n6236) );
  OR U6850 ( .A(n6237), .B(n6236), .Z(n6238) );
  NAND U6851 ( .A(n6239), .B(n6238), .Z(n6240) );
  NANDN U6852 ( .A(n6241), .B(n6240), .Z(n6242) );
  NAND U6853 ( .A(n6243), .B(n6242), .Z(n6244) );
  NANDN U6854 ( .A(n6245), .B(n6244), .Z(n6246) );
  AND U6855 ( .A(n6247), .B(n6246), .Z(n6248) );
  OR U6856 ( .A(n6249), .B(n6248), .Z(n6250) );
  NAND U6857 ( .A(n6251), .B(n6250), .Z(n6252) );
  NANDN U6858 ( .A(n6253), .B(n6252), .Z(n6254) );
  NAND U6859 ( .A(n6255), .B(n6254), .Z(n6256) );
  NANDN U6860 ( .A(n6257), .B(n6256), .Z(n6258) );
  AND U6861 ( .A(n6259), .B(n6258), .Z(n6260) );
  OR U6862 ( .A(n6261), .B(n6260), .Z(n6262) );
  NAND U6863 ( .A(n6263), .B(n6262), .Z(n6264) );
  NANDN U6864 ( .A(n6265), .B(n6264), .Z(n6266) );
  NAND U6865 ( .A(n6267), .B(n6266), .Z(n6268) );
  NANDN U6866 ( .A(n6269), .B(n6268), .Z(n6270) );
  AND U6867 ( .A(n6271), .B(n6270), .Z(n6272) );
  OR U6868 ( .A(n6273), .B(n6272), .Z(n6274) );
  NAND U6869 ( .A(n6275), .B(n6274), .Z(n6276) );
  NANDN U6870 ( .A(n6277), .B(n6276), .Z(n6278) );
  NAND U6871 ( .A(n6279), .B(n6278), .Z(n6280) );
  NANDN U6872 ( .A(n6281), .B(n6280), .Z(n6282) );
  AND U6873 ( .A(n6283), .B(n6282), .Z(n6284) );
  OR U6874 ( .A(n6285), .B(n6284), .Z(n6286) );
  NAND U6875 ( .A(n6287), .B(n6286), .Z(n6288) );
  NANDN U6876 ( .A(n6289), .B(n6288), .Z(n6290) );
  NAND U6877 ( .A(n6291), .B(n6290), .Z(n6292) );
  NANDN U6878 ( .A(n6293), .B(n6292), .Z(n6294) );
  AND U6879 ( .A(n6295), .B(n6294), .Z(n6296) );
  OR U6880 ( .A(n6297), .B(n6296), .Z(n6298) );
  NAND U6881 ( .A(n6299), .B(n6298), .Z(n6300) );
  NANDN U6882 ( .A(n6301), .B(n6300), .Z(n6302) );
  NAND U6883 ( .A(n6303), .B(n6302), .Z(n6304) );
  NANDN U6884 ( .A(n6305), .B(n6304), .Z(n6306) );
  AND U6885 ( .A(n6307), .B(n6306), .Z(n6308) );
  OR U6886 ( .A(n6309), .B(n6308), .Z(n6310) );
  NAND U6887 ( .A(n6311), .B(n6310), .Z(n6312) );
  NANDN U6888 ( .A(n6313), .B(n6312), .Z(n6314) );
  NAND U6889 ( .A(n6315), .B(n6314), .Z(n6316) );
  NANDN U6890 ( .A(n6317), .B(n6316), .Z(n6318) );
  AND U6891 ( .A(n6319), .B(n6318), .Z(n6320) );
  OR U6892 ( .A(n6321), .B(n6320), .Z(n6322) );
  NAND U6893 ( .A(n6323), .B(n6322), .Z(n6324) );
  NANDN U6894 ( .A(n6325), .B(n6324), .Z(n6326) );
  NAND U6895 ( .A(n6327), .B(n6326), .Z(n6328) );
  NANDN U6896 ( .A(n6329), .B(n6328), .Z(n6330) );
  AND U6897 ( .A(n6331), .B(n6330), .Z(n6332) );
  OR U6898 ( .A(n6333), .B(n6332), .Z(n6334) );
  NAND U6899 ( .A(n6335), .B(n6334), .Z(n6336) );
  NANDN U6900 ( .A(n6337), .B(n6336), .Z(n6338) );
  NAND U6901 ( .A(n6339), .B(n6338), .Z(n6340) );
  NANDN U6902 ( .A(n6341), .B(n6340), .Z(n6342) );
  AND U6903 ( .A(n6343), .B(n6342), .Z(n6344) );
  OR U6904 ( .A(n6345), .B(n6344), .Z(n6346) );
  NAND U6905 ( .A(n6347), .B(n6346), .Z(n6348) );
  NANDN U6906 ( .A(n6349), .B(n6348), .Z(n6350) );
  NAND U6907 ( .A(n6351), .B(n6350), .Z(n6352) );
  NANDN U6908 ( .A(n6353), .B(n6352), .Z(n6354) );
  AND U6909 ( .A(n6355), .B(n6354), .Z(n6356) );
  OR U6910 ( .A(n6357), .B(n6356), .Z(n6358) );
  NAND U6911 ( .A(n6359), .B(n6358), .Z(n6360) );
  NANDN U6912 ( .A(n6361), .B(n6360), .Z(n6362) );
  NAND U6913 ( .A(n6363), .B(n6362), .Z(n6364) );
  NANDN U6914 ( .A(n6365), .B(n6364), .Z(n6366) );
  AND U6915 ( .A(n6367), .B(n6366), .Z(n6368) );
  OR U6916 ( .A(n6369), .B(n6368), .Z(n6370) );
  NAND U6917 ( .A(n6371), .B(n6370), .Z(n6372) );
  NANDN U6918 ( .A(n6373), .B(n6372), .Z(n6374) );
  NAND U6919 ( .A(n6375), .B(n6374), .Z(n6376) );
  NANDN U6920 ( .A(n6377), .B(n6376), .Z(n6378) );
  AND U6921 ( .A(n6379), .B(n6378), .Z(n6380) );
  OR U6922 ( .A(n6381), .B(n6380), .Z(n6382) );
  NAND U6923 ( .A(n6383), .B(n6382), .Z(n6384) );
  NANDN U6924 ( .A(n6385), .B(n6384), .Z(n6386) );
  NAND U6925 ( .A(n6387), .B(n6386), .Z(n6388) );
  NANDN U6926 ( .A(n6389), .B(n6388), .Z(n6390) );
  AND U6927 ( .A(n6391), .B(n6390), .Z(n6392) );
  OR U6928 ( .A(n6393), .B(n6392), .Z(n6394) );
  NAND U6929 ( .A(n6395), .B(n6394), .Z(n6396) );
  NANDN U6930 ( .A(n6397), .B(n6396), .Z(n6398) );
  NAND U6931 ( .A(n6399), .B(n6398), .Z(n6400) );
  NANDN U6932 ( .A(n6401), .B(n6400), .Z(n6402) );
  AND U6933 ( .A(n6403), .B(n6402), .Z(n6404) );
  OR U6934 ( .A(n6405), .B(n6404), .Z(n6406) );
  NAND U6935 ( .A(n6407), .B(n6406), .Z(n6408) );
  NANDN U6936 ( .A(n6409), .B(n6408), .Z(n6410) );
  NAND U6937 ( .A(n6411), .B(n6410), .Z(n6412) );
  NANDN U6938 ( .A(n6413), .B(n6412), .Z(n6414) );
  AND U6939 ( .A(n6415), .B(n6414), .Z(n6416) );
  OR U6940 ( .A(n6417), .B(n6416), .Z(n6418) );
  NAND U6941 ( .A(n6419), .B(n6418), .Z(n6420) );
  NANDN U6942 ( .A(n6421), .B(n6420), .Z(n6422) );
  NAND U6943 ( .A(n6423), .B(n6422), .Z(n6424) );
  NANDN U6944 ( .A(n6425), .B(n6424), .Z(n6426) );
  AND U6945 ( .A(n6427), .B(n6426), .Z(n6428) );
  OR U6946 ( .A(n6429), .B(n6428), .Z(n6430) );
  NAND U6947 ( .A(n6431), .B(n6430), .Z(n6432) );
  NANDN U6948 ( .A(n6433), .B(n6432), .Z(n6434) );
  NAND U6949 ( .A(n6435), .B(n6434), .Z(n6436) );
  NANDN U6950 ( .A(n6437), .B(n6436), .Z(n6438) );
  AND U6951 ( .A(n6439), .B(n6438), .Z(n6440) );
  OR U6952 ( .A(n6441), .B(n6440), .Z(n6442) );
  NAND U6953 ( .A(n6443), .B(n6442), .Z(n6444) );
  NANDN U6954 ( .A(n6445), .B(n6444), .Z(n6446) );
  NAND U6955 ( .A(n6447), .B(n6446), .Z(n6448) );
  NANDN U6956 ( .A(n6449), .B(n6448), .Z(n6450) );
  AND U6957 ( .A(n6451), .B(n6450), .Z(n6452) );
  OR U6958 ( .A(n6453), .B(n6452), .Z(n6454) );
  NAND U6959 ( .A(n6455), .B(n6454), .Z(n6456) );
  NANDN U6960 ( .A(n6457), .B(n6456), .Z(n6458) );
  NAND U6961 ( .A(n6459), .B(n6458), .Z(n6460) );
  NANDN U6962 ( .A(n6461), .B(n6460), .Z(n6462) );
  AND U6963 ( .A(n6463), .B(n6462), .Z(n6464) );
  OR U6964 ( .A(n6465), .B(n6464), .Z(n6466) );
  NAND U6965 ( .A(n6467), .B(n6466), .Z(n6468) );
  NANDN U6966 ( .A(n6469), .B(n6468), .Z(n6470) );
  NAND U6967 ( .A(n6471), .B(n6470), .Z(n6472) );
  NANDN U6968 ( .A(n6473), .B(n6472), .Z(n6474) );
  AND U6969 ( .A(n6475), .B(n6474), .Z(n6476) );
  OR U6970 ( .A(n6477), .B(n6476), .Z(n6478) );
  NAND U6971 ( .A(n6479), .B(n6478), .Z(n6480) );
  NANDN U6972 ( .A(n6481), .B(n6480), .Z(n6482) );
  NAND U6973 ( .A(n6483), .B(n6482), .Z(n6484) );
  NANDN U6974 ( .A(n6485), .B(n6484), .Z(n6486) );
  AND U6975 ( .A(n6487), .B(n6486), .Z(n6488) );
  OR U6976 ( .A(n6489), .B(n6488), .Z(n6490) );
  NAND U6977 ( .A(n6491), .B(n6490), .Z(n6492) );
  NANDN U6978 ( .A(n6493), .B(n6492), .Z(n6494) );
  NAND U6979 ( .A(n6495), .B(n6494), .Z(n6496) );
  NANDN U6980 ( .A(n6497), .B(n6496), .Z(n6498) );
  AND U6981 ( .A(n6499), .B(n6498), .Z(n6500) );
  OR U6982 ( .A(n6501), .B(n6500), .Z(n6502) );
  NAND U6983 ( .A(n6503), .B(n6502), .Z(n6504) );
  NANDN U6984 ( .A(n6505), .B(n6504), .Z(n6506) );
  NAND U6985 ( .A(n6507), .B(n6506), .Z(n6508) );
  NANDN U6986 ( .A(n6509), .B(n6508), .Z(n6510) );
  AND U6987 ( .A(n6511), .B(n6510), .Z(n6512) );
  OR U6988 ( .A(n6513), .B(n6512), .Z(n6514) );
  NAND U6989 ( .A(n6515), .B(n6514), .Z(n6516) );
  NANDN U6990 ( .A(n6517), .B(n6516), .Z(n6518) );
  NAND U6991 ( .A(n6519), .B(n6518), .Z(n6520) );
  NANDN U6992 ( .A(n6521), .B(n6520), .Z(n6522) );
  AND U6993 ( .A(n6523), .B(n6522), .Z(n6524) );
  OR U6994 ( .A(n6525), .B(n6524), .Z(n6526) );
  NAND U6995 ( .A(n6527), .B(n6526), .Z(n6528) );
  NANDN U6996 ( .A(n6529), .B(n6528), .Z(n6530) );
  NAND U6997 ( .A(n6531), .B(n6530), .Z(n6532) );
  NANDN U6998 ( .A(n6533), .B(n6532), .Z(n6534) );
  AND U6999 ( .A(n6535), .B(n6534), .Z(n6536) );
  OR U7000 ( .A(n6537), .B(n6536), .Z(n6538) );
  NAND U7001 ( .A(n6539), .B(n6538), .Z(n6540) );
  NANDN U7002 ( .A(n6541), .B(n6540), .Z(n6542) );
  NAND U7003 ( .A(n6543), .B(n6542), .Z(n6544) );
  NANDN U7004 ( .A(n6545), .B(n6544), .Z(n6546) );
  AND U7005 ( .A(n6547), .B(n6546), .Z(n6548) );
  OR U7006 ( .A(n6549), .B(n6548), .Z(n6550) );
  NAND U7007 ( .A(n6551), .B(n6550), .Z(n6552) );
  NANDN U7008 ( .A(n6553), .B(n6552), .Z(n6554) );
  NAND U7009 ( .A(n6555), .B(n6554), .Z(n6556) );
  NAND U7010 ( .A(n6557), .B(n6556), .Z(n6559) );
  ANDN U7011 ( .B(n6559), .A(n6558), .Z(n6560) );
  OR U7012 ( .A(n6561), .B(n6560), .Z(n6562) );
  NAND U7013 ( .A(n6563), .B(n6562), .Z(n6564) );
  NANDN U7014 ( .A(n6565), .B(n6564), .Z(n6566) );
  NAND U7015 ( .A(n6567), .B(n6566), .Z(n6568) );
  NANDN U7016 ( .A(n6569), .B(n6568), .Z(n6570) );
  AND U7017 ( .A(n6571), .B(n6570), .Z(n6572) );
  OR U7018 ( .A(n6573), .B(n6572), .Z(n6574) );
  NAND U7019 ( .A(n6575), .B(n6574), .Z(n6576) );
  NANDN U7020 ( .A(n6577), .B(n6576), .Z(n6578) );
  NAND U7021 ( .A(n6579), .B(n6578), .Z(n6580) );
  NANDN U7022 ( .A(n6581), .B(n6580), .Z(n6582) );
  AND U7023 ( .A(n6583), .B(n6582), .Z(n6584) );
  OR U7024 ( .A(n6585), .B(n6584), .Z(n6586) );
  NAND U7025 ( .A(n6587), .B(n6586), .Z(n6588) );
  NANDN U7026 ( .A(n6589), .B(n6588), .Z(n6590) );
  NAND U7027 ( .A(n6591), .B(n6590), .Z(n6592) );
  NANDN U7028 ( .A(n6593), .B(n6592), .Z(n6594) );
  AND U7029 ( .A(n6595), .B(n6594), .Z(n6596) );
  OR U7030 ( .A(n6597), .B(n6596), .Z(n6598) );
  NAND U7031 ( .A(n6599), .B(n6598), .Z(n6600) );
  NANDN U7032 ( .A(n6601), .B(n6600), .Z(n6602) );
  NAND U7033 ( .A(n6603), .B(n6602), .Z(n6604) );
  NANDN U7034 ( .A(n6605), .B(n6604), .Z(n6606) );
  AND U7035 ( .A(n6607), .B(n6606), .Z(n6608) );
  OR U7036 ( .A(n6609), .B(n6608), .Z(n6610) );
  NAND U7037 ( .A(n6611), .B(n6610), .Z(n6612) );
  NANDN U7038 ( .A(n6613), .B(n6612), .Z(n6614) );
  NAND U7039 ( .A(n6615), .B(n6614), .Z(n6616) );
  NANDN U7040 ( .A(n6617), .B(n6616), .Z(n6618) );
  AND U7041 ( .A(n6619), .B(n6618), .Z(n6620) );
  OR U7042 ( .A(n6621), .B(n6620), .Z(n6622) );
  NAND U7043 ( .A(n6623), .B(n6622), .Z(n6624) );
  NANDN U7044 ( .A(n6625), .B(n6624), .Z(n6626) );
  NAND U7045 ( .A(n6627), .B(n6626), .Z(n6628) );
  NANDN U7046 ( .A(n6629), .B(n6628), .Z(n6630) );
  AND U7047 ( .A(n6631), .B(n6630), .Z(n6632) );
  OR U7048 ( .A(n6633), .B(n6632), .Z(n6634) );
  NAND U7049 ( .A(n6635), .B(n6634), .Z(n6636) );
  NANDN U7050 ( .A(n6637), .B(n6636), .Z(n6638) );
  NAND U7051 ( .A(n6639), .B(n6638), .Z(n6640) );
  NANDN U7052 ( .A(n6641), .B(n6640), .Z(n6642) );
  AND U7053 ( .A(n6643), .B(n6642), .Z(n6644) );
  OR U7054 ( .A(n6645), .B(n6644), .Z(n6646) );
  NAND U7055 ( .A(n6647), .B(n6646), .Z(n6648) );
  NANDN U7056 ( .A(n6649), .B(n6648), .Z(n6650) );
  NAND U7057 ( .A(n6651), .B(n6650), .Z(n6652) );
  NANDN U7058 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U7059 ( .A(n6655), .B(n6654), .Z(n6656) );
  OR U7060 ( .A(n6657), .B(n6656), .Z(n6658) );
  NAND U7061 ( .A(n6659), .B(n6658), .Z(n6660) );
  NANDN U7062 ( .A(n6661), .B(n6660), .Z(n6662) );
  NAND U7063 ( .A(n6663), .B(n6662), .Z(n6664) );
  NANDN U7064 ( .A(n6665), .B(n6664), .Z(n6666) );
  AND U7065 ( .A(n6667), .B(n6666), .Z(n6668) );
  OR U7066 ( .A(n6669), .B(n6668), .Z(n6670) );
  NAND U7067 ( .A(n6671), .B(n6670), .Z(n6672) );
  NANDN U7068 ( .A(n6673), .B(n6672), .Z(n6674) );
  NAND U7069 ( .A(n6675), .B(n6674), .Z(n6676) );
  NANDN U7070 ( .A(n6677), .B(n6676), .Z(n6678) );
  AND U7071 ( .A(n6679), .B(n6678), .Z(n6680) );
  OR U7072 ( .A(n6681), .B(n6680), .Z(n6682) );
  NAND U7073 ( .A(n6683), .B(n6682), .Z(n6684) );
  NANDN U7074 ( .A(n6685), .B(n6684), .Z(n6686) );
  NAND U7075 ( .A(n6687), .B(n6686), .Z(n6688) );
  NANDN U7076 ( .A(n6689), .B(n6688), .Z(n6690) );
  AND U7077 ( .A(n6691), .B(n6690), .Z(n6692) );
  OR U7078 ( .A(n6693), .B(n6692), .Z(n6694) );
  NAND U7079 ( .A(n6695), .B(n6694), .Z(n6696) );
  NAND U7080 ( .A(n6716), .B(n6715), .Z(n6717) );
  NANDN U7081 ( .A(n6718), .B(n6717), .Z(n6719) );
  AND U7082 ( .A(n6720), .B(n6719), .Z(n6721) );
  OR U7083 ( .A(n6722), .B(n6721), .Z(n6723) );
  NAND U7084 ( .A(n6724), .B(n6723), .Z(n6725) );
  NANDN U7085 ( .A(n6726), .B(n6725), .Z(n6727) );
  NAND U7086 ( .A(n6728), .B(n6727), .Z(n6729) );
  NANDN U7087 ( .A(n6730), .B(n6729), .Z(n6731) );
  AND U7088 ( .A(n6732), .B(n6731), .Z(n6733) );
  OR U7089 ( .A(n6734), .B(n6733), .Z(n6735) );
  NAND U7090 ( .A(n6736), .B(n6735), .Z(n6737) );
  NANDN U7091 ( .A(n6738), .B(n6737), .Z(n6739) );
  NAND U7092 ( .A(n6740), .B(n6739), .Z(n6741) );
  NANDN U7093 ( .A(n6742), .B(n6741), .Z(n6743) );
  AND U7094 ( .A(n6744), .B(n6743), .Z(n6745) );
  OR U7095 ( .A(n6746), .B(n6745), .Z(n6747) );
  NAND U7096 ( .A(n6748), .B(n6747), .Z(n6749) );
  NANDN U7097 ( .A(n6750), .B(n6749), .Z(n6751) );
  NAND U7098 ( .A(n6752), .B(n6751), .Z(n6753) );
  NANDN U7099 ( .A(n6754), .B(n6753), .Z(n6755) );
  AND U7100 ( .A(n6756), .B(n6755), .Z(n6757) );
  OR U7101 ( .A(n6758), .B(n6757), .Z(n6759) );
  NAND U7102 ( .A(n6760), .B(n6759), .Z(n6761) );
  NANDN U7103 ( .A(n6762), .B(n6761), .Z(n6763) );
  NAND U7104 ( .A(n6764), .B(n6763), .Z(n6765) );
  NANDN U7105 ( .A(n6766), .B(n6765), .Z(n6767) );
  AND U7106 ( .A(n6768), .B(n6767), .Z(n6769) );
  OR U7107 ( .A(n6770), .B(n6769), .Z(n6771) );
  NAND U7108 ( .A(n6772), .B(n6771), .Z(n6773) );
  NANDN U7109 ( .A(n6774), .B(n6773), .Z(n6775) );
  NAND U7110 ( .A(n6776), .B(n6775), .Z(n6777) );
  NANDN U7111 ( .A(n6778), .B(n6777), .Z(n6779) );
  AND U7112 ( .A(n6780), .B(n6779), .Z(n6781) );
  OR U7113 ( .A(n6782), .B(n6781), .Z(n6783) );
  NAND U7114 ( .A(n6784), .B(n6783), .Z(n6785) );
  NANDN U7115 ( .A(n6786), .B(n6785), .Z(n6787) );
  NAND U7116 ( .A(n6788), .B(n6787), .Z(n6789) );
  NANDN U7117 ( .A(n6790), .B(n6789), .Z(n6791) );
  AND U7118 ( .A(n6792), .B(n6791), .Z(n6793) );
  OR U7119 ( .A(n6794), .B(n6793), .Z(n6795) );
  NAND U7120 ( .A(n6796), .B(n6795), .Z(n6797) );
  NANDN U7121 ( .A(n6798), .B(n6797), .Z(n6799) );
  NAND U7122 ( .A(n6800), .B(n6799), .Z(n6801) );
  NANDN U7123 ( .A(n6802), .B(n6801), .Z(n6803) );
  AND U7124 ( .A(n6804), .B(n6803), .Z(n6805) );
  OR U7125 ( .A(n6806), .B(n6805), .Z(n6807) );
  NAND U7126 ( .A(n6808), .B(n6807), .Z(n6809) );
  NANDN U7127 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND U7128 ( .A(n6812), .B(n6811), .Z(n6813) );
  NANDN U7129 ( .A(n6814), .B(n6813), .Z(n6815) );
  AND U7130 ( .A(n6816), .B(n6815), .Z(n6817) );
  OR U7131 ( .A(n6818), .B(n6817), .Z(n6819) );
  NAND U7132 ( .A(n6820), .B(n6819), .Z(n6821) );
  NANDN U7133 ( .A(n6822), .B(n6821), .Z(n6823) );
  NAND U7134 ( .A(n6824), .B(n6823), .Z(n6825) );
  NANDN U7135 ( .A(n6826), .B(n6825), .Z(n6827) );
  AND U7136 ( .A(n6828), .B(n6827), .Z(n6829) );
  OR U7137 ( .A(n6830), .B(n6829), .Z(n6831) );
  NAND U7138 ( .A(n6832), .B(n6831), .Z(n6833) );
  NANDN U7139 ( .A(n6834), .B(n6833), .Z(n6835) );
  NAND U7140 ( .A(n6836), .B(n6835), .Z(n6837) );
  NANDN U7141 ( .A(n6838), .B(n6837), .Z(n6840) );
  ANDN U7142 ( .B(n6840), .A(n6839), .Z(n6841) );
  OR U7143 ( .A(n6842), .B(n6841), .Z(n6843) );
  NAND U7144 ( .A(n6844), .B(n6843), .Z(n6845) );
  NANDN U7145 ( .A(n6846), .B(n6845), .Z(n6847) );
  NAND U7146 ( .A(n6848), .B(n6847), .Z(n6849) );
  NANDN U7147 ( .A(n6850), .B(n6849), .Z(n6851) );
  AND U7148 ( .A(n6852), .B(n6851), .Z(n6853) );
  OR U7149 ( .A(n6854), .B(n6853), .Z(n6855) );
  NAND U7150 ( .A(n6856), .B(n6855), .Z(n6857) );
  NANDN U7151 ( .A(n6858), .B(n6857), .Z(n6859) );
  NAND U7152 ( .A(n6860), .B(n6859), .Z(n6861) );
  NANDN U7153 ( .A(n6862), .B(n6861), .Z(n6863) );
  AND U7154 ( .A(n6864), .B(n6863), .Z(n6865) );
  OR U7155 ( .A(n6866), .B(n6865), .Z(n6867) );
  NAND U7156 ( .A(n6868), .B(n6867), .Z(n6869) );
  NANDN U7157 ( .A(n6870), .B(n6869), .Z(n6871) );
  NAND U7158 ( .A(n6872), .B(n6871), .Z(n6873) );
  NANDN U7159 ( .A(n6874), .B(n6873), .Z(n6875) );
  AND U7160 ( .A(n6876), .B(n6875), .Z(n6877) );
  OR U7161 ( .A(n6878), .B(n6877), .Z(n6879) );
  NAND U7162 ( .A(n6880), .B(n6879), .Z(n6881) );
  NANDN U7163 ( .A(n6882), .B(n6881), .Z(n6883) );
  NAND U7164 ( .A(n6884), .B(n6883), .Z(n6885) );
  NANDN U7165 ( .A(n6886), .B(n6885), .Z(n6887) );
  AND U7166 ( .A(n6888), .B(n6887), .Z(n6889) );
  OR U7167 ( .A(n6890), .B(n6889), .Z(n6891) );
  NAND U7168 ( .A(n6892), .B(n6891), .Z(n6893) );
  NANDN U7169 ( .A(n6894), .B(n6893), .Z(n6895) );
  NAND U7170 ( .A(n6896), .B(n6895), .Z(n6897) );
  NANDN U7171 ( .A(n6898), .B(n6897), .Z(n6899) );
  AND U7172 ( .A(n6900), .B(n6899), .Z(n6901) );
  OR U7173 ( .A(n6902), .B(n6901), .Z(n6903) );
  NAND U7174 ( .A(n6904), .B(n6903), .Z(n6905) );
  NANDN U7175 ( .A(n6906), .B(n6905), .Z(n6907) );
  NAND U7176 ( .A(n6908), .B(n6907), .Z(n6909) );
  NANDN U7177 ( .A(n6910), .B(n6909), .Z(n6911) );
  AND U7178 ( .A(n6912), .B(n6911), .Z(n6913) );
  OR U7179 ( .A(n6914), .B(n6913), .Z(n6915) );
  NAND U7180 ( .A(n6916), .B(n6915), .Z(n6917) );
  NANDN U7181 ( .A(n6918), .B(n6917), .Z(n6919) );
  NAND U7182 ( .A(n6920), .B(n6919), .Z(n6921) );
  NANDN U7183 ( .A(n6922), .B(n6921), .Z(n6923) );
  AND U7184 ( .A(n6924), .B(n6923), .Z(n6925) );
  OR U7185 ( .A(n6926), .B(n6925), .Z(n6927) );
  NAND U7186 ( .A(n6928), .B(n6927), .Z(n6929) );
  NANDN U7187 ( .A(n6930), .B(n6929), .Z(n6931) );
  NAND U7188 ( .A(n6932), .B(n6931), .Z(n6933) );
  NANDN U7189 ( .A(n6934), .B(n6933), .Z(n6935) );
  AND U7190 ( .A(n6936), .B(n6935), .Z(n6937) );
  OR U7191 ( .A(n6938), .B(n6937), .Z(n6939) );
  NAND U7192 ( .A(n6940), .B(n6939), .Z(n6941) );
  NANDN U7193 ( .A(n6942), .B(n6941), .Z(n6943) );
  NAND U7194 ( .A(n6944), .B(n6943), .Z(n6945) );
  NANDN U7195 ( .A(n6946), .B(n6945), .Z(n6947) );
  AND U7196 ( .A(n6948), .B(n6947), .Z(n6949) );
  OR U7197 ( .A(n6950), .B(n6949), .Z(n6951) );
  NAND U7198 ( .A(n6952), .B(n6951), .Z(n6953) );
  NANDN U7199 ( .A(n6954), .B(n6953), .Z(n6955) );
  NAND U7200 ( .A(n6956), .B(n6955), .Z(n6957) );
  NANDN U7201 ( .A(n6958), .B(n6957), .Z(n6959) );
  AND U7202 ( .A(n6960), .B(n6959), .Z(n6961) );
  OR U7203 ( .A(n6962), .B(n6961), .Z(n6963) );
  NAND U7204 ( .A(n6964), .B(n6963), .Z(n6965) );
  NANDN U7205 ( .A(n6966), .B(n6965), .Z(n6967) );
  NAND U7206 ( .A(n6968), .B(n6967), .Z(n6969) );
  NANDN U7207 ( .A(n6970), .B(n6969), .Z(n6971) );
  AND U7208 ( .A(n6972), .B(n6971), .Z(n6973) );
  OR U7209 ( .A(n6974), .B(n6973), .Z(n6975) );
  NAND U7210 ( .A(n6976), .B(n6975), .Z(n6977) );
  NANDN U7211 ( .A(n6978), .B(n6977), .Z(n6979) );
  NAND U7212 ( .A(n6980), .B(n6979), .Z(n6981) );
  NANDN U7213 ( .A(n6982), .B(n6981), .Z(n6983) );
  AND U7214 ( .A(n6984), .B(n6983), .Z(n6985) );
  OR U7215 ( .A(n6986), .B(n6985), .Z(n6987) );
  NAND U7216 ( .A(n6988), .B(n6987), .Z(n6989) );
  NANDN U7217 ( .A(n6990), .B(n6989), .Z(n6991) );
  NAND U7218 ( .A(n6992), .B(n6991), .Z(n6993) );
  NANDN U7219 ( .A(n6994), .B(n6993), .Z(n6995) );
  AND U7220 ( .A(n6996), .B(n6995), .Z(n6997) );
  OR U7221 ( .A(n6998), .B(n6997), .Z(n6999) );
  NAND U7222 ( .A(n7000), .B(n6999), .Z(n7001) );
  NANDN U7223 ( .A(n7002), .B(n7001), .Z(n7003) );
  NAND U7224 ( .A(n7004), .B(n7003), .Z(n7005) );
  NANDN U7225 ( .A(n7006), .B(n7005), .Z(n7007) );
  AND U7226 ( .A(n7008), .B(n7007), .Z(n7009) );
  OR U7227 ( .A(n7010), .B(n7009), .Z(n7011) );
  NAND U7228 ( .A(n7012), .B(n7011), .Z(n7013) );
  NANDN U7229 ( .A(n7014), .B(n7013), .Z(n7015) );
  NAND U7230 ( .A(n7016), .B(n7015), .Z(n7017) );
  NANDN U7231 ( .A(n7018), .B(n7017), .Z(n7019) );
  AND U7232 ( .A(n7020), .B(n7019), .Z(n7021) );
  OR U7233 ( .A(n7022), .B(n7021), .Z(n7023) );
  NAND U7234 ( .A(n7024), .B(n7023), .Z(n7025) );
  NANDN U7235 ( .A(n7026), .B(n7025), .Z(n7027) );
  NAND U7236 ( .A(n7028), .B(n7027), .Z(n7029) );
  NANDN U7237 ( .A(n7030), .B(n7029), .Z(n7031) );
  AND U7238 ( .A(n7032), .B(n7031), .Z(n7033) );
  OR U7239 ( .A(n7034), .B(n7033), .Z(n7035) );
  IV U7240 ( .A(n7070), .Z(n7071) );
  AND U7241 ( .A(n7072), .B(n7071), .Z(n7074) );
  NANDN U7242 ( .A(n7074), .B(n7073), .Z(n7075) );
  NAND U7243 ( .A(n7076), .B(n7075), .Z(n7077) );
  NANDN U7244 ( .A(n7078), .B(n7077), .Z(n7079) );
  NAND U7245 ( .A(n7080), .B(n7079), .Z(n7081) );
  NANDN U7246 ( .A(n7082), .B(n7081), .Z(n7083) );
  AND U7247 ( .A(n7084), .B(n7083), .Z(n7087) );
  IV U7248 ( .A(n7085), .Z(n7086) );
  NANDN U7249 ( .A(n7087), .B(n7086), .Z(n7089) );
  AND U7250 ( .A(n7089), .B(n7088), .Z(n7090) );
  OR U7251 ( .A(n7091), .B(n7090), .Z(n7092) );
  AND U7252 ( .A(n7093), .B(n7092), .Z(n7094) );
  ANDN U7253 ( .B(n7095), .A(n7094), .Z(n7096) );
  NANDN U7254 ( .A(n7097), .B(n7096), .Z(n7098) );
  NAND U7255 ( .A(n7099), .B(n7098), .Z(n7100) );
  NAND U7256 ( .A(n7101), .B(n7100), .Z(n7104) );
  IV U7257 ( .A(n7102), .Z(n7103) );
  AND U7258 ( .A(n7104), .B(n7103), .Z(n7106) );
  OR U7259 ( .A(n7106), .B(n7105), .Z(n7107) );
  NAND U7260 ( .A(n7108), .B(n7107), .Z(n7109) );
  NANDN U7261 ( .A(n7110), .B(n7109), .Z(n7111) );
  NAND U7262 ( .A(n7112), .B(n7111), .Z(n7113) );
  NANDN U7263 ( .A(n7114), .B(n7113), .Z(n7115) );
  AND U7264 ( .A(n7116), .B(n7115), .Z(n7117) );
  OR U7265 ( .A(n7118), .B(n7117), .Z(n7119) );
  NAND U7266 ( .A(n7120), .B(n7119), .Z(n7121) );
  NANDN U7267 ( .A(n7122), .B(n7121), .Z(n7125) );
  IV U7268 ( .A(n7123), .Z(n7124) );
  AND U7269 ( .A(n7125), .B(n7124), .Z(n7127) );
  NAND U7270 ( .A(n7127), .B(n7126), .Z(n7128) );
  NAND U7271 ( .A(n7129), .B(n7128), .Z(n7131) );
  OR U7272 ( .A(n7131), .B(n7130), .Z(n7132) );
  NAND U7273 ( .A(n7133), .B(n7132), .Z(n7134) );
  NAND U7274 ( .A(n7135), .B(n7134), .Z(n7136) );
  NAND U7275 ( .A(n7137), .B(n7136), .Z(n7138) );
  NANDN U7276 ( .A(n7139), .B(n7138), .Z(n7142) );
  IV U7277 ( .A(n7140), .Z(n7141) );
  AND U7278 ( .A(n7142), .B(n7141), .Z(n7144) );
  OR U7279 ( .A(n7144), .B(n7143), .Z(n7145) );
  NAND U7280 ( .A(n7146), .B(n7145), .Z(n7147) );
  NANDN U7281 ( .A(n7148), .B(n7147), .Z(n7149) );
  NAND U7282 ( .A(n7150), .B(n7149), .Z(n7151) );
  NANDN U7283 ( .A(n7152), .B(n7151), .Z(n7155) );
  IV U7284 ( .A(n7153), .Z(n7154) );
  AND U7285 ( .A(n7155), .B(n7154), .Z(n7157) );
  NANDN U7286 ( .A(n7157), .B(n7156), .Z(n7158) );
  NAND U7287 ( .A(n7159), .B(n7158), .Z(n7160) );
  NAND U7288 ( .A(n7161), .B(n7160), .Z(n7163) );
  NAND U7289 ( .A(n7163), .B(n7162), .Z(n7164) );
  NANDN U7290 ( .A(n7165), .B(n7164), .Z(n7168) );
  IV U7291 ( .A(n7166), .Z(n7167) );
  AND U7292 ( .A(n7168), .B(n7167), .Z(n7170) );
  NAND U7293 ( .A(n7170), .B(n7169), .Z(n7171) );
  NAND U7294 ( .A(n7172), .B(n7171), .Z(n7174) );
  OR U7295 ( .A(n7174), .B(n7173), .Z(n7177) );
  IV U7296 ( .A(n7175), .Z(n7176) );
  AND U7297 ( .A(n7177), .B(n7176), .Z(n7179) );
  OR U7298 ( .A(n7179), .B(n7178), .Z(n7180) );
  AND U7299 ( .A(n7181), .B(n7180), .Z(n7183) );
  NANDN U7300 ( .A(n7183), .B(n7182), .Z(n7184) );
  NANDN U7301 ( .A(n7185), .B(n7184), .Z(n7186) );
  NAND U7302 ( .A(n7187), .B(n7186), .Z(n7188) );
  NANDN U7303 ( .A(n7189), .B(n7188), .Z(n7190) );
  AND U7304 ( .A(n7191), .B(n7190), .Z(n7192) );
  OR U7305 ( .A(n7193), .B(n7192), .Z(n7194) );
  NAND U7306 ( .A(n7195), .B(n7194), .Z(n7196) );
  NAND U7307 ( .A(n7197), .B(n7196), .Z(n7198) );
  NAND U7308 ( .A(n7199), .B(n7198), .Z(n7200) );
  NANDN U7309 ( .A(n7201), .B(n7200), .Z(n7202) );
  NANDN U7310 ( .A(n7203), .B(n7202), .Z(n7205) );
  IV U7311 ( .A(n7206), .Z(n7207) );
  NANDN U7312 ( .A(n7239), .B(n7238), .Z(n7242) );
  IV U7313 ( .A(n7240), .Z(n7241) );
  AND U7314 ( .A(n7242), .B(n7241), .Z(n7243) );
  NAND U7315 ( .A(n7244), .B(n7243), .Z(n7245) );
  NAND U7316 ( .A(n7246), .B(n7245), .Z(n7248) );
  OR U7317 ( .A(n7248), .B(n7247), .Z(n7249) );
  NAND U7318 ( .A(n7250), .B(n7249), .Z(n7251) );
  NANDN U7319 ( .A(n7252), .B(n7251), .Z(n7253) );
  AND U7320 ( .A(n7254), .B(n7253), .Z(n7255) );
  OR U7321 ( .A(n7256), .B(n7255), .Z(n7257) );
  NAND U7322 ( .A(n7258), .B(n7257), .Z(n7259) );
  NAND U7323 ( .A(n7260), .B(n7259), .Z(n7261) );
  AND U7324 ( .A(n7262), .B(n7261), .Z(n7263) );
  NAND U7325 ( .A(n7264), .B(n7263), .Z(n7265) );
  NANDN U7326 ( .A(n7266), .B(n7265), .Z(n7268) );
  AND U7327 ( .A(n7268), .B(n7267), .Z(n7271) );
  IV U7328 ( .A(n7269), .Z(n7270) );
  NAND U7329 ( .A(n7286), .B(n7285), .Z(n7287) );
  NANDN U7330 ( .A(n7288), .B(n7287), .Z(n7289) );
  AND U7331 ( .A(n7290), .B(n7289), .Z(n7292) );
  NANDN U7332 ( .A(n7292), .B(n7291), .Z(n7293) );
  AND U7333 ( .A(n7294), .B(n7293), .Z(n7296) );
  NANDN U7334 ( .A(n7296), .B(n7295), .Z(n7297) );
  NAND U7335 ( .A(n7298), .B(n7297), .Z(n7299) );
  NANDN U7336 ( .A(n7300), .B(n7299), .Z(n7301) );
  NAND U7337 ( .A(n7302), .B(n7301), .Z(n7305) );
  IV U7338 ( .A(n7303), .Z(n7304) );
  AND U7339 ( .A(n7305), .B(n7304), .Z(n7307) );
  OR U7340 ( .A(n7307), .B(n7306), .Z(n7308) );
  NANDN U7341 ( .A(n7309), .B(n7308), .Z(n7310) );
  NAND U7342 ( .A(n7311), .B(n7310), .Z(n7313) );
  AND U7343 ( .A(n7313), .B(n7312), .Z(n7314) );
  NAND U7344 ( .A(n7315), .B(n7314), .Z(n7316) );
  NAND U7345 ( .A(n7317), .B(n7316), .Z(n7318) );
  NAND U7346 ( .A(n7319), .B(n7318), .Z(n7320) );
endmodule

