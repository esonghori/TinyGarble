
module mult_N64_CC32 ( clk, rst, a, b, c );
  input [63:0] a;
  input [1:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479;
  wire   [63:2] swire;
  wire   [127:64] sreg;

  DFF \sreg_reg[64]  ( .D(swire[2]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[3]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[96]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[97]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[98]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[99]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[100]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[101]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[102]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[103]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[104]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[105]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[106]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[107]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[108]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[109]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[110]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[111]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[112]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[113]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[114]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[115]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[116]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[117]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[118]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[119]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[120]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[121]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[122]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[123]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[124]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[125]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[3]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[2]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U5 ( .A(n1), .B(n2), .Z(swire[9]) );
  XNOR U6 ( .A(n3), .B(n4), .Z(swire[8]) );
  XNOR U7 ( .A(n5), .B(n6), .Z(swire[7]) );
  XNOR U8 ( .A(n7), .B(n8), .Z(swire[6]) );
  XOR U9 ( .A(n9), .B(n10), .Z(swire[63]) );
  AND U10 ( .A(a[63]), .B(b[0]), .Z(n10) );
  AND U11 ( .A(b[1]), .B(a[62]), .Z(n9) );
  XOR U12 ( .A(n11), .B(n12), .Z(swire[62]) );
  AND U13 ( .A(a[62]), .B(b[0]), .Z(n12) );
  AND U14 ( .A(b[1]), .B(a[61]), .Z(n11) );
  XOR U15 ( .A(n13), .B(n14), .Z(swire[61]) );
  XOR U16 ( .A(sreg[125]), .B(n15), .Z(n14) );
  AND U17 ( .A(b[1]), .B(a[60]), .Z(n15) );
  AND U18 ( .A(a[61]), .B(b[0]), .Z(n13) );
  XOR U19 ( .A(n16), .B(n17), .Z(swire[60]) );
  XOR U20 ( .A(sreg[124]), .B(n18), .Z(n17) );
  AND U21 ( .A(b[1]), .B(a[59]), .Z(n18) );
  AND U22 ( .A(a[60]), .B(b[0]), .Z(n16) );
  XNOR U23 ( .A(n19), .B(n20), .Z(swire[5]) );
  XOR U24 ( .A(n21), .B(n22), .Z(swire[59]) );
  XOR U25 ( .A(sreg[123]), .B(n23), .Z(n22) );
  XOR U26 ( .A(n23), .B(n24), .Z(n21) );
  XOR U27 ( .A(n25), .B(n26), .Z(n24) );
  AND U28 ( .A(a[59]), .B(b[0]), .Z(n26) );
  AND U29 ( .A(b[1]), .B(a[58]), .Z(n25) );
  XOR U30 ( .A(n27), .B(n28), .Z(n23) );
  ANDN U31 ( .B(n29), .A(n30), .Z(n27) );
  XNOR U32 ( .A(n29), .B(n30), .Z(swire[58]) );
  XOR U33 ( .A(sreg[122]), .B(n31), .Z(n30) );
  XOR U34 ( .A(n31), .B(n32), .Z(n29) );
  XOR U35 ( .A(n33), .B(n34), .Z(n32) );
  NAND U36 ( .A(b[0]), .B(a[58]), .Z(n34) );
  AND U37 ( .A(b[1]), .B(a[57]), .Z(n33) );
  IV U38 ( .A(n28), .Z(n31) );
  XOR U39 ( .A(n35), .B(n36), .Z(n28) );
  ANDN U40 ( .B(n37), .A(n38), .Z(n35) );
  XNOR U41 ( .A(n37), .B(n38), .Z(swire[57]) );
  XOR U42 ( .A(sreg[121]), .B(n39), .Z(n38) );
  XOR U43 ( .A(n39), .B(n40), .Z(n37) );
  XOR U44 ( .A(n41), .B(n42), .Z(n40) );
  NAND U45 ( .A(b[0]), .B(a[57]), .Z(n42) );
  AND U46 ( .A(b[1]), .B(a[56]), .Z(n41) );
  IV U47 ( .A(n36), .Z(n39) );
  XOR U48 ( .A(n43), .B(n44), .Z(n36) );
  ANDN U49 ( .B(n45), .A(n46), .Z(n43) );
  XNOR U50 ( .A(n45), .B(n46), .Z(swire[56]) );
  XOR U51 ( .A(sreg[120]), .B(n47), .Z(n46) );
  XOR U52 ( .A(n47), .B(n48), .Z(n45) );
  XOR U53 ( .A(n49), .B(n50), .Z(n48) );
  NAND U54 ( .A(b[0]), .B(a[56]), .Z(n50) );
  AND U55 ( .A(b[1]), .B(a[55]), .Z(n49) );
  IV U56 ( .A(n44), .Z(n47) );
  XOR U57 ( .A(n51), .B(n52), .Z(n44) );
  ANDN U58 ( .B(n53), .A(n54), .Z(n51) );
  XNOR U59 ( .A(n53), .B(n54), .Z(swire[55]) );
  XOR U60 ( .A(sreg[119]), .B(n55), .Z(n54) );
  XOR U61 ( .A(n55), .B(n56), .Z(n53) );
  XOR U62 ( .A(n57), .B(n58), .Z(n56) );
  NAND U63 ( .A(b[0]), .B(a[55]), .Z(n58) );
  AND U64 ( .A(b[1]), .B(a[54]), .Z(n57) );
  IV U65 ( .A(n52), .Z(n55) );
  XOR U66 ( .A(n59), .B(n60), .Z(n52) );
  ANDN U67 ( .B(n61), .A(n62), .Z(n59) );
  XNOR U68 ( .A(n61), .B(n62), .Z(swire[54]) );
  XOR U69 ( .A(sreg[118]), .B(n63), .Z(n62) );
  XOR U70 ( .A(n63), .B(n64), .Z(n61) );
  XOR U71 ( .A(n65), .B(n66), .Z(n64) );
  NAND U72 ( .A(b[0]), .B(a[54]), .Z(n66) );
  AND U73 ( .A(b[1]), .B(a[53]), .Z(n65) );
  IV U74 ( .A(n60), .Z(n63) );
  XOR U75 ( .A(n67), .B(n68), .Z(n60) );
  ANDN U76 ( .B(n69), .A(n70), .Z(n67) );
  XNOR U77 ( .A(n69), .B(n70), .Z(swire[53]) );
  XOR U78 ( .A(sreg[117]), .B(n71), .Z(n70) );
  XOR U79 ( .A(n71), .B(n72), .Z(n69) );
  XOR U80 ( .A(n73), .B(n74), .Z(n72) );
  NAND U81 ( .A(b[0]), .B(a[53]), .Z(n74) );
  AND U82 ( .A(b[1]), .B(a[52]), .Z(n73) );
  IV U83 ( .A(n68), .Z(n71) );
  XOR U84 ( .A(n75), .B(n76), .Z(n68) );
  ANDN U85 ( .B(n77), .A(n78), .Z(n75) );
  XNOR U86 ( .A(n77), .B(n78), .Z(swire[52]) );
  XOR U87 ( .A(sreg[116]), .B(n79), .Z(n78) );
  XOR U88 ( .A(n79), .B(n80), .Z(n77) );
  XOR U89 ( .A(n81), .B(n82), .Z(n80) );
  NAND U90 ( .A(b[0]), .B(a[52]), .Z(n82) );
  AND U91 ( .A(b[1]), .B(a[51]), .Z(n81) );
  IV U92 ( .A(n76), .Z(n79) );
  XOR U93 ( .A(n83), .B(n84), .Z(n76) );
  ANDN U94 ( .B(n85), .A(n86), .Z(n83) );
  XNOR U95 ( .A(n85), .B(n86), .Z(swire[51]) );
  XOR U96 ( .A(sreg[115]), .B(n87), .Z(n86) );
  XOR U97 ( .A(n87), .B(n88), .Z(n85) );
  XOR U98 ( .A(n89), .B(n90), .Z(n88) );
  NAND U99 ( .A(b[0]), .B(a[51]), .Z(n90) );
  AND U100 ( .A(b[1]), .B(a[50]), .Z(n89) );
  IV U101 ( .A(n84), .Z(n87) );
  XOR U102 ( .A(n91), .B(n92), .Z(n84) );
  ANDN U103 ( .B(n93), .A(n94), .Z(n91) );
  XNOR U104 ( .A(n93), .B(n94), .Z(swire[50]) );
  XOR U105 ( .A(sreg[114]), .B(n95), .Z(n94) );
  XOR U106 ( .A(n95), .B(n96), .Z(n93) );
  XOR U107 ( .A(n97), .B(n98), .Z(n96) );
  NAND U108 ( .A(b[0]), .B(a[50]), .Z(n98) );
  AND U109 ( .A(b[1]), .B(a[49]), .Z(n97) );
  IV U110 ( .A(n92), .Z(n95) );
  XOR U111 ( .A(n99), .B(n100), .Z(n92) );
  ANDN U112 ( .B(n101), .A(n102), .Z(n99) );
  XNOR U113 ( .A(n103), .B(n104), .Z(swire[4]) );
  XNOR U114 ( .A(n101), .B(n102), .Z(swire[49]) );
  XOR U115 ( .A(sreg[113]), .B(n105), .Z(n102) );
  XOR U116 ( .A(n105), .B(n106), .Z(n101) );
  XOR U117 ( .A(n107), .B(n108), .Z(n106) );
  NAND U118 ( .A(b[0]), .B(a[49]), .Z(n108) );
  AND U119 ( .A(b[1]), .B(a[48]), .Z(n107) );
  IV U120 ( .A(n100), .Z(n105) );
  XOR U121 ( .A(n109), .B(n110), .Z(n100) );
  ANDN U122 ( .B(n111), .A(n112), .Z(n109) );
  XNOR U123 ( .A(n111), .B(n112), .Z(swire[48]) );
  XOR U124 ( .A(sreg[112]), .B(n113), .Z(n112) );
  XOR U125 ( .A(n113), .B(n114), .Z(n111) );
  XOR U126 ( .A(n115), .B(n116), .Z(n114) );
  NAND U127 ( .A(b[0]), .B(a[48]), .Z(n116) );
  AND U128 ( .A(b[1]), .B(a[47]), .Z(n115) );
  IV U129 ( .A(n110), .Z(n113) );
  XOR U130 ( .A(n117), .B(n118), .Z(n110) );
  ANDN U131 ( .B(n119), .A(n120), .Z(n117) );
  XNOR U132 ( .A(n119), .B(n120), .Z(swire[47]) );
  XOR U133 ( .A(sreg[111]), .B(n121), .Z(n120) );
  XOR U134 ( .A(n121), .B(n122), .Z(n119) );
  XOR U135 ( .A(n123), .B(n124), .Z(n122) );
  NAND U136 ( .A(b[0]), .B(a[47]), .Z(n124) );
  AND U137 ( .A(b[1]), .B(a[46]), .Z(n123) );
  IV U138 ( .A(n118), .Z(n121) );
  XOR U139 ( .A(n125), .B(n126), .Z(n118) );
  ANDN U140 ( .B(n127), .A(n128), .Z(n125) );
  XNOR U141 ( .A(n127), .B(n128), .Z(swire[46]) );
  XOR U142 ( .A(sreg[110]), .B(n129), .Z(n128) );
  XOR U143 ( .A(n129), .B(n130), .Z(n127) );
  XOR U144 ( .A(n131), .B(n132), .Z(n130) );
  NAND U145 ( .A(b[0]), .B(a[46]), .Z(n132) );
  AND U146 ( .A(b[1]), .B(a[45]), .Z(n131) );
  IV U147 ( .A(n126), .Z(n129) );
  XOR U148 ( .A(n133), .B(n134), .Z(n126) );
  ANDN U149 ( .B(n135), .A(n136), .Z(n133) );
  XNOR U150 ( .A(n135), .B(n136), .Z(swire[45]) );
  XOR U151 ( .A(sreg[109]), .B(n137), .Z(n136) );
  XOR U152 ( .A(n137), .B(n138), .Z(n135) );
  XOR U153 ( .A(n139), .B(n140), .Z(n138) );
  NAND U154 ( .A(b[0]), .B(a[45]), .Z(n140) );
  AND U155 ( .A(b[1]), .B(a[44]), .Z(n139) );
  IV U156 ( .A(n134), .Z(n137) );
  XOR U157 ( .A(n141), .B(n142), .Z(n134) );
  ANDN U158 ( .B(n143), .A(n144), .Z(n141) );
  XNOR U159 ( .A(n143), .B(n144), .Z(swire[44]) );
  XOR U160 ( .A(sreg[108]), .B(n145), .Z(n144) );
  XOR U161 ( .A(n145), .B(n146), .Z(n143) );
  XOR U162 ( .A(n147), .B(n148), .Z(n146) );
  NAND U163 ( .A(b[0]), .B(a[44]), .Z(n148) );
  AND U164 ( .A(b[1]), .B(a[43]), .Z(n147) );
  IV U165 ( .A(n142), .Z(n145) );
  XOR U166 ( .A(n149), .B(n150), .Z(n142) );
  ANDN U167 ( .B(n151), .A(n152), .Z(n149) );
  XNOR U168 ( .A(n151), .B(n152), .Z(swire[43]) );
  XOR U169 ( .A(sreg[107]), .B(n153), .Z(n152) );
  XOR U170 ( .A(n153), .B(n154), .Z(n151) );
  XOR U171 ( .A(n155), .B(n156), .Z(n154) );
  NAND U172 ( .A(b[0]), .B(a[43]), .Z(n156) );
  AND U173 ( .A(b[1]), .B(a[42]), .Z(n155) );
  IV U174 ( .A(n150), .Z(n153) );
  XOR U175 ( .A(n157), .B(n158), .Z(n150) );
  ANDN U176 ( .B(n159), .A(n160), .Z(n157) );
  XNOR U177 ( .A(n159), .B(n160), .Z(swire[42]) );
  XOR U178 ( .A(sreg[106]), .B(n161), .Z(n160) );
  XOR U179 ( .A(n161), .B(n162), .Z(n159) );
  XOR U180 ( .A(n163), .B(n164), .Z(n162) );
  NAND U181 ( .A(b[0]), .B(a[42]), .Z(n164) );
  AND U182 ( .A(b[1]), .B(a[41]), .Z(n163) );
  IV U183 ( .A(n158), .Z(n161) );
  XOR U184 ( .A(n165), .B(n166), .Z(n158) );
  ANDN U185 ( .B(n167), .A(n168), .Z(n165) );
  XNOR U186 ( .A(n167), .B(n168), .Z(swire[41]) );
  XOR U187 ( .A(sreg[105]), .B(n169), .Z(n168) );
  XOR U188 ( .A(n169), .B(n170), .Z(n167) );
  XOR U189 ( .A(n171), .B(n172), .Z(n170) );
  NAND U190 ( .A(b[0]), .B(a[41]), .Z(n172) );
  AND U191 ( .A(b[1]), .B(a[40]), .Z(n171) );
  IV U192 ( .A(n166), .Z(n169) );
  XOR U193 ( .A(n173), .B(n174), .Z(n166) );
  ANDN U194 ( .B(n175), .A(n176), .Z(n173) );
  XNOR U195 ( .A(n175), .B(n176), .Z(swire[40]) );
  XOR U196 ( .A(sreg[104]), .B(n177), .Z(n176) );
  XOR U197 ( .A(n177), .B(n178), .Z(n175) );
  XOR U198 ( .A(n179), .B(n180), .Z(n178) );
  NAND U199 ( .A(b[0]), .B(a[40]), .Z(n180) );
  AND U200 ( .A(b[1]), .B(a[39]), .Z(n179) );
  IV U201 ( .A(n174), .Z(n177) );
  XOR U202 ( .A(n181), .B(n182), .Z(n174) );
  ANDN U203 ( .B(n183), .A(n184), .Z(n181) );
  XNOR U204 ( .A(n185), .B(n186), .Z(swire[3]) );
  XNOR U205 ( .A(n183), .B(n184), .Z(swire[39]) );
  XOR U206 ( .A(sreg[103]), .B(n187), .Z(n184) );
  XOR U207 ( .A(n187), .B(n188), .Z(n183) );
  XOR U208 ( .A(n189), .B(n190), .Z(n188) );
  NAND U209 ( .A(b[0]), .B(a[39]), .Z(n190) );
  AND U210 ( .A(b[1]), .B(a[38]), .Z(n189) );
  IV U211 ( .A(n182), .Z(n187) );
  XOR U212 ( .A(n191), .B(n192), .Z(n182) );
  ANDN U213 ( .B(n193), .A(n194), .Z(n191) );
  XNOR U214 ( .A(n193), .B(n194), .Z(swire[38]) );
  XOR U215 ( .A(sreg[102]), .B(n195), .Z(n194) );
  XOR U216 ( .A(n195), .B(n196), .Z(n193) );
  XOR U217 ( .A(n197), .B(n198), .Z(n196) );
  NAND U218 ( .A(b[0]), .B(a[38]), .Z(n198) );
  AND U219 ( .A(b[1]), .B(a[37]), .Z(n197) );
  IV U220 ( .A(n192), .Z(n195) );
  XOR U221 ( .A(n199), .B(n200), .Z(n192) );
  ANDN U222 ( .B(n201), .A(n202), .Z(n199) );
  XNOR U223 ( .A(n201), .B(n202), .Z(swire[37]) );
  XOR U224 ( .A(sreg[101]), .B(n203), .Z(n202) );
  XOR U225 ( .A(n203), .B(n204), .Z(n201) );
  XOR U226 ( .A(n205), .B(n206), .Z(n204) );
  NAND U227 ( .A(b[0]), .B(a[37]), .Z(n206) );
  AND U228 ( .A(b[1]), .B(a[36]), .Z(n205) );
  IV U229 ( .A(n200), .Z(n203) );
  XOR U230 ( .A(n207), .B(n208), .Z(n200) );
  ANDN U231 ( .B(n209), .A(n210), .Z(n207) );
  XNOR U232 ( .A(n209), .B(n210), .Z(swire[36]) );
  XOR U233 ( .A(sreg[100]), .B(n211), .Z(n210) );
  XOR U234 ( .A(n211), .B(n212), .Z(n209) );
  XOR U235 ( .A(n213), .B(n214), .Z(n212) );
  NAND U236 ( .A(b[0]), .B(a[36]), .Z(n214) );
  AND U237 ( .A(b[1]), .B(a[35]), .Z(n213) );
  IV U238 ( .A(n208), .Z(n211) );
  XOR U239 ( .A(n215), .B(n216), .Z(n208) );
  ANDN U240 ( .B(n217), .A(n218), .Z(n215) );
  XNOR U241 ( .A(n217), .B(n218), .Z(swire[35]) );
  XOR U242 ( .A(sreg[99]), .B(n219), .Z(n218) );
  XOR U243 ( .A(n219), .B(n220), .Z(n217) );
  XOR U244 ( .A(n221), .B(n222), .Z(n220) );
  NAND U245 ( .A(b[0]), .B(a[35]), .Z(n222) );
  AND U246 ( .A(b[1]), .B(a[34]), .Z(n221) );
  IV U247 ( .A(n216), .Z(n219) );
  XOR U248 ( .A(n223), .B(n224), .Z(n216) );
  ANDN U249 ( .B(n225), .A(n226), .Z(n223) );
  XNOR U250 ( .A(n225), .B(n226), .Z(swire[34]) );
  XOR U251 ( .A(sreg[98]), .B(n227), .Z(n226) );
  XOR U252 ( .A(n227), .B(n228), .Z(n225) );
  XOR U253 ( .A(n229), .B(n230), .Z(n228) );
  NAND U254 ( .A(b[0]), .B(a[34]), .Z(n230) );
  AND U255 ( .A(b[1]), .B(a[33]), .Z(n229) );
  IV U256 ( .A(n224), .Z(n227) );
  XOR U257 ( .A(n231), .B(n232), .Z(n224) );
  ANDN U258 ( .B(n233), .A(n234), .Z(n231) );
  XNOR U259 ( .A(n233), .B(n234), .Z(swire[33]) );
  XOR U260 ( .A(sreg[97]), .B(n235), .Z(n234) );
  XOR U261 ( .A(n235), .B(n236), .Z(n233) );
  XOR U262 ( .A(n237), .B(n238), .Z(n236) );
  NAND U263 ( .A(b[0]), .B(a[33]), .Z(n238) );
  AND U264 ( .A(b[1]), .B(a[32]), .Z(n237) );
  IV U265 ( .A(n232), .Z(n235) );
  XOR U266 ( .A(n239), .B(n240), .Z(n232) );
  ANDN U267 ( .B(n241), .A(n242), .Z(n239) );
  XNOR U268 ( .A(n241), .B(n242), .Z(swire[32]) );
  XOR U269 ( .A(sreg[96]), .B(n243), .Z(n242) );
  XOR U270 ( .A(n243), .B(n244), .Z(n241) );
  XOR U271 ( .A(n245), .B(n246), .Z(n244) );
  NAND U272 ( .A(b[0]), .B(a[32]), .Z(n246) );
  AND U273 ( .A(b[1]), .B(a[31]), .Z(n245) );
  IV U274 ( .A(n240), .Z(n243) );
  XOR U275 ( .A(n247), .B(n248), .Z(n240) );
  ANDN U276 ( .B(n249), .A(n250), .Z(n247) );
  XNOR U277 ( .A(n249), .B(n250), .Z(swire[31]) );
  XOR U278 ( .A(sreg[95]), .B(n251), .Z(n250) );
  XOR U279 ( .A(n251), .B(n252), .Z(n249) );
  XOR U280 ( .A(n253), .B(n254), .Z(n252) );
  NAND U281 ( .A(b[0]), .B(a[31]), .Z(n254) );
  AND U282 ( .A(b[1]), .B(a[30]), .Z(n253) );
  IV U283 ( .A(n248), .Z(n251) );
  XOR U284 ( .A(n255), .B(n256), .Z(n248) );
  ANDN U285 ( .B(n257), .A(n258), .Z(n255) );
  XNOR U286 ( .A(n257), .B(n258), .Z(swire[30]) );
  XOR U287 ( .A(sreg[94]), .B(n259), .Z(n258) );
  XOR U288 ( .A(n259), .B(n260), .Z(n257) );
  XOR U289 ( .A(n261), .B(n262), .Z(n260) );
  NAND U290 ( .A(b[0]), .B(a[30]), .Z(n262) );
  AND U291 ( .A(b[1]), .B(a[29]), .Z(n261) );
  IV U292 ( .A(n256), .Z(n259) );
  XOR U293 ( .A(n263), .B(n264), .Z(n256) );
  ANDN U294 ( .B(n265), .A(n266), .Z(n263) );
  XNOR U295 ( .A(n267), .B(n268), .Z(swire[2]) );
  XNOR U296 ( .A(n265), .B(n266), .Z(swire[29]) );
  XOR U297 ( .A(sreg[93]), .B(n269), .Z(n266) );
  XOR U298 ( .A(n269), .B(n270), .Z(n265) );
  XOR U299 ( .A(n271), .B(n272), .Z(n270) );
  NAND U300 ( .A(b[0]), .B(a[29]), .Z(n272) );
  AND U301 ( .A(b[1]), .B(a[28]), .Z(n271) );
  IV U302 ( .A(n264), .Z(n269) );
  XOR U303 ( .A(n273), .B(n274), .Z(n264) );
  ANDN U304 ( .B(n275), .A(n276), .Z(n273) );
  XNOR U305 ( .A(n275), .B(n276), .Z(swire[28]) );
  XOR U306 ( .A(sreg[92]), .B(n277), .Z(n276) );
  XOR U307 ( .A(n277), .B(n278), .Z(n275) );
  XOR U308 ( .A(n279), .B(n280), .Z(n278) );
  NAND U309 ( .A(b[0]), .B(a[28]), .Z(n280) );
  AND U310 ( .A(b[1]), .B(a[27]), .Z(n279) );
  IV U311 ( .A(n274), .Z(n277) );
  XOR U312 ( .A(n281), .B(n282), .Z(n274) );
  ANDN U313 ( .B(n283), .A(n284), .Z(n281) );
  XNOR U314 ( .A(n283), .B(n284), .Z(swire[27]) );
  XOR U315 ( .A(sreg[91]), .B(n285), .Z(n284) );
  XOR U316 ( .A(n285), .B(n286), .Z(n283) );
  XOR U317 ( .A(n287), .B(n288), .Z(n286) );
  NAND U318 ( .A(b[0]), .B(a[27]), .Z(n288) );
  AND U319 ( .A(b[1]), .B(a[26]), .Z(n287) );
  IV U320 ( .A(n282), .Z(n285) );
  XOR U321 ( .A(n289), .B(n290), .Z(n282) );
  ANDN U322 ( .B(n291), .A(n292), .Z(n289) );
  XNOR U323 ( .A(n291), .B(n292), .Z(swire[26]) );
  XOR U324 ( .A(sreg[90]), .B(n293), .Z(n292) );
  XOR U325 ( .A(n293), .B(n294), .Z(n291) );
  XOR U326 ( .A(n295), .B(n296), .Z(n294) );
  NAND U327 ( .A(b[0]), .B(a[26]), .Z(n296) );
  AND U328 ( .A(b[1]), .B(a[25]), .Z(n295) );
  IV U329 ( .A(n290), .Z(n293) );
  XOR U330 ( .A(n297), .B(n298), .Z(n290) );
  ANDN U331 ( .B(n299), .A(n300), .Z(n297) );
  XNOR U332 ( .A(n299), .B(n300), .Z(swire[25]) );
  XOR U333 ( .A(sreg[89]), .B(n301), .Z(n300) );
  XOR U334 ( .A(n301), .B(n302), .Z(n299) );
  XOR U335 ( .A(n303), .B(n304), .Z(n302) );
  NAND U336 ( .A(b[0]), .B(a[25]), .Z(n304) );
  AND U337 ( .A(b[1]), .B(a[24]), .Z(n303) );
  IV U338 ( .A(n298), .Z(n301) );
  XOR U339 ( .A(n305), .B(n306), .Z(n298) );
  ANDN U340 ( .B(n307), .A(n308), .Z(n305) );
  XNOR U341 ( .A(n307), .B(n308), .Z(swire[24]) );
  XOR U342 ( .A(sreg[88]), .B(n309), .Z(n308) );
  XOR U343 ( .A(n309), .B(n310), .Z(n307) );
  XOR U344 ( .A(n311), .B(n312), .Z(n310) );
  NAND U345 ( .A(b[0]), .B(a[24]), .Z(n312) );
  AND U346 ( .A(b[1]), .B(a[23]), .Z(n311) );
  IV U347 ( .A(n306), .Z(n309) );
  XOR U348 ( .A(n313), .B(n314), .Z(n306) );
  ANDN U349 ( .B(n315), .A(n316), .Z(n313) );
  XNOR U350 ( .A(n315), .B(n316), .Z(swire[23]) );
  XOR U351 ( .A(sreg[87]), .B(n317), .Z(n316) );
  XOR U352 ( .A(n317), .B(n318), .Z(n315) );
  XOR U353 ( .A(n319), .B(n320), .Z(n318) );
  NAND U354 ( .A(b[0]), .B(a[23]), .Z(n320) );
  AND U355 ( .A(b[1]), .B(a[22]), .Z(n319) );
  IV U356 ( .A(n314), .Z(n317) );
  XOR U357 ( .A(n321), .B(n322), .Z(n314) );
  ANDN U358 ( .B(n323), .A(n324), .Z(n321) );
  XNOR U359 ( .A(n323), .B(n324), .Z(swire[22]) );
  XOR U360 ( .A(sreg[86]), .B(n325), .Z(n324) );
  XOR U361 ( .A(n325), .B(n326), .Z(n323) );
  XOR U362 ( .A(n327), .B(n328), .Z(n326) );
  NAND U363 ( .A(b[0]), .B(a[22]), .Z(n328) );
  AND U364 ( .A(b[1]), .B(a[21]), .Z(n327) );
  IV U365 ( .A(n322), .Z(n325) );
  XOR U366 ( .A(n329), .B(n330), .Z(n322) );
  ANDN U367 ( .B(n331), .A(n332), .Z(n329) );
  XNOR U368 ( .A(n331), .B(n332), .Z(swire[21]) );
  XOR U369 ( .A(sreg[85]), .B(n333), .Z(n332) );
  XOR U370 ( .A(n333), .B(n334), .Z(n331) );
  XOR U371 ( .A(n335), .B(n336), .Z(n334) );
  NAND U372 ( .A(b[0]), .B(a[21]), .Z(n336) );
  AND U373 ( .A(b[1]), .B(a[20]), .Z(n335) );
  IV U374 ( .A(n330), .Z(n333) );
  XOR U375 ( .A(n337), .B(n338), .Z(n330) );
  ANDN U376 ( .B(n339), .A(n340), .Z(n337) );
  XNOR U377 ( .A(n339), .B(n340), .Z(swire[20]) );
  XOR U378 ( .A(sreg[84]), .B(n341), .Z(n340) );
  XOR U379 ( .A(n341), .B(n342), .Z(n339) );
  XOR U380 ( .A(n343), .B(n344), .Z(n342) );
  NAND U381 ( .A(b[0]), .B(a[20]), .Z(n344) );
  AND U382 ( .A(b[1]), .B(a[19]), .Z(n343) );
  IV U383 ( .A(n338), .Z(n341) );
  XOR U384 ( .A(n345), .B(n346), .Z(n338) );
  ANDN U385 ( .B(n347), .A(n348), .Z(n345) );
  XNOR U386 ( .A(n347), .B(n348), .Z(swire[19]) );
  XOR U387 ( .A(sreg[83]), .B(n349), .Z(n348) );
  XOR U388 ( .A(n349), .B(n350), .Z(n347) );
  XOR U389 ( .A(n351), .B(n352), .Z(n350) );
  NAND U390 ( .A(b[0]), .B(a[19]), .Z(n352) );
  AND U391 ( .A(b[1]), .B(a[18]), .Z(n351) );
  IV U392 ( .A(n346), .Z(n349) );
  XOR U393 ( .A(n353), .B(n354), .Z(n346) );
  ANDN U394 ( .B(n355), .A(n356), .Z(n353) );
  XNOR U395 ( .A(n355), .B(n356), .Z(swire[18]) );
  XOR U396 ( .A(sreg[82]), .B(n357), .Z(n356) );
  XOR U397 ( .A(n357), .B(n358), .Z(n355) );
  XOR U398 ( .A(n359), .B(n360), .Z(n358) );
  NAND U399 ( .A(b[0]), .B(a[18]), .Z(n360) );
  AND U400 ( .A(b[1]), .B(a[17]), .Z(n359) );
  IV U401 ( .A(n354), .Z(n357) );
  XOR U402 ( .A(n361), .B(n362), .Z(n354) );
  ANDN U403 ( .B(n363), .A(n364), .Z(n361) );
  XNOR U404 ( .A(n363), .B(n364), .Z(swire[17]) );
  XOR U405 ( .A(sreg[81]), .B(n365), .Z(n364) );
  XOR U406 ( .A(n365), .B(n366), .Z(n363) );
  XOR U407 ( .A(n367), .B(n368), .Z(n366) );
  NAND U408 ( .A(b[0]), .B(a[17]), .Z(n368) );
  AND U409 ( .A(b[1]), .B(a[16]), .Z(n367) );
  IV U410 ( .A(n362), .Z(n365) );
  XOR U411 ( .A(n369), .B(n370), .Z(n362) );
  ANDN U412 ( .B(n371), .A(n372), .Z(n369) );
  XNOR U413 ( .A(n371), .B(n372), .Z(swire[16]) );
  XOR U414 ( .A(sreg[80]), .B(n373), .Z(n372) );
  XOR U415 ( .A(n373), .B(n374), .Z(n371) );
  XOR U416 ( .A(n375), .B(n376), .Z(n374) );
  NAND U417 ( .A(b[0]), .B(a[16]), .Z(n376) );
  AND U418 ( .A(b[1]), .B(a[15]), .Z(n375) );
  IV U419 ( .A(n370), .Z(n373) );
  XOR U420 ( .A(n377), .B(n378), .Z(n370) );
  ANDN U421 ( .B(n379), .A(n380), .Z(n377) );
  XNOR U422 ( .A(n379), .B(n380), .Z(swire[15]) );
  XOR U423 ( .A(sreg[79]), .B(n381), .Z(n380) );
  XOR U424 ( .A(n381), .B(n382), .Z(n379) );
  XOR U425 ( .A(n383), .B(n384), .Z(n382) );
  NAND U426 ( .A(b[0]), .B(a[15]), .Z(n384) );
  AND U427 ( .A(b[1]), .B(a[14]), .Z(n383) );
  IV U428 ( .A(n378), .Z(n381) );
  XOR U429 ( .A(n385), .B(n386), .Z(n378) );
  ANDN U430 ( .B(n387), .A(n388), .Z(n385) );
  XNOR U431 ( .A(n387), .B(n388), .Z(swire[14]) );
  XOR U432 ( .A(sreg[78]), .B(n389), .Z(n388) );
  XOR U433 ( .A(n389), .B(n390), .Z(n387) );
  XOR U434 ( .A(n391), .B(n392), .Z(n390) );
  NAND U435 ( .A(b[0]), .B(a[14]), .Z(n392) );
  AND U436 ( .A(b[1]), .B(a[13]), .Z(n391) );
  IV U437 ( .A(n386), .Z(n389) );
  XOR U438 ( .A(n393), .B(n394), .Z(n386) );
  ANDN U439 ( .B(n395), .A(n396), .Z(n393) );
  XNOR U440 ( .A(n395), .B(n396), .Z(swire[13]) );
  XOR U441 ( .A(sreg[77]), .B(n397), .Z(n396) );
  XOR U442 ( .A(n397), .B(n398), .Z(n395) );
  XOR U443 ( .A(n399), .B(n400), .Z(n398) );
  NAND U444 ( .A(b[0]), .B(a[13]), .Z(n400) );
  AND U445 ( .A(b[1]), .B(a[12]), .Z(n399) );
  IV U446 ( .A(n394), .Z(n397) );
  XOR U447 ( .A(n401), .B(n402), .Z(n394) );
  ANDN U448 ( .B(n403), .A(n404), .Z(n401) );
  XNOR U449 ( .A(n403), .B(n404), .Z(swire[12]) );
  XOR U450 ( .A(sreg[76]), .B(n405), .Z(n404) );
  XOR U451 ( .A(n405), .B(n406), .Z(n403) );
  XOR U452 ( .A(n407), .B(n408), .Z(n406) );
  NAND U453 ( .A(b[0]), .B(a[12]), .Z(n408) );
  AND U454 ( .A(b[1]), .B(a[11]), .Z(n407) );
  IV U455 ( .A(n402), .Z(n405) );
  XOR U456 ( .A(n409), .B(n410), .Z(n402) );
  ANDN U457 ( .B(n411), .A(n412), .Z(n409) );
  XNOR U458 ( .A(n411), .B(n412), .Z(swire[11]) );
  XOR U459 ( .A(sreg[75]), .B(n413), .Z(n412) );
  XOR U460 ( .A(n413), .B(n414), .Z(n411) );
  XOR U461 ( .A(n415), .B(n416), .Z(n414) );
  NAND U462 ( .A(b[0]), .B(a[11]), .Z(n416) );
  AND U463 ( .A(b[1]), .B(a[10]), .Z(n415) );
  IV U464 ( .A(n410), .Z(n413) );
  XOR U465 ( .A(n417), .B(n418), .Z(n410) );
  ANDN U466 ( .B(n419), .A(n420), .Z(n417) );
  XNOR U467 ( .A(n419), .B(n420), .Z(swire[10]) );
  XOR U468 ( .A(sreg[74]), .B(n421), .Z(n420) );
  XOR U469 ( .A(n421), .B(n422), .Z(n419) );
  XOR U470 ( .A(n423), .B(n424), .Z(n422) );
  NAND U471 ( .A(b[0]), .B(a[10]), .Z(n424) );
  AND U472 ( .A(a[9]), .B(b[1]), .Z(n423) );
  IV U473 ( .A(n418), .Z(n421) );
  XOR U474 ( .A(n425), .B(n426), .Z(n418) );
  ANDN U475 ( .B(n2), .A(n1), .Z(n425) );
  XOR U476 ( .A(sreg[73]), .B(n427), .Z(n1) );
  XOR U477 ( .A(n427), .B(n428), .Z(n2) );
  XOR U478 ( .A(n429), .B(n430), .Z(n428) );
  NAND U479 ( .A(b[1]), .B(a[8]), .Z(n430) );
  AND U480 ( .A(b[0]), .B(a[9]), .Z(n429) );
  IV U481 ( .A(n426), .Z(n427) );
  XOR U482 ( .A(n431), .B(n432), .Z(n426) );
  ANDN U483 ( .B(n3), .A(n4), .Z(n431) );
  XOR U484 ( .A(sreg[72]), .B(n433), .Z(n4) );
  XOR U485 ( .A(n433), .B(n434), .Z(n3) );
  XOR U486 ( .A(n435), .B(n436), .Z(n434) );
  NAND U487 ( .A(a[7]), .B(b[1]), .Z(n436) );
  AND U488 ( .A(a[8]), .B(b[0]), .Z(n435) );
  IV U489 ( .A(n432), .Z(n433) );
  XOR U490 ( .A(n437), .B(n438), .Z(n432) );
  ANDN U491 ( .B(n5), .A(n6), .Z(n437) );
  XOR U492 ( .A(sreg[71]), .B(n439), .Z(n6) );
  XOR U493 ( .A(n439), .B(n440), .Z(n5) );
  XOR U494 ( .A(n441), .B(n442), .Z(n440) );
  NAND U495 ( .A(b[1]), .B(a[6]), .Z(n442) );
  AND U496 ( .A(a[7]), .B(b[0]), .Z(n441) );
  IV U497 ( .A(n438), .Z(n439) );
  XOR U498 ( .A(n443), .B(n444), .Z(n438) );
  ANDN U499 ( .B(n7), .A(n8), .Z(n443) );
  XOR U500 ( .A(sreg[70]), .B(n445), .Z(n8) );
  XOR U501 ( .A(n445), .B(n446), .Z(n7) );
  XOR U502 ( .A(n447), .B(n448), .Z(n446) );
  NAND U503 ( .A(b[1]), .B(a[5]), .Z(n448) );
  AND U504 ( .A(b[0]), .B(a[6]), .Z(n447) );
  IV U505 ( .A(n444), .Z(n445) );
  XOR U506 ( .A(n449), .B(n450), .Z(n444) );
  ANDN U507 ( .B(n19), .A(n20), .Z(n449) );
  XOR U508 ( .A(sreg[69]), .B(n451), .Z(n20) );
  XOR U509 ( .A(n451), .B(n452), .Z(n19) );
  XOR U510 ( .A(n453), .B(n454), .Z(n452) );
  NAND U511 ( .A(b[1]), .B(a[4]), .Z(n454) );
  AND U512 ( .A(b[0]), .B(a[5]), .Z(n453) );
  IV U513 ( .A(n450), .Z(n451) );
  XOR U514 ( .A(n455), .B(n456), .Z(n450) );
  ANDN U515 ( .B(n103), .A(n104), .Z(n455) );
  XOR U516 ( .A(sreg[68]), .B(n457), .Z(n104) );
  XOR U517 ( .A(n457), .B(n458), .Z(n103) );
  XOR U518 ( .A(n459), .B(n460), .Z(n458) );
  NAND U519 ( .A(b[1]), .B(a[3]), .Z(n460) );
  AND U520 ( .A(b[0]), .B(a[4]), .Z(n459) );
  IV U521 ( .A(n456), .Z(n457) );
  XOR U522 ( .A(n461), .B(n462), .Z(n456) );
  ANDN U523 ( .B(n185), .A(n186), .Z(n461) );
  XOR U524 ( .A(sreg[67]), .B(n463), .Z(n186) );
  XOR U525 ( .A(n463), .B(n464), .Z(n185) );
  XOR U526 ( .A(n465), .B(n466), .Z(n464) );
  NAND U527 ( .A(b[1]), .B(a[2]), .Z(n466) );
  AND U528 ( .A(b[0]), .B(a[3]), .Z(n465) );
  IV U529 ( .A(n462), .Z(n463) );
  XNOR U530 ( .A(n467), .B(n468), .Z(n462) );
  ANDN U531 ( .B(n267), .A(n268), .Z(n467) );
  XOR U532 ( .A(sreg[66]), .B(n468), .Z(n268) );
  XOR U533 ( .A(n468), .B(n469), .Z(n267) );
  XOR U534 ( .A(n470), .B(n471), .Z(n469) );
  NAND U535 ( .A(b[1]), .B(a[1]), .Z(n471) );
  AND U536 ( .A(b[0]), .B(a[2]), .Z(n470) );
  XOR U537 ( .A(n472), .B(n473), .Z(n468) );
  NAND U538 ( .A(n474), .B(n475), .Z(n473) );
  XOR U539 ( .A(n474), .B(n475), .Z(c[63]) );
  XOR U540 ( .A(sreg[65]), .B(n472), .Z(n475) );
  XNOR U541 ( .A(n472), .B(n476), .Z(n474) );
  XOR U542 ( .A(n477), .B(n478), .Z(n476) );
  NAND U543 ( .A(b[0]), .B(a[1]), .Z(n478) );
  AND U544 ( .A(b[1]), .B(a[0]), .Z(n477) );
  ANDN U545 ( .B(sreg[64]), .A(n479), .Z(n472) );
  XNOR U546 ( .A(sreg[64]), .B(n479), .Z(c[62]) );
  NAND U547 ( .A(a[0]), .B(b[0]), .Z(n479) );
endmodule

