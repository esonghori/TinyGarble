
module Control ( opcode, rs_index, rt_index, rd_index, imm_out, alu_func, 
        shift_func, mult_func, branch_func, a_source_out, b_source_out, 
        c_source_out, pc_source_out, mem_source_out );
  input [31:0] opcode;
  output [4:0] rs_index;
  output [4:0] rt_index;
  output [4:0] rd_index;
  output [15:0] imm_out;
  output [3:0] alu_func;
  output [1:0] shift_func;
  output [3:0] mult_func;
  output [2:0] branch_func;
  output [1:0] a_source_out;
  output [1:0] b_source_out;
  output [2:0] c_source_out;
  output [1:0] pc_source_out;
  output [3:0] mem_source_out;
  wire   n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949;
  assign a_source_out[1] = 1'b0;
  assign imm_out[15] = opcode[15];
  assign imm_out[14] = opcode[14];
  assign imm_out[13] = opcode[13];
  assign imm_out[12] = opcode[12];
  assign imm_out[11] = opcode[11];
  assign imm_out[10] = opcode[10];
  assign imm_out[9] = opcode[9];
  assign imm_out[8] = opcode[8];
  assign imm_out[7] = opcode[7];
  assign imm_out[6] = opcode[6];
  assign imm_out[5] = opcode[5];
  assign imm_out[4] = opcode[4];
  assign imm_out[3] = opcode[3];
  assign imm_out[2] = opcode[2];
  assign imm_out[1] = opcode[1];
  assign imm_out[0] = opcode[0];

  ANDN U545 ( .B(n503), .A(n504), .Z(shift_func[1]) );
  AND U546 ( .A(n503), .B(n505), .Z(shift_func[0]) );
  AND U547 ( .A(n506), .B(n507), .Z(n505) );
  NANDN U548 ( .A(n508), .B(n509), .Z(n507) );
  NAND U549 ( .A(imm_out[1]), .B(imm_out[0]), .Z(n509) );
  NAND U550 ( .A(n510), .B(n511), .Z(rt_index[4]) );
  NAND U551 ( .A(n512), .B(opcode[20]), .Z(n511) );
  AND U552 ( .A(n513), .B(n514), .Z(n510) );
  NAND U553 ( .A(n515), .B(n506), .Z(n514) );
  NAND U554 ( .A(n516), .B(n517), .Z(n515) );
  NAND U555 ( .A(n518), .B(n519), .Z(n517) );
  NAND U556 ( .A(n520), .B(n521), .Z(n519) );
  NAND U557 ( .A(imm_out[1]), .B(opcode[20]), .Z(n521) );
  NANDN U558 ( .A(n522), .B(opcode[20]), .Z(n520) );
  AND U559 ( .A(n523), .B(n524), .Z(n516) );
  NAND U560 ( .A(n525), .B(n526), .Z(n524) );
  NAND U561 ( .A(n527), .B(n528), .Z(n526) );
  NAND U562 ( .A(n529), .B(opcode[20]), .Z(n528) );
  NAND U563 ( .A(opcode[19]), .B(opcode[20]), .Z(n527) );
  NAND U564 ( .A(n530), .B(opcode[20]), .Z(n523) );
  NAND U565 ( .A(n531), .B(n532), .Z(n513) );
  NAND U566 ( .A(n533), .B(n534), .Z(n531) );
  NAND U567 ( .A(n535), .B(opcode[20]), .Z(n534) );
  NAND U568 ( .A(n536), .B(opcode[20]), .Z(n533) );
  NAND U569 ( .A(n537), .B(n538), .Z(rt_index[3]) );
  NAND U570 ( .A(opcode[19]), .B(n512), .Z(n538) );
  AND U571 ( .A(n539), .B(n540), .Z(n537) );
  NAND U572 ( .A(n541), .B(n506), .Z(n540) );
  NAND U573 ( .A(n542), .B(n543), .Z(n541) );
  NAND U574 ( .A(n518), .B(n544), .Z(n543) );
  NAND U575 ( .A(n545), .B(n546), .Z(n544) );
  NAND U576 ( .A(imm_out[1]), .B(opcode[19]), .Z(n546) );
  OR U577 ( .A(n522), .B(n547), .Z(n545) );
  AND U578 ( .A(n548), .B(n549), .Z(n542) );
  NAND U579 ( .A(opcode[19]), .B(n525), .Z(n549) );
  NAND U580 ( .A(opcode[19]), .B(n530), .Z(n548) );
  NAND U581 ( .A(n550), .B(n532), .Z(n539) );
  NAND U582 ( .A(n551), .B(n552), .Z(n550) );
  NAND U583 ( .A(opcode[19]), .B(n535), .Z(n552) );
  NAND U584 ( .A(opcode[19]), .B(n536), .Z(n551) );
  NAND U585 ( .A(n553), .B(n554), .Z(rt_index[2]) );
  NAND U586 ( .A(n512), .B(opcode[18]), .Z(n554) );
  AND U587 ( .A(n555), .B(n556), .Z(n553) );
  NAND U588 ( .A(n557), .B(n506), .Z(n556) );
  NAND U589 ( .A(n558), .B(n559), .Z(n557) );
  NAND U590 ( .A(n518), .B(n560), .Z(n559) );
  NAND U591 ( .A(n561), .B(n562), .Z(n560) );
  NAND U592 ( .A(imm_out[1]), .B(opcode[18]), .Z(n562) );
  NANDN U593 ( .A(n522), .B(opcode[18]), .Z(n561) );
  AND U594 ( .A(n563), .B(n564), .Z(n558) );
  NAND U595 ( .A(n525), .B(opcode[18]), .Z(n564) );
  NAND U596 ( .A(n530), .B(opcode[18]), .Z(n563) );
  NAND U597 ( .A(n565), .B(n532), .Z(n555) );
  NAND U598 ( .A(n566), .B(n567), .Z(n565) );
  NAND U599 ( .A(n535), .B(opcode[18]), .Z(n567) );
  NAND U600 ( .A(n536), .B(opcode[18]), .Z(n566) );
  NAND U601 ( .A(n568), .B(n569), .Z(rt_index[1]) );
  NAND U602 ( .A(n512), .B(opcode[17]), .Z(n569) );
  AND U603 ( .A(n570), .B(n571), .Z(n568) );
  NAND U604 ( .A(n572), .B(n506), .Z(n571) );
  NAND U605 ( .A(n573), .B(n574), .Z(n572) );
  NAND U606 ( .A(n518), .B(n575), .Z(n574) );
  NAND U607 ( .A(n576), .B(n577), .Z(n575) );
  NAND U608 ( .A(imm_out[1]), .B(opcode[17]), .Z(n577) );
  NANDN U609 ( .A(n522), .B(opcode[17]), .Z(n576) );
  AND U610 ( .A(n578), .B(n579), .Z(n573) );
  NAND U611 ( .A(n525), .B(opcode[17]), .Z(n579) );
  NAND U612 ( .A(n530), .B(opcode[17]), .Z(n578) );
  NAND U613 ( .A(n580), .B(n532), .Z(n570) );
  NAND U614 ( .A(n581), .B(n582), .Z(n580) );
  NAND U615 ( .A(n535), .B(opcode[17]), .Z(n582) );
  NAND U616 ( .A(n536), .B(opcode[17]), .Z(n581) );
  NAND U617 ( .A(n583), .B(n584), .Z(rt_index[0]) );
  NAND U618 ( .A(n512), .B(opcode[16]), .Z(n584) );
  AND U619 ( .A(n585), .B(n586), .Z(n583) );
  NAND U620 ( .A(n587), .B(n506), .Z(n586) );
  NAND U621 ( .A(n588), .B(n589), .Z(n587) );
  NAND U622 ( .A(n518), .B(n590), .Z(n589) );
  NAND U623 ( .A(n591), .B(n592), .Z(n590) );
  NAND U624 ( .A(imm_out[1]), .B(opcode[16]), .Z(n592) );
  NANDN U625 ( .A(n522), .B(opcode[16]), .Z(n591) );
  AND U626 ( .A(n593), .B(n594), .Z(n588) );
  NAND U627 ( .A(n525), .B(n595), .Z(n594) );
  NAND U628 ( .A(n596), .B(n597), .Z(n595) );
  NAND U629 ( .A(n529), .B(opcode[16]), .Z(n597) );
  IV U630 ( .A(n598), .Z(n529) );
  NAND U631 ( .A(opcode[19]), .B(opcode[16]), .Z(n596) );
  NAND U632 ( .A(opcode[16]), .B(n530), .Z(n593) );
  NANDN U633 ( .A(n599), .B(n600), .Z(n530) );
  IV U634 ( .A(n601), .Z(n599) );
  NAND U635 ( .A(n602), .B(n532), .Z(n585) );
  NAND U636 ( .A(n603), .B(n604), .Z(n602) );
  NAND U637 ( .A(n535), .B(opcode[16]), .Z(n604) );
  NAND U638 ( .A(opcode[16]), .B(n536), .Z(n603) );
  NAND U639 ( .A(n605), .B(n606), .Z(rs_index[4]) );
  ANDN U640 ( .B(n607), .A(opcode[25]), .Z(n605) );
  NAND U641 ( .A(n608), .B(n609), .Z(n607) );
  MUX U642 ( .IN0(opcode[20]), .IN1(imm_out[15]), .SEL(n610), .F(n609) );
  NAND U643 ( .A(n611), .B(n612), .Z(rs_index[3]) );
  NAND U644 ( .A(n608), .B(n613), .Z(n612) );
  MUX U645 ( .IN0(opcode[19]), .IN1(imm_out[14]), .SEL(n610), .F(n613) );
  ANDN U646 ( .B(n606), .A(opcode[24]), .Z(n611) );
  NAND U647 ( .A(n614), .B(n615), .Z(rs_index[2]) );
  NAND U648 ( .A(n616), .B(n506), .Z(n615) );
  NAND U649 ( .A(n610), .B(n617), .Z(n616) );
  NAND U650 ( .A(n618), .B(n619), .Z(n617) );
  AND U651 ( .A(n620), .B(n518), .Z(n618) );
  AND U652 ( .A(n621), .B(n622), .Z(n614) );
  NAND U653 ( .A(n623), .B(n532), .Z(n622) );
  NAND U654 ( .A(n624), .B(n625), .Z(n623) );
  NAND U655 ( .A(n518), .B(n626), .Z(n625) );
  NAND U656 ( .A(n627), .B(n628), .Z(n626) );
  NAND U657 ( .A(n629), .B(n630), .Z(n628) );
  MUX U658 ( .IN0(opcode[18]), .IN1(imm_out[13]), .SEL(n610), .F(n629) );
  NAND U659 ( .A(opcode[23]), .B(n535), .Z(n627) );
  NANDN U660 ( .A(n631), .B(n632), .Z(n535) );
  NAND U661 ( .A(opcode[23]), .B(n536), .Z(n624) );
  NAND U662 ( .A(n633), .B(n634), .Z(n536) );
  AND U663 ( .A(n635), .B(n636), .Z(n634) );
  NAND U664 ( .A(opcode[23]), .B(n512), .Z(n621) );
  NAND U665 ( .A(n637), .B(n638), .Z(n512) );
  AND U666 ( .A(n639), .B(n640), .Z(n637) );
  IV U667 ( .A(opcode[29]), .Z(n639) );
  NAND U668 ( .A(n641), .B(n642), .Z(rs_index[1]) );
  NAND U669 ( .A(n608), .B(n643), .Z(n642) );
  MUX U670 ( .IN0(opcode[17]), .IN1(imm_out[12]), .SEL(n610), .F(n643) );
  ANDN U671 ( .B(n606), .A(opcode[22]), .Z(n641) );
  NAND U672 ( .A(n644), .B(n645), .Z(rs_index[0]) );
  NAND U673 ( .A(n608), .B(n646), .Z(n645) );
  MUX U674 ( .IN0(opcode[16]), .IN1(imm_out[11]), .SEL(n610), .F(n646) );
  ANDN U675 ( .B(n606), .A(opcode[21]), .Z(n644) );
  NAND U676 ( .A(n647), .B(n648), .Z(n606) );
  AND U677 ( .A(n620), .B(n619), .Z(n647) );
  NAND U678 ( .A(n649), .B(n650), .Z(rd_index[4]) );
  AND U679 ( .A(n651), .B(n652), .Z(n650) );
  NAND U680 ( .A(opcode[20]), .B(n653), .Z(n652) );
  NAND U681 ( .A(n654), .B(n506), .Z(n651) );
  NAND U682 ( .A(n655), .B(n656), .Z(n654) );
  AND U683 ( .A(n657), .B(n658), .Z(n655) );
  NAND U684 ( .A(n518), .B(n659), .Z(n658) );
  NAND U685 ( .A(n660), .B(n661), .Z(n659) );
  AND U686 ( .A(n662), .B(n663), .Z(n661) );
  NAND U687 ( .A(n664), .B(n665), .Z(n663) );
  AND U688 ( .A(n666), .B(imm_out[15]), .Z(n664) );
  AND U689 ( .A(n667), .B(n668), .Z(n662) );
  NAND U690 ( .A(n669), .B(imm_out[15]), .Z(n668) );
  NANDN U691 ( .A(n670), .B(imm_out[15]), .Z(n667) );
  AND U692 ( .A(n671), .B(n672), .Z(n660) );
  NANDN U693 ( .A(n673), .B(n674), .Z(n672) );
  AND U694 ( .A(n675), .B(imm_out[15]), .Z(n674) );
  NANDN U695 ( .A(n676), .B(n677), .Z(n671) );
  AND U696 ( .A(n619), .B(imm_out[15]), .Z(n677) );
  AND U697 ( .A(n678), .B(n679), .Z(n649) );
  NAND U698 ( .A(n608), .B(n680), .Z(n679) );
  MUX U699 ( .IN0(imm_out[15]), .IN1(opcode[20]), .SEL(n610), .F(n680) );
  NAND U700 ( .A(n681), .B(n682), .Z(n678) );
  AND U701 ( .A(n683), .B(opcode[20]), .Z(n682) );
  NAND U702 ( .A(n684), .B(n685), .Z(rd_index[3]) );
  AND U703 ( .A(n686), .B(n687), .Z(n685) );
  NAND U704 ( .A(opcode[19]), .B(n653), .Z(n687) );
  NAND U705 ( .A(n688), .B(n506), .Z(n686) );
  NAND U706 ( .A(n689), .B(n690), .Z(n688) );
  NAND U707 ( .A(n518), .B(n691), .Z(n690) );
  NAND U708 ( .A(n692), .B(n693), .Z(n691) );
  AND U709 ( .A(n694), .B(n695), .Z(n693) );
  NAND U710 ( .A(n696), .B(imm_out[14]), .Z(n695) );
  AND U711 ( .A(n697), .B(n698), .Z(n694) );
  NAND U712 ( .A(n669), .B(imm_out[14]), .Z(n698) );
  NANDN U713 ( .A(n670), .B(imm_out[14]), .Z(n697) );
  AND U714 ( .A(n699), .B(n700), .Z(n692) );
  NAND U715 ( .A(n701), .B(imm_out[14]), .Z(n700) );
  NAND U716 ( .A(n702), .B(n619), .Z(n699) );
  NANDN U717 ( .A(n620), .B(n703), .Z(n702) );
  NANDN U718 ( .A(n676), .B(imm_out[14]), .Z(n703) );
  AND U719 ( .A(n704), .B(n705), .Z(n684) );
  NAND U720 ( .A(n608), .B(n706), .Z(n705) );
  MUX U721 ( .IN0(imm_out[14]), .IN1(opcode[19]), .SEL(n610), .F(n706) );
  NAND U722 ( .A(n681), .B(n707), .Z(n704) );
  AND U723 ( .A(n683), .B(opcode[19]), .Z(n707) );
  NAND U724 ( .A(n708), .B(n709), .Z(rd_index[2]) );
  AND U725 ( .A(n710), .B(n711), .Z(n709) );
  NAND U726 ( .A(opcode[18]), .B(n653), .Z(n711) );
  NAND U727 ( .A(n712), .B(n506), .Z(n710) );
  NAND U728 ( .A(n689), .B(n713), .Z(n712) );
  NAND U729 ( .A(n518), .B(n714), .Z(n713) );
  NAND U730 ( .A(n715), .B(n716), .Z(n714) );
  AND U731 ( .A(n717), .B(n718), .Z(n716) );
  NAND U732 ( .A(n696), .B(imm_out[13]), .Z(n718) );
  AND U733 ( .A(n719), .B(n720), .Z(n717) );
  NAND U734 ( .A(n669), .B(imm_out[13]), .Z(n720) );
  NANDN U735 ( .A(n670), .B(imm_out[13]), .Z(n719) );
  AND U736 ( .A(n721), .B(n722), .Z(n715) );
  NAND U737 ( .A(n701), .B(imm_out[13]), .Z(n722) );
  NAND U738 ( .A(n723), .B(n619), .Z(n721) );
  NANDN U739 ( .A(n620), .B(n724), .Z(n723) );
  NANDN U740 ( .A(n676), .B(imm_out[13]), .Z(n724) );
  AND U741 ( .A(n725), .B(n726), .Z(n708) );
  NAND U742 ( .A(n608), .B(n727), .Z(n726) );
  MUX U743 ( .IN0(imm_out[13]), .IN1(opcode[18]), .SEL(n610), .F(n727) );
  NAND U744 ( .A(n681), .B(n728), .Z(n725) );
  AND U745 ( .A(n683), .B(opcode[18]), .Z(n728) );
  NAND U746 ( .A(n729), .B(n730), .Z(rd_index[1]) );
  AND U747 ( .A(n731), .B(n732), .Z(n730) );
  NAND U748 ( .A(opcode[17]), .B(n653), .Z(n732) );
  NAND U749 ( .A(n733), .B(n506), .Z(n731) );
  NAND U750 ( .A(n689), .B(n734), .Z(n733) );
  NAND U751 ( .A(n518), .B(n735), .Z(n734) );
  NAND U752 ( .A(n736), .B(n737), .Z(n735) );
  AND U753 ( .A(n738), .B(n739), .Z(n737) );
  NAND U754 ( .A(n696), .B(imm_out[12]), .Z(n739) );
  AND U755 ( .A(n740), .B(n741), .Z(n738) );
  NAND U756 ( .A(n669), .B(imm_out[12]), .Z(n741) );
  NANDN U757 ( .A(n670), .B(imm_out[12]), .Z(n740) );
  AND U758 ( .A(n742), .B(n743), .Z(n736) );
  NAND U759 ( .A(n701), .B(imm_out[12]), .Z(n743) );
  NAND U760 ( .A(n744), .B(n619), .Z(n742) );
  NANDN U761 ( .A(n620), .B(n745), .Z(n744) );
  NANDN U762 ( .A(n676), .B(imm_out[12]), .Z(n745) );
  AND U763 ( .A(n746), .B(n747), .Z(n729) );
  NAND U764 ( .A(n608), .B(n748), .Z(n747) );
  MUX U765 ( .IN0(imm_out[12]), .IN1(opcode[17]), .SEL(n610), .F(n748) );
  NAND U766 ( .A(n681), .B(n749), .Z(n746) );
  AND U767 ( .A(n683), .B(opcode[17]), .Z(n749) );
  NAND U768 ( .A(n750), .B(n751), .Z(rd_index[0]) );
  AND U769 ( .A(n752), .B(n753), .Z(n751) );
  NAND U770 ( .A(opcode[16]), .B(n653), .Z(n753) );
  NAND U771 ( .A(n754), .B(n506), .Z(n752) );
  NAND U772 ( .A(n689), .B(n755), .Z(n754) );
  NAND U773 ( .A(n518), .B(n756), .Z(n755) );
  NAND U774 ( .A(n757), .B(n758), .Z(n756) );
  AND U775 ( .A(n759), .B(n760), .Z(n758) );
  NAND U776 ( .A(n696), .B(imm_out[11]), .Z(n760) );
  AND U777 ( .A(n665), .B(n666), .Z(n696) );
  OR U778 ( .A(n761), .B(n762), .Z(n666) );
  AND U779 ( .A(n763), .B(n764), .Z(n759) );
  NAND U780 ( .A(n669), .B(imm_out[11]), .Z(n764) );
  NANDN U781 ( .A(n670), .B(imm_out[11]), .Z(n763) );
  NAND U782 ( .A(n765), .B(n766), .Z(n670) );
  NANDN U783 ( .A(n508), .B(n767), .Z(n765) );
  ANDN U784 ( .B(n767), .A(imm_out[0]), .Z(n508) );
  AND U785 ( .A(n768), .B(n769), .Z(n757) );
  NAND U786 ( .A(n701), .B(imm_out[11]), .Z(n769) );
  ANDN U787 ( .B(n675), .A(n673), .Z(n701) );
  NAND U788 ( .A(n770), .B(imm_out[11]), .Z(n768) );
  ANDN U789 ( .B(n619), .A(n676), .Z(n770) );
  AND U790 ( .A(n771), .B(n772), .Z(n750) );
  NAND U791 ( .A(n608), .B(n773), .Z(n772) );
  MUX U792 ( .IN0(imm_out[11]), .IN1(opcode[16]), .SEL(n610), .F(n773) );
  IV U793 ( .A(opcode[23]), .Z(n610) );
  ANDN U794 ( .B(n518), .A(n774), .Z(n608) );
  NAND U795 ( .A(n532), .B(n630), .Z(n774) );
  ANDN U796 ( .B(n632), .A(n631), .Z(n630) );
  NAND U797 ( .A(n681), .B(n775), .Z(n771) );
  AND U798 ( .A(n683), .B(opcode[16]), .Z(n775) );
  AND U799 ( .A(n506), .B(n776), .Z(pc_source_out[1]) );
  NAND U800 ( .A(n777), .B(n778), .Z(n776) );
  ANDN U801 ( .B(n779), .A(n780), .Z(n777) );
  AND U802 ( .A(n506), .B(n781), .Z(pc_source_out[0]) );
  NANDN U803 ( .A(n780), .B(n601), .Z(n781) );
  NOR U804 ( .A(n782), .B(n783), .Z(n780) );
  AND U805 ( .A(n784), .B(n785), .Z(mult_func[3]) );
  AND U806 ( .A(n648), .B(imm_out[1]), .Z(n785) );
  AND U807 ( .A(n506), .B(n518), .Z(n648) );
  ANDN U808 ( .B(n786), .A(n787), .Z(n784) );
  AND U809 ( .A(n506), .B(n788), .Z(mult_func[2]) );
  AND U810 ( .A(n789), .B(n518), .Z(n788) );
  NAND U811 ( .A(n790), .B(n791), .Z(n789) );
  NAND U812 ( .A(n792), .B(n665), .Z(n791) );
  ANDN U813 ( .B(imm_out[0]), .A(n793), .Z(n792) );
  NAND U814 ( .A(n794), .B(n786), .Z(n790) );
  NANDN U815 ( .A(n795), .B(n796), .Z(n794) );
  AND U816 ( .A(n506), .B(n797), .Z(mult_func[1]) );
  AND U817 ( .A(n798), .B(n518), .Z(n797) );
  NAND U818 ( .A(n799), .B(n800), .Z(n798) );
  NAND U819 ( .A(n801), .B(n665), .Z(n800) );
  NANDN U820 ( .A(n761), .B(n802), .Z(n801) );
  IV U821 ( .A(n803), .Z(n802) );
  ANDN U822 ( .B(n804), .A(n793), .Z(n761) );
  NAND U823 ( .A(n805), .B(n786), .Z(n799) );
  NAND U824 ( .A(n806), .B(n796), .Z(n805) );
  NANDN U825 ( .A(n807), .B(imm_out[0]), .Z(n806) );
  AND U826 ( .A(n506), .B(n808), .Z(mult_func[0]) );
  AND U827 ( .A(n809), .B(n518), .Z(n808) );
  NAND U828 ( .A(n810), .B(n811), .Z(n809) );
  NAND U829 ( .A(n675), .B(n665), .Z(n811) );
  AND U830 ( .A(n812), .B(imm_out[4]), .Z(n665) );
  ANDN U831 ( .B(n813), .A(imm_out[5]), .Z(n812) );
  IV U832 ( .A(imm_out[3]), .Z(n813) );
  OR U833 ( .A(n762), .B(n803), .Z(n675) );
  NAND U834 ( .A(n786), .B(n795), .Z(n810) );
  AND U835 ( .A(n814), .B(imm_out[0]), .Z(n795) );
  AND U836 ( .A(n815), .B(imm_out[4]), .Z(n786) );
  ANDN U837 ( .B(imm_out[3]), .A(imm_out[5]), .Z(n815) );
  NAND U838 ( .A(n816), .B(n817), .Z(mem_source_out[3]) );
  NAND U839 ( .A(n681), .B(n818), .Z(n817) );
  NAND U840 ( .A(n819), .B(n600), .Z(n818) );
  NANDN U841 ( .A(n820), .B(n821), .Z(n816) );
  NAND U842 ( .A(n822), .B(n823), .Z(mem_source_out[2]) );
  NAND U843 ( .A(n824), .B(n821), .Z(n823) );
  NAND U844 ( .A(n657), .B(n825), .Z(n824) );
  NAND U845 ( .A(n681), .B(n826), .Z(n822) );
  NAND U846 ( .A(n827), .B(n828), .Z(n826) );
  AND U847 ( .A(n657), .B(n829), .Z(n828) );
  ANDN U848 ( .B(n825), .A(n830), .Z(n827) );
  ANDN U849 ( .B(n681), .A(n820), .Z(mem_source_out[1]) );
  ANDN U850 ( .B(n636), .A(n518), .Z(n820) );
  NAND U851 ( .A(n831), .B(n832), .Z(c_source_out[2]) );
  NAND U852 ( .A(n833), .B(n506), .Z(n832) );
  NAND U853 ( .A(n689), .B(n834), .Z(n833) );
  NAND U854 ( .A(n835), .B(n619), .Z(n834) );
  AND U855 ( .A(n836), .B(n518), .Z(n835) );
  NANDN U856 ( .A(n620), .B(n676), .Z(n836) );
  AND U857 ( .A(n656), .B(n657), .Z(n689) );
  NANDN U858 ( .A(n837), .B(n838), .Z(n656) );
  AND U859 ( .A(n598), .B(n525), .Z(n838) );
  NAND U860 ( .A(n839), .B(n653), .Z(n831) );
  AND U861 ( .A(n683), .B(n681), .Z(c_source_out[1]) );
  NAND U862 ( .A(n840), .B(n841), .Z(c_source_out[0]) );
  AND U863 ( .A(n638), .B(n635), .Z(n841) );
  AND U864 ( .A(n842), .B(n843), .Z(n840) );
  NAND U865 ( .A(n844), .B(n506), .Z(n843) );
  NAND U866 ( .A(n845), .B(n846), .Z(n844) );
  AND U867 ( .A(n847), .B(n848), .Z(n846) );
  NAND U868 ( .A(n525), .B(n849), .Z(n848) );
  NANDN U869 ( .A(n837), .B(n598), .Z(n849) );
  NAND U870 ( .A(n547), .B(opcode[20]), .Z(n837) );
  AND U871 ( .A(n850), .B(n851), .Z(n845) );
  NAND U872 ( .A(n518), .B(n852), .Z(n851) );
  NAND U873 ( .A(n853), .B(n522), .Z(n852) );
  AND U874 ( .A(n796), .B(n767), .Z(n853) );
  NAND U875 ( .A(n854), .B(n855), .Z(branch_func[2]) );
  AND U876 ( .A(n856), .B(n857), .Z(n855) );
  AND U877 ( .A(n782), .B(n635), .Z(n856) );
  AND U878 ( .A(n858), .B(n859), .Z(n854) );
  AND U879 ( .A(n657), .B(n860), .Z(n859) );
  NAND U880 ( .A(n525), .B(n861), .Z(n860) );
  NAND U881 ( .A(n862), .B(n863), .Z(n861) );
  ANDN U882 ( .B(n547), .A(opcode[18]), .Z(n863) );
  NOR U883 ( .A(opcode[16]), .B(opcode[17]), .Z(n862) );
  NAND U884 ( .A(n864), .B(n865), .Z(branch_func[1]) );
  AND U885 ( .A(n825), .B(n866), .Z(n865) );
  AND U886 ( .A(n867), .B(n868), .Z(n866) );
  ANDN U887 ( .B(n782), .A(n869), .Z(n825) );
  ANDN U888 ( .B(n858), .A(n870), .Z(n864) );
  NAND U889 ( .A(n871), .B(n872), .Z(branch_func[0]) );
  ANDN U890 ( .B(n873), .A(n830), .Z(n872) );
  AND U891 ( .A(n867), .B(n635), .Z(n873) );
  AND U892 ( .A(n858), .B(n874), .Z(n871) );
  AND U893 ( .A(n868), .B(n875), .Z(n874) );
  NAND U894 ( .A(n518), .B(n876), .Z(n875) );
  NAND U895 ( .A(n767), .B(n522), .Z(n876) );
  AND U896 ( .A(n877), .B(imm_out[3]), .Z(n522) );
  ANDN U897 ( .B(n673), .A(imm_out[4]), .Z(n877) );
  NAND U898 ( .A(n525), .B(n878), .Z(n868) );
  NAND U899 ( .A(n547), .B(n598), .Z(n878) );
  AND U900 ( .A(n842), .B(n879), .Z(n858) );
  AND U901 ( .A(n638), .B(n640), .Z(n879) );
  IV U902 ( .A(n681), .Z(n640) );
  NAND U903 ( .A(opcode[30]), .B(opcode[31]), .Z(n638) );
  NOR U904 ( .A(opcode[29]), .B(n532), .Z(n842) );
  NAND U905 ( .A(n880), .B(n881), .Z(b_source_out[1]) );
  ANDN U906 ( .B(n882), .A(mem_source_out[0]), .Z(n880) );
  NAND U907 ( .A(n883), .B(n653), .Z(n882) );
  NAND U908 ( .A(n857), .B(n819), .Z(n883) );
  AND U909 ( .A(n653), .B(n884), .Z(b_source_out[0]) );
  NANDN U910 ( .A(n870), .B(n847), .Z(n884) );
  AND U911 ( .A(n885), .B(n886), .Z(alu_func[3]) );
  AND U912 ( .A(n887), .B(imm_out[0]), .Z(n886) );
  ANDN U913 ( .B(n518), .A(n504), .Z(n887) );
  NAND U914 ( .A(imm_out[1]), .B(n506), .Z(n504) );
  AND U915 ( .A(n669), .B(imm_out[2]), .Z(n885) );
  NAND U916 ( .A(n888), .B(n889), .Z(alu_func[2]) );
  NAND U917 ( .A(n890), .B(n506), .Z(n889) );
  NAND U918 ( .A(n891), .B(n778), .Z(n890) );
  AND U919 ( .A(n779), .B(n892), .Z(n891) );
  NAND U920 ( .A(n518), .B(n893), .Z(n892) );
  NAND U921 ( .A(n894), .B(n895), .Z(n893) );
  NANDN U922 ( .A(n673), .B(n762), .Z(n895) );
  ANDN U923 ( .B(imm_out[1]), .A(n787), .Z(n762) );
  AND U924 ( .A(n783), .B(n896), .Z(n894) );
  NAND U925 ( .A(n897), .B(n669), .Z(n896) );
  NANDN U926 ( .A(n620), .B(n898), .Z(n897) );
  ANDN U927 ( .B(n899), .A(n900), .Z(n888) );
  NAND U928 ( .A(n901), .B(n653), .Z(n899) );
  NAND U929 ( .A(n847), .B(n850), .Z(n901) );
  ANDN U930 ( .B(n829), .A(n869), .Z(n850) );
  NAND U931 ( .A(n902), .B(n903), .Z(alu_func[1]) );
  NAND U932 ( .A(n904), .B(n653), .Z(n903) );
  OR U933 ( .A(n870), .B(n830), .Z(n904) );
  NAND U934 ( .A(n829), .B(n657), .Z(n870) );
  NAND U935 ( .A(n905), .B(n506), .Z(n902) );
  NAND U936 ( .A(n906), .B(n600), .Z(n905) );
  NAND U937 ( .A(n518), .B(n907), .Z(n906) );
  NANDN U938 ( .A(n908), .B(n909), .Z(n907) );
  NAND U939 ( .A(n910), .B(n669), .Z(n909) );
  NAND U940 ( .A(n898), .B(n807), .Z(n910) );
  NANDN U941 ( .A(imm_out[0]), .B(imm_out[2]), .Z(n898) );
  NAND U942 ( .A(n911), .B(n912), .Z(alu_func[0]) );
  ANDN U943 ( .B(n913), .A(n900), .Z(n912) );
  AND U944 ( .A(n914), .B(n915), .Z(n900) );
  AND U945 ( .A(n632), .B(n518), .Z(n915) );
  NOR U946 ( .A(opcode[21]), .B(opcode[22]), .Z(n632) );
  ANDN U947 ( .B(n532), .A(n631), .Z(n914) );
  OR U948 ( .A(opcode[25]), .B(opcode[24]), .Z(n631) );
  AND U949 ( .A(n916), .B(opcode[30]), .Z(n532) );
  NOR U950 ( .A(opcode[29]), .B(opcode[31]), .Z(n916) );
  ANDN U951 ( .B(n881), .A(mem_source_out[0]), .Z(n913) );
  ANDN U952 ( .B(n821), .A(n917), .Z(mem_source_out[0]) );
  AND U953 ( .A(n819), .B(n601), .Z(n917) );
  AND U954 ( .A(n918), .B(opcode[29]), .Z(n821) );
  NAND U955 ( .A(n681), .B(n683), .Z(n881) );
  NAND U956 ( .A(n819), .B(n633), .Z(n683) );
  ANDN U957 ( .B(n601), .A(n919), .Z(n633) );
  NANDN U958 ( .A(n830), .B(n600), .Z(n919) );
  AND U959 ( .A(n867), .B(n829), .Z(n600) );
  AND U960 ( .A(n657), .B(n857), .Z(n601) );
  IV U961 ( .A(n869), .Z(n857) );
  NOR U962 ( .A(opcode[26]), .B(n920), .Z(n869) );
  ANDN U963 ( .B(n918), .A(opcode[29]), .Z(n681) );
  ANDN U964 ( .B(opcode[31]), .A(opcode[30]), .Z(n918) );
  AND U965 ( .A(n921), .B(n922), .Z(n911) );
  NAND U966 ( .A(n923), .B(n506), .Z(n922) );
  NAND U967 ( .A(n924), .B(n778), .Z(n923) );
  AND U968 ( .A(n925), .B(n847), .Z(n778) );
  AND U969 ( .A(n829), .B(n635), .Z(n925) );
  IV U970 ( .A(n839), .Z(n635) );
  AND U971 ( .A(n926), .B(opcode[27]), .Z(n839) );
  AND U972 ( .A(opcode[26]), .B(opcode[28]), .Z(n926) );
  OR U973 ( .A(opcode[26]), .B(n927), .Z(n829) );
  AND U974 ( .A(n779), .B(n928), .Z(n924) );
  NAND U975 ( .A(n518), .B(n929), .Z(n928) );
  NAND U976 ( .A(n930), .B(n931), .Z(n929) );
  NAND U977 ( .A(n932), .B(n669), .Z(n931) );
  AND U978 ( .A(n933), .B(imm_out[5]), .Z(n669) );
  NOR U979 ( .A(imm_out[3]), .B(imm_out[4]), .Z(n933) );
  NANDN U980 ( .A(n934), .B(n793), .Z(n932) );
  MUX U981 ( .IN0(n935), .IN1(n767), .SEL(imm_out[0]), .F(n934) );
  AND U982 ( .A(imm_out[1]), .B(imm_out[2]), .Z(n935) );
  ANDN U983 ( .B(n783), .A(n908), .Z(n930) );
  ANDN U984 ( .B(n803), .A(n673), .Z(n908) );
  NAND U985 ( .A(n936), .B(imm_out[5]), .Z(n673) );
  ANDN U986 ( .B(imm_out[3]), .A(imm_out[4]), .Z(n936) );
  ANDN U987 ( .B(imm_out[0]), .A(n807), .Z(n803) );
  NAND U988 ( .A(n937), .B(n619), .Z(n783) );
  AND U989 ( .A(n938), .B(imm_out[3]), .Z(n619) );
  NAND U990 ( .A(n939), .B(n796), .Z(n937) );
  OR U991 ( .A(n793), .B(imm_out[0]), .Z(n796) );
  ANDN U992 ( .B(n676), .A(n620), .Z(n939) );
  ANDN U993 ( .B(n767), .A(n814), .Z(n620) );
  NANDN U994 ( .A(n793), .B(imm_out[0]), .Z(n676) );
  NAND U995 ( .A(n767), .B(n814), .Z(n793) );
  IV U996 ( .A(imm_out[1]), .Z(n767) );
  IV U997 ( .A(n782), .Z(n518) );
  NAND U998 ( .A(n940), .B(n598), .Z(n779) );
  NOR U999 ( .A(opcode[17]), .B(opcode[18]), .Z(n598) );
  AND U1000 ( .A(n547), .B(n525), .Z(n940) );
  IV U1001 ( .A(opcode[19]), .Z(n547) );
  NAND U1002 ( .A(n941), .B(n653), .Z(n921) );
  AND U1003 ( .A(n942), .B(opcode[29]), .Z(n653) );
  NAND U1004 ( .A(n943), .B(n819), .Z(n941) );
  AND U1005 ( .A(n782), .B(n636), .Z(n819) );
  IV U1006 ( .A(n525), .Z(n636) );
  AND U1007 ( .A(n944), .B(opcode[26]), .Z(n525) );
  AND U1008 ( .A(n657), .B(n847), .Z(n943) );
  ANDN U1009 ( .B(n867), .A(n830), .Z(n847) );
  AND U1010 ( .A(n945), .B(opcode[27]), .Z(n830) );
  NOR U1011 ( .A(n946), .B(opcode[26]), .Z(n945) );
  NANDN U1012 ( .A(n927), .B(opcode[26]), .Z(n867) );
  NAND U1013 ( .A(opcode[28]), .B(n947), .Z(n927) );
  NANDN U1014 ( .A(n920), .B(opcode[26]), .Z(n657) );
  NAND U1015 ( .A(opcode[27]), .B(n946), .Z(n920) );
  AND U1016 ( .A(n503), .B(n948), .Z(a_source_out[0]) );
  AND U1017 ( .A(n506), .B(n949), .Z(n948) );
  NAND U1018 ( .A(n787), .B(n807), .Z(n949) );
  NAND U1019 ( .A(imm_out[1]), .B(n814), .Z(n807) );
  NAND U1020 ( .A(n804), .B(n814), .Z(n787) );
  IV U1021 ( .A(imm_out[2]), .Z(n814) );
  IV U1022 ( .A(imm_out[0]), .Z(n804) );
  ANDN U1023 ( .B(n942), .A(opcode[29]), .Z(n506) );
  NOR U1024 ( .A(opcode[31]), .B(opcode[30]), .Z(n942) );
  ANDN U1025 ( .B(n766), .A(n782), .Z(n503) );
  NANDN U1026 ( .A(opcode[26]), .B(n944), .Z(n782) );
  AND U1027 ( .A(n947), .B(n946), .Z(n944) );
  IV U1028 ( .A(opcode[28]), .Z(n946) );
  IV U1029 ( .A(opcode[27]), .Z(n947) );
  ANDN U1030 ( .B(n938), .A(imm_out[3]), .Z(n766) );
  NOR U1031 ( .A(imm_out[4]), .B(imm_out[5]), .Z(n938) );
endmodule

