
module modmult_step_N256_1 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N4, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871;
  assign N4 = y[0];

  XNOR U2 ( .A(n3962), .B(n3963), .Z(n1) );
  NAND U3 ( .A(n1), .B(n2322), .Z(n2) );
  NAND U4 ( .A(n2), .B(n3087), .Z(n3) );
  NAND U5 ( .A(n[97]), .B(n3958), .Z(n4) );
  XOR U6 ( .A(n3958), .B(n[97]), .Z(n5) );
  NAND U7 ( .A(n5), .B(n3), .Z(n6) );
  NAND U8 ( .A(n4), .B(n6), .Z(n7) );
  NAND U9 ( .A(n[98]), .B(n3954), .Z(n8) );
  XOR U10 ( .A(n3954), .B(n[98]), .Z(n9) );
  NAND U11 ( .A(n9), .B(n7), .Z(n10) );
  NAND U12 ( .A(n8), .B(n10), .Z(n11) );
  NANDN U13 ( .A(n5344), .B(n3950), .Z(n12) );
  XOR U14 ( .A(n3950), .B(n[99]), .Z(n13) );
  NAND U15 ( .A(n13), .B(n11), .Z(n14) );
  NAND U16 ( .A(n12), .B(n14), .Z(n15) );
  NAND U17 ( .A(n[100]), .B(n3946), .Z(n16) );
  XOR U18 ( .A(n3946), .B(n[100]), .Z(n17) );
  NAND U19 ( .A(n17), .B(n15), .Z(n18) );
  NAND U20 ( .A(n16), .B(n18), .Z(n2323) );
  XOR U21 ( .A(n3369), .B(n[242]), .Z(n19) );
  NANDN U22 ( .A(n3366), .B(n19), .Z(n20) );
  NAND U23 ( .A(n3369), .B(n[242]), .Z(n21) );
  AND U24 ( .A(n20), .B(n21), .Z(n3362) );
  NAND U25 ( .A(n6456), .B(n5257), .Z(n22) );
  XOR U26 ( .A(n5257), .B(n6456), .Z(n23) );
  NANDN U27 ( .A(n5260), .B(n23), .Z(n24) );
  NAND U28 ( .A(n22), .B(n24), .Z(n3383) );
  XOR U29 ( .A(n3512), .B(n[205]), .Z(n25) );
  NANDN U30 ( .A(n3509), .B(n25), .Z(n26) );
  NAND U31 ( .A(n3512), .B(n[205]), .Z(n27) );
  AND U32 ( .A(n26), .B(n27), .Z(n3504) );
  XOR U33 ( .A(n3726), .B(n[150]), .Z(n28) );
  NANDN U34 ( .A(n3723), .B(n28), .Z(n29) );
  NAND U35 ( .A(n3726), .B(n[150]), .Z(n30) );
  AND U36 ( .A(n29), .B(n30), .Z(n3719) );
  XOR U37 ( .A(n3373), .B(n[241]), .Z(n31) );
  NANDN U38 ( .A(n3370), .B(n31), .Z(n32) );
  NAND U39 ( .A(n3373), .B(n[241]), .Z(n33) );
  AND U40 ( .A(n32), .B(n33), .Z(n3366) );
  NAND U41 ( .A(n6449), .B(n3387), .Z(n34) );
  XOR U42 ( .A(n3387), .B(n6449), .Z(n35) );
  NANDN U43 ( .A(n3390), .B(n35), .Z(n36) );
  NAND U44 ( .A(n34), .B(n36), .Z(n5257) );
  XOR U45 ( .A(n5233), .B(n[230]), .Z(n37) );
  NANDN U46 ( .A(n5230), .B(n37), .Z(n38) );
  NAND U47 ( .A(n5233), .B(n[230]), .Z(n39) );
  AND U48 ( .A(n38), .B(n39), .Z(n3408) );
  XOR U49 ( .A(n3447), .B(n[221]), .Z(n40) );
  NANDN U50 ( .A(n3444), .B(n40), .Z(n41) );
  NAND U51 ( .A(n3447), .B(n[221]), .Z(n42) );
  AND U52 ( .A(n41), .B(n42), .Z(n3440) );
  XOR U53 ( .A(n3463), .B(n[216]), .Z(n43) );
  NANDN U54 ( .A(n3460), .B(n43), .Z(n44) );
  NAND U55 ( .A(n3463), .B(n[216]), .Z(n45) );
  AND U56 ( .A(n44), .B(n45), .Z(n5175) );
  XOR U57 ( .A(n3484), .B(n[211]), .Z(n46) );
  NANDN U58 ( .A(n3481), .B(n46), .Z(n47) );
  NAND U59 ( .A(n3484), .B(n[211]), .Z(n48) );
  AND U60 ( .A(n47), .B(n48), .Z(n3477) );
  XOR U61 ( .A(n3542), .B(n[198]), .Z(n49) );
  NANDN U62 ( .A(n3539), .B(n49), .Z(n50) );
  NAND U63 ( .A(n3542), .B(n[198]), .Z(n51) );
  AND U64 ( .A(n50), .B(n51), .Z(n3534) );
  XOR U65 ( .A(n3560), .B(n[194]), .Z(n52) );
  NANDN U66 ( .A(n3557), .B(n52), .Z(n53) );
  NAND U67 ( .A(n3560), .B(n[194]), .Z(n54) );
  AND U68 ( .A(n53), .B(n54), .Z(n3551) );
  XOR U69 ( .A(n3615), .B(n[180]), .Z(n55) );
  NANDN U70 ( .A(n3612), .B(n55), .Z(n56) );
  NAND U71 ( .A(n3615), .B(n[180]), .Z(n57) );
  AND U72 ( .A(n56), .B(n57), .Z(n3608) );
  XOR U73 ( .A(n3685), .B(n[163]), .Z(n58) );
  NANDN U74 ( .A(n3682), .B(n58), .Z(n59) );
  NAND U75 ( .A(n3685), .B(n[163]), .Z(n60) );
  AND U76 ( .A(n59), .B(n60), .Z(n3678) );
  XOR U77 ( .A(n3734), .B(n3731), .Z(n61) );
  NAND U78 ( .A(n61), .B(n[148]), .Z(n62) );
  NAND U79 ( .A(n3734), .B(n3731), .Z(n63) );
  AND U80 ( .A(n62), .B(n63), .Z(n3727) );
  XOR U81 ( .A(n3773), .B(n[139]), .Z(n64) );
  NANDN U82 ( .A(n3770), .B(n64), .Z(n65) );
  NAND U83 ( .A(n3773), .B(n[139]), .Z(n66) );
  AND U84 ( .A(n65), .B(n66), .Z(n3765) );
  XOR U85 ( .A(n3785), .B(n[136]), .Z(n67) );
  NANDN U86 ( .A(n3782), .B(n67), .Z(n68) );
  NAND U87 ( .A(n3785), .B(n[136]), .Z(n69) );
  AND U88 ( .A(n68), .B(n69), .Z(n3778) );
  XOR U89 ( .A(n3920), .B(n[106]), .Z(n70) );
  NANDN U90 ( .A(n3917), .B(n70), .Z(n71) );
  NAND U91 ( .A(n3920), .B(n[106]), .Z(n72) );
  AND U92 ( .A(n71), .B(n72), .Z(n3913) );
  NAND U93 ( .A(n5344), .B(n3947), .Z(n73) );
  XOR U94 ( .A(n3947), .B(n5344), .Z(n74) );
  NANDN U95 ( .A(n3950), .B(n74), .Z(n75) );
  NAND U96 ( .A(n73), .B(n75), .Z(n3943) );
  XOR U97 ( .A(n4010), .B(n[84]), .Z(n76) );
  NANDN U98 ( .A(n4007), .B(n76), .Z(n77) );
  NAND U99 ( .A(n4010), .B(n[84]), .Z(n78) );
  AND U100 ( .A(n77), .B(n78), .Z(n4003) );
  XOR U101 ( .A(n4032), .B(n[79]), .Z(n79) );
  NANDN U102 ( .A(n4029), .B(n79), .Z(n80) );
  NAND U103 ( .A(n4032), .B(n[79]), .Z(n81) );
  AND U104 ( .A(n80), .B(n81), .Z(n4024) );
  XOR U105 ( .A(n3331), .B(n[251]), .Z(n82) );
  NANDN U106 ( .A(n3328), .B(n82), .Z(n83) );
  NAND U107 ( .A(n3331), .B(n[251]), .Z(n84) );
  AND U108 ( .A(n83), .B(n84), .Z(n3323) );
  XOR U109 ( .A(n3403), .B(n[233]), .Z(n85) );
  NANDN U110 ( .A(n3400), .B(n85), .Z(n86) );
  NAND U111 ( .A(n3403), .B(n[233]), .Z(n87) );
  AND U112 ( .A(n86), .B(n87), .Z(n3395) );
  XOR U113 ( .A(n3503), .B(n3500), .Z(n88) );
  NAND U114 ( .A(n88), .B(n[207]), .Z(n89) );
  NAND U115 ( .A(n3503), .B(n3500), .Z(n90) );
  AND U116 ( .A(n89), .B(n90), .Z(n3495) );
  XOR U117 ( .A(n3702), .B(n3699), .Z(n91) );
  NAND U118 ( .A(n91), .B(n[159]), .Z(n92) );
  NAND U119 ( .A(n3702), .B(n3699), .Z(n93) );
  AND U120 ( .A(n92), .B(n93), .Z(n3694) );
  XOR U121 ( .A(n4209), .B(n[34]), .Z(n94) );
  NANDN U122 ( .A(n4206), .B(n94), .Z(n95) );
  NAND U123 ( .A(n4209), .B(n[34]), .Z(n96) );
  AND U124 ( .A(n95), .B(n96), .Z(n4428) );
  NAND U125 ( .A(n4399), .B(n4398), .Z(n97) );
  XOR U126 ( .A(n4398), .B(n4399), .Z(n98) );
  NANDN U127 ( .A(n2879), .B(n98), .Z(n99) );
  NAND U128 ( .A(n97), .B(n99), .Z(n4403) );
  NAND U129 ( .A(n[1]), .B(n4296), .Z(n100) );
  XOR U130 ( .A(n4296), .B(n[1]), .Z(n101) );
  NANDN U131 ( .A(n4299), .B(n101), .Z(n102) );
  NAND U132 ( .A(n100), .B(n102), .Z(n4300) );
  XOR U133 ( .A(n5928), .B(n5929), .Z(n103) );
  NANDN U134 ( .A(n5927), .B(n103), .Z(n104) );
  NAND U135 ( .A(n5928), .B(n5929), .Z(n105) );
  AND U136 ( .A(n104), .B(n105), .Z(n5933) );
  NAND U137 ( .A(n5621), .B(n5620), .Z(n106) );
  XOR U138 ( .A(n5620), .B(n5621), .Z(n107) );
  NANDN U139 ( .A(n5622), .B(n107), .Z(n108) );
  NAND U140 ( .A(n106), .B(n108), .Z(n5624) );
  XOR U141 ( .A(n[3]), .B(n6676), .Z(n109) );
  NAND U142 ( .A(n109), .B(n6673), .Z(n110) );
  NAND U143 ( .A(n[3]), .B(n6676), .Z(n111) );
  AND U144 ( .A(n110), .B(n111), .Z(n6726) );
  XOR U145 ( .A(n3394), .B(n[235]), .Z(n112) );
  NANDN U146 ( .A(n3391), .B(n112), .Z(n113) );
  NAND U147 ( .A(n3394), .B(n[235]), .Z(n114) );
  AND U148 ( .A(n113), .B(n114), .Z(n3387) );
  XOR U149 ( .A(n4073), .B(n[69]), .Z(n115) );
  NANDN U150 ( .A(n4070), .B(n115), .Z(n116) );
  NAND U151 ( .A(n4073), .B(n[69]), .Z(n117) );
  AND U152 ( .A(n116), .B(n117), .Z(n4066) );
  XOR U153 ( .A(n3343), .B(n3340), .Z(n118) );
  NAND U154 ( .A(n118), .B(n[248]), .Z(n119) );
  NAND U155 ( .A(n3343), .B(n3340), .Z(n120) );
  AND U156 ( .A(n119), .B(n120), .Z(n3336) );
  XOR U157 ( .A(n3423), .B(n[227]), .Z(n121) );
  NANDN U158 ( .A(n3420), .B(n121), .Z(n122) );
  NAND U159 ( .A(n3423), .B(n[227]), .Z(n123) );
  AND U160 ( .A(n122), .B(n123), .Z(n3416) );
  XOR U161 ( .A(n3435), .B(n[224]), .Z(n124) );
  NANDN U162 ( .A(n3432), .B(n124), .Z(n125) );
  NAND U163 ( .A(n3435), .B(n[224]), .Z(n126) );
  AND U164 ( .A(n125), .B(n126), .Z(n3428) );
  XOR U165 ( .A(n3451), .B(n[220]), .Z(n127) );
  NANDN U166 ( .A(n3448), .B(n127), .Z(n128) );
  NAND U167 ( .A(n3451), .B(n[220]), .Z(n129) );
  AND U168 ( .A(n128), .B(n129), .Z(n3444) );
  XOR U169 ( .A(n5178), .B(n[217]), .Z(n130) );
  NANDN U170 ( .A(n5175), .B(n130), .Z(n131) );
  NAND U171 ( .A(n5178), .B(n[217]), .Z(n132) );
  AND U172 ( .A(n131), .B(n132), .Z(n3456) );
  XOR U173 ( .A(n3471), .B(n3468), .Z(n133) );
  NAND U174 ( .A(n133), .B(n[214]), .Z(n134) );
  NAND U175 ( .A(n3471), .B(n3468), .Z(n135) );
  AND U176 ( .A(n134), .B(n135), .Z(n3464) );
  NAND U177 ( .A(n6268), .B(n3485), .Z(n136) );
  XOR U178 ( .A(n3485), .B(n6268), .Z(n137) );
  NANDN U179 ( .A(n2874), .B(n137), .Z(n138) );
  NAND U180 ( .A(n136), .B(n138), .Z(n3481) );
  XOR U181 ( .A(n3546), .B(n[197]), .Z(n139) );
  NANDN U182 ( .A(n3543), .B(n139), .Z(n140) );
  NAND U183 ( .A(n3546), .B(n[197]), .Z(n141) );
  AND U184 ( .A(n140), .B(n141), .Z(n3539) );
  XOR U185 ( .A(n3564), .B(n[193]), .Z(n142) );
  NANDN U186 ( .A(n3561), .B(n142), .Z(n143) );
  NAND U187 ( .A(n3564), .B(n[193]), .Z(n144) );
  AND U188 ( .A(n143), .B(n144), .Z(n3557) );
  XOR U189 ( .A(n3577), .B(n2875), .Z(n145) );
  NANDN U190 ( .A(n3581), .B(n145), .Z(n146) );
  NAND U191 ( .A(n3577), .B(n2875), .Z(n147) );
  AND U192 ( .A(n146), .B(n147), .Z(n3573) );
  XOR U193 ( .A(n3594), .B(n[186]), .Z(n148) );
  NANDN U194 ( .A(n3591), .B(n148), .Z(n149) );
  NAND U195 ( .A(n3594), .B(n[186]), .Z(n150) );
  AND U196 ( .A(n149), .B(n150), .Z(n3587) );
  XOR U197 ( .A(n3607), .B(n[182]), .Z(n151) );
  NANDN U198 ( .A(n3604), .B(n151), .Z(n152) );
  NAND U199 ( .A(n3607), .B(n[182]), .Z(n153) );
  AND U200 ( .A(n152), .B(n153), .Z(n3599) );
  XOR U201 ( .A(n5026), .B(n[179]), .Z(n154) );
  NANDN U202 ( .A(n5023), .B(n154), .Z(n155) );
  NAND U203 ( .A(n5026), .B(n[179]), .Z(n156) );
  AND U204 ( .A(n155), .B(n156), .Z(n3612) );
  XOR U205 ( .A(n3625), .B(n3628), .Z(n157) );
  NANDN U206 ( .A(n6025), .B(n157), .Z(n158) );
  NAND U207 ( .A(n3625), .B(n3628), .Z(n159) );
  AND U208 ( .A(n158), .B(n159), .Z(n3620) );
  XOR U209 ( .A(n3689), .B(n[162]), .Z(n160) );
  NANDN U210 ( .A(n3686), .B(n160), .Z(n161) );
  NAND U211 ( .A(n3689), .B(n[162]), .Z(n162) );
  AND U212 ( .A(n161), .B(n162), .Z(n3682) );
  XOR U213 ( .A(n3764), .B(n3761), .Z(n163) );
  NAND U214 ( .A(n163), .B(n[141]), .Z(n164) );
  NAND U215 ( .A(n3764), .B(n3761), .Z(n165) );
  AND U216 ( .A(n164), .B(n165), .Z(n3757) );
  XOR U217 ( .A(n3781), .B(n[137]), .Z(n166) );
  NANDN U218 ( .A(n3778), .B(n166), .Z(n167) );
  NAND U219 ( .A(n3781), .B(n[137]), .Z(n168) );
  AND U220 ( .A(n167), .B(n168), .Z(n3774) );
  XOR U221 ( .A(n3793), .B(n3790), .Z(n169) );
  NAND U222 ( .A(n169), .B(n[134]), .Z(n170) );
  NAND U223 ( .A(n3793), .B(n3790), .Z(n171) );
  AND U224 ( .A(n170), .B(n171), .Z(n3786) );
  XOR U225 ( .A(n3823), .B(n[127]), .Z(n172) );
  NANDN U226 ( .A(n3820), .B(n172), .Z(n173) );
  NAND U227 ( .A(n3823), .B(n[127]), .Z(n174) );
  AND U228 ( .A(n173), .B(n174), .Z(n3816) );
  XOR U229 ( .A(n3916), .B(n[107]), .Z(n175) );
  NANDN U230 ( .A(n3913), .B(n175), .Z(n176) );
  NAND U231 ( .A(n3916), .B(n[107]), .Z(n177) );
  AND U232 ( .A(n176), .B(n177), .Z(n3908) );
  XOR U233 ( .A(n3928), .B(n3925), .Z(n178) );
  NAND U234 ( .A(n178), .B(n[104]), .Z(n179) );
  NAND U235 ( .A(n3928), .B(n3925), .Z(n180) );
  AND U236 ( .A(n179), .B(n180), .Z(n3921) );
  XOR U237 ( .A(n3958), .B(n3955), .Z(n181) );
  NAND U238 ( .A(n181), .B(n[97]), .Z(n182) );
  NAND U239 ( .A(n3958), .B(n3955), .Z(n183) );
  AND U240 ( .A(n182), .B(n183), .Z(n3951) );
  XOR U241 ( .A(n3993), .B(n3990), .Z(n184) );
  NAND U242 ( .A(n184), .B(n[88]), .Z(n185) );
  NAND U243 ( .A(n3993), .B(n3990), .Z(n186) );
  AND U244 ( .A(n185), .B(n186), .Z(n3986) );
  XOR U245 ( .A(n4014), .B(n[83]), .Z(n187) );
  NANDN U246 ( .A(n4011), .B(n187), .Z(n188) );
  NAND U247 ( .A(n4014), .B(n[83]), .Z(n189) );
  AND U248 ( .A(n188), .B(n189), .Z(n4007) );
  XOR U249 ( .A(n4057), .B(n[73]), .Z(n190) );
  NANDN U250 ( .A(n4054), .B(n190), .Z(n191) );
  NAND U251 ( .A(n4057), .B(n[73]), .Z(n192) );
  AND U252 ( .A(n191), .B(n192), .Z(n4050) );
  XOR U253 ( .A(n4086), .B(n[66]), .Z(n193) );
  NAND U254 ( .A(n193), .B(n4083), .Z(n194) );
  NAND U255 ( .A(n4086), .B(n[66]), .Z(n195) );
  AND U256 ( .A(n194), .B(n195), .Z(n4079) );
  ANDN U257 ( .B(n[46]), .A(n4174), .Z(n2989) );
  XOR U258 ( .A(n3322), .B(n3319), .Z(n196) );
  NAND U259 ( .A(n196), .B(n[253]), .Z(n197) );
  NAND U260 ( .A(n3322), .B(n3319), .Z(n198) );
  AND U261 ( .A(n197), .B(n198), .Z(n3315) );
  XOR U262 ( .A(n3365), .B(n[243]), .Z(n199) );
  NANDN U263 ( .A(n3362), .B(n199), .Z(n200) );
  NAND U264 ( .A(n3365), .B(n[243]), .Z(n201) );
  AND U265 ( .A(n200), .B(n201), .Z(n3357) );
  XOR U266 ( .A(n3386), .B(n[238]), .Z(n202) );
  NANDN U267 ( .A(n3383), .B(n202), .Z(n203) );
  NAND U268 ( .A(n3386), .B(n[238]), .Z(n204) );
  AND U269 ( .A(n203), .B(n204), .Z(n3378) );
  XOR U270 ( .A(n3407), .B(n3404), .Z(n205) );
  NAND U271 ( .A(n205), .B(n[232]), .Z(n206) );
  NAND U272 ( .A(n3407), .B(n3404), .Z(n207) );
  AND U273 ( .A(n206), .B(n207), .Z(n3400) );
  XOR U274 ( .A(n3516), .B(n3513), .Z(n208) );
  NAND U275 ( .A(n208), .B(n[204]), .Z(n209) );
  NAND U276 ( .A(n3516), .B(n3513), .Z(n210) );
  AND U277 ( .A(n209), .B(n210), .Z(n3509) );
  XOR U278 ( .A(n3659), .B(n3656), .Z(n211) );
  NAND U279 ( .A(n211), .B(n[169]), .Z(n212) );
  NAND U280 ( .A(n3659), .B(n3656), .Z(n213) );
  AND U281 ( .A(n212), .B(n213), .Z(n3651) );
  XOR U282 ( .A(n3718), .B(n3715), .Z(n214) );
  NAND U283 ( .A(n214), .B(n[152]), .Z(n215) );
  NAND U284 ( .A(n3718), .B(n3715), .Z(n216) );
  AND U285 ( .A(n215), .B(n216), .Z(n4909) );
  XOR U286 ( .A(n3730), .B(n[149]), .Z(n217) );
  NANDN U287 ( .A(n3727), .B(n217), .Z(n218) );
  NAND U288 ( .A(n3730), .B(n[149]), .Z(n219) );
  AND U289 ( .A(n218), .B(n219), .Z(n3723) );
  XOR U290 ( .A(n3836), .B(n3833), .Z(n220) );
  NAND U291 ( .A(n220), .B(n[124]), .Z(n221) );
  NAND U292 ( .A(n3836), .B(n3833), .Z(n222) );
  AND U293 ( .A(n221), .B(n222), .Z(n3828) );
  XOR U294 ( .A(n3946), .B(n[100]), .Z(n223) );
  NANDN U295 ( .A(n3943), .B(n223), .Z(n224) );
  NAND U296 ( .A(n3946), .B(n[100]), .Z(n225) );
  AND U297 ( .A(n224), .B(n225), .Z(n3938) );
  XOR U298 ( .A(n4045), .B(n[76]), .Z(n226) );
  NANDN U299 ( .A(n4042), .B(n226), .Z(n227) );
  NAND U300 ( .A(n4045), .B(n[76]), .Z(n228) );
  AND U301 ( .A(n227), .B(n228), .Z(n4037) );
  NAND U302 ( .A(n4432), .B(n4428), .Z(n229) );
  XOR U303 ( .A(n4428), .B(n4432), .Z(n230) );
  NANDN U304 ( .A(n4431), .B(n230), .Z(n231) );
  NAND U305 ( .A(n229), .B(n231), .Z(n4202) );
  XOR U306 ( .A(n4217), .B(n4214), .Z(n232) );
  NAND U307 ( .A(n232), .B(n[32]), .Z(n233) );
  NAND U308 ( .A(n4217), .B(n4214), .Z(n234) );
  AND U309 ( .A(n233), .B(n234), .Z(n4210) );
  XOR U310 ( .A(n[28]), .B(n6613), .Z(n235) );
  NAND U311 ( .A(n235), .B(n6610), .Z(n236) );
  NAND U312 ( .A(n[28]), .B(n6613), .Z(n237) );
  AND U313 ( .A(n236), .B(n237), .Z(n6614) );
  XOR U314 ( .A(n4230), .B(n[26]), .Z(n238) );
  NANDN U315 ( .A(n4227), .B(n238), .Z(n239) );
  NAND U316 ( .A(n4230), .B(n[26]), .Z(n240) );
  AND U317 ( .A(n239), .B(n240), .Z(n4398) );
  XNOR U318 ( .A(n6544), .B(n4239), .Z(n241) );
  NANDN U319 ( .A(n4387), .B(n6473), .Z(n242) );
  XOR U320 ( .A(n6473), .B(n[23]), .Z(n243) );
  NAND U321 ( .A(n243), .B(n6537), .Z(n244) );
  NAND U322 ( .A(n242), .B(n244), .Z(n245) );
  NAND U323 ( .A(n241), .B(n245), .Z(n246) );
  NANDN U324 ( .A(n4239), .B(n6544), .Z(n247) );
  AND U325 ( .A(n246), .B(n247), .Z(n6595) );
  NANDN U326 ( .A(n4358), .B(n5918), .Z(n248) );
  XOR U327 ( .A(n5918), .B(n[15]), .Z(n249) );
  NAND U328 ( .A(n249), .B(n5978), .Z(n250) );
  NAND U329 ( .A(n248), .B(n250), .Z(n251) );
  XNOR U330 ( .A(n5985), .B(n4266), .Z(n252) );
  NAND U331 ( .A(n252), .B(n251), .Z(n253) );
  NANDN U332 ( .A(n4266), .B(n5985), .Z(n254) );
  AND U333 ( .A(n253), .B(n254), .Z(n6054) );
  NAND U334 ( .A(n6439), .B(n6438), .Z(n255) );
  XOR U335 ( .A(n6438), .B(n6439), .Z(n256) );
  NANDN U336 ( .A(n6440), .B(n256), .Z(n257) );
  NAND U337 ( .A(n255), .B(n257), .Z(n6445) );
  NAND U338 ( .A(n6250), .B(n6251), .Z(n258) );
  XOR U339 ( .A(n6251), .B(n6250), .Z(n259) );
  NANDN U340 ( .A(n6249), .B(n259), .Z(n260) );
  NAND U341 ( .A(n258), .B(n260), .Z(n6253) );
  XOR U342 ( .A(n5924), .B(n5925), .Z(n261) );
  NANDN U343 ( .A(n5923), .B(n261), .Z(n262) );
  NAND U344 ( .A(n5924), .B(n5925), .Z(n263) );
  AND U345 ( .A(n262), .B(n263), .Z(n5927) );
  NAND U346 ( .A(n5616), .B(n5617), .Z(n264) );
  XOR U347 ( .A(n5617), .B(n5616), .Z(n265) );
  NANDN U348 ( .A(n5618), .B(n265), .Z(n266) );
  NAND U349 ( .A(n264), .B(n266), .Z(n5620) );
  XOR U350 ( .A(n6810), .B(n6812), .Z(n267) );
  NAND U351 ( .A(n267), .B(n6809), .Z(n268) );
  NAND U352 ( .A(n6810), .B(n6812), .Z(n269) );
  AND U353 ( .A(n268), .B(n269), .Z(n6816) );
  XOR U354 ( .A(n6776), .B(n6773), .Z(n270) );
  NANDN U355 ( .A(n6774), .B(n270), .Z(n271) );
  NAND U356 ( .A(n6776), .B(n6773), .Z(n272) );
  AND U357 ( .A(n271), .B(n272), .Z(n6778) );
  XOR U358 ( .A(n6731), .B(n6730), .Z(n273) );
  NAND U359 ( .A(n273), .B(n6733), .Z(n274) );
  NAND U360 ( .A(n6731), .B(n6730), .Z(n275) );
  AND U361 ( .A(n274), .B(n275), .Z(n6735) );
  XOR U362 ( .A(n[44]), .B(n6705), .Z(n276) );
  NAND U363 ( .A(n276), .B(n6702), .Z(n277) );
  NAND U364 ( .A(n[44]), .B(n6705), .Z(n278) );
  AND U365 ( .A(n277), .B(n278), .Z(n6706) );
  NAND U366 ( .A(n6615), .B(n6619), .Z(n279) );
  XOR U367 ( .A(n6619), .B(n6615), .Z(n280) );
  NANDN U368 ( .A(n6616), .B(n280), .Z(n281) );
  NAND U369 ( .A(n279), .B(n281), .Z(n6673) );
  XOR U370 ( .A(n3377), .B(n3374), .Z(n282) );
  NAND U371 ( .A(n282), .B(n[240]), .Z(n283) );
  NAND U372 ( .A(n3377), .B(n3374), .Z(n284) );
  AND U373 ( .A(n283), .B(n284), .Z(n3370) );
  NAND U374 ( .A(n3399), .B(n3395), .Z(n285) );
  XOR U375 ( .A(n3395), .B(n3399), .Z(n286) );
  NANDN U376 ( .A(n2872), .B(n286), .Z(n287) );
  NAND U377 ( .A(n285), .B(n287), .Z(n3391) );
  XOR U378 ( .A(n3415), .B(n[229]), .Z(n288) );
  NANDN U379 ( .A(n3412), .B(n288), .Z(n289) );
  NAND U380 ( .A(n3415), .B(n[229]), .Z(n290) );
  AND U381 ( .A(n289), .B(n290), .Z(n5230) );
  XOR U382 ( .A(n3427), .B(n3424), .Z(n291) );
  NAND U383 ( .A(n291), .B(n[226]), .Z(n292) );
  NAND U384 ( .A(n3427), .B(n3424), .Z(n293) );
  AND U385 ( .A(n292), .B(n293), .Z(n3420) );
  XOR U386 ( .A(n3439), .B(n3436), .Z(n294) );
  NAND U387 ( .A(n294), .B(n[223]), .Z(n295) );
  NAND U388 ( .A(n3439), .B(n3436), .Z(n296) );
  AND U389 ( .A(n295), .B(n296), .Z(n3432) );
  XOR U390 ( .A(n3455), .B(n3452), .Z(n297) );
  NAND U391 ( .A(n297), .B(n[219]), .Z(n298) );
  NAND U392 ( .A(n3455), .B(n3452), .Z(n299) );
  AND U393 ( .A(n298), .B(n299), .Z(n3448) );
  XOR U394 ( .A(n3467), .B(n[215]), .Z(n300) );
  NANDN U395 ( .A(n3464), .B(n300), .Z(n301) );
  NAND U396 ( .A(n3467), .B(n[215]), .Z(n302) );
  AND U397 ( .A(n301), .B(n302), .Z(n3460) );
  XOR U398 ( .A(n3480), .B(n[212]), .Z(n303) );
  NANDN U399 ( .A(n3477), .B(n303), .Z(n304) );
  NAND U400 ( .A(n3480), .B(n[212]), .Z(n305) );
  AND U401 ( .A(n304), .B(n305), .Z(n3472) );
  XOR U402 ( .A(n3489), .B(n3492), .Z(n306) );
  NANDN U403 ( .A(n6256), .B(n306), .Z(n307) );
  NAND U404 ( .A(n3489), .B(n3492), .Z(n308) );
  AND U405 ( .A(n307), .B(n308), .Z(n3485) );
  XOR U406 ( .A(n3524), .B(n3521), .Z(n309) );
  NAND U407 ( .A(n309), .B(n[202]), .Z(n310) );
  NAND U408 ( .A(n3524), .B(n3521), .Z(n311) );
  AND U409 ( .A(n310), .B(n311), .Z(n3517) );
  XOR U410 ( .A(n3537), .B(n[199]), .Z(n312) );
  NANDN U411 ( .A(n3534), .B(n312), .Z(n313) );
  NAND U412 ( .A(n3537), .B(n[199]), .Z(n314) );
  AND U413 ( .A(n313), .B(n314), .Z(n3530) );
  XOR U414 ( .A(n3547), .B(n3550), .Z(n315) );
  NANDN U415 ( .A(n6166), .B(n315), .Z(n316) );
  NAND U416 ( .A(n3547), .B(n3550), .Z(n317) );
  AND U417 ( .A(n316), .B(n317), .Z(n3543) );
  XOR U418 ( .A(n3568), .B(n3565), .Z(n318) );
  NAND U419 ( .A(n318), .B(n[192]), .Z(n319) );
  NAND U420 ( .A(n3568), .B(n3565), .Z(n320) );
  AND U421 ( .A(n319), .B(n320), .Z(n3561) );
  XOR U422 ( .A(n5054), .B(n5051), .Z(n321) );
  NAND U423 ( .A(n321), .B(n[185]), .Z(n322) );
  NAND U424 ( .A(n5054), .B(n5051), .Z(n323) );
  AND U425 ( .A(n322), .B(n323), .Z(n3591) );
  XOR U426 ( .A(n3611), .B(n[181]), .Z(n324) );
  NANDN U427 ( .A(n3608), .B(n324), .Z(n325) );
  NAND U428 ( .A(n3611), .B(n[181]), .Z(n326) );
  AND U429 ( .A(n325), .B(n326), .Z(n3604) );
  XOR U430 ( .A(n3616), .B(n3619), .Z(n327) );
  NANDN U431 ( .A(n6039), .B(n327), .Z(n328) );
  NAND U432 ( .A(n3616), .B(n3619), .Z(n329) );
  AND U433 ( .A(n328), .B(n329), .Z(n5023) );
  XOR U434 ( .A(n3636), .B(n3633), .Z(n330) );
  NAND U435 ( .A(n330), .B(n[174]), .Z(n331) );
  NAND U436 ( .A(n3636), .B(n3633), .Z(n332) );
  AND U437 ( .A(n331), .B(n332), .Z(n3629) );
  XOR U438 ( .A(n3693), .B(n3690), .Z(n333) );
  NAND U439 ( .A(n333), .B(n[161]), .Z(n334) );
  NAND U440 ( .A(n3693), .B(n3690), .Z(n335) );
  AND U441 ( .A(n334), .B(n335), .Z(n3686) );
  XOR U442 ( .A(n4926), .B(n4923), .Z(n336) );
  NAND U443 ( .A(n336), .B(n[155]), .Z(n337) );
  NAND U444 ( .A(n4926), .B(n4923), .Z(n338) );
  AND U445 ( .A(n337), .B(n338), .Z(n3707) );
  XOR U446 ( .A(n3743), .B(n3740), .Z(n339) );
  NAND U447 ( .A(n339), .B(n[146]), .Z(n340) );
  NAND U448 ( .A(n3743), .B(n3740), .Z(n341) );
  AND U449 ( .A(n340), .B(n341), .Z(n3735) );
  XOR U450 ( .A(n3756), .B(n[143]), .Z(n342) );
  NANDN U451 ( .A(n3753), .B(n342), .Z(n343) );
  NAND U452 ( .A(n3756), .B(n[143]), .Z(n344) );
  AND U453 ( .A(n343), .B(n344), .Z(n3748) );
  XOR U454 ( .A(n3777), .B(n[138]), .Z(n345) );
  NANDN U455 ( .A(n3774), .B(n345), .Z(n346) );
  NAND U456 ( .A(n3777), .B(n[138]), .Z(n347) );
  AND U457 ( .A(n346), .B(n347), .Z(n3770) );
  XOR U458 ( .A(n3789), .B(n[135]), .Z(n348) );
  NANDN U459 ( .A(n3786), .B(n348), .Z(n349) );
  NAND U460 ( .A(n3789), .B(n[135]), .Z(n350) );
  AND U461 ( .A(n349), .B(n350), .Z(n3782) );
  XOR U462 ( .A(n3802), .B(n3799), .Z(n351) );
  NAND U463 ( .A(n351), .B(n[132]), .Z(n352) );
  NAND U464 ( .A(n3802), .B(n3799), .Z(n353) );
  AND U465 ( .A(n352), .B(n353), .Z(n3794) );
  XOR U466 ( .A(n3815), .B(n3812), .Z(n354) );
  NAND U467 ( .A(n354), .B(n[129]), .Z(n355) );
  NAND U468 ( .A(n3815), .B(n3812), .Z(n356) );
  AND U469 ( .A(n355), .B(n356), .Z(n3807) );
  XOR U470 ( .A(n3827), .B(n3824), .Z(n357) );
  NAND U471 ( .A(n357), .B(n[126]), .Z(n358) );
  NAND U472 ( .A(n3827), .B(n3824), .Z(n359) );
  AND U473 ( .A(n358), .B(n359), .Z(n3820) );
  XOR U474 ( .A(n3924), .B(n[105]), .Z(n360) );
  NANDN U475 ( .A(n3921), .B(n360), .Z(n361) );
  NAND U476 ( .A(n3924), .B(n[105]), .Z(n362) );
  AND U477 ( .A(n361), .B(n362), .Z(n3917) );
  XOR U478 ( .A(n3937), .B(n3934), .Z(n363) );
  NAND U479 ( .A(n363), .B(n[102]), .Z(n364) );
  NAND U480 ( .A(n3937), .B(n3934), .Z(n365) );
  AND U481 ( .A(n364), .B(n365), .Z(n3929) );
  XOR U482 ( .A(n3985), .B(n3982), .Z(n366) );
  NAND U483 ( .A(n366), .B(n[90]), .Z(n367) );
  NAND U484 ( .A(n3985), .B(n3982), .Z(n368) );
  AND U485 ( .A(n367), .B(n368), .Z(n3978) );
  XOR U486 ( .A(n4002), .B(n3999), .Z(n369) );
  NAND U487 ( .A(n369), .B(n[86]), .Z(n370) );
  NAND U488 ( .A(n4002), .B(n3999), .Z(n371) );
  AND U489 ( .A(n370), .B(n371), .Z(n3994) );
  XOR U490 ( .A(n4018), .B(n4015), .Z(n372) );
  NAND U491 ( .A(n372), .B(n[82]), .Z(n373) );
  NAND U492 ( .A(n4018), .B(n4015), .Z(n374) );
  AND U493 ( .A(n373), .B(n374), .Z(n4011) );
  XOR U494 ( .A(n4049), .B(n[75]), .Z(n375) );
  NANDN U495 ( .A(n4046), .B(n375), .Z(n376) );
  NAND U496 ( .A(n4049), .B(n[75]), .Z(n377) );
  AND U497 ( .A(n376), .B(n377), .Z(n4042) );
  XOR U498 ( .A(n4062), .B(n4065), .Z(n378) );
  NANDN U499 ( .A(n5390), .B(n378), .Z(n379) );
  NAND U500 ( .A(n4062), .B(n4065), .Z(n380) );
  AND U501 ( .A(n379), .B(n380), .Z(n4058) );
  XOR U502 ( .A(n4099), .B(n4096), .Z(n381) );
  NAND U503 ( .A(n381), .B(n[63]), .Z(n382) );
  NAND U504 ( .A(n4099), .B(n4096), .Z(n383) );
  AND U505 ( .A(n382), .B(n383), .Z(n4092) );
  NAND U506 ( .A(n[57]), .B(n4126), .Z(n384) );
  XOR U507 ( .A(n4126), .B(n[57]), .Z(n385) );
  NANDN U508 ( .A(n4123), .B(n385), .Z(n386) );
  NAND U509 ( .A(n384), .B(n386), .Z(n4119) );
  XOR U510 ( .A(n4153), .B(n4150), .Z(n387) );
  NAND U511 ( .A(n387), .B(n[51]), .Z(n388) );
  NAND U512 ( .A(n4153), .B(n4150), .Z(n389) );
  AND U513 ( .A(n388), .B(n389), .Z(n4146) );
  XOR U514 ( .A(n3335), .B(n3332), .Z(n390) );
  NAND U515 ( .A(n390), .B(n[250]), .Z(n391) );
  NAND U516 ( .A(n3335), .B(n3332), .Z(n392) );
  AND U517 ( .A(n391), .B(n392), .Z(n3328) );
  NAND U518 ( .A(n2856), .B(n2855), .Z(n393) );
  NAND U519 ( .A(n[251]), .B(n3331), .Z(n394) );
  NAND U520 ( .A(n393), .B(n394), .Z(n395) );
  XNOR U521 ( .A(n3327), .B(n3326), .Z(n396) );
  NAND U522 ( .A(n396), .B(n395), .Z(n397) );
  NAND U523 ( .A(n397), .B(n3300), .Z(n398) );
  NAND U524 ( .A(n[253]), .B(n3322), .Z(n399) );
  XOR U525 ( .A(n3322), .B(n[253]), .Z(n400) );
  NAND U526 ( .A(n400), .B(n398), .Z(n401) );
  NAND U527 ( .A(n399), .B(n401), .Z(n402) );
  XNOR U528 ( .A(n6582), .B(n3318), .Z(n403) );
  NAND U529 ( .A(n403), .B(n402), .Z(n404) );
  AND U530 ( .A(n3303), .B(n404), .Z(n405) );
  NANDN U531 ( .A(n405), .B(n3308), .Z(n406) );
  XNOR U532 ( .A(n3308), .B(n405), .Z(n407) );
  NAND U533 ( .A(n407), .B(n[255]), .Z(n408) );
  NAND U534 ( .A(n406), .B(n408), .Z(n409) );
  ANDN U535 ( .B(n409), .A(n3313), .Z(n410) );
  NANDN U536 ( .A(n3312), .B(n410), .Z(n523) );
  NANDN U537 ( .A(n6457), .B(n[237]), .Z(n6459) );
  XOR U538 ( .A(n3954), .B(n[98]), .Z(n411) );
  NANDN U539 ( .A(n3951), .B(n411), .Z(n412) );
  NAND U540 ( .A(n3954), .B(n[98]), .Z(n413) );
  AND U541 ( .A(n412), .B(n413), .Z(n3947) );
  XOR U542 ( .A(n4036), .B(n4033), .Z(n414) );
  NAND U543 ( .A(n414), .B(n[78]), .Z(n415) );
  NAND U544 ( .A(n4036), .B(n4033), .Z(n416) );
  AND U545 ( .A(n415), .B(n416), .Z(n4029) );
  XOR U546 ( .A(n4082), .B(n[67]), .Z(n417) );
  NANDN U547 ( .A(n4079), .B(n417), .Z(n418) );
  NAND U548 ( .A(n4082), .B(n[67]), .Z(n419) );
  AND U549 ( .A(n418), .B(n419), .Z(n4074) );
  XOR U550 ( .A(n4474), .B(n[45]), .Z(n420) );
  NANDN U551 ( .A(n4471), .B(n420), .Z(n421) );
  NAND U552 ( .A(n4474), .B(n[45]), .Z(n422) );
  AND U553 ( .A(n421), .B(n422), .Z(n4171) );
  XOR U554 ( .A(n4213), .B(n[33]), .Z(n423) );
  NANDN U555 ( .A(n4210), .B(n423), .Z(n424) );
  NAND U556 ( .A(n4213), .B(n[33]), .Z(n425) );
  AND U557 ( .A(n424), .B(n425), .Z(n4206) );
  XOR U558 ( .A(n4234), .B(n4231), .Z(n426) );
  NAND U559 ( .A(n426), .B(n[25]), .Z(n427) );
  NAND U560 ( .A(n4234), .B(n4231), .Z(n428) );
  AND U561 ( .A(n427), .B(n428), .Z(n4227) );
  XOR U562 ( .A(n5716), .B(n5719), .Z(n429) );
  NAND U563 ( .A(n429), .B(n[12]), .Z(n430) );
  NAND U564 ( .A(n5716), .B(n5719), .Z(n431) );
  AND U565 ( .A(n430), .B(n431), .Z(n5782) );
  XOR U566 ( .A(n6505), .B(n6504), .Z(n432) );
  NANDN U567 ( .A(n6503), .B(n432), .Z(n433) );
  NAND U568 ( .A(n6505), .B(n6504), .Z(n434) );
  AND U569 ( .A(n433), .B(n434), .Z(n6510) );
  XOR U570 ( .A(n6474), .B(n6475), .Z(n435) );
  NAND U571 ( .A(n435), .B(n6476), .Z(n436) );
  NAND U572 ( .A(n6474), .B(n6475), .Z(n437) );
  AND U573 ( .A(n436), .B(n437), .Z(n6479) );
  XOR U574 ( .A(n6436), .B(n6435), .Z(n438) );
  NANDN U575 ( .A(n6434), .B(n438), .Z(n439) );
  NAND U576 ( .A(n6436), .B(n6435), .Z(n440) );
  AND U577 ( .A(n439), .B(n440), .Z(n6438) );
  NAND U578 ( .A(n6302), .B(n6303), .Z(n441) );
  XOR U579 ( .A(n6303), .B(n6302), .Z(n442) );
  NANDN U580 ( .A(n6304), .B(n442), .Z(n443) );
  NAND U581 ( .A(n441), .B(n443), .Z(n6307) );
  XOR U582 ( .A(n6254), .B(n6255), .Z(n444) );
  NANDN U583 ( .A(n6253), .B(n444), .Z(n445) );
  NAND U584 ( .A(n6254), .B(n6255), .Z(n446) );
  AND U585 ( .A(n445), .B(n446), .Z(n6274) );
  XOR U586 ( .A(n6239), .B(n6240), .Z(n447) );
  NAND U587 ( .A(n447), .B(n6241), .Z(n448) );
  NAND U588 ( .A(n6239), .B(n6240), .Z(n449) );
  AND U589 ( .A(n448), .B(n449), .Z(n6244) );
  XOR U590 ( .A(n6130), .B(n6131), .Z(n450) );
  NAND U591 ( .A(n450), .B(n6132), .Z(n451) );
  NAND U592 ( .A(n6130), .B(n6131), .Z(n452) );
  AND U593 ( .A(n451), .B(n452), .Z(n6139) );
  NAND U594 ( .A(n5995), .B(n5993), .Z(n453) );
  NANDN U595 ( .A(n5995), .B(n5994), .Z(n454) );
  NANDN U596 ( .A(n5996), .B(n454), .Z(n455) );
  NAND U597 ( .A(n453), .B(n455), .Z(n6002) );
  NAND U598 ( .A(n5919), .B(n5920), .Z(n456) );
  XOR U599 ( .A(n5920), .B(n5919), .Z(n457) );
  NAND U600 ( .A(n457), .B(n5921), .Z(n458) );
  NAND U601 ( .A(n456), .B(n458), .Z(n5925) );
  XOR U602 ( .A(n5881), .B(n5880), .Z(n459) );
  NANDN U603 ( .A(n5879), .B(n459), .Z(n460) );
  NAND U604 ( .A(n5881), .B(n5880), .Z(n461) );
  AND U605 ( .A(n460), .B(n461), .Z(n5885) );
  XOR U606 ( .A(n5863), .B(n5862), .Z(n462) );
  NANDN U607 ( .A(n5861), .B(n462), .Z(n463) );
  NAND U608 ( .A(n5863), .B(n5862), .Z(n464) );
  AND U609 ( .A(n463), .B(n464), .Z(n5868) );
  NAND U610 ( .A(n5796), .B(n5797), .Z(n465) );
  XOR U611 ( .A(n5797), .B(n5796), .Z(n466) );
  NANDN U612 ( .A(n5798), .B(n466), .Z(n467) );
  NAND U613 ( .A(n465), .B(n467), .Z(n5803) );
  XOR U614 ( .A(n5696), .B(n5695), .Z(n468) );
  NANDN U615 ( .A(n5694), .B(n468), .Z(n469) );
  NAND U616 ( .A(n5696), .B(n5695), .Z(n470) );
  AND U617 ( .A(n469), .B(n470), .Z(n5699) );
  XOR U618 ( .A(n5666), .B(n5667), .Z(n471) );
  NAND U619 ( .A(n471), .B(n5668), .Z(n472) );
  NAND U620 ( .A(n5666), .B(n5667), .Z(n473) );
  AND U621 ( .A(n472), .B(n473), .Z(n5671) );
  NAND U622 ( .A(n5625), .B(n5624), .Z(n474) );
  XOR U623 ( .A(n5624), .B(n5625), .Z(n475) );
  NANDN U624 ( .A(n5626), .B(n475), .Z(n476) );
  NAND U625 ( .A(n474), .B(n476), .Z(n5629) );
  NAND U626 ( .A(n5612), .B(n5613), .Z(n477) );
  XOR U627 ( .A(n5613), .B(n5612), .Z(n478) );
  NAND U628 ( .A(n478), .B(n5614), .Z(n479) );
  NAND U629 ( .A(n477), .B(n479), .Z(n5617) );
  XOR U630 ( .A(n5569), .B(n5568), .Z(n480) );
  NANDN U631 ( .A(n5567), .B(n480), .Z(n481) );
  NAND U632 ( .A(n5569), .B(n5568), .Z(n482) );
  AND U633 ( .A(n481), .B(n482), .Z(n5572) );
  XOR U634 ( .A(n5551), .B(n5552), .Z(n483) );
  NAND U635 ( .A(n483), .B(n5553), .Z(n484) );
  NAND U636 ( .A(n5551), .B(n5552), .Z(n485) );
  AND U637 ( .A(n484), .B(n485), .Z(n5556) );
  XOR U638 ( .A(n6862), .B(n6859), .Z(n486) );
  NANDN U639 ( .A(n6860), .B(n486), .Z(n487) );
  NAND U640 ( .A(n6862), .B(n6859), .Z(n488) );
  AND U641 ( .A(n487), .B(n488), .Z(n6864) );
  XOR U642 ( .A(n6804), .B(n6806), .Z(n489) );
  NAND U643 ( .A(n489), .B(n6803), .Z(n490) );
  NAND U644 ( .A(n6804), .B(n6806), .Z(n491) );
  AND U645 ( .A(n490), .B(n491), .Z(n6807) );
  XOR U646 ( .A(n6770), .B(n6767), .Z(n492) );
  NANDN U647 ( .A(n6768), .B(n492), .Z(n493) );
  NAND U648 ( .A(n6770), .B(n6767), .Z(n494) );
  AND U649 ( .A(n493), .B(n494), .Z(n6772) );
  XOR U650 ( .A(n6741), .B(n6738), .Z(n495) );
  NANDN U651 ( .A(n6739), .B(n495), .Z(n496) );
  NAND U652 ( .A(n6741), .B(n6738), .Z(n497) );
  AND U653 ( .A(n496), .B(n497), .Z(n6743) );
  NAND U654 ( .A(n6723), .B(n6725), .Z(n498) );
  XOR U655 ( .A(n6725), .B(n6723), .Z(n499) );
  NAND U656 ( .A(n499), .B(n6722), .Z(n500) );
  NAND U657 ( .A(n498), .B(n500), .Z(n6730) );
  NAND U658 ( .A(n6698), .B(n6701), .Z(n501) );
  XOR U659 ( .A(n6701), .B(n6698), .Z(n502) );
  NANDN U660 ( .A(n4463), .B(n502), .Z(n503) );
  NAND U661 ( .A(n501), .B(n503), .Z(n6702) );
  NANDN U662 ( .A(n4416), .B(n6630), .Z(n504) );
  XOR U663 ( .A(n6630), .B(n[31]), .Z(n505) );
  NAND U664 ( .A(n505), .B(n6633), .Z(n506) );
  NAND U665 ( .A(n504), .B(n506), .Z(n507) );
  XOR U666 ( .A(n[32]), .B(n6640), .Z(n508) );
  NAND U667 ( .A(n508), .B(n507), .Z(n509) );
  NAND U668 ( .A(n[32]), .B(n6640), .Z(n510) );
  AND U669 ( .A(n509), .B(n510), .Z(n6641) );
  NAND U670 ( .A(n6606), .B(n6609), .Z(n511) );
  XOR U671 ( .A(n6609), .B(n6606), .Z(n512) );
  NANDN U672 ( .A(n4399), .B(n512), .Z(n513) );
  NAND U673 ( .A(n511), .B(n513), .Z(n6610) );
  XOR U674 ( .A(n[21]), .B(n6334), .Z(n514) );
  NAND U675 ( .A(n514), .B(n6331), .Z(n515) );
  NAND U676 ( .A(n[21]), .B(n6334), .Z(n516) );
  AND U677 ( .A(n515), .B(n516), .Z(n6403) );
  XOR U678 ( .A(n6867), .B(n6871), .Z(n517) );
  NANDN U679 ( .A(n6868), .B(n517), .Z(n518) );
  NAND U680 ( .A(n6867), .B(n6871), .Z(n519) );
  AND U681 ( .A(n518), .B(n519), .Z(n5595) );
  NAND U682 ( .A(n6195), .B(n[1]), .Z(n520) );
  XOR U683 ( .A(n[1]), .B(n6195), .Z(n521) );
  NANDN U684 ( .A(n6198), .B(n521), .Z(n522) );
  NAND U685 ( .A(n520), .B(n522), .Z(n6615) );
  IV U686 ( .A(n523), .Z(n524) );
  IV U687 ( .A(n6814), .Z(n525) );
  AND U688 ( .A(N4), .B(xregN_1), .Z(n2880) );
  IV U689 ( .A(n[254]), .Z(n6582) );
  NAND U690 ( .A(y[253]), .B(zin[252]), .Z(n1281) );
  XOR U691 ( .A(zin[252]), .B(y[253]), .Z(n1279) );
  NAND U692 ( .A(y[252]), .B(zin[251]), .Z(n1278) );
  XOR U693 ( .A(zin[251]), .B(y[252]), .Z(n1276) );
  NAND U694 ( .A(y[251]), .B(zin[250]), .Z(n1275) );
  XOR U695 ( .A(zin[250]), .B(y[251]), .Z(n1273) );
  NAND U696 ( .A(y[250]), .B(zin[249]), .Z(n1272) );
  XOR U697 ( .A(zin[249]), .B(y[250]), .Z(n1270) );
  NAND U698 ( .A(y[249]), .B(zin[248]), .Z(n1269) );
  XOR U699 ( .A(zin[248]), .B(y[249]), .Z(n1267) );
  NAND U700 ( .A(y[248]), .B(zin[247]), .Z(n1266) );
  XOR U701 ( .A(zin[247]), .B(y[248]), .Z(n1264) );
  NAND U702 ( .A(y[247]), .B(zin[246]), .Z(n1263) );
  XOR U703 ( .A(zin[246]), .B(y[247]), .Z(n1261) );
  NAND U704 ( .A(y[246]), .B(zin[245]), .Z(n1260) );
  XOR U705 ( .A(zin[245]), .B(y[246]), .Z(n1258) );
  NAND U706 ( .A(y[245]), .B(zin[244]), .Z(n1257) );
  XOR U707 ( .A(zin[244]), .B(y[245]), .Z(n1255) );
  NAND U708 ( .A(y[244]), .B(zin[243]), .Z(n1254) );
  XOR U709 ( .A(zin[243]), .B(y[244]), .Z(n1252) );
  NAND U710 ( .A(y[243]), .B(zin[242]), .Z(n1251) );
  XOR U711 ( .A(zin[242]), .B(y[243]), .Z(n1249) );
  NAND U712 ( .A(y[242]), .B(zin[241]), .Z(n1248) );
  XOR U713 ( .A(zin[241]), .B(y[242]), .Z(n1246) );
  NAND U714 ( .A(y[241]), .B(zin[240]), .Z(n1245) );
  XOR U715 ( .A(zin[240]), .B(y[241]), .Z(n1243) );
  NAND U716 ( .A(y[240]), .B(zin[239]), .Z(n1242) );
  XOR U717 ( .A(zin[239]), .B(y[240]), .Z(n1240) );
  NAND U718 ( .A(y[239]), .B(zin[238]), .Z(n1239) );
  XOR U719 ( .A(zin[238]), .B(y[239]), .Z(n1237) );
  NAND U720 ( .A(y[238]), .B(zin[237]), .Z(n1236) );
  XOR U721 ( .A(zin[237]), .B(y[238]), .Z(n1234) );
  NAND U722 ( .A(y[237]), .B(zin[236]), .Z(n1233) );
  XOR U723 ( .A(zin[236]), .B(y[237]), .Z(n1231) );
  NAND U724 ( .A(y[236]), .B(zin[235]), .Z(n1230) );
  XOR U725 ( .A(zin[235]), .B(y[236]), .Z(n1228) );
  NAND U726 ( .A(y[235]), .B(zin[234]), .Z(n1227) );
  XOR U727 ( .A(zin[234]), .B(y[235]), .Z(n1225) );
  NAND U728 ( .A(y[234]), .B(zin[233]), .Z(n1224) );
  XOR U729 ( .A(zin[233]), .B(y[234]), .Z(n1222) );
  NAND U730 ( .A(y[233]), .B(zin[232]), .Z(n1221) );
  XOR U731 ( .A(zin[232]), .B(y[233]), .Z(n1219) );
  NAND U732 ( .A(y[232]), .B(zin[231]), .Z(n1218) );
  XOR U733 ( .A(zin[231]), .B(y[232]), .Z(n1216) );
  NAND U734 ( .A(y[231]), .B(zin[230]), .Z(n1215) );
  XOR U735 ( .A(zin[230]), .B(y[231]), .Z(n1213) );
  NAND U736 ( .A(y[230]), .B(zin[229]), .Z(n1212) );
  XOR U737 ( .A(zin[229]), .B(y[230]), .Z(n1210) );
  NAND U738 ( .A(y[229]), .B(zin[228]), .Z(n1209) );
  XOR U739 ( .A(zin[228]), .B(y[229]), .Z(n1207) );
  NAND U740 ( .A(y[228]), .B(zin[227]), .Z(n1206) );
  XOR U741 ( .A(zin[227]), .B(y[228]), .Z(n1204) );
  NAND U742 ( .A(y[227]), .B(zin[226]), .Z(n1203) );
  XOR U743 ( .A(zin[226]), .B(y[227]), .Z(n1201) );
  NAND U744 ( .A(y[226]), .B(zin[225]), .Z(n1200) );
  XOR U745 ( .A(zin[225]), .B(y[226]), .Z(n1198) );
  NAND U746 ( .A(y[225]), .B(zin[224]), .Z(n1197) );
  XOR U747 ( .A(zin[224]), .B(y[225]), .Z(n1195) );
  NAND U748 ( .A(y[224]), .B(zin[223]), .Z(n1194) );
  XOR U749 ( .A(zin[223]), .B(y[224]), .Z(n1192) );
  NAND U750 ( .A(y[223]), .B(zin[222]), .Z(n1191) );
  XOR U751 ( .A(zin[222]), .B(y[223]), .Z(n1189) );
  NAND U752 ( .A(y[222]), .B(zin[221]), .Z(n1188) );
  XOR U753 ( .A(zin[221]), .B(y[222]), .Z(n1186) );
  NAND U754 ( .A(y[221]), .B(zin[220]), .Z(n1185) );
  XOR U755 ( .A(zin[220]), .B(y[221]), .Z(n1183) );
  NAND U756 ( .A(y[220]), .B(zin[219]), .Z(n1182) );
  XOR U757 ( .A(zin[219]), .B(y[220]), .Z(n1180) );
  NAND U758 ( .A(y[219]), .B(zin[218]), .Z(n1179) );
  XOR U759 ( .A(zin[218]), .B(y[219]), .Z(n1177) );
  NAND U760 ( .A(y[218]), .B(zin[217]), .Z(n1176) );
  XOR U761 ( .A(zin[217]), .B(y[218]), .Z(n1174) );
  NAND U762 ( .A(y[217]), .B(zin[216]), .Z(n1173) );
  XOR U763 ( .A(zin[216]), .B(y[217]), .Z(n1171) );
  NAND U764 ( .A(y[216]), .B(zin[215]), .Z(n1170) );
  XOR U765 ( .A(zin[215]), .B(y[216]), .Z(n1168) );
  NAND U766 ( .A(y[215]), .B(zin[214]), .Z(n1167) );
  XOR U767 ( .A(zin[214]), .B(y[215]), .Z(n1165) );
  NAND U768 ( .A(y[214]), .B(zin[213]), .Z(n1164) );
  XOR U769 ( .A(zin[213]), .B(y[214]), .Z(n1162) );
  NAND U770 ( .A(y[213]), .B(zin[212]), .Z(n1161) );
  XOR U771 ( .A(zin[212]), .B(y[213]), .Z(n1159) );
  NAND U772 ( .A(y[212]), .B(zin[211]), .Z(n1158) );
  XOR U773 ( .A(zin[211]), .B(y[212]), .Z(n1156) );
  NAND U774 ( .A(y[211]), .B(zin[210]), .Z(n1155) );
  XOR U775 ( .A(zin[210]), .B(y[211]), .Z(n1153) );
  NAND U776 ( .A(y[210]), .B(zin[209]), .Z(n1152) );
  XOR U777 ( .A(zin[209]), .B(y[210]), .Z(n1150) );
  NAND U778 ( .A(y[209]), .B(zin[208]), .Z(n1149) );
  XOR U779 ( .A(zin[208]), .B(y[209]), .Z(n1147) );
  NAND U780 ( .A(y[208]), .B(zin[207]), .Z(n1146) );
  XOR U781 ( .A(zin[207]), .B(y[208]), .Z(n1144) );
  NAND U782 ( .A(y[207]), .B(zin[206]), .Z(n1143) );
  XOR U783 ( .A(zin[206]), .B(y[207]), .Z(n1141) );
  NAND U784 ( .A(y[206]), .B(zin[205]), .Z(n1140) );
  XOR U785 ( .A(zin[205]), .B(y[206]), .Z(n1138) );
  NAND U786 ( .A(y[205]), .B(zin[204]), .Z(n1137) );
  XOR U787 ( .A(zin[204]), .B(y[205]), .Z(n1135) );
  NAND U788 ( .A(y[204]), .B(zin[203]), .Z(n1134) );
  XOR U789 ( .A(zin[203]), .B(y[204]), .Z(n1132) );
  NAND U790 ( .A(y[203]), .B(zin[202]), .Z(n1131) );
  XOR U791 ( .A(zin[202]), .B(y[203]), .Z(n1129) );
  NAND U792 ( .A(y[202]), .B(zin[201]), .Z(n1128) );
  XOR U793 ( .A(zin[201]), .B(y[202]), .Z(n1126) );
  NAND U794 ( .A(y[201]), .B(zin[200]), .Z(n1125) );
  XOR U795 ( .A(zin[200]), .B(y[201]), .Z(n1123) );
  NAND U796 ( .A(y[200]), .B(zin[199]), .Z(n1122) );
  XOR U797 ( .A(zin[199]), .B(y[200]), .Z(n1120) );
  NAND U798 ( .A(y[199]), .B(zin[198]), .Z(n1119) );
  XOR U799 ( .A(zin[198]), .B(y[199]), .Z(n1117) );
  NAND U800 ( .A(y[198]), .B(zin[197]), .Z(n1116) );
  XOR U801 ( .A(zin[197]), .B(y[198]), .Z(n1114) );
  NAND U802 ( .A(y[197]), .B(zin[196]), .Z(n1113) );
  XOR U803 ( .A(zin[196]), .B(y[197]), .Z(n1111) );
  NAND U804 ( .A(y[196]), .B(zin[195]), .Z(n1110) );
  XOR U805 ( .A(zin[195]), .B(y[196]), .Z(n1108) );
  NAND U806 ( .A(y[195]), .B(zin[194]), .Z(n1107) );
  XOR U807 ( .A(zin[194]), .B(y[195]), .Z(n1105) );
  NAND U808 ( .A(y[194]), .B(zin[193]), .Z(n1104) );
  XOR U809 ( .A(zin[193]), .B(y[194]), .Z(n1102) );
  NAND U810 ( .A(y[193]), .B(zin[192]), .Z(n1101) );
  XOR U811 ( .A(zin[192]), .B(y[193]), .Z(n1099) );
  NAND U812 ( .A(y[192]), .B(zin[191]), .Z(n1098) );
  XOR U813 ( .A(zin[191]), .B(y[192]), .Z(n1096) );
  NAND U814 ( .A(y[191]), .B(zin[190]), .Z(n1095) );
  XOR U815 ( .A(zin[190]), .B(y[191]), .Z(n1093) );
  NAND U816 ( .A(y[190]), .B(zin[189]), .Z(n1092) );
  XOR U817 ( .A(zin[189]), .B(y[190]), .Z(n1090) );
  NAND U818 ( .A(y[189]), .B(zin[188]), .Z(n1089) );
  XOR U819 ( .A(zin[188]), .B(y[189]), .Z(n1087) );
  NAND U820 ( .A(y[188]), .B(zin[187]), .Z(n1086) );
  XOR U821 ( .A(zin[187]), .B(y[188]), .Z(n1084) );
  NAND U822 ( .A(y[187]), .B(zin[186]), .Z(n1083) );
  XOR U823 ( .A(zin[186]), .B(y[187]), .Z(n1081) );
  NAND U824 ( .A(y[186]), .B(zin[185]), .Z(n1080) );
  XOR U825 ( .A(zin[185]), .B(y[186]), .Z(n1078) );
  NAND U826 ( .A(y[185]), .B(zin[184]), .Z(n1077) );
  XOR U827 ( .A(zin[184]), .B(y[185]), .Z(n1075) );
  NAND U828 ( .A(y[184]), .B(zin[183]), .Z(n1074) );
  XOR U829 ( .A(zin[183]), .B(y[184]), .Z(n1072) );
  NAND U830 ( .A(y[183]), .B(zin[182]), .Z(n1071) );
  XOR U831 ( .A(zin[182]), .B(y[183]), .Z(n1069) );
  NAND U832 ( .A(y[182]), .B(zin[181]), .Z(n1068) );
  XOR U833 ( .A(zin[181]), .B(y[182]), .Z(n1066) );
  NAND U834 ( .A(y[181]), .B(zin[180]), .Z(n1065) );
  XOR U835 ( .A(zin[180]), .B(y[181]), .Z(n1063) );
  NAND U836 ( .A(y[180]), .B(zin[179]), .Z(n1062) );
  XOR U837 ( .A(zin[179]), .B(y[180]), .Z(n1060) );
  NAND U838 ( .A(y[179]), .B(zin[178]), .Z(n1059) );
  XOR U839 ( .A(zin[178]), .B(y[179]), .Z(n1057) );
  NAND U840 ( .A(y[178]), .B(zin[177]), .Z(n1056) );
  XOR U841 ( .A(zin[177]), .B(y[178]), .Z(n1054) );
  NAND U842 ( .A(y[177]), .B(zin[176]), .Z(n1053) );
  XOR U843 ( .A(zin[176]), .B(y[177]), .Z(n1051) );
  NAND U844 ( .A(y[176]), .B(zin[175]), .Z(n1050) );
  XOR U845 ( .A(zin[175]), .B(y[176]), .Z(n1048) );
  NAND U846 ( .A(y[175]), .B(zin[174]), .Z(n1047) );
  XOR U847 ( .A(zin[174]), .B(y[175]), .Z(n1045) );
  NAND U848 ( .A(y[174]), .B(zin[173]), .Z(n1044) );
  XOR U849 ( .A(zin[173]), .B(y[174]), .Z(n1042) );
  NAND U850 ( .A(y[173]), .B(zin[172]), .Z(n1041) );
  XOR U851 ( .A(zin[172]), .B(y[173]), .Z(n1039) );
  NAND U852 ( .A(y[172]), .B(zin[171]), .Z(n1038) );
  XOR U853 ( .A(zin[171]), .B(y[172]), .Z(n1036) );
  NAND U854 ( .A(y[171]), .B(zin[170]), .Z(n1035) );
  XOR U855 ( .A(zin[170]), .B(y[171]), .Z(n1033) );
  NAND U856 ( .A(y[170]), .B(zin[169]), .Z(n1032) );
  XOR U857 ( .A(zin[169]), .B(y[170]), .Z(n1030) );
  NAND U858 ( .A(y[169]), .B(zin[168]), .Z(n1029) );
  XOR U859 ( .A(zin[168]), .B(y[169]), .Z(n1027) );
  NAND U860 ( .A(y[168]), .B(zin[167]), .Z(n1026) );
  XOR U861 ( .A(zin[167]), .B(y[168]), .Z(n1024) );
  NAND U862 ( .A(y[167]), .B(zin[166]), .Z(n1023) );
  XOR U863 ( .A(zin[166]), .B(y[167]), .Z(n1021) );
  NAND U864 ( .A(y[166]), .B(zin[165]), .Z(n1020) );
  XOR U865 ( .A(zin[165]), .B(y[166]), .Z(n1018) );
  NAND U866 ( .A(y[165]), .B(zin[164]), .Z(n1017) );
  XOR U867 ( .A(zin[164]), .B(y[165]), .Z(n1015) );
  NAND U868 ( .A(y[164]), .B(zin[163]), .Z(n1014) );
  XOR U869 ( .A(zin[163]), .B(y[164]), .Z(n1012) );
  NAND U870 ( .A(y[163]), .B(zin[162]), .Z(n1011) );
  XOR U871 ( .A(zin[162]), .B(y[163]), .Z(n1009) );
  NAND U872 ( .A(y[162]), .B(zin[161]), .Z(n1008) );
  XOR U873 ( .A(zin[161]), .B(y[162]), .Z(n1006) );
  NAND U874 ( .A(y[161]), .B(zin[160]), .Z(n1005) );
  XOR U875 ( .A(zin[160]), .B(y[161]), .Z(n1003) );
  NAND U876 ( .A(y[160]), .B(zin[159]), .Z(n1002) );
  XOR U877 ( .A(zin[159]), .B(y[160]), .Z(n1000) );
  NAND U878 ( .A(y[159]), .B(zin[158]), .Z(n999) );
  XOR U879 ( .A(zin[158]), .B(y[159]), .Z(n997) );
  NAND U880 ( .A(y[158]), .B(zin[157]), .Z(n996) );
  XOR U881 ( .A(zin[157]), .B(y[158]), .Z(n994) );
  NAND U882 ( .A(y[157]), .B(zin[156]), .Z(n993) );
  XOR U883 ( .A(zin[156]), .B(y[157]), .Z(n991) );
  NAND U884 ( .A(y[156]), .B(zin[155]), .Z(n990) );
  XOR U885 ( .A(zin[155]), .B(y[156]), .Z(n988) );
  NAND U886 ( .A(y[155]), .B(zin[154]), .Z(n987) );
  XOR U887 ( .A(zin[154]), .B(y[155]), .Z(n985) );
  NAND U888 ( .A(y[154]), .B(zin[153]), .Z(n984) );
  XOR U889 ( .A(zin[153]), .B(y[154]), .Z(n982) );
  NAND U890 ( .A(y[153]), .B(zin[152]), .Z(n981) );
  XOR U891 ( .A(zin[152]), .B(y[153]), .Z(n979) );
  NAND U892 ( .A(y[152]), .B(zin[151]), .Z(n978) );
  XOR U893 ( .A(zin[151]), .B(y[152]), .Z(n976) );
  NAND U894 ( .A(y[151]), .B(zin[150]), .Z(n975) );
  XOR U895 ( .A(zin[150]), .B(y[151]), .Z(n973) );
  NAND U896 ( .A(y[150]), .B(zin[149]), .Z(n972) );
  XOR U897 ( .A(zin[149]), .B(y[150]), .Z(n970) );
  NAND U898 ( .A(y[149]), .B(zin[148]), .Z(n969) );
  XOR U899 ( .A(zin[148]), .B(y[149]), .Z(n967) );
  NAND U900 ( .A(y[148]), .B(zin[147]), .Z(n966) );
  XOR U901 ( .A(zin[147]), .B(y[148]), .Z(n964) );
  NAND U902 ( .A(y[147]), .B(zin[146]), .Z(n963) );
  XOR U903 ( .A(zin[146]), .B(y[147]), .Z(n961) );
  NAND U904 ( .A(y[146]), .B(zin[145]), .Z(n960) );
  XOR U905 ( .A(zin[145]), .B(y[146]), .Z(n958) );
  NAND U906 ( .A(y[145]), .B(zin[144]), .Z(n957) );
  XOR U907 ( .A(zin[144]), .B(y[145]), .Z(n955) );
  NAND U908 ( .A(y[144]), .B(zin[143]), .Z(n954) );
  XOR U909 ( .A(zin[143]), .B(y[144]), .Z(n952) );
  NAND U910 ( .A(y[143]), .B(zin[142]), .Z(n951) );
  XOR U911 ( .A(zin[142]), .B(y[143]), .Z(n949) );
  NAND U912 ( .A(y[142]), .B(zin[141]), .Z(n948) );
  XOR U913 ( .A(zin[141]), .B(y[142]), .Z(n946) );
  NAND U914 ( .A(y[141]), .B(zin[140]), .Z(n945) );
  XOR U915 ( .A(zin[140]), .B(y[141]), .Z(n943) );
  NAND U916 ( .A(y[140]), .B(zin[139]), .Z(n942) );
  XOR U917 ( .A(zin[139]), .B(y[140]), .Z(n940) );
  NAND U918 ( .A(y[139]), .B(zin[138]), .Z(n939) );
  XOR U919 ( .A(zin[138]), .B(y[139]), .Z(n937) );
  NAND U920 ( .A(y[138]), .B(zin[137]), .Z(n936) );
  XOR U921 ( .A(zin[137]), .B(y[138]), .Z(n934) );
  NAND U922 ( .A(y[137]), .B(zin[136]), .Z(n933) );
  XOR U923 ( .A(zin[136]), .B(y[137]), .Z(n931) );
  NAND U924 ( .A(y[136]), .B(zin[135]), .Z(n930) );
  XOR U925 ( .A(zin[135]), .B(y[136]), .Z(n928) );
  NAND U926 ( .A(y[135]), .B(zin[134]), .Z(n927) );
  XOR U927 ( .A(zin[134]), .B(y[135]), .Z(n925) );
  NAND U928 ( .A(y[134]), .B(zin[133]), .Z(n924) );
  XOR U929 ( .A(zin[133]), .B(y[134]), .Z(n922) );
  NAND U930 ( .A(y[133]), .B(zin[132]), .Z(n921) );
  XOR U931 ( .A(zin[132]), .B(y[133]), .Z(n919) );
  NAND U932 ( .A(y[132]), .B(zin[131]), .Z(n918) );
  XOR U933 ( .A(zin[131]), .B(y[132]), .Z(n916) );
  NAND U934 ( .A(y[131]), .B(zin[130]), .Z(n915) );
  XOR U935 ( .A(zin[130]), .B(y[131]), .Z(n913) );
  NAND U936 ( .A(y[130]), .B(zin[129]), .Z(n912) );
  XOR U937 ( .A(zin[129]), .B(y[130]), .Z(n910) );
  NAND U938 ( .A(y[129]), .B(zin[128]), .Z(n909) );
  XOR U939 ( .A(zin[128]), .B(y[129]), .Z(n907) );
  NAND U940 ( .A(y[128]), .B(zin[127]), .Z(n906) );
  XOR U941 ( .A(zin[127]), .B(y[128]), .Z(n904) );
  NAND U942 ( .A(y[127]), .B(zin[126]), .Z(n903) );
  XOR U943 ( .A(zin[126]), .B(y[127]), .Z(n901) );
  NAND U944 ( .A(y[126]), .B(zin[125]), .Z(n900) );
  XOR U945 ( .A(zin[125]), .B(y[126]), .Z(n898) );
  NAND U946 ( .A(y[125]), .B(zin[124]), .Z(n897) );
  XOR U947 ( .A(zin[124]), .B(y[125]), .Z(n895) );
  NAND U948 ( .A(y[124]), .B(zin[123]), .Z(n894) );
  XOR U949 ( .A(zin[123]), .B(y[124]), .Z(n892) );
  NAND U950 ( .A(y[123]), .B(zin[122]), .Z(n891) );
  XOR U951 ( .A(zin[122]), .B(y[123]), .Z(n889) );
  NAND U952 ( .A(y[122]), .B(zin[121]), .Z(n888) );
  XOR U953 ( .A(zin[121]), .B(y[122]), .Z(n886) );
  NAND U954 ( .A(y[121]), .B(zin[120]), .Z(n885) );
  XOR U955 ( .A(zin[120]), .B(y[121]), .Z(n883) );
  NAND U956 ( .A(y[120]), .B(zin[119]), .Z(n882) );
  XOR U957 ( .A(zin[119]), .B(y[120]), .Z(n880) );
  NAND U958 ( .A(y[119]), .B(zin[118]), .Z(n879) );
  XOR U959 ( .A(zin[118]), .B(y[119]), .Z(n877) );
  NAND U960 ( .A(y[118]), .B(zin[117]), .Z(n876) );
  XOR U961 ( .A(zin[117]), .B(y[118]), .Z(n874) );
  NAND U962 ( .A(y[117]), .B(zin[116]), .Z(n873) );
  XOR U963 ( .A(zin[116]), .B(y[117]), .Z(n871) );
  NAND U964 ( .A(y[116]), .B(zin[115]), .Z(n870) );
  XOR U965 ( .A(zin[115]), .B(y[116]), .Z(n868) );
  NAND U966 ( .A(y[115]), .B(zin[114]), .Z(n867) );
  XOR U967 ( .A(zin[114]), .B(y[115]), .Z(n865) );
  NAND U968 ( .A(y[114]), .B(zin[113]), .Z(n864) );
  XOR U969 ( .A(zin[113]), .B(y[114]), .Z(n862) );
  NAND U970 ( .A(y[113]), .B(zin[112]), .Z(n861) );
  XOR U971 ( .A(zin[112]), .B(y[113]), .Z(n859) );
  NAND U972 ( .A(y[112]), .B(zin[111]), .Z(n858) );
  XOR U973 ( .A(zin[111]), .B(y[112]), .Z(n856) );
  NAND U974 ( .A(y[111]), .B(zin[110]), .Z(n855) );
  XOR U975 ( .A(zin[110]), .B(y[111]), .Z(n853) );
  NAND U976 ( .A(y[110]), .B(zin[109]), .Z(n852) );
  XOR U977 ( .A(zin[109]), .B(y[110]), .Z(n850) );
  NAND U978 ( .A(y[109]), .B(zin[108]), .Z(n849) );
  XOR U979 ( .A(zin[108]), .B(y[109]), .Z(n847) );
  NAND U980 ( .A(y[108]), .B(zin[107]), .Z(n846) );
  XOR U981 ( .A(zin[107]), .B(y[108]), .Z(n844) );
  NAND U982 ( .A(y[107]), .B(zin[106]), .Z(n843) );
  XOR U983 ( .A(zin[106]), .B(y[107]), .Z(n841) );
  NAND U984 ( .A(y[106]), .B(zin[105]), .Z(n840) );
  XOR U985 ( .A(zin[105]), .B(y[106]), .Z(n838) );
  NAND U986 ( .A(y[105]), .B(zin[104]), .Z(n837) );
  XOR U987 ( .A(zin[104]), .B(y[105]), .Z(n835) );
  NAND U988 ( .A(y[104]), .B(zin[103]), .Z(n834) );
  XOR U989 ( .A(zin[103]), .B(y[104]), .Z(n832) );
  NAND U990 ( .A(y[103]), .B(zin[102]), .Z(n831) );
  XOR U991 ( .A(zin[102]), .B(y[103]), .Z(n829) );
  NAND U992 ( .A(y[102]), .B(zin[101]), .Z(n828) );
  XOR U993 ( .A(zin[101]), .B(y[102]), .Z(n826) );
  NAND U994 ( .A(y[101]), .B(zin[100]), .Z(n825) );
  XOR U995 ( .A(zin[100]), .B(y[101]), .Z(n823) );
  NAND U996 ( .A(y[100]), .B(zin[99]), .Z(n822) );
  XOR U997 ( .A(zin[99]), .B(y[100]), .Z(n820) );
  NAND U998 ( .A(zin[98]), .B(y[99]), .Z(n819) );
  XOR U999 ( .A(y[99]), .B(zin[98]), .Z(n817) );
  NAND U1000 ( .A(y[98]), .B(zin[97]), .Z(n816) );
  XOR U1001 ( .A(zin[97]), .B(y[98]), .Z(n814) );
  NAND U1002 ( .A(y[97]), .B(zin[96]), .Z(n813) );
  XOR U1003 ( .A(zin[96]), .B(y[97]), .Z(n811) );
  NAND U1004 ( .A(y[96]), .B(zin[95]), .Z(n810) );
  XOR U1005 ( .A(zin[95]), .B(y[96]), .Z(n808) );
  NAND U1006 ( .A(y[95]), .B(zin[94]), .Z(n807) );
  XOR U1007 ( .A(zin[94]), .B(y[95]), .Z(n805) );
  NAND U1008 ( .A(y[94]), .B(zin[93]), .Z(n804) );
  XOR U1009 ( .A(zin[93]), .B(y[94]), .Z(n802) );
  NAND U1010 ( .A(y[93]), .B(zin[92]), .Z(n801) );
  XOR U1011 ( .A(zin[92]), .B(y[93]), .Z(n799) );
  NAND U1012 ( .A(y[92]), .B(zin[91]), .Z(n798) );
  XOR U1013 ( .A(zin[91]), .B(y[92]), .Z(n796) );
  NAND U1014 ( .A(y[91]), .B(zin[90]), .Z(n795) );
  XOR U1015 ( .A(zin[90]), .B(y[91]), .Z(n793) );
  NAND U1016 ( .A(y[90]), .B(zin[89]), .Z(n792) );
  XOR U1017 ( .A(zin[89]), .B(y[90]), .Z(n790) );
  NAND U1018 ( .A(y[89]), .B(zin[88]), .Z(n789) );
  XOR U1019 ( .A(zin[88]), .B(y[89]), .Z(n787) );
  NAND U1020 ( .A(y[88]), .B(zin[87]), .Z(n786) );
  XOR U1021 ( .A(zin[87]), .B(y[88]), .Z(n784) );
  NAND U1022 ( .A(y[87]), .B(zin[86]), .Z(n783) );
  XOR U1023 ( .A(zin[86]), .B(y[87]), .Z(n781) );
  NAND U1024 ( .A(y[86]), .B(zin[85]), .Z(n780) );
  XOR U1025 ( .A(zin[85]), .B(y[86]), .Z(n778) );
  NAND U1026 ( .A(y[85]), .B(zin[84]), .Z(n777) );
  XOR U1027 ( .A(zin[84]), .B(y[85]), .Z(n775) );
  NAND U1028 ( .A(y[84]), .B(zin[83]), .Z(n774) );
  XOR U1029 ( .A(zin[83]), .B(y[84]), .Z(n772) );
  NAND U1030 ( .A(y[83]), .B(zin[82]), .Z(n771) );
  XOR U1031 ( .A(zin[82]), .B(y[83]), .Z(n769) );
  NAND U1032 ( .A(y[82]), .B(zin[81]), .Z(n768) );
  XOR U1033 ( .A(zin[81]), .B(y[82]), .Z(n766) );
  NAND U1034 ( .A(y[81]), .B(zin[80]), .Z(n765) );
  XOR U1035 ( .A(zin[80]), .B(y[81]), .Z(n763) );
  NAND U1036 ( .A(y[80]), .B(zin[79]), .Z(n762) );
  XOR U1037 ( .A(zin[79]), .B(y[80]), .Z(n760) );
  NAND U1038 ( .A(y[79]), .B(zin[78]), .Z(n759) );
  XOR U1039 ( .A(zin[78]), .B(y[79]), .Z(n757) );
  NAND U1040 ( .A(y[78]), .B(zin[77]), .Z(n756) );
  XOR U1041 ( .A(zin[77]), .B(y[78]), .Z(n754) );
  NAND U1042 ( .A(y[77]), .B(zin[76]), .Z(n753) );
  XOR U1043 ( .A(zin[76]), .B(y[77]), .Z(n751) );
  NAND U1044 ( .A(y[76]), .B(zin[75]), .Z(n750) );
  XOR U1045 ( .A(zin[75]), .B(y[76]), .Z(n748) );
  NAND U1046 ( .A(y[75]), .B(zin[74]), .Z(n747) );
  XOR U1047 ( .A(zin[74]), .B(y[75]), .Z(n745) );
  NAND U1048 ( .A(y[74]), .B(zin[73]), .Z(n744) );
  XOR U1049 ( .A(zin[73]), .B(y[74]), .Z(n742) );
  NAND U1050 ( .A(y[73]), .B(zin[72]), .Z(n741) );
  XOR U1051 ( .A(zin[72]), .B(y[73]), .Z(n739) );
  NAND U1052 ( .A(y[72]), .B(zin[71]), .Z(n738) );
  XOR U1053 ( .A(zin[71]), .B(y[72]), .Z(n736) );
  NAND U1054 ( .A(y[71]), .B(zin[70]), .Z(n735) );
  XOR U1055 ( .A(zin[70]), .B(y[71]), .Z(n733) );
  NAND U1056 ( .A(y[70]), .B(zin[69]), .Z(n732) );
  XOR U1057 ( .A(zin[69]), .B(y[70]), .Z(n730) );
  NAND U1058 ( .A(y[69]), .B(zin[68]), .Z(n729) );
  XOR U1059 ( .A(zin[68]), .B(y[69]), .Z(n727) );
  NAND U1060 ( .A(y[68]), .B(zin[67]), .Z(n726) );
  XOR U1061 ( .A(zin[67]), .B(y[68]), .Z(n724) );
  NAND U1062 ( .A(y[67]), .B(zin[66]), .Z(n723) );
  XOR U1063 ( .A(zin[66]), .B(y[67]), .Z(n721) );
  NAND U1064 ( .A(y[66]), .B(zin[65]), .Z(n720) );
  XOR U1065 ( .A(zin[65]), .B(y[66]), .Z(n718) );
  NAND U1066 ( .A(y[65]), .B(zin[64]), .Z(n717) );
  XOR U1067 ( .A(zin[64]), .B(y[65]), .Z(n715) );
  NAND U1068 ( .A(y[64]), .B(zin[63]), .Z(n714) );
  XOR U1069 ( .A(zin[63]), .B(y[64]), .Z(n712) );
  NAND U1070 ( .A(y[63]), .B(zin[62]), .Z(n711) );
  XOR U1071 ( .A(zin[62]), .B(y[63]), .Z(n709) );
  NAND U1072 ( .A(y[62]), .B(zin[61]), .Z(n708) );
  XOR U1073 ( .A(zin[61]), .B(y[62]), .Z(n706) );
  NAND U1074 ( .A(y[61]), .B(zin[60]), .Z(n705) );
  XOR U1075 ( .A(zin[60]), .B(y[61]), .Z(n703) );
  NAND U1076 ( .A(y[60]), .B(zin[59]), .Z(n702) );
  XOR U1077 ( .A(zin[59]), .B(y[60]), .Z(n700) );
  NAND U1078 ( .A(y[59]), .B(zin[58]), .Z(n699) );
  XOR U1079 ( .A(zin[58]), .B(y[59]), .Z(n697) );
  NAND U1080 ( .A(y[58]), .B(zin[57]), .Z(n696) );
  XOR U1081 ( .A(zin[57]), .B(y[58]), .Z(n694) );
  NAND U1082 ( .A(y[57]), .B(zin[56]), .Z(n693) );
  XOR U1083 ( .A(zin[56]), .B(y[57]), .Z(n691) );
  NAND U1084 ( .A(y[56]), .B(zin[55]), .Z(n690) );
  XOR U1085 ( .A(zin[55]), .B(y[56]), .Z(n688) );
  NAND U1086 ( .A(y[55]), .B(zin[54]), .Z(n687) );
  XOR U1087 ( .A(zin[54]), .B(y[55]), .Z(n685) );
  NAND U1088 ( .A(y[54]), .B(zin[53]), .Z(n684) );
  XOR U1089 ( .A(zin[53]), .B(y[54]), .Z(n682) );
  NAND U1090 ( .A(y[53]), .B(zin[52]), .Z(n681) );
  XOR U1091 ( .A(zin[52]), .B(y[53]), .Z(n679) );
  NAND U1092 ( .A(y[52]), .B(zin[51]), .Z(n678) );
  XOR U1093 ( .A(zin[51]), .B(y[52]), .Z(n676) );
  NAND U1094 ( .A(y[51]), .B(zin[50]), .Z(n675) );
  XOR U1095 ( .A(zin[50]), .B(y[51]), .Z(n673) );
  NAND U1096 ( .A(y[50]), .B(zin[49]), .Z(n672) );
  XOR U1097 ( .A(zin[49]), .B(y[50]), .Z(n670) );
  NAND U1098 ( .A(y[49]), .B(zin[48]), .Z(n669) );
  XOR U1099 ( .A(zin[48]), .B(y[49]), .Z(n667) );
  NAND U1100 ( .A(y[48]), .B(zin[47]), .Z(n666) );
  XOR U1101 ( .A(zin[47]), .B(y[48]), .Z(n664) );
  NAND U1102 ( .A(y[47]), .B(zin[46]), .Z(n663) );
  XOR U1103 ( .A(zin[46]), .B(y[47]), .Z(n661) );
  NAND U1104 ( .A(y[46]), .B(zin[45]), .Z(n660) );
  XOR U1105 ( .A(zin[45]), .B(y[46]), .Z(n658) );
  NAND U1106 ( .A(y[45]), .B(zin[44]), .Z(n657) );
  XOR U1107 ( .A(zin[44]), .B(y[45]), .Z(n655) );
  NAND U1108 ( .A(y[44]), .B(zin[43]), .Z(n654) );
  XOR U1109 ( .A(zin[43]), .B(y[44]), .Z(n652) );
  NAND U1110 ( .A(y[43]), .B(zin[42]), .Z(n651) );
  XOR U1111 ( .A(zin[42]), .B(y[43]), .Z(n649) );
  NAND U1112 ( .A(y[42]), .B(zin[41]), .Z(n648) );
  XOR U1113 ( .A(zin[41]), .B(y[42]), .Z(n646) );
  NAND U1114 ( .A(y[41]), .B(zin[40]), .Z(n645) );
  XOR U1115 ( .A(zin[40]), .B(y[41]), .Z(n643) );
  NAND U1116 ( .A(y[40]), .B(zin[39]), .Z(n642) );
  XOR U1117 ( .A(zin[39]), .B(y[40]), .Z(n640) );
  NAND U1118 ( .A(y[39]), .B(zin[38]), .Z(n639) );
  XOR U1119 ( .A(zin[38]), .B(y[39]), .Z(n637) );
  NAND U1120 ( .A(y[38]), .B(zin[37]), .Z(n636) );
  XOR U1121 ( .A(zin[37]), .B(y[38]), .Z(n634) );
  NAND U1122 ( .A(y[37]), .B(zin[36]), .Z(n633) );
  XOR U1123 ( .A(zin[36]), .B(y[37]), .Z(n631) );
  NAND U1124 ( .A(y[36]), .B(zin[35]), .Z(n630) );
  XOR U1125 ( .A(zin[35]), .B(y[36]), .Z(n628) );
  NAND U1126 ( .A(y[35]), .B(zin[34]), .Z(n627) );
  XOR U1127 ( .A(zin[34]), .B(y[35]), .Z(n625) );
  NAND U1128 ( .A(y[34]), .B(zin[33]), .Z(n624) );
  XOR U1129 ( .A(zin[33]), .B(y[34]), .Z(n622) );
  NAND U1130 ( .A(y[33]), .B(zin[32]), .Z(n621) );
  XOR U1131 ( .A(zin[32]), .B(y[33]), .Z(n619) );
  NAND U1132 ( .A(y[32]), .B(zin[31]), .Z(n618) );
  XOR U1133 ( .A(zin[31]), .B(y[32]), .Z(n616) );
  NAND U1134 ( .A(y[31]), .B(zin[30]), .Z(n615) );
  XOR U1135 ( .A(zin[30]), .B(y[31]), .Z(n613) );
  NAND U1136 ( .A(y[30]), .B(zin[29]), .Z(n612) );
  XOR U1137 ( .A(zin[29]), .B(y[30]), .Z(n610) );
  NAND U1138 ( .A(y[29]), .B(zin[28]), .Z(n609) );
  XOR U1139 ( .A(zin[28]), .B(y[29]), .Z(n607) );
  NAND U1140 ( .A(y[28]), .B(zin[27]), .Z(n606) );
  XOR U1141 ( .A(zin[27]), .B(y[28]), .Z(n604) );
  NAND U1142 ( .A(y[27]), .B(zin[26]), .Z(n603) );
  XOR U1143 ( .A(zin[26]), .B(y[27]), .Z(n601) );
  NAND U1144 ( .A(y[26]), .B(zin[25]), .Z(n600) );
  XOR U1145 ( .A(zin[25]), .B(y[26]), .Z(n598) );
  NAND U1146 ( .A(y[25]), .B(zin[24]), .Z(n597) );
  XOR U1147 ( .A(zin[24]), .B(y[25]), .Z(n595) );
  NAND U1148 ( .A(y[24]), .B(zin[23]), .Z(n594) );
  XOR U1149 ( .A(zin[23]), .B(y[24]), .Z(n592) );
  NAND U1150 ( .A(y[23]), .B(zin[22]), .Z(n591) );
  XOR U1151 ( .A(zin[22]), .B(y[23]), .Z(n589) );
  NAND U1152 ( .A(y[22]), .B(zin[21]), .Z(n588) );
  XOR U1153 ( .A(zin[21]), .B(y[22]), .Z(n586) );
  NAND U1154 ( .A(y[21]), .B(zin[20]), .Z(n585) );
  XOR U1155 ( .A(zin[20]), .B(y[21]), .Z(n583) );
  NAND U1156 ( .A(y[20]), .B(zin[19]), .Z(n582) );
  XOR U1157 ( .A(zin[19]), .B(y[20]), .Z(n580) );
  NAND U1158 ( .A(y[19]), .B(zin[18]), .Z(n579) );
  XOR U1159 ( .A(zin[18]), .B(y[19]), .Z(n577) );
  NAND U1160 ( .A(y[18]), .B(zin[17]), .Z(n576) );
  XOR U1161 ( .A(zin[17]), .B(y[18]), .Z(n574) );
  NAND U1162 ( .A(y[17]), .B(zin[16]), .Z(n573) );
  XOR U1163 ( .A(zin[16]), .B(y[17]), .Z(n571) );
  NAND U1164 ( .A(y[16]), .B(zin[15]), .Z(n570) );
  XOR U1165 ( .A(zin[15]), .B(y[16]), .Z(n568) );
  NAND U1166 ( .A(y[15]), .B(zin[14]), .Z(n567) );
  XOR U1167 ( .A(zin[14]), .B(y[15]), .Z(n565) );
  NAND U1168 ( .A(y[14]), .B(zin[13]), .Z(n564) );
  XOR U1169 ( .A(zin[13]), .B(y[14]), .Z(n562) );
  NAND U1170 ( .A(y[13]), .B(zin[12]), .Z(n561) );
  XOR U1171 ( .A(zin[12]), .B(y[13]), .Z(n559) );
  NAND U1172 ( .A(y[12]), .B(zin[11]), .Z(n558) );
  XOR U1173 ( .A(zin[11]), .B(y[12]), .Z(n556) );
  NAND U1174 ( .A(y[11]), .B(zin[10]), .Z(n555) );
  XOR U1175 ( .A(zin[10]), .B(y[11]), .Z(n553) );
  NAND U1176 ( .A(y[10]), .B(zin[9]), .Z(n552) );
  XOR U1177 ( .A(zin[9]), .B(y[10]), .Z(n550) );
  NAND U1178 ( .A(y[9]), .B(zin[8]), .Z(n549) );
  NAND U1179 ( .A(y[8]), .B(zin[7]), .Z(n546) );
  XOR U1180 ( .A(zin[7]), .B(y[8]), .Z(n544) );
  NAND U1181 ( .A(y[7]), .B(zin[6]), .Z(n543) );
  XOR U1182 ( .A(zin[6]), .B(y[7]), .Z(n541) );
  NAND U1183 ( .A(y[6]), .B(zin[5]), .Z(n540) );
  XOR U1184 ( .A(zin[5]), .B(y[6]), .Z(n538) );
  NAND U1185 ( .A(y[5]), .B(zin[4]), .Z(n537) );
  XOR U1186 ( .A(zin[4]), .B(y[5]), .Z(n535) );
  NAND U1187 ( .A(y[4]), .B(zin[3]), .Z(n534) );
  XOR U1188 ( .A(zin[3]), .B(y[4]), .Z(n532) );
  NAND U1189 ( .A(y[3]), .B(zin[2]), .Z(n531) );
  XOR U1190 ( .A(zin[2]), .B(y[3]), .Z(n529) );
  NAND U1191 ( .A(y[2]), .B(zin[1]), .Z(n528) );
  NAND U1192 ( .A(zin[0]), .B(y[1]), .Z(n2003) );
  XOR U1193 ( .A(zin[1]), .B(y[2]), .Z(n526) );
  NANDN U1194 ( .A(n2003), .B(n526), .Z(n527) );
  NAND U1195 ( .A(n528), .B(n527), .Z(n2000) );
  NAND U1196 ( .A(n529), .B(n2000), .Z(n530) );
  NAND U1197 ( .A(n531), .B(n530), .Z(n1997) );
  NAND U1198 ( .A(n532), .B(n1997), .Z(n533) );
  NAND U1199 ( .A(n534), .B(n533), .Z(n2019) );
  NAND U1200 ( .A(n535), .B(n2019), .Z(n536) );
  NAND U1201 ( .A(n537), .B(n536), .Z(n1994) );
  NAND U1202 ( .A(n538), .B(n1994), .Z(n539) );
  NAND U1203 ( .A(n540), .B(n539), .Z(n1991) );
  NAND U1204 ( .A(n541), .B(n1991), .Z(n542) );
  NAND U1205 ( .A(n543), .B(n542), .Z(n2028) );
  NAND U1206 ( .A(n544), .B(n2028), .Z(n545) );
  AND U1207 ( .A(n546), .B(n545), .Z(n2033) );
  XOR U1208 ( .A(zin[8]), .B(y[9]), .Z(n547) );
  NANDN U1209 ( .A(n2033), .B(n547), .Z(n548) );
  NAND U1210 ( .A(n549), .B(n548), .Z(n2036) );
  NAND U1211 ( .A(n550), .B(n2036), .Z(n551) );
  NAND U1212 ( .A(n552), .B(n551), .Z(n1988) );
  NAND U1213 ( .A(n553), .B(n1988), .Z(n554) );
  NAND U1214 ( .A(n555), .B(n554), .Z(n1984) );
  NAND U1215 ( .A(n556), .B(n1984), .Z(n557) );
  NAND U1216 ( .A(n558), .B(n557), .Z(n1981) );
  NAND U1217 ( .A(n559), .B(n1981), .Z(n560) );
  NAND U1218 ( .A(n561), .B(n560), .Z(n2050) );
  NAND U1219 ( .A(n562), .B(n2050), .Z(n563) );
  NAND U1220 ( .A(n564), .B(n563), .Z(n1978) );
  NAND U1221 ( .A(n565), .B(n1978), .Z(n566) );
  NAND U1222 ( .A(n567), .B(n566), .Z(n1975) );
  NAND U1223 ( .A(n568), .B(n1975), .Z(n569) );
  NAND U1224 ( .A(n570), .B(n569), .Z(n1972) );
  NAND U1225 ( .A(n571), .B(n1972), .Z(n572) );
  NAND U1226 ( .A(n573), .B(n572), .Z(n1969) );
  NAND U1227 ( .A(n574), .B(n1969), .Z(n575) );
  NAND U1228 ( .A(n576), .B(n575), .Z(n1966) );
  NAND U1229 ( .A(n577), .B(n1966), .Z(n578) );
  NAND U1230 ( .A(n579), .B(n578), .Z(n1963) );
  NAND U1231 ( .A(n580), .B(n1963), .Z(n581) );
  NAND U1232 ( .A(n582), .B(n581), .Z(n1960) );
  NAND U1233 ( .A(n583), .B(n1960), .Z(n584) );
  NAND U1234 ( .A(n585), .B(n584), .Z(n1957) );
  NAND U1235 ( .A(n586), .B(n1957), .Z(n587) );
  NAND U1236 ( .A(n588), .B(n587), .Z(n1954) );
  NAND U1237 ( .A(n589), .B(n1954), .Z(n590) );
  NAND U1238 ( .A(n591), .B(n590), .Z(n1951) );
  NAND U1239 ( .A(n592), .B(n1951), .Z(n593) );
  NAND U1240 ( .A(n594), .B(n593), .Z(n1948) );
  NAND U1241 ( .A(n595), .B(n1948), .Z(n596) );
  NAND U1242 ( .A(n597), .B(n596), .Z(n1945) );
  NAND U1243 ( .A(n598), .B(n1945), .Z(n599) );
  NAND U1244 ( .A(n600), .B(n599), .Z(n1942) );
  NAND U1245 ( .A(n601), .B(n1942), .Z(n602) );
  NAND U1246 ( .A(n603), .B(n602), .Z(n1939) );
  NAND U1247 ( .A(n604), .B(n1939), .Z(n605) );
  NAND U1248 ( .A(n606), .B(n605), .Z(n1936) );
  NAND U1249 ( .A(n607), .B(n1936), .Z(n608) );
  NAND U1250 ( .A(n609), .B(n608), .Z(n1933) );
  NAND U1251 ( .A(n610), .B(n1933), .Z(n611) );
  NAND U1252 ( .A(n612), .B(n611), .Z(n1930) );
  NAND U1253 ( .A(n613), .B(n1930), .Z(n614) );
  NAND U1254 ( .A(n615), .B(n614), .Z(n1927) );
  NAND U1255 ( .A(n616), .B(n1927), .Z(n617) );
  NAND U1256 ( .A(n618), .B(n617), .Z(n1924) );
  NAND U1257 ( .A(n619), .B(n1924), .Z(n620) );
  NAND U1258 ( .A(n621), .B(n620), .Z(n1921) );
  NAND U1259 ( .A(n622), .B(n1921), .Z(n623) );
  NAND U1260 ( .A(n624), .B(n623), .Z(n2119) );
  NAND U1261 ( .A(n625), .B(n2119), .Z(n626) );
  NAND U1262 ( .A(n627), .B(n626), .Z(n1918) );
  NAND U1263 ( .A(n628), .B(n1918), .Z(n629) );
  NAND U1264 ( .A(n630), .B(n629), .Z(n1915) );
  NAND U1265 ( .A(n631), .B(n1915), .Z(n632) );
  NAND U1266 ( .A(n633), .B(n632), .Z(n1912) );
  NAND U1267 ( .A(n634), .B(n1912), .Z(n635) );
  NAND U1268 ( .A(n636), .B(n635), .Z(n2134) );
  NAND U1269 ( .A(n637), .B(n2134), .Z(n638) );
  NAND U1270 ( .A(n639), .B(n638), .Z(n1909) );
  NAND U1271 ( .A(n640), .B(n1909), .Z(n641) );
  NAND U1272 ( .A(n642), .B(n641), .Z(n1906) );
  NAND U1273 ( .A(n643), .B(n1906), .Z(n644) );
  NAND U1274 ( .A(n645), .B(n644), .Z(n1903) );
  NAND U1275 ( .A(n646), .B(n1903), .Z(n647) );
  NAND U1276 ( .A(n648), .B(n647), .Z(n1900) );
  NAND U1277 ( .A(n649), .B(n1900), .Z(n650) );
  NAND U1278 ( .A(n651), .B(n650), .Z(n1897) );
  NAND U1279 ( .A(n652), .B(n1897), .Z(n653) );
  NAND U1280 ( .A(n654), .B(n653), .Z(n2149) );
  NAND U1281 ( .A(n655), .B(n2149), .Z(n656) );
  NAND U1282 ( .A(n657), .B(n656), .Z(n1894) );
  NAND U1283 ( .A(n658), .B(n1894), .Z(n659) );
  NAND U1284 ( .A(n660), .B(n659), .Z(n1891) );
  NAND U1285 ( .A(n661), .B(n1891), .Z(n662) );
  NAND U1286 ( .A(n663), .B(n662), .Z(n1888) );
  NAND U1287 ( .A(n664), .B(n1888), .Z(n665) );
  NAND U1288 ( .A(n666), .B(n665), .Z(n1885) );
  NAND U1289 ( .A(n667), .B(n1885), .Z(n668) );
  NAND U1290 ( .A(n669), .B(n668), .Z(n1882) );
  NAND U1291 ( .A(n670), .B(n1882), .Z(n671) );
  NAND U1292 ( .A(n672), .B(n671), .Z(n2167) );
  NAND U1293 ( .A(n673), .B(n2167), .Z(n674) );
  NAND U1294 ( .A(n675), .B(n674), .Z(n1879) );
  NAND U1295 ( .A(n676), .B(n1879), .Z(n677) );
  NAND U1296 ( .A(n678), .B(n677), .Z(n1876) );
  NAND U1297 ( .A(n679), .B(n1876), .Z(n680) );
  NAND U1298 ( .A(n681), .B(n680), .Z(n1873) );
  NAND U1299 ( .A(n682), .B(n1873), .Z(n683) );
  NAND U1300 ( .A(n684), .B(n683), .Z(n1870) );
  NAND U1301 ( .A(n685), .B(n1870), .Z(n686) );
  NAND U1302 ( .A(n687), .B(n686), .Z(n1867) );
  NAND U1303 ( .A(n688), .B(n1867), .Z(n689) );
  NAND U1304 ( .A(n690), .B(n689), .Z(n2186) );
  NAND U1305 ( .A(n691), .B(n2186), .Z(n692) );
  NAND U1306 ( .A(n693), .B(n692), .Z(n1861) );
  NAND U1307 ( .A(n694), .B(n1861), .Z(n695) );
  NAND U1308 ( .A(n696), .B(n695), .Z(n1864) );
  NAND U1309 ( .A(n697), .B(n1864), .Z(n698) );
  NAND U1310 ( .A(n699), .B(n698), .Z(n2197) );
  NAND U1311 ( .A(n700), .B(n2197), .Z(n701) );
  NAND U1312 ( .A(n702), .B(n701), .Z(n1858) );
  NAND U1313 ( .A(n703), .B(n1858), .Z(n704) );
  NAND U1314 ( .A(n705), .B(n704), .Z(n1855) );
  NAND U1315 ( .A(n706), .B(n1855), .Z(n707) );
  NAND U1316 ( .A(n708), .B(n707), .Z(n2206) );
  NAND U1317 ( .A(n709), .B(n2206), .Z(n710) );
  NAND U1318 ( .A(n711), .B(n710), .Z(n1852) );
  NAND U1319 ( .A(n712), .B(n1852), .Z(n713) );
  NAND U1320 ( .A(n714), .B(n713), .Z(n1849) );
  NAND U1321 ( .A(n715), .B(n1849), .Z(n716) );
  NAND U1322 ( .A(n717), .B(n716), .Z(n1846) );
  NAND U1323 ( .A(n718), .B(n1846), .Z(n719) );
  NAND U1324 ( .A(n720), .B(n719), .Z(n1839) );
  NAND U1325 ( .A(n721), .B(n1839), .Z(n722) );
  NAND U1326 ( .A(n723), .B(n722), .Z(n1842) );
  NAND U1327 ( .A(n724), .B(n1842), .Z(n725) );
  NAND U1328 ( .A(n726), .B(n725), .Z(n1836) );
  NAND U1329 ( .A(n727), .B(n1836), .Z(n728) );
  NAND U1330 ( .A(n729), .B(n728), .Z(n1833) );
  NAND U1331 ( .A(n730), .B(n1833), .Z(n731) );
  NAND U1332 ( .A(n732), .B(n731), .Z(n1830) );
  NAND U1333 ( .A(n733), .B(n1830), .Z(n734) );
  NAND U1334 ( .A(n735), .B(n734), .Z(n1827) );
  NAND U1335 ( .A(n736), .B(n1827), .Z(n737) );
  NAND U1336 ( .A(n738), .B(n737), .Z(n1824) );
  NAND U1337 ( .A(n739), .B(n1824), .Z(n740) );
  NAND U1338 ( .A(n741), .B(n740), .Z(n1821) );
  NAND U1339 ( .A(n742), .B(n1821), .Z(n743) );
  NAND U1340 ( .A(n744), .B(n743), .Z(n1818) );
  NAND U1341 ( .A(n745), .B(n1818), .Z(n746) );
  NAND U1342 ( .A(n747), .B(n746), .Z(n1815) );
  NAND U1343 ( .A(n748), .B(n1815), .Z(n749) );
  NAND U1344 ( .A(n750), .B(n749), .Z(n1812) );
  NAND U1345 ( .A(n751), .B(n1812), .Z(n752) );
  NAND U1346 ( .A(n753), .B(n752), .Z(n1809) );
  NAND U1347 ( .A(n754), .B(n1809), .Z(n755) );
  NAND U1348 ( .A(n756), .B(n755), .Z(n1806) );
  NAND U1349 ( .A(n757), .B(n1806), .Z(n758) );
  NAND U1350 ( .A(n759), .B(n758), .Z(n1803) );
  NAND U1351 ( .A(n760), .B(n1803), .Z(n761) );
  NAND U1352 ( .A(n762), .B(n761), .Z(n1800) );
  NAND U1353 ( .A(n763), .B(n1800), .Z(n764) );
  NAND U1354 ( .A(n765), .B(n764), .Z(n1797) );
  NAND U1355 ( .A(n766), .B(n1797), .Z(n767) );
  NAND U1356 ( .A(n768), .B(n767), .Z(n1794) );
  NAND U1357 ( .A(n769), .B(n1794), .Z(n770) );
  NAND U1358 ( .A(n771), .B(n770), .Z(n1791) );
  NAND U1359 ( .A(n772), .B(n1791), .Z(n773) );
  NAND U1360 ( .A(n774), .B(n773), .Z(n1788) );
  NAND U1361 ( .A(n775), .B(n1788), .Z(n776) );
  NAND U1362 ( .A(n777), .B(n776), .Z(n1785) );
  NAND U1363 ( .A(n778), .B(n1785), .Z(n779) );
  NAND U1364 ( .A(n780), .B(n779), .Z(n1782) );
  NAND U1365 ( .A(n781), .B(n1782), .Z(n782) );
  NAND U1366 ( .A(n783), .B(n782), .Z(n1779) );
  NAND U1367 ( .A(n784), .B(n1779), .Z(n785) );
  NAND U1368 ( .A(n786), .B(n785), .Z(n1776) );
  NAND U1369 ( .A(n787), .B(n1776), .Z(n788) );
  NAND U1370 ( .A(n789), .B(n788), .Z(n1773) );
  NAND U1371 ( .A(n790), .B(n1773), .Z(n791) );
  NAND U1372 ( .A(n792), .B(n791), .Z(n1770) );
  NAND U1373 ( .A(n793), .B(n1770), .Z(n794) );
  NAND U1374 ( .A(n795), .B(n794), .Z(n1767) );
  NAND U1375 ( .A(n796), .B(n1767), .Z(n797) );
  NAND U1376 ( .A(n798), .B(n797), .Z(n1764) );
  NAND U1377 ( .A(n799), .B(n1764), .Z(n800) );
  NAND U1378 ( .A(n801), .B(n800), .Z(n1761) );
  NAND U1379 ( .A(n802), .B(n1761), .Z(n803) );
  NAND U1380 ( .A(n804), .B(n803), .Z(n1758) );
  NAND U1381 ( .A(n805), .B(n1758), .Z(n806) );
  NAND U1382 ( .A(n807), .B(n806), .Z(n1755) );
  NAND U1383 ( .A(n808), .B(n1755), .Z(n809) );
  NAND U1384 ( .A(n810), .B(n809), .Z(n1752) );
  NAND U1385 ( .A(n811), .B(n1752), .Z(n812) );
  NAND U1386 ( .A(n813), .B(n812), .Z(n1749) );
  NAND U1387 ( .A(n814), .B(n1749), .Z(n815) );
  NAND U1388 ( .A(n816), .B(n815), .Z(n1746) );
  NAND U1389 ( .A(n817), .B(n1746), .Z(n818) );
  NAND U1390 ( .A(n819), .B(n818), .Z(n1743) );
  NAND U1391 ( .A(n820), .B(n1743), .Z(n821) );
  NAND U1392 ( .A(n822), .B(n821), .Z(n1740) );
  NAND U1393 ( .A(n823), .B(n1740), .Z(n824) );
  NAND U1394 ( .A(n825), .B(n824), .Z(n1737) );
  NAND U1395 ( .A(n826), .B(n1737), .Z(n827) );
  NAND U1396 ( .A(n828), .B(n827), .Z(n1734) );
  NAND U1397 ( .A(n829), .B(n1734), .Z(n830) );
  NAND U1398 ( .A(n831), .B(n830), .Z(n1731) );
  NAND U1399 ( .A(n832), .B(n1731), .Z(n833) );
  NAND U1400 ( .A(n834), .B(n833), .Z(n1728) );
  NAND U1401 ( .A(n835), .B(n1728), .Z(n836) );
  NAND U1402 ( .A(n837), .B(n836), .Z(n1725) );
  NAND U1403 ( .A(n838), .B(n1725), .Z(n839) );
  NAND U1404 ( .A(n840), .B(n839), .Z(n1722) );
  NAND U1405 ( .A(n841), .B(n1722), .Z(n842) );
  NAND U1406 ( .A(n843), .B(n842), .Z(n1719) );
  NAND U1407 ( .A(n844), .B(n1719), .Z(n845) );
  NAND U1408 ( .A(n846), .B(n845), .Z(n1716) );
  NAND U1409 ( .A(n847), .B(n1716), .Z(n848) );
  NAND U1410 ( .A(n849), .B(n848), .Z(n1713) );
  NAND U1411 ( .A(n850), .B(n1713), .Z(n851) );
  NAND U1412 ( .A(n852), .B(n851), .Z(n1710) );
  NAND U1413 ( .A(n853), .B(n1710), .Z(n854) );
  NAND U1414 ( .A(n855), .B(n854), .Z(n1707) );
  NAND U1415 ( .A(n856), .B(n1707), .Z(n857) );
  NAND U1416 ( .A(n858), .B(n857), .Z(n1704) );
  NAND U1417 ( .A(n859), .B(n1704), .Z(n860) );
  NAND U1418 ( .A(n861), .B(n860), .Z(n1701) );
  NAND U1419 ( .A(n862), .B(n1701), .Z(n863) );
  NAND U1420 ( .A(n864), .B(n863), .Z(n1698) );
  NAND U1421 ( .A(n865), .B(n1698), .Z(n866) );
  NAND U1422 ( .A(n867), .B(n866), .Z(n1695) );
  NAND U1423 ( .A(n868), .B(n1695), .Z(n869) );
  NAND U1424 ( .A(n870), .B(n869), .Z(n1692) );
  NAND U1425 ( .A(n871), .B(n1692), .Z(n872) );
  NAND U1426 ( .A(n873), .B(n872), .Z(n1689) );
  NAND U1427 ( .A(n874), .B(n1689), .Z(n875) );
  NAND U1428 ( .A(n876), .B(n875), .Z(n1686) );
  NAND U1429 ( .A(n877), .B(n1686), .Z(n878) );
  NAND U1430 ( .A(n879), .B(n878), .Z(n1683) );
  NAND U1431 ( .A(n880), .B(n1683), .Z(n881) );
  NAND U1432 ( .A(n882), .B(n881), .Z(n1680) );
  NAND U1433 ( .A(n883), .B(n1680), .Z(n884) );
  NAND U1434 ( .A(n885), .B(n884), .Z(n1677) );
  NAND U1435 ( .A(n886), .B(n1677), .Z(n887) );
  NAND U1436 ( .A(n888), .B(n887), .Z(n1674) );
  NAND U1437 ( .A(n889), .B(n1674), .Z(n890) );
  NAND U1438 ( .A(n891), .B(n890), .Z(n1671) );
  NAND U1439 ( .A(n892), .B(n1671), .Z(n893) );
  NAND U1440 ( .A(n894), .B(n893), .Z(n1668) );
  NAND U1441 ( .A(n895), .B(n1668), .Z(n896) );
  NAND U1442 ( .A(n897), .B(n896), .Z(n1665) );
  NAND U1443 ( .A(n898), .B(n1665), .Z(n899) );
  NAND U1444 ( .A(n900), .B(n899), .Z(n1662) );
  NAND U1445 ( .A(n901), .B(n1662), .Z(n902) );
  NAND U1446 ( .A(n903), .B(n902), .Z(n1659) );
  NAND U1447 ( .A(n904), .B(n1659), .Z(n905) );
  NAND U1448 ( .A(n906), .B(n905), .Z(n1656) );
  NAND U1449 ( .A(n907), .B(n1656), .Z(n908) );
  NAND U1450 ( .A(n909), .B(n908), .Z(n1653) );
  NAND U1451 ( .A(n910), .B(n1653), .Z(n911) );
  NAND U1452 ( .A(n912), .B(n911), .Z(n1650) );
  NAND U1453 ( .A(n913), .B(n1650), .Z(n914) );
  NAND U1454 ( .A(n915), .B(n914), .Z(n1647) );
  NAND U1455 ( .A(n916), .B(n1647), .Z(n917) );
  NAND U1456 ( .A(n918), .B(n917), .Z(n1644) );
  NAND U1457 ( .A(n919), .B(n1644), .Z(n920) );
  NAND U1458 ( .A(n921), .B(n920), .Z(n1641) );
  NAND U1459 ( .A(n922), .B(n1641), .Z(n923) );
  NAND U1460 ( .A(n924), .B(n923), .Z(n1638) );
  NAND U1461 ( .A(n925), .B(n1638), .Z(n926) );
  NAND U1462 ( .A(n927), .B(n926), .Z(n1635) );
  NAND U1463 ( .A(n928), .B(n1635), .Z(n929) );
  NAND U1464 ( .A(n930), .B(n929), .Z(n1632) );
  NAND U1465 ( .A(n931), .B(n1632), .Z(n932) );
  NAND U1466 ( .A(n933), .B(n932), .Z(n1629) );
  NAND U1467 ( .A(n934), .B(n1629), .Z(n935) );
  NAND U1468 ( .A(n936), .B(n935), .Z(n1626) );
  NAND U1469 ( .A(n937), .B(n1626), .Z(n938) );
  NAND U1470 ( .A(n939), .B(n938), .Z(n1623) );
  NAND U1471 ( .A(n940), .B(n1623), .Z(n941) );
  NAND U1472 ( .A(n942), .B(n941), .Z(n1620) );
  NAND U1473 ( .A(n943), .B(n1620), .Z(n944) );
  NAND U1474 ( .A(n945), .B(n944), .Z(n1617) );
  NAND U1475 ( .A(n946), .B(n1617), .Z(n947) );
  NAND U1476 ( .A(n948), .B(n947), .Z(n1614) );
  NAND U1477 ( .A(n949), .B(n1614), .Z(n950) );
  NAND U1478 ( .A(n951), .B(n950), .Z(n1611) );
  NAND U1479 ( .A(n952), .B(n1611), .Z(n953) );
  NAND U1480 ( .A(n954), .B(n953), .Z(n1608) );
  NAND U1481 ( .A(n955), .B(n1608), .Z(n956) );
  NAND U1482 ( .A(n957), .B(n956), .Z(n1605) );
  NAND U1483 ( .A(n958), .B(n1605), .Z(n959) );
  NAND U1484 ( .A(n960), .B(n959), .Z(n1602) );
  NAND U1485 ( .A(n961), .B(n1602), .Z(n962) );
  NAND U1486 ( .A(n963), .B(n962), .Z(n1599) );
  NAND U1487 ( .A(n964), .B(n1599), .Z(n965) );
  NAND U1488 ( .A(n966), .B(n965), .Z(n1596) );
  NAND U1489 ( .A(n967), .B(n1596), .Z(n968) );
  NAND U1490 ( .A(n969), .B(n968), .Z(n1593) );
  NAND U1491 ( .A(n970), .B(n1593), .Z(n971) );
  NAND U1492 ( .A(n972), .B(n971), .Z(n1590) );
  NAND U1493 ( .A(n973), .B(n1590), .Z(n974) );
  NAND U1494 ( .A(n975), .B(n974), .Z(n1587) );
  NAND U1495 ( .A(n976), .B(n1587), .Z(n977) );
  NAND U1496 ( .A(n978), .B(n977), .Z(n1584) );
  NAND U1497 ( .A(n979), .B(n1584), .Z(n980) );
  NAND U1498 ( .A(n981), .B(n980), .Z(n1581) );
  NAND U1499 ( .A(n982), .B(n1581), .Z(n983) );
  NAND U1500 ( .A(n984), .B(n983), .Z(n1578) );
  NAND U1501 ( .A(n985), .B(n1578), .Z(n986) );
  NAND U1502 ( .A(n987), .B(n986), .Z(n1575) );
  NAND U1503 ( .A(n988), .B(n1575), .Z(n989) );
  NAND U1504 ( .A(n990), .B(n989), .Z(n1572) );
  NAND U1505 ( .A(n991), .B(n1572), .Z(n992) );
  NAND U1506 ( .A(n993), .B(n992), .Z(n1569) );
  NAND U1507 ( .A(n994), .B(n1569), .Z(n995) );
  NAND U1508 ( .A(n996), .B(n995), .Z(n1566) );
  NAND U1509 ( .A(n997), .B(n1566), .Z(n998) );
  NAND U1510 ( .A(n999), .B(n998), .Z(n1563) );
  NAND U1511 ( .A(n1000), .B(n1563), .Z(n1001) );
  NAND U1512 ( .A(n1002), .B(n1001), .Z(n1560) );
  NAND U1513 ( .A(n1003), .B(n1560), .Z(n1004) );
  NAND U1514 ( .A(n1005), .B(n1004), .Z(n1557) );
  NAND U1515 ( .A(n1006), .B(n1557), .Z(n1007) );
  NAND U1516 ( .A(n1008), .B(n1007), .Z(n1554) );
  NAND U1517 ( .A(n1009), .B(n1554), .Z(n1010) );
  NAND U1518 ( .A(n1011), .B(n1010), .Z(n1551) );
  NAND U1519 ( .A(n1012), .B(n1551), .Z(n1013) );
  NAND U1520 ( .A(n1014), .B(n1013), .Z(n1548) );
  NAND U1521 ( .A(n1015), .B(n1548), .Z(n1016) );
  NAND U1522 ( .A(n1017), .B(n1016), .Z(n1545) );
  NAND U1523 ( .A(n1018), .B(n1545), .Z(n1019) );
  NAND U1524 ( .A(n1020), .B(n1019), .Z(n1542) );
  NAND U1525 ( .A(n1021), .B(n1542), .Z(n1022) );
  NAND U1526 ( .A(n1023), .B(n1022), .Z(n1539) );
  NAND U1527 ( .A(n1024), .B(n1539), .Z(n1025) );
  NAND U1528 ( .A(n1026), .B(n1025), .Z(n1536) );
  NAND U1529 ( .A(n1027), .B(n1536), .Z(n1028) );
  NAND U1530 ( .A(n1029), .B(n1028), .Z(n1533) );
  NAND U1531 ( .A(n1030), .B(n1533), .Z(n1031) );
  NAND U1532 ( .A(n1032), .B(n1031), .Z(n1530) );
  NAND U1533 ( .A(n1033), .B(n1530), .Z(n1034) );
  NAND U1534 ( .A(n1035), .B(n1034), .Z(n1527) );
  NAND U1535 ( .A(n1036), .B(n1527), .Z(n1037) );
  NAND U1536 ( .A(n1038), .B(n1037), .Z(n1524) );
  NAND U1537 ( .A(n1039), .B(n1524), .Z(n1040) );
  NAND U1538 ( .A(n1041), .B(n1040), .Z(n1521) );
  NAND U1539 ( .A(n1042), .B(n1521), .Z(n1043) );
  NAND U1540 ( .A(n1044), .B(n1043), .Z(n1518) );
  NAND U1541 ( .A(n1045), .B(n1518), .Z(n1046) );
  NAND U1542 ( .A(n1047), .B(n1046), .Z(n1515) );
  NAND U1543 ( .A(n1048), .B(n1515), .Z(n1049) );
  NAND U1544 ( .A(n1050), .B(n1049), .Z(n1512) );
  NAND U1545 ( .A(n1051), .B(n1512), .Z(n1052) );
  NAND U1546 ( .A(n1053), .B(n1052), .Z(n1509) );
  NAND U1547 ( .A(n1054), .B(n1509), .Z(n1055) );
  NAND U1548 ( .A(n1056), .B(n1055), .Z(n1506) );
  NAND U1549 ( .A(n1057), .B(n1506), .Z(n1058) );
  NAND U1550 ( .A(n1059), .B(n1058), .Z(n1503) );
  NAND U1551 ( .A(n1060), .B(n1503), .Z(n1061) );
  NAND U1552 ( .A(n1062), .B(n1061), .Z(n1500) );
  NAND U1553 ( .A(n1063), .B(n1500), .Z(n1064) );
  NAND U1554 ( .A(n1065), .B(n1064), .Z(n1497) );
  NAND U1555 ( .A(n1066), .B(n1497), .Z(n1067) );
  NAND U1556 ( .A(n1068), .B(n1067), .Z(n1494) );
  NAND U1557 ( .A(n1069), .B(n1494), .Z(n1070) );
  NAND U1558 ( .A(n1071), .B(n1070), .Z(n1491) );
  NAND U1559 ( .A(n1072), .B(n1491), .Z(n1073) );
  NAND U1560 ( .A(n1074), .B(n1073), .Z(n1488) );
  NAND U1561 ( .A(n1075), .B(n1488), .Z(n1076) );
  NAND U1562 ( .A(n1077), .B(n1076), .Z(n1485) );
  NAND U1563 ( .A(n1078), .B(n1485), .Z(n1079) );
  NAND U1564 ( .A(n1080), .B(n1079), .Z(n1482) );
  NAND U1565 ( .A(n1081), .B(n1482), .Z(n1082) );
  NAND U1566 ( .A(n1083), .B(n1082), .Z(n1479) );
  NAND U1567 ( .A(n1084), .B(n1479), .Z(n1085) );
  NAND U1568 ( .A(n1086), .B(n1085), .Z(n1476) );
  NAND U1569 ( .A(n1087), .B(n1476), .Z(n1088) );
  NAND U1570 ( .A(n1089), .B(n1088), .Z(n1473) );
  NAND U1571 ( .A(n1090), .B(n1473), .Z(n1091) );
  NAND U1572 ( .A(n1092), .B(n1091), .Z(n1470) );
  NAND U1573 ( .A(n1093), .B(n1470), .Z(n1094) );
  NAND U1574 ( .A(n1095), .B(n1094), .Z(n1467) );
  NAND U1575 ( .A(n1096), .B(n1467), .Z(n1097) );
  NAND U1576 ( .A(n1098), .B(n1097), .Z(n1464) );
  NAND U1577 ( .A(n1099), .B(n1464), .Z(n1100) );
  NAND U1578 ( .A(n1101), .B(n1100), .Z(n1461) );
  NAND U1579 ( .A(n1102), .B(n1461), .Z(n1103) );
  NAND U1580 ( .A(n1104), .B(n1103), .Z(n1458) );
  NAND U1581 ( .A(n1105), .B(n1458), .Z(n1106) );
  NAND U1582 ( .A(n1107), .B(n1106), .Z(n1455) );
  NAND U1583 ( .A(n1108), .B(n1455), .Z(n1109) );
  NAND U1584 ( .A(n1110), .B(n1109), .Z(n1452) );
  NAND U1585 ( .A(n1111), .B(n1452), .Z(n1112) );
  NAND U1586 ( .A(n1113), .B(n1112), .Z(n1449) );
  NAND U1587 ( .A(n1114), .B(n1449), .Z(n1115) );
  NAND U1588 ( .A(n1116), .B(n1115), .Z(n1446) );
  NAND U1589 ( .A(n1117), .B(n1446), .Z(n1118) );
  NAND U1590 ( .A(n1119), .B(n1118), .Z(n1443) );
  NAND U1591 ( .A(n1120), .B(n1443), .Z(n1121) );
  NAND U1592 ( .A(n1122), .B(n1121), .Z(n1440) );
  NAND U1593 ( .A(n1123), .B(n1440), .Z(n1124) );
  NAND U1594 ( .A(n1125), .B(n1124), .Z(n1437) );
  NAND U1595 ( .A(n1126), .B(n1437), .Z(n1127) );
  NAND U1596 ( .A(n1128), .B(n1127), .Z(n1434) );
  NAND U1597 ( .A(n1129), .B(n1434), .Z(n1130) );
  NAND U1598 ( .A(n1131), .B(n1130), .Z(n1431) );
  NAND U1599 ( .A(n1132), .B(n1431), .Z(n1133) );
  NAND U1600 ( .A(n1134), .B(n1133), .Z(n1428) );
  NAND U1601 ( .A(n1135), .B(n1428), .Z(n1136) );
  NAND U1602 ( .A(n1137), .B(n1136), .Z(n1425) );
  NAND U1603 ( .A(n1138), .B(n1425), .Z(n1139) );
  NAND U1604 ( .A(n1140), .B(n1139), .Z(n1422) );
  NAND U1605 ( .A(n1141), .B(n1422), .Z(n1142) );
  NAND U1606 ( .A(n1143), .B(n1142), .Z(n1419) );
  NAND U1607 ( .A(n1144), .B(n1419), .Z(n1145) );
  NAND U1608 ( .A(n1146), .B(n1145), .Z(n1416) );
  NAND U1609 ( .A(n1147), .B(n1416), .Z(n1148) );
  NAND U1610 ( .A(n1149), .B(n1148), .Z(n1413) );
  NAND U1611 ( .A(n1150), .B(n1413), .Z(n1151) );
  NAND U1612 ( .A(n1152), .B(n1151), .Z(n1410) );
  NAND U1613 ( .A(n1153), .B(n1410), .Z(n1154) );
  NAND U1614 ( .A(n1155), .B(n1154), .Z(n1407) );
  NAND U1615 ( .A(n1156), .B(n1407), .Z(n1157) );
  NAND U1616 ( .A(n1158), .B(n1157), .Z(n1404) );
  NAND U1617 ( .A(n1159), .B(n1404), .Z(n1160) );
  NAND U1618 ( .A(n1161), .B(n1160), .Z(n1401) );
  NAND U1619 ( .A(n1162), .B(n1401), .Z(n1163) );
  NAND U1620 ( .A(n1164), .B(n1163), .Z(n1398) );
  NAND U1621 ( .A(n1165), .B(n1398), .Z(n1166) );
  NAND U1622 ( .A(n1167), .B(n1166), .Z(n1395) );
  NAND U1623 ( .A(n1168), .B(n1395), .Z(n1169) );
  NAND U1624 ( .A(n1170), .B(n1169), .Z(n1392) );
  NAND U1625 ( .A(n1171), .B(n1392), .Z(n1172) );
  NAND U1626 ( .A(n1173), .B(n1172), .Z(n1389) );
  NAND U1627 ( .A(n1174), .B(n1389), .Z(n1175) );
  NAND U1628 ( .A(n1176), .B(n1175), .Z(n1386) );
  NAND U1629 ( .A(n1177), .B(n1386), .Z(n1178) );
  NAND U1630 ( .A(n1179), .B(n1178), .Z(n1383) );
  NAND U1631 ( .A(n1180), .B(n1383), .Z(n1181) );
  NAND U1632 ( .A(n1182), .B(n1181), .Z(n1380) );
  NAND U1633 ( .A(n1183), .B(n1380), .Z(n1184) );
  NAND U1634 ( .A(n1185), .B(n1184), .Z(n1377) );
  NAND U1635 ( .A(n1186), .B(n1377), .Z(n1187) );
  NAND U1636 ( .A(n1188), .B(n1187), .Z(n1374) );
  NAND U1637 ( .A(n1189), .B(n1374), .Z(n1190) );
  NAND U1638 ( .A(n1191), .B(n1190), .Z(n1371) );
  NAND U1639 ( .A(n1192), .B(n1371), .Z(n1193) );
  NAND U1640 ( .A(n1194), .B(n1193), .Z(n1368) );
  NAND U1641 ( .A(n1195), .B(n1368), .Z(n1196) );
  NAND U1642 ( .A(n1197), .B(n1196), .Z(n1365) );
  NAND U1643 ( .A(n1198), .B(n1365), .Z(n1199) );
  NAND U1644 ( .A(n1200), .B(n1199), .Z(n1362) );
  NAND U1645 ( .A(n1201), .B(n1362), .Z(n1202) );
  NAND U1646 ( .A(n1203), .B(n1202), .Z(n1359) );
  NAND U1647 ( .A(n1204), .B(n1359), .Z(n1205) );
  NAND U1648 ( .A(n1206), .B(n1205), .Z(n1356) );
  NAND U1649 ( .A(n1207), .B(n1356), .Z(n1208) );
  NAND U1650 ( .A(n1209), .B(n1208), .Z(n1353) );
  NAND U1651 ( .A(n1210), .B(n1353), .Z(n1211) );
  NAND U1652 ( .A(n1212), .B(n1211), .Z(n1350) );
  NAND U1653 ( .A(n1213), .B(n1350), .Z(n1214) );
  NAND U1654 ( .A(n1215), .B(n1214), .Z(n1347) );
  NAND U1655 ( .A(n1216), .B(n1347), .Z(n1217) );
  NAND U1656 ( .A(n1218), .B(n1217), .Z(n1344) );
  NAND U1657 ( .A(n1219), .B(n1344), .Z(n1220) );
  NAND U1658 ( .A(n1221), .B(n1220), .Z(n1341) );
  NAND U1659 ( .A(n1222), .B(n1341), .Z(n1223) );
  NAND U1660 ( .A(n1224), .B(n1223), .Z(n1338) );
  NAND U1661 ( .A(n1225), .B(n1338), .Z(n1226) );
  NAND U1662 ( .A(n1227), .B(n1226), .Z(n1335) );
  NAND U1663 ( .A(n1228), .B(n1335), .Z(n1229) );
  NAND U1664 ( .A(n1230), .B(n1229), .Z(n1332) );
  NAND U1665 ( .A(n1231), .B(n1332), .Z(n1232) );
  NAND U1666 ( .A(n1233), .B(n1232), .Z(n1329) );
  NAND U1667 ( .A(n1234), .B(n1329), .Z(n1235) );
  NAND U1668 ( .A(n1236), .B(n1235), .Z(n1326) );
  NAND U1669 ( .A(n1237), .B(n1326), .Z(n1238) );
  NAND U1670 ( .A(n1239), .B(n1238), .Z(n1323) );
  NAND U1671 ( .A(n1240), .B(n1323), .Z(n1241) );
  NAND U1672 ( .A(n1242), .B(n1241), .Z(n1320) );
  NAND U1673 ( .A(n1243), .B(n1320), .Z(n1244) );
  NAND U1674 ( .A(n1245), .B(n1244), .Z(n1317) );
  NAND U1675 ( .A(n1246), .B(n1317), .Z(n1247) );
  NAND U1676 ( .A(n1248), .B(n1247), .Z(n1314) );
  NAND U1677 ( .A(n1249), .B(n1314), .Z(n1250) );
  NAND U1678 ( .A(n1251), .B(n1250), .Z(n1311) );
  NAND U1679 ( .A(n1252), .B(n1311), .Z(n1253) );
  NAND U1680 ( .A(n1254), .B(n1253), .Z(n1308) );
  NAND U1681 ( .A(n1255), .B(n1308), .Z(n1256) );
  NAND U1682 ( .A(n1257), .B(n1256), .Z(n1305) );
  NAND U1683 ( .A(n1258), .B(n1305), .Z(n1259) );
  NAND U1684 ( .A(n1260), .B(n1259), .Z(n1302) );
  NAND U1685 ( .A(n1261), .B(n1302), .Z(n1262) );
  NAND U1686 ( .A(n1263), .B(n1262), .Z(n1299) );
  NAND U1687 ( .A(n1264), .B(n1299), .Z(n1265) );
  NAND U1688 ( .A(n1266), .B(n1265), .Z(n1296) );
  NAND U1689 ( .A(n1267), .B(n1296), .Z(n1268) );
  NAND U1690 ( .A(n1269), .B(n1268), .Z(n1293) );
  NAND U1691 ( .A(n1270), .B(n1293), .Z(n1271) );
  NAND U1692 ( .A(n1272), .B(n1271), .Z(n1290) );
  NAND U1693 ( .A(n1273), .B(n1290), .Z(n1274) );
  NAND U1694 ( .A(n1275), .B(n1274), .Z(n1287) );
  NAND U1695 ( .A(n1276), .B(n1287), .Z(n1277) );
  NAND U1696 ( .A(n1278), .B(n1277), .Z(n1284) );
  NAND U1697 ( .A(n1279), .B(n1284), .Z(n1280) );
  NAND U1698 ( .A(n1281), .B(n1280), .Z(n2857) );
  XOR U1699 ( .A(y[254]), .B(n2857), .Z(n1282) );
  IV U1700 ( .A(xregN_1), .Z(n2868) );
  ANDN U1701 ( .B(n1282), .A(n2868), .Z(n1283) );
  XNOR U1702 ( .A(zin[253]), .B(n1283), .Z(n3318) );
  NANDN U1703 ( .A(n6582), .B(n3318), .Z(n3303) );
  XOR U1704 ( .A(y[253]), .B(n1284), .Z(n1285) );
  ANDN U1705 ( .B(n1285), .A(n2868), .Z(n1286) );
  XNOR U1706 ( .A(zin[252]), .B(n1286), .Z(n3322) );
  IV U1707 ( .A(n[252]), .Z(n3327) );
  XOR U1708 ( .A(y[252]), .B(n1287), .Z(n1288) );
  ANDN U1709 ( .B(n1288), .A(n2868), .Z(n1289) );
  XNOR U1710 ( .A(zin[251]), .B(n1289), .Z(n3326) );
  NANDN U1711 ( .A(n3327), .B(n3326), .Z(n3300) );
  XOR U1712 ( .A(y[251]), .B(n1290), .Z(n1291) );
  ANDN U1713 ( .B(n1291), .A(n2868), .Z(n1292) );
  XNOR U1714 ( .A(zin[250]), .B(n1292), .Z(n3331) );
  XOR U1715 ( .A(n3331), .B(n[251]), .Z(n2856) );
  XOR U1716 ( .A(y[250]), .B(n1293), .Z(n1294) );
  ANDN U1717 ( .B(n1294), .A(n2868), .Z(n1295) );
  XNOR U1718 ( .A(zin[249]), .B(n1295), .Z(n3335) );
  NAND U1719 ( .A(n3335), .B(n[250]), .Z(n2854) );
  XOR U1720 ( .A(n[250]), .B(n3335), .Z(n2852) );
  IV U1721 ( .A(n[249]), .Z(n6534) );
  XOR U1722 ( .A(y[249]), .B(n1296), .Z(n1297) );
  ANDN U1723 ( .B(n1297), .A(n2868), .Z(n1298) );
  XNOR U1724 ( .A(zin[248]), .B(n1298), .Z(n3339) );
  NANDN U1725 ( .A(n6534), .B(n3339), .Z(n3297) );
  XNOR U1726 ( .A(n6534), .B(n3339), .Z(n2849) );
  XOR U1727 ( .A(y[248]), .B(n1299), .Z(n1300) );
  ANDN U1728 ( .B(n1300), .A(n2868), .Z(n1301) );
  XNOR U1729 ( .A(zin[247]), .B(n1301), .Z(n3343) );
  NAND U1730 ( .A(n3343), .B(n[248]), .Z(n2847) );
  XOR U1731 ( .A(n[248]), .B(n3343), .Z(n2845) );
  IV U1732 ( .A(n[247]), .Z(n3348) );
  XOR U1733 ( .A(y[247]), .B(n1302), .Z(n1303) );
  ANDN U1734 ( .B(n1303), .A(n2868), .Z(n1304) );
  XNOR U1735 ( .A(zin[246]), .B(n1304), .Z(n3347) );
  NANDN U1736 ( .A(n3348), .B(n3347), .Z(n3294) );
  XNOR U1737 ( .A(n3348), .B(n3347), .Z(n2842) );
  IV U1738 ( .A(n[246]), .Z(n6514) );
  XOR U1739 ( .A(y[246]), .B(n1305), .Z(n1306) );
  ANDN U1740 ( .B(n1306), .A(n2868), .Z(n1307) );
  XNOR U1741 ( .A(zin[245]), .B(n1307), .Z(n3352) );
  NANDN U1742 ( .A(n6514), .B(n3352), .Z(n3291) );
  XNOR U1743 ( .A(n3352), .B(n6514), .Z(n2839) );
  XOR U1744 ( .A(y[245]), .B(n1308), .Z(n1309) );
  ANDN U1745 ( .B(n1309), .A(n2868), .Z(n1310) );
  XNOR U1746 ( .A(zin[244]), .B(n1310), .Z(n3356) );
  NAND U1747 ( .A(n[245]), .B(n3356), .Z(n3288) );
  XOR U1748 ( .A(n[245]), .B(n3356), .Z(n2836) );
  IV U1749 ( .A(n[244]), .Z(n3361) );
  XOR U1750 ( .A(y[244]), .B(n1311), .Z(n1312) );
  ANDN U1751 ( .B(n1312), .A(n2868), .Z(n1313) );
  XNOR U1752 ( .A(zin[243]), .B(n1313), .Z(n3360) );
  NANDN U1753 ( .A(n3361), .B(n3360), .Z(n3285) );
  XNOR U1754 ( .A(n3360), .B(n3361), .Z(n2833) );
  XOR U1755 ( .A(y[243]), .B(n1314), .Z(n1315) );
  ANDN U1756 ( .B(n1315), .A(n2868), .Z(n1316) );
  XNOR U1757 ( .A(zin[242]), .B(n1316), .Z(n3365) );
  NAND U1758 ( .A(n[243]), .B(n3365), .Z(n2831) );
  XOR U1759 ( .A(n3365), .B(n[243]), .Z(n2829) );
  XOR U1760 ( .A(y[242]), .B(n1317), .Z(n1318) );
  ANDN U1761 ( .B(n1318), .A(n2868), .Z(n1319) );
  XNOR U1762 ( .A(zin[241]), .B(n1319), .Z(n3369) );
  NAND U1763 ( .A(n3369), .B(n[242]), .Z(n2827) );
  XOR U1764 ( .A(n[242]), .B(n3369), .Z(n2825) );
  XOR U1765 ( .A(y[241]), .B(n1320), .Z(n1321) );
  ANDN U1766 ( .B(n1321), .A(n2868), .Z(n1322) );
  XNOR U1767 ( .A(zin[240]), .B(n1322), .Z(n3373) );
  NAND U1768 ( .A(n[241]), .B(n3373), .Z(n2823) );
  XOR U1769 ( .A(n3373), .B(n[241]), .Z(n2821) );
  XOR U1770 ( .A(y[240]), .B(n1323), .Z(n1324) );
  ANDN U1771 ( .B(n1324), .A(n2868), .Z(n1325) );
  XNOR U1772 ( .A(zin[239]), .B(n1325), .Z(n3377) );
  NAND U1773 ( .A(n3377), .B(n[240]), .Z(n2819) );
  XOR U1774 ( .A(n[240]), .B(n3377), .Z(n2817) );
  IV U1775 ( .A(n[239]), .Z(n3382) );
  XOR U1776 ( .A(y[239]), .B(n1326), .Z(n1327) );
  ANDN U1777 ( .B(n1327), .A(n2868), .Z(n1328) );
  XNOR U1778 ( .A(zin[238]), .B(n1328), .Z(n3381) );
  NANDN U1779 ( .A(n3382), .B(n3381), .Z(n3282) );
  XNOR U1780 ( .A(n3382), .B(n3381), .Z(n2814) );
  XOR U1781 ( .A(y[238]), .B(n1329), .Z(n1330) );
  ANDN U1782 ( .B(n1330), .A(n2868), .Z(n1331) );
  XNOR U1783 ( .A(zin[237]), .B(n1331), .Z(n3386) );
  NAND U1784 ( .A(n3386), .B(n[238]), .Z(n2812) );
  XOR U1785 ( .A(n[238]), .B(n3386), .Z(n2810) );
  IV U1786 ( .A(n[237]), .Z(n6456) );
  XOR U1787 ( .A(y[237]), .B(n1332), .Z(n1333) );
  ANDN U1788 ( .B(n1333), .A(n2868), .Z(n1334) );
  XNOR U1789 ( .A(zin[236]), .B(n1334), .Z(n5260) );
  NANDN U1790 ( .A(n6456), .B(n5260), .Z(n2808) );
  XNOR U1791 ( .A(n5260), .B(n6456), .Z(n2806) );
  IV U1792 ( .A(n[236]), .Z(n6449) );
  XOR U1793 ( .A(y[236]), .B(n1335), .Z(n1336) );
  ANDN U1794 ( .B(n1336), .A(n2868), .Z(n1337) );
  XNOR U1795 ( .A(zin[235]), .B(n1337), .Z(n3390) );
  NANDN U1796 ( .A(n6449), .B(n3390), .Z(n2804) );
  XNOR U1797 ( .A(n6449), .B(n3390), .Z(n2802) );
  XOR U1798 ( .A(y[235]), .B(n1338), .Z(n1339) );
  ANDN U1799 ( .B(n1339), .A(n2868), .Z(n1340) );
  XNOR U1800 ( .A(zin[234]), .B(n1340), .Z(n3394) );
  NAND U1801 ( .A(n[235]), .B(n3394), .Z(n2800) );
  XOR U1802 ( .A(n3394), .B(n[235]), .Z(n2798) );
  IV U1803 ( .A(n[234]), .Z(n3399) );
  XOR U1804 ( .A(y[234]), .B(n1341), .Z(n1342) );
  ANDN U1805 ( .B(n1342), .A(n2868), .Z(n1343) );
  XOR U1806 ( .A(zin[233]), .B(n1343), .Z(n3398) );
  IV U1807 ( .A(n3398), .Z(n2872) );
  NANDN U1808 ( .A(n3399), .B(n2872), .Z(n2796) );
  XNOR U1809 ( .A(n3398), .B(n[234]), .Z(n2794) );
  XOR U1810 ( .A(y[233]), .B(n1344), .Z(n1345) );
  ANDN U1811 ( .B(n1345), .A(n2868), .Z(n1346) );
  XNOR U1812 ( .A(zin[232]), .B(n1346), .Z(n3403) );
  NAND U1813 ( .A(n[233]), .B(n3403), .Z(n2792) );
  XOR U1814 ( .A(n3403), .B(n[233]), .Z(n2790) );
  XOR U1815 ( .A(y[232]), .B(n1347), .Z(n1348) );
  ANDN U1816 ( .B(n1348), .A(n2868), .Z(n1349) );
  XNOR U1817 ( .A(zin[231]), .B(n1349), .Z(n3407) );
  NAND U1818 ( .A(n3407), .B(n[232]), .Z(n2788) );
  XOR U1819 ( .A(n[232]), .B(n3407), .Z(n2786) );
  IV U1820 ( .A(n[231]), .Z(n6413) );
  XOR U1821 ( .A(y[231]), .B(n1350), .Z(n1351) );
  ANDN U1822 ( .B(n1351), .A(n2868), .Z(n1352) );
  XNOR U1823 ( .A(zin[230]), .B(n1352), .Z(n3411) );
  NANDN U1824 ( .A(n6413), .B(n3411), .Z(n3279) );
  XNOR U1825 ( .A(n6413), .B(n3411), .Z(n2783) );
  XOR U1826 ( .A(y[230]), .B(n1353), .Z(n1354) );
  ANDN U1827 ( .B(n1354), .A(n2868), .Z(n1355) );
  XNOR U1828 ( .A(zin[229]), .B(n1355), .Z(n5233) );
  NAND U1829 ( .A(n5233), .B(n[230]), .Z(n2781) );
  XOR U1830 ( .A(n[230]), .B(n5233), .Z(n2779) );
  XOR U1831 ( .A(y[229]), .B(n1356), .Z(n1357) );
  ANDN U1832 ( .B(n1357), .A(n2868), .Z(n1358) );
  XNOR U1833 ( .A(zin[228]), .B(n1358), .Z(n3415) );
  NAND U1834 ( .A(n[229]), .B(n3415), .Z(n2777) );
  XOR U1835 ( .A(n3415), .B(n[229]), .Z(n2775) );
  XOR U1836 ( .A(y[228]), .B(n1359), .Z(n1360) );
  ANDN U1837 ( .B(n1360), .A(n2868), .Z(n1361) );
  XOR U1838 ( .A(zin[227]), .B(n1361), .Z(n2873) );
  NANDN U1839 ( .A(n2873), .B(n[228]), .Z(n2773) );
  XNOR U1840 ( .A(n[228]), .B(n2873), .Z(n2771) );
  XOR U1841 ( .A(y[227]), .B(n1362), .Z(n1363) );
  ANDN U1842 ( .B(n1363), .A(n2868), .Z(n1364) );
  XNOR U1843 ( .A(zin[226]), .B(n1364), .Z(n3423) );
  NAND U1844 ( .A(n[227]), .B(n3423), .Z(n2769) );
  XOR U1845 ( .A(n3423), .B(n[227]), .Z(n2767) );
  XOR U1846 ( .A(y[226]), .B(n1365), .Z(n1366) );
  ANDN U1847 ( .B(n1366), .A(n2868), .Z(n1367) );
  XNOR U1848 ( .A(zin[225]), .B(n1367), .Z(n3427) );
  NAND U1849 ( .A(n3427), .B(n[226]), .Z(n2765) );
  XOR U1850 ( .A(n[226]), .B(n3427), .Z(n2763) );
  IV U1851 ( .A(n[225]), .Z(n6376) );
  XOR U1852 ( .A(y[225]), .B(n1368), .Z(n1369) );
  ANDN U1853 ( .B(n1369), .A(n2868), .Z(n1370) );
  XNOR U1854 ( .A(zin[224]), .B(n1370), .Z(n3431) );
  NANDN U1855 ( .A(n6376), .B(n3431), .Z(n3273) );
  XNOR U1856 ( .A(n6376), .B(n3431), .Z(n2760) );
  XOR U1857 ( .A(y[224]), .B(n1371), .Z(n1372) );
  ANDN U1858 ( .B(n1372), .A(n2868), .Z(n1373) );
  XNOR U1859 ( .A(zin[223]), .B(n1373), .Z(n3435) );
  NAND U1860 ( .A(n3435), .B(n[224]), .Z(n2758) );
  XOR U1861 ( .A(n[224]), .B(n3435), .Z(n2756) );
  XOR U1862 ( .A(y[223]), .B(n1374), .Z(n1375) );
  ANDN U1863 ( .B(n1375), .A(n2868), .Z(n1376) );
  XNOR U1864 ( .A(zin[222]), .B(n1376), .Z(n3439) );
  NAND U1865 ( .A(n[223]), .B(n3439), .Z(n2754) );
  XOR U1866 ( .A(n3439), .B(n[223]), .Z(n2752) );
  IV U1867 ( .A(n[222]), .Z(n6357) );
  XOR U1868 ( .A(y[222]), .B(n1377), .Z(n1378) );
  ANDN U1869 ( .B(n1378), .A(n2868), .Z(n1379) );
  XNOR U1870 ( .A(zin[221]), .B(n1379), .Z(n3443) );
  NANDN U1871 ( .A(n6357), .B(n3443), .Z(n3270) );
  XNOR U1872 ( .A(n3443), .B(n6357), .Z(n2749) );
  XOR U1873 ( .A(y[221]), .B(n1380), .Z(n1381) );
  ANDN U1874 ( .B(n1381), .A(n2868), .Z(n1382) );
  XNOR U1875 ( .A(zin[220]), .B(n1382), .Z(n3447) );
  NAND U1876 ( .A(n[221]), .B(n3447), .Z(n2747) );
  XOR U1877 ( .A(n3447), .B(n[221]), .Z(n2745) );
  XOR U1878 ( .A(y[220]), .B(n1383), .Z(n1384) );
  ANDN U1879 ( .B(n1384), .A(n2868), .Z(n1385) );
  XNOR U1880 ( .A(zin[219]), .B(n1385), .Z(n3451) );
  NAND U1881 ( .A(n3451), .B(n[220]), .Z(n2743) );
  XOR U1882 ( .A(n[220]), .B(n3451), .Z(n2741) );
  XOR U1883 ( .A(y[219]), .B(n1386), .Z(n1387) );
  ANDN U1884 ( .B(n1387), .A(n2868), .Z(n1388) );
  XNOR U1885 ( .A(zin[218]), .B(n1388), .Z(n3455) );
  NAND U1886 ( .A(n[219]), .B(n3455), .Z(n2739) );
  XOR U1887 ( .A(n3455), .B(n[219]), .Z(n2737) );
  IV U1888 ( .A(n[218]), .Z(n6317) );
  XOR U1889 ( .A(y[218]), .B(n1389), .Z(n1390) );
  ANDN U1890 ( .B(n1390), .A(n2868), .Z(n1391) );
  XNOR U1891 ( .A(zin[217]), .B(n1391), .Z(n3459) );
  NANDN U1892 ( .A(n6317), .B(n3459), .Z(n3267) );
  XNOR U1893 ( .A(n3459), .B(n6317), .Z(n2734) );
  XOR U1894 ( .A(y[217]), .B(n1392), .Z(n1393) );
  ANDN U1895 ( .B(n1393), .A(n2868), .Z(n1394) );
  XNOR U1896 ( .A(zin[216]), .B(n1394), .Z(n5178) );
  NAND U1897 ( .A(n[217]), .B(n5178), .Z(n2732) );
  XOR U1898 ( .A(n5178), .B(n[217]), .Z(n2730) );
  XOR U1899 ( .A(y[216]), .B(n1395), .Z(n1396) );
  ANDN U1900 ( .B(n1396), .A(n2868), .Z(n1397) );
  XNOR U1901 ( .A(zin[215]), .B(n1397), .Z(n3463) );
  NAND U1902 ( .A(n3463), .B(n[216]), .Z(n2728) );
  XOR U1903 ( .A(n[216]), .B(n3463), .Z(n2726) );
  XOR U1904 ( .A(y[215]), .B(n1398), .Z(n1399) );
  ANDN U1905 ( .B(n1399), .A(n2868), .Z(n1400) );
  XNOR U1906 ( .A(zin[214]), .B(n1400), .Z(n3467) );
  NAND U1907 ( .A(n[215]), .B(n3467), .Z(n2724) );
  XOR U1908 ( .A(n3467), .B(n[215]), .Z(n2722) );
  XOR U1909 ( .A(y[214]), .B(n1401), .Z(n1402) );
  ANDN U1910 ( .B(n1402), .A(n2868), .Z(n1403) );
  XNOR U1911 ( .A(zin[213]), .B(n1403), .Z(n3471) );
  NAND U1912 ( .A(n3471), .B(n[214]), .Z(n2720) );
  XOR U1913 ( .A(n[214]), .B(n3471), .Z(n2718) );
  IV U1914 ( .A(n[213]), .Z(n3476) );
  XOR U1915 ( .A(y[213]), .B(n1404), .Z(n1405) );
  ANDN U1916 ( .B(n1405), .A(n2868), .Z(n1406) );
  XNOR U1917 ( .A(zin[212]), .B(n1406), .Z(n3475) );
  NANDN U1918 ( .A(n3476), .B(n3475), .Z(n3264) );
  XNOR U1919 ( .A(n3476), .B(n3475), .Z(n2715) );
  XOR U1920 ( .A(y[212]), .B(n1407), .Z(n1408) );
  ANDN U1921 ( .B(n1408), .A(n2868), .Z(n1409) );
  XNOR U1922 ( .A(zin[211]), .B(n1409), .Z(n3480) );
  NAND U1923 ( .A(n3480), .B(n[212]), .Z(n2713) );
  XOR U1924 ( .A(n[212]), .B(n3480), .Z(n2711) );
  XOR U1925 ( .A(y[211]), .B(n1410), .Z(n1411) );
  ANDN U1926 ( .B(n1411), .A(n2868), .Z(n1412) );
  XNOR U1927 ( .A(zin[210]), .B(n1412), .Z(n3484) );
  NAND U1928 ( .A(n[211]), .B(n3484), .Z(n2709) );
  XOR U1929 ( .A(n3484), .B(n[211]), .Z(n2707) );
  XOR U1930 ( .A(y[210]), .B(n1413), .Z(n1414) );
  ANDN U1931 ( .B(n1414), .A(n2868), .Z(n1415) );
  XOR U1932 ( .A(zin[209]), .B(n1415), .Z(n3488) );
  NANDN U1933 ( .A(n3488), .B(n[210]), .Z(n2705) );
  IV U1934 ( .A(n[210]), .Z(n6268) );
  IV U1935 ( .A(n3488), .Z(n2874) );
  XNOR U1936 ( .A(n6268), .B(n2874), .Z(n2703) );
  IV U1937 ( .A(n[209]), .Z(n6256) );
  XOR U1938 ( .A(y[209]), .B(n1416), .Z(n1417) );
  ANDN U1939 ( .B(n1417), .A(n2868), .Z(n1418) );
  XNOR U1940 ( .A(zin[208]), .B(n1418), .Z(n3492) );
  NANDN U1941 ( .A(n6256), .B(n3492), .Z(n2701) );
  XNOR U1942 ( .A(n3492), .B(n6256), .Z(n2699) );
  IV U1943 ( .A(n[208]), .Z(n3499) );
  XOR U1944 ( .A(y[208]), .B(n1419), .Z(n1420) );
  ANDN U1945 ( .B(n1420), .A(n2868), .Z(n1421) );
  XNOR U1946 ( .A(zin[207]), .B(n1421), .Z(n3498) );
  NANDN U1947 ( .A(n3499), .B(n3498), .Z(n3261) );
  XNOR U1948 ( .A(n3498), .B(n3499), .Z(n2696) );
  XOR U1949 ( .A(y[207]), .B(n1422), .Z(n1423) );
  ANDN U1950 ( .B(n1423), .A(n2868), .Z(n1424) );
  XNOR U1951 ( .A(zin[206]), .B(n1424), .Z(n3503) );
  NAND U1952 ( .A(n[207]), .B(n3503), .Z(n2694) );
  XOR U1953 ( .A(n3503), .B(n[207]), .Z(n2692) );
  IV U1954 ( .A(n[206]), .Z(n3508) );
  XOR U1955 ( .A(y[206]), .B(n1425), .Z(n1426) );
  ANDN U1956 ( .B(n1426), .A(n2868), .Z(n1427) );
  XNOR U1957 ( .A(zin[205]), .B(n1427), .Z(n3507) );
  NANDN U1958 ( .A(n3508), .B(n3507), .Z(n3258) );
  XNOR U1959 ( .A(n3507), .B(n3508), .Z(n2689) );
  XOR U1960 ( .A(y[205]), .B(n1428), .Z(n1429) );
  ANDN U1961 ( .B(n1429), .A(n2868), .Z(n1430) );
  XNOR U1962 ( .A(zin[204]), .B(n1430), .Z(n3512) );
  NAND U1963 ( .A(n[205]), .B(n3512), .Z(n2687) );
  XOR U1964 ( .A(n3512), .B(n[205]), .Z(n2685) );
  XOR U1965 ( .A(y[204]), .B(n1431), .Z(n1432) );
  ANDN U1966 ( .B(n1432), .A(n2868), .Z(n1433) );
  XNOR U1967 ( .A(zin[203]), .B(n1433), .Z(n3516) );
  NAND U1968 ( .A(n3516), .B(n[204]), .Z(n2683) );
  XOR U1969 ( .A(n[204]), .B(n3516), .Z(n2681) );
  IV U1970 ( .A(n[203]), .Z(n6225) );
  XOR U1971 ( .A(y[203]), .B(n1434), .Z(n1435) );
  ANDN U1972 ( .B(n1435), .A(n2868), .Z(n1436) );
  XNOR U1973 ( .A(zin[202]), .B(n1436), .Z(n3520) );
  NANDN U1974 ( .A(n6225), .B(n3520), .Z(n3255) );
  XNOR U1975 ( .A(n6225), .B(n3520), .Z(n2678) );
  XOR U1976 ( .A(y[202]), .B(n1437), .Z(n1438) );
  ANDN U1977 ( .B(n1438), .A(n2868), .Z(n1439) );
  XNOR U1978 ( .A(zin[201]), .B(n1439), .Z(n3524) );
  NAND U1979 ( .A(n3524), .B(n[202]), .Z(n2676) );
  XOR U1980 ( .A(n[202]), .B(n3524), .Z(n2674) );
  IV U1981 ( .A(n[201]), .Z(n3529) );
  XOR U1982 ( .A(y[201]), .B(n1440), .Z(n1441) );
  ANDN U1983 ( .B(n1441), .A(n2868), .Z(n1442) );
  XNOR U1984 ( .A(zin[200]), .B(n1442), .Z(n3528) );
  NANDN U1985 ( .A(n3529), .B(n3528), .Z(n3252) );
  XNOR U1986 ( .A(n3529), .B(n3528), .Z(n2671) );
  IV U1987 ( .A(n[200]), .Z(n6199) );
  XOR U1988 ( .A(y[200]), .B(n1443), .Z(n1444) );
  ANDN U1989 ( .B(n1444), .A(n2868), .Z(n1445) );
  XNOR U1990 ( .A(zin[199]), .B(n1445), .Z(n3533) );
  NANDN U1991 ( .A(n6199), .B(n3533), .Z(n3249) );
  XNOR U1992 ( .A(n3533), .B(n6199), .Z(n2668) );
  XOR U1993 ( .A(y[199]), .B(n1446), .Z(n1447) );
  ANDN U1994 ( .B(n1447), .A(n2868), .Z(n1448) );
  XNOR U1995 ( .A(zin[198]), .B(n1448), .Z(n3537) );
  NAND U1996 ( .A(n[199]), .B(n3537), .Z(n2666) );
  XOR U1997 ( .A(n3537), .B(n[199]), .Z(n2664) );
  XOR U1998 ( .A(y[198]), .B(n1449), .Z(n1450) );
  ANDN U1999 ( .B(n1450), .A(n2868), .Z(n1451) );
  XNOR U2000 ( .A(zin[197]), .B(n1451), .Z(n3542) );
  NAND U2001 ( .A(n[198]), .B(n3542), .Z(n2662) );
  XOR U2002 ( .A(n3542), .B(n[198]), .Z(n2660) );
  XOR U2003 ( .A(y[197]), .B(n1452), .Z(n1453) );
  ANDN U2004 ( .B(n1453), .A(n2868), .Z(n1454) );
  XNOR U2005 ( .A(zin[196]), .B(n1454), .Z(n3546) );
  NAND U2006 ( .A(n[197]), .B(n3546), .Z(n2658) );
  XOR U2007 ( .A(n3546), .B(n[197]), .Z(n2656) );
  IV U2008 ( .A(n[196]), .Z(n6166) );
  XOR U2009 ( .A(y[196]), .B(n1455), .Z(n1456) );
  ANDN U2010 ( .B(n1456), .A(n2868), .Z(n1457) );
  XNOR U2011 ( .A(zin[195]), .B(n1457), .Z(n3550) );
  NANDN U2012 ( .A(n6166), .B(n3550), .Z(n2654) );
  XNOR U2013 ( .A(n3550), .B(n6166), .Z(n2652) );
  IV U2014 ( .A(n[195]), .Z(n3556) );
  XOR U2015 ( .A(y[195]), .B(n1458), .Z(n1459) );
  ANDN U2016 ( .B(n1459), .A(n2868), .Z(n1460) );
  XNOR U2017 ( .A(zin[194]), .B(n1460), .Z(n3554) );
  NANDN U2018 ( .A(n3556), .B(n3554), .Z(n3246) );
  XNOR U2019 ( .A(n3554), .B(n3556), .Z(n2649) );
  XOR U2020 ( .A(y[194]), .B(n1461), .Z(n1462) );
  ANDN U2021 ( .B(n1462), .A(n2868), .Z(n1463) );
  XNOR U2022 ( .A(zin[193]), .B(n1463), .Z(n3560) );
  NAND U2023 ( .A(n[194]), .B(n3560), .Z(n2647) );
  XOR U2024 ( .A(n3560), .B(n[194]), .Z(n2645) );
  XOR U2025 ( .A(y[193]), .B(n1464), .Z(n1465) );
  ANDN U2026 ( .B(n1465), .A(n2868), .Z(n1466) );
  XNOR U2027 ( .A(zin[192]), .B(n1466), .Z(n3564) );
  NAND U2028 ( .A(n[193]), .B(n3564), .Z(n2643) );
  XOR U2029 ( .A(n3564), .B(n[193]), .Z(n2641) );
  XOR U2030 ( .A(y[192]), .B(n1467), .Z(n1468) );
  ANDN U2031 ( .B(n1468), .A(n2868), .Z(n1469) );
  XNOR U2032 ( .A(zin[191]), .B(n1469), .Z(n3568) );
  NAND U2033 ( .A(n3568), .B(n[192]), .Z(n2639) );
  XOR U2034 ( .A(n[192]), .B(n3568), .Z(n2637) );
  XOR U2035 ( .A(y[191]), .B(n1470), .Z(n1471) );
  ANDN U2036 ( .B(n1471), .A(n2868), .Z(n1472) );
  XNOR U2037 ( .A(zin[190]), .B(n1472), .Z(n3572) );
  NAND U2038 ( .A(n[191]), .B(n3572), .Z(n3243) );
  XOR U2039 ( .A(n[191]), .B(n3572), .Z(n2634) );
  IV U2040 ( .A(n[190]), .Z(n6135) );
  XOR U2041 ( .A(y[190]), .B(n1473), .Z(n1474) );
  ANDN U2042 ( .B(n1474), .A(n2868), .Z(n1475) );
  XNOR U2043 ( .A(zin[189]), .B(n1475), .Z(n3576) );
  NANDN U2044 ( .A(n6135), .B(n3576), .Z(n3240) );
  XNOR U2045 ( .A(n3576), .B(n6135), .Z(n2631) );
  IV U2046 ( .A(n[189]), .Z(n3581) );
  XOR U2047 ( .A(y[189]), .B(n1476), .Z(n1477) );
  ANDN U2048 ( .B(n1477), .A(n2868), .Z(n1478) );
  XOR U2049 ( .A(zin[188]), .B(n1478), .Z(n3580) );
  IV U2050 ( .A(n3580), .Z(n2875) );
  NANDN U2051 ( .A(n3581), .B(n2875), .Z(n2629) );
  XNOR U2052 ( .A(n3580), .B(n[189]), .Z(n2627) );
  IV U2053 ( .A(n[188]), .Z(n3586) );
  XOR U2054 ( .A(y[188]), .B(n1479), .Z(n1480) );
  ANDN U2055 ( .B(n1480), .A(n2868), .Z(n1481) );
  XNOR U2056 ( .A(zin[187]), .B(n1481), .Z(n3585) );
  NANDN U2057 ( .A(n3586), .B(n3585), .Z(n3237) );
  XNOR U2058 ( .A(n3586), .B(n3585), .Z(n2624) );
  IV U2059 ( .A(n[187]), .Z(n6106) );
  XOR U2060 ( .A(y[187]), .B(n1482), .Z(n1483) );
  ANDN U2061 ( .B(n1483), .A(n2868), .Z(n1484) );
  XNOR U2062 ( .A(zin[186]), .B(n1484), .Z(n3590) );
  NANDN U2063 ( .A(n6106), .B(n3590), .Z(n3234) );
  XNOR U2064 ( .A(n6106), .B(n3590), .Z(n2621) );
  XOR U2065 ( .A(y[186]), .B(n1485), .Z(n1486) );
  ANDN U2066 ( .B(n1486), .A(n2868), .Z(n1487) );
  XNOR U2067 ( .A(zin[185]), .B(n1487), .Z(n3594) );
  NAND U2068 ( .A(n3594), .B(n[186]), .Z(n2619) );
  XOR U2069 ( .A(n[186]), .B(n3594), .Z(n2617) );
  XOR U2070 ( .A(y[185]), .B(n1488), .Z(n1489) );
  ANDN U2071 ( .B(n1489), .A(n2868), .Z(n1490) );
  XNOR U2072 ( .A(zin[184]), .B(n1490), .Z(n5054) );
  NAND U2073 ( .A(n[185]), .B(n5054), .Z(n2615) );
  XOR U2074 ( .A(n5054), .B(n[185]), .Z(n2613) );
  IV U2075 ( .A(n[184]), .Z(n6086) );
  XOR U2076 ( .A(y[184]), .B(n1491), .Z(n1492) );
  ANDN U2077 ( .B(n1492), .A(n2868), .Z(n1493) );
  XNOR U2078 ( .A(zin[183]), .B(n1493), .Z(n3598) );
  NANDN U2079 ( .A(n6086), .B(n3598), .Z(n3231) );
  XNOR U2080 ( .A(n3598), .B(n6086), .Z(n2610) );
  IV U2081 ( .A(n[183]), .Z(n3603) );
  XOR U2082 ( .A(y[183]), .B(n1494), .Z(n1495) );
  ANDN U2083 ( .B(n1495), .A(n2868), .Z(n1496) );
  XNOR U2084 ( .A(zin[182]), .B(n1496), .Z(n3602) );
  NANDN U2085 ( .A(n3603), .B(n3602), .Z(n3228) );
  XNOR U2086 ( .A(n3603), .B(n3602), .Z(n2607) );
  XOR U2087 ( .A(y[182]), .B(n1497), .Z(n1498) );
  ANDN U2088 ( .B(n1498), .A(n2868), .Z(n1499) );
  XNOR U2089 ( .A(zin[181]), .B(n1499), .Z(n3607) );
  NAND U2090 ( .A(n[182]), .B(n3607), .Z(n2605) );
  XOR U2091 ( .A(n3607), .B(n[182]), .Z(n2603) );
  XOR U2092 ( .A(y[181]), .B(n1500), .Z(n1501) );
  ANDN U2093 ( .B(n1501), .A(n2868), .Z(n1502) );
  XNOR U2094 ( .A(zin[180]), .B(n1502), .Z(n3611) );
  NAND U2095 ( .A(n3611), .B(n[181]), .Z(n2601) );
  XOR U2096 ( .A(n[181]), .B(n3611), .Z(n2599) );
  XOR U2097 ( .A(y[180]), .B(n1503), .Z(n1504) );
  ANDN U2098 ( .B(n1504), .A(n2868), .Z(n1505) );
  XNOR U2099 ( .A(zin[179]), .B(n1505), .Z(n3615) );
  NAND U2100 ( .A(n[180]), .B(n3615), .Z(n2597) );
  XOR U2101 ( .A(n3615), .B(n[180]), .Z(n2595) );
  XOR U2102 ( .A(y[179]), .B(n1506), .Z(n1507) );
  ANDN U2103 ( .B(n1507), .A(n2868), .Z(n1508) );
  XNOR U2104 ( .A(zin[178]), .B(n1508), .Z(n5026) );
  NAND U2105 ( .A(n[179]), .B(n5026), .Z(n2593) );
  XOR U2106 ( .A(n5026), .B(n[179]), .Z(n2591) );
  IV U2107 ( .A(n[178]), .Z(n6039) );
  XOR U2108 ( .A(y[178]), .B(n1509), .Z(n1510) );
  ANDN U2109 ( .B(n1510), .A(n2868), .Z(n1511) );
  XNOR U2110 ( .A(zin[177]), .B(n1511), .Z(n3619) );
  NANDN U2111 ( .A(n6039), .B(n3619), .Z(n2589) );
  XNOR U2112 ( .A(n3619), .B(n6039), .Z(n2587) );
  IV U2113 ( .A(n[177]), .Z(n6042) );
  XOR U2114 ( .A(y[177]), .B(n1512), .Z(n1513) );
  ANDN U2115 ( .B(n1513), .A(n2868), .Z(n1514) );
  XNOR U2116 ( .A(zin[176]), .B(n1514), .Z(n3623) );
  NANDN U2117 ( .A(n6042), .B(n3623), .Z(n3225) );
  XNOR U2118 ( .A(n3623), .B(n6042), .Z(n2584) );
  IV U2119 ( .A(n[176]), .Z(n6025) );
  XOR U2120 ( .A(y[176]), .B(n1515), .Z(n1516) );
  ANDN U2121 ( .B(n1516), .A(n2868), .Z(n1517) );
  XNOR U2122 ( .A(zin[175]), .B(n1517), .Z(n3628) );
  NANDN U2123 ( .A(n6025), .B(n3628), .Z(n2582) );
  XNOR U2124 ( .A(n3628), .B(n6025), .Z(n2580) );
  IV U2125 ( .A(n[175]), .Z(n6024) );
  XOR U2126 ( .A(y[175]), .B(n1518), .Z(n1519) );
  ANDN U2127 ( .B(n1519), .A(n2868), .Z(n1520) );
  XNOR U2128 ( .A(zin[174]), .B(n1520), .Z(n3632) );
  NANDN U2129 ( .A(n6024), .B(n3632), .Z(n3222) );
  XNOR U2130 ( .A(n6024), .B(n3632), .Z(n2577) );
  XOR U2131 ( .A(y[174]), .B(n1521), .Z(n1522) );
  ANDN U2132 ( .B(n1522), .A(n2868), .Z(n1523) );
  XNOR U2133 ( .A(zin[173]), .B(n1523), .Z(n3636) );
  NAND U2134 ( .A(n[174]), .B(n3636), .Z(n2575) );
  XOR U2135 ( .A(n3636), .B(n[174]), .Z(n2573) );
  IV U2136 ( .A(n[173]), .Z(n3641) );
  XOR U2137 ( .A(y[173]), .B(n1524), .Z(n1525) );
  ANDN U2138 ( .B(n1525), .A(n2868), .Z(n1526) );
  XNOR U2139 ( .A(zin[172]), .B(n1526), .Z(n3640) );
  NANDN U2140 ( .A(n3641), .B(n3640), .Z(n3219) );
  XNOR U2141 ( .A(n3640), .B(n3641), .Z(n2570) );
  IV U2142 ( .A(n[172]), .Z(n3646) );
  XOR U2143 ( .A(y[172]), .B(n1527), .Z(n1528) );
  ANDN U2144 ( .B(n1528), .A(n2868), .Z(n1529) );
  XNOR U2145 ( .A(zin[171]), .B(n1529), .Z(n3645) );
  NANDN U2146 ( .A(n3646), .B(n3645), .Z(n3216) );
  XNOR U2147 ( .A(n3646), .B(n3645), .Z(n2567) );
  IV U2148 ( .A(n[171]), .Z(n5998) );
  XOR U2149 ( .A(y[171]), .B(n1530), .Z(n1531) );
  ANDN U2150 ( .B(n1531), .A(n2868), .Z(n1532) );
  XNOR U2151 ( .A(zin[170]), .B(n1532), .Z(n3650) );
  NANDN U2152 ( .A(n5998), .B(n3650), .Z(n3213) );
  XNOR U2153 ( .A(n3650), .B(n5998), .Z(n2564) );
  IV U2154 ( .A(n[170]), .Z(n3655) );
  XOR U2155 ( .A(y[170]), .B(n1533), .Z(n1534) );
  ANDN U2156 ( .B(n1534), .A(n2868), .Z(n1535) );
  XNOR U2157 ( .A(zin[169]), .B(n1535), .Z(n3654) );
  NANDN U2158 ( .A(n3655), .B(n3654), .Z(n3210) );
  XNOR U2159 ( .A(n3655), .B(n3654), .Z(n2561) );
  XOR U2160 ( .A(y[169]), .B(n1536), .Z(n1537) );
  ANDN U2161 ( .B(n1537), .A(n2868), .Z(n1538) );
  XNOR U2162 ( .A(zin[168]), .B(n1538), .Z(n3659) );
  NAND U2163 ( .A(n3659), .B(n[169]), .Z(n2559) );
  XOR U2164 ( .A(n[169]), .B(n3659), .Z(n2557) );
  IV U2165 ( .A(n[168]), .Z(n3664) );
  XOR U2166 ( .A(y[168]), .B(n1539), .Z(n1540) );
  ANDN U2167 ( .B(n1540), .A(n2868), .Z(n1541) );
  XNOR U2168 ( .A(zin[167]), .B(n1541), .Z(n3663) );
  NANDN U2169 ( .A(n3664), .B(n3663), .Z(n3207) );
  XNOR U2170 ( .A(n3664), .B(n3663), .Z(n2554) );
  XOR U2171 ( .A(y[167]), .B(n1542), .Z(n1543) );
  ANDN U2172 ( .B(n1543), .A(n2868), .Z(n1544) );
  XNOR U2173 ( .A(zin[166]), .B(n1544), .Z(n3668) );
  NAND U2174 ( .A(n[167]), .B(n3668), .Z(n3204) );
  XOR U2175 ( .A(n[167]), .B(n3668), .Z(n2551) );
  IV U2176 ( .A(n[166]), .Z(n3673) );
  XOR U2177 ( .A(y[166]), .B(n1545), .Z(n1546) );
  ANDN U2178 ( .B(n1546), .A(n2868), .Z(n1547) );
  XNOR U2179 ( .A(zin[165]), .B(n1547), .Z(n3672) );
  NANDN U2180 ( .A(n3673), .B(n3672), .Z(n3201) );
  XNOR U2181 ( .A(n3672), .B(n3673), .Z(n2548) );
  XOR U2182 ( .A(y[165]), .B(n1548), .Z(n1549) );
  ANDN U2183 ( .B(n1549), .A(n2868), .Z(n1550) );
  XNOR U2184 ( .A(zin[164]), .B(n1550), .Z(n3677) );
  NAND U2185 ( .A(n[165]), .B(n3677), .Z(n3198) );
  XOR U2186 ( .A(n[165]), .B(n3677), .Z(n2545) );
  IV U2187 ( .A(n[164]), .Z(n5943) );
  XOR U2188 ( .A(y[164]), .B(n1551), .Z(n1552) );
  ANDN U2189 ( .B(n1552), .A(n2868), .Z(n1553) );
  XNOR U2190 ( .A(zin[163]), .B(n1553), .Z(n3681) );
  NANDN U2191 ( .A(n5943), .B(n3681), .Z(n3195) );
  XNOR U2192 ( .A(n3681), .B(n5943), .Z(n2542) );
  XOR U2193 ( .A(y[163]), .B(n1554), .Z(n1555) );
  ANDN U2194 ( .B(n1555), .A(n2868), .Z(n1556) );
  XNOR U2195 ( .A(zin[162]), .B(n1556), .Z(n3685) );
  NAND U2196 ( .A(n[163]), .B(n3685), .Z(n2540) );
  XOR U2197 ( .A(n3685), .B(n[163]), .Z(n2538) );
  XOR U2198 ( .A(y[162]), .B(n1557), .Z(n1558) );
  ANDN U2199 ( .B(n1558), .A(n2868), .Z(n1559) );
  XNOR U2200 ( .A(zin[161]), .B(n1559), .Z(n3689) );
  NAND U2201 ( .A(n3689), .B(n[162]), .Z(n2536) );
  XOR U2202 ( .A(n[162]), .B(n3689), .Z(n2534) );
  XOR U2203 ( .A(y[161]), .B(n1560), .Z(n1561) );
  ANDN U2204 ( .B(n1561), .A(n2868), .Z(n1562) );
  XNOR U2205 ( .A(zin[160]), .B(n1562), .Z(n3693) );
  NAND U2206 ( .A(n[161]), .B(n3693), .Z(n2532) );
  XOR U2207 ( .A(n3693), .B(n[161]), .Z(n2530) );
  IV U2208 ( .A(n[160]), .Z(n3698) );
  XOR U2209 ( .A(y[160]), .B(n1563), .Z(n1564) );
  ANDN U2210 ( .B(n1564), .A(n2868), .Z(n1565) );
  XNOR U2211 ( .A(zin[159]), .B(n1565), .Z(n3697) );
  NANDN U2212 ( .A(n3698), .B(n3697), .Z(n3192) );
  XNOR U2213 ( .A(n3697), .B(n3698), .Z(n2527) );
  XOR U2214 ( .A(y[159]), .B(n1566), .Z(n1567) );
  ANDN U2215 ( .B(n1567), .A(n2868), .Z(n1568) );
  XNOR U2216 ( .A(zin[158]), .B(n1568), .Z(n3702) );
  NAND U2217 ( .A(n[159]), .B(n3702), .Z(n2525) );
  XOR U2218 ( .A(n3702), .B(n[159]), .Z(n2523) );
  IV U2219 ( .A(n[158]), .Z(n5903) );
  XOR U2220 ( .A(y[158]), .B(n1569), .Z(n1570) );
  ANDN U2221 ( .B(n1570), .A(n2868), .Z(n1571) );
  XNOR U2222 ( .A(zin[157]), .B(n1571), .Z(n3706) );
  NANDN U2223 ( .A(n5903), .B(n3706), .Z(n3189) );
  XNOR U2224 ( .A(n3706), .B(n5903), .Z(n2520) );
  IV U2225 ( .A(n[157]), .Z(n4939) );
  XOR U2226 ( .A(y[157]), .B(n1572), .Z(n1573) );
  ANDN U2227 ( .B(n1573), .A(n2868), .Z(n1574) );
  XNOR U2228 ( .A(zin[156]), .B(n1574), .Z(n4937) );
  NANDN U2229 ( .A(n4939), .B(n4937), .Z(n3186) );
  XNOR U2230 ( .A(n4939), .B(n4937), .Z(n2517) );
  IV U2231 ( .A(n[156]), .Z(n5889) );
  XOR U2232 ( .A(y[156]), .B(n1575), .Z(n1576) );
  ANDN U2233 ( .B(n1576), .A(n2868), .Z(n1577) );
  XNOR U2234 ( .A(zin[155]), .B(n1577), .Z(n3710) );
  NANDN U2235 ( .A(n5889), .B(n3710), .Z(n3183) );
  XNOR U2236 ( .A(n3710), .B(n5889), .Z(n2514) );
  XOR U2237 ( .A(y[155]), .B(n1578), .Z(n1579) );
  ANDN U2238 ( .B(n1579), .A(n2868), .Z(n1580) );
  XNOR U2239 ( .A(zin[154]), .B(n1580), .Z(n4926) );
  NAND U2240 ( .A(n[155]), .B(n4926), .Z(n2512) );
  XOR U2241 ( .A(n4926), .B(n[155]), .Z(n2510) );
  XOR U2242 ( .A(y[154]), .B(n1581), .Z(n1582) );
  ANDN U2243 ( .B(n1582), .A(n2868), .Z(n1583) );
  XNOR U2244 ( .A(zin[153]), .B(n1583), .Z(n3714) );
  NAND U2245 ( .A(n[154]), .B(n3714), .Z(n3180) );
  XOR U2246 ( .A(n[154]), .B(n3714), .Z(n2507) );
  IV U2247 ( .A(n[153]), .Z(n4910) );
  XOR U2248 ( .A(y[153]), .B(n1584), .Z(n1585) );
  ANDN U2249 ( .B(n1585), .A(n2868), .Z(n1586) );
  XNOR U2250 ( .A(zin[152]), .B(n1586), .Z(n4913) );
  NANDN U2251 ( .A(n4910), .B(n4913), .Z(n3177) );
  XNOR U2252 ( .A(n4910), .B(n4913), .Z(n2504) );
  XOR U2253 ( .A(y[152]), .B(n1587), .Z(n1588) );
  ANDN U2254 ( .B(n1588), .A(n2868), .Z(n1589) );
  XNOR U2255 ( .A(zin[151]), .B(n1589), .Z(n3718) );
  NAND U2256 ( .A(n[152]), .B(n3718), .Z(n2502) );
  XOR U2257 ( .A(n3718), .B(n[152]), .Z(n2500) );
  XOR U2258 ( .A(y[151]), .B(n1590), .Z(n1591) );
  ANDN U2259 ( .B(n1591), .A(n2868), .Z(n1592) );
  XNOR U2260 ( .A(zin[150]), .B(n1592), .Z(n3722) );
  NAND U2261 ( .A(n[151]), .B(n3722), .Z(n3174) );
  XOR U2262 ( .A(n[151]), .B(n3722), .Z(n2497) );
  XOR U2263 ( .A(y[150]), .B(n1593), .Z(n1594) );
  ANDN U2264 ( .B(n1594), .A(n2868), .Z(n1595) );
  XNOR U2265 ( .A(zin[149]), .B(n1595), .Z(n3726) );
  NAND U2266 ( .A(n3726), .B(n[150]), .Z(n2495) );
  XOR U2267 ( .A(n[150]), .B(n3726), .Z(n2493) );
  XOR U2268 ( .A(y[149]), .B(n1596), .Z(n1597) );
  ANDN U2269 ( .B(n1597), .A(n2868), .Z(n1598) );
  XNOR U2270 ( .A(zin[148]), .B(n1598), .Z(n3730) );
  NAND U2271 ( .A(n[149]), .B(n3730), .Z(n2491) );
  XOR U2272 ( .A(n3730), .B(n[149]), .Z(n2489) );
  XOR U2273 ( .A(y[148]), .B(n1599), .Z(n1600) );
  ANDN U2274 ( .B(n1600), .A(n2868), .Z(n1601) );
  XNOR U2275 ( .A(zin[147]), .B(n1601), .Z(n3734) );
  NAND U2276 ( .A(n3734), .B(n[148]), .Z(n2487) );
  XOR U2277 ( .A(n[148]), .B(n3734), .Z(n2485) );
  IV U2278 ( .A(n[147]), .Z(n3739) );
  XOR U2279 ( .A(y[147]), .B(n1602), .Z(n1603) );
  ANDN U2280 ( .B(n1603), .A(n2868), .Z(n1604) );
  XNOR U2281 ( .A(zin[146]), .B(n1604), .Z(n3738) );
  NANDN U2282 ( .A(n3739), .B(n3738), .Z(n3171) );
  XNOR U2283 ( .A(n3739), .B(n3738), .Z(n2482) );
  XOR U2284 ( .A(y[146]), .B(n1605), .Z(n1606) );
  ANDN U2285 ( .B(n1606), .A(n2868), .Z(n1607) );
  XNOR U2286 ( .A(zin[145]), .B(n1607), .Z(n3743) );
  NAND U2287 ( .A(n[146]), .B(n3743), .Z(n2480) );
  XOR U2288 ( .A(n3743), .B(n[146]), .Z(n2478) );
  XOR U2289 ( .A(y[145]), .B(n1608), .Z(n1609) );
  ANDN U2290 ( .B(n1609), .A(n2868), .Z(n1610) );
  XNOR U2291 ( .A(zin[144]), .B(n1610), .Z(n3747) );
  NAND U2292 ( .A(n[145]), .B(n3747), .Z(n3168) );
  XOR U2293 ( .A(n[145]), .B(n3747), .Z(n2475) );
  IV U2294 ( .A(n[144]), .Z(n3752) );
  XOR U2295 ( .A(y[144]), .B(n1611), .Z(n1612) );
  ANDN U2296 ( .B(n1612), .A(n2868), .Z(n1613) );
  XNOR U2297 ( .A(zin[143]), .B(n1613), .Z(n3751) );
  NANDN U2298 ( .A(n3752), .B(n3751), .Z(n3165) );
  XNOR U2299 ( .A(n3752), .B(n3751), .Z(n2472) );
  XOR U2300 ( .A(y[143]), .B(n1614), .Z(n1615) );
  ANDN U2301 ( .B(n1615), .A(n2868), .Z(n1616) );
  XNOR U2302 ( .A(zin[142]), .B(n1616), .Z(n3756) );
  NAND U2303 ( .A(n[143]), .B(n3756), .Z(n2470) );
  XOR U2304 ( .A(n3756), .B(n[143]), .Z(n2468) );
  XOR U2305 ( .A(y[142]), .B(n1617), .Z(n1618) );
  ANDN U2306 ( .B(n1618), .A(n2868), .Z(n1619) );
  XOR U2307 ( .A(zin[141]), .B(n1619), .Z(n2876) );
  NANDN U2308 ( .A(n2876), .B(n[142]), .Z(n2466) );
  XNOR U2309 ( .A(n[142]), .B(n2876), .Z(n2464) );
  XOR U2310 ( .A(y[141]), .B(n1620), .Z(n1621) );
  ANDN U2311 ( .B(n1621), .A(n2868), .Z(n1622) );
  XNOR U2312 ( .A(zin[140]), .B(n1622), .Z(n3764) );
  NAND U2313 ( .A(n[141]), .B(n3764), .Z(n2462) );
  XOR U2314 ( .A(n3764), .B(n[141]), .Z(n2460) );
  IV U2315 ( .A(n[140]), .Z(n3769) );
  XOR U2316 ( .A(y[140]), .B(n1623), .Z(n1624) );
  ANDN U2317 ( .B(n1624), .A(n2868), .Z(n1625) );
  XNOR U2318 ( .A(zin[139]), .B(n1625), .Z(n3768) );
  NANDN U2319 ( .A(n3769), .B(n3768), .Z(n3159) );
  XNOR U2320 ( .A(n3768), .B(n3769), .Z(n2457) );
  XOR U2321 ( .A(y[139]), .B(n1626), .Z(n1627) );
  ANDN U2322 ( .B(n1627), .A(n2868), .Z(n1628) );
  XNOR U2323 ( .A(zin[138]), .B(n1628), .Z(n3773) );
  NAND U2324 ( .A(n[139]), .B(n3773), .Z(n2455) );
  XOR U2325 ( .A(n3773), .B(n[139]), .Z(n2453) );
  XOR U2326 ( .A(y[138]), .B(n1629), .Z(n1630) );
  ANDN U2327 ( .B(n1630), .A(n2868), .Z(n1631) );
  XNOR U2328 ( .A(zin[137]), .B(n1631), .Z(n3777) );
  NAND U2329 ( .A(n3777), .B(n[138]), .Z(n2451) );
  XOR U2330 ( .A(n[138]), .B(n3777), .Z(n2449) );
  XOR U2331 ( .A(y[137]), .B(n1632), .Z(n1633) );
  ANDN U2332 ( .B(n1633), .A(n2868), .Z(n1634) );
  XNOR U2333 ( .A(zin[136]), .B(n1634), .Z(n3781) );
  NAND U2334 ( .A(n[137]), .B(n3781), .Z(n2447) );
  XOR U2335 ( .A(n3781), .B(n[137]), .Z(n2445) );
  XOR U2336 ( .A(y[136]), .B(n1635), .Z(n1636) );
  ANDN U2337 ( .B(n1636), .A(n2868), .Z(n1637) );
  XNOR U2338 ( .A(zin[135]), .B(n1637), .Z(n3785) );
  NAND U2339 ( .A(n3785), .B(n[136]), .Z(n2443) );
  XOR U2340 ( .A(n[136]), .B(n3785), .Z(n2441) );
  XOR U2341 ( .A(y[135]), .B(n1638), .Z(n1639) );
  ANDN U2342 ( .B(n1639), .A(n2868), .Z(n1640) );
  XNOR U2343 ( .A(zin[134]), .B(n1640), .Z(n3789) );
  NAND U2344 ( .A(n[135]), .B(n3789), .Z(n2439) );
  XOR U2345 ( .A(n3789), .B(n[135]), .Z(n2437) );
  XOR U2346 ( .A(y[134]), .B(n1641), .Z(n1642) );
  ANDN U2347 ( .B(n1642), .A(n2868), .Z(n1643) );
  XNOR U2348 ( .A(zin[133]), .B(n1643), .Z(n3793) );
  NAND U2349 ( .A(n[134]), .B(n3793), .Z(n2435) );
  XOR U2350 ( .A(n3793), .B(n[134]), .Z(n2433) );
  IV U2351 ( .A(n[133]), .Z(n3798) );
  XOR U2352 ( .A(y[133]), .B(n1644), .Z(n1645) );
  ANDN U2353 ( .B(n1645), .A(n2868), .Z(n1646) );
  XNOR U2354 ( .A(zin[132]), .B(n1646), .Z(n3797) );
  NANDN U2355 ( .A(n3798), .B(n3797), .Z(n3156) );
  XNOR U2356 ( .A(n3797), .B(n3798), .Z(n2430) );
  XOR U2357 ( .A(y[132]), .B(n1647), .Z(n1648) );
  ANDN U2358 ( .B(n1648), .A(n2868), .Z(n1649) );
  XNOR U2359 ( .A(zin[131]), .B(n1649), .Z(n3802) );
  NAND U2360 ( .A(n[132]), .B(n3802), .Z(n2428) );
  XOR U2361 ( .A(n3802), .B(n[132]), .Z(n2426) );
  XOR U2362 ( .A(y[131]), .B(n1650), .Z(n1651) );
  ANDN U2363 ( .B(n1651), .A(n2868), .Z(n1652) );
  XNOR U2364 ( .A(zin[130]), .B(n1652), .Z(n3806) );
  NAND U2365 ( .A(n[131]), .B(n3806), .Z(n3153) );
  XOR U2366 ( .A(n[131]), .B(n3806), .Z(n2423) );
  IV U2367 ( .A(n[130]), .Z(n3811) );
  XOR U2368 ( .A(y[130]), .B(n1653), .Z(n1654) );
  ANDN U2369 ( .B(n1654), .A(n2868), .Z(n1655) );
  XNOR U2370 ( .A(zin[129]), .B(n1655), .Z(n3810) );
  NANDN U2371 ( .A(n3811), .B(n3810), .Z(n3150) );
  XNOR U2372 ( .A(n3810), .B(n3811), .Z(n2420) );
  XOR U2373 ( .A(y[129]), .B(n1656), .Z(n1657) );
  ANDN U2374 ( .B(n1657), .A(n2868), .Z(n1658) );
  XNOR U2375 ( .A(zin[128]), .B(n1658), .Z(n3815) );
  NAND U2376 ( .A(n[129]), .B(n3815), .Z(n2418) );
  XOR U2377 ( .A(n3815), .B(n[129]), .Z(n2416) );
  XOR U2378 ( .A(y[128]), .B(n1659), .Z(n1660) );
  ANDN U2379 ( .B(n1660), .A(n2868), .Z(n1661) );
  XNOR U2380 ( .A(zin[127]), .B(n1661), .Z(n3819) );
  NAND U2381 ( .A(n[128]), .B(n3819), .Z(n3147) );
  XOR U2382 ( .A(n[128]), .B(n3819), .Z(n2413) );
  XOR U2383 ( .A(y[127]), .B(n1662), .Z(n1663) );
  ANDN U2384 ( .B(n1663), .A(n2868), .Z(n1664) );
  XNOR U2385 ( .A(zin[126]), .B(n1664), .Z(n3823) );
  NAND U2386 ( .A(n3823), .B(n[127]), .Z(n2411) );
  XOR U2387 ( .A(n[127]), .B(n3823), .Z(n2409) );
  XOR U2388 ( .A(y[126]), .B(n1665), .Z(n1666) );
  ANDN U2389 ( .B(n1666), .A(n2868), .Z(n1667) );
  XNOR U2390 ( .A(zin[125]), .B(n1667), .Z(n3827) );
  NAND U2391 ( .A(n[126]), .B(n3827), .Z(n2407) );
  XOR U2392 ( .A(n3827), .B(n[126]), .Z(n2405) );
  IV U2393 ( .A(n[125]), .Z(n3832) );
  XOR U2394 ( .A(y[125]), .B(n1668), .Z(n1669) );
  ANDN U2395 ( .B(n1669), .A(n2868), .Z(n1670) );
  XNOR U2396 ( .A(zin[124]), .B(n1670), .Z(n3831) );
  NANDN U2397 ( .A(n3832), .B(n3831), .Z(n3144) );
  XNOR U2398 ( .A(n3831), .B(n3832), .Z(n2402) );
  XOR U2399 ( .A(y[124]), .B(n1671), .Z(n1672) );
  ANDN U2400 ( .B(n1672), .A(n2868), .Z(n1673) );
  XNOR U2401 ( .A(zin[123]), .B(n1673), .Z(n3836) );
  NAND U2402 ( .A(n[124]), .B(n3836), .Z(n2400) );
  XOR U2403 ( .A(n3836), .B(n[124]), .Z(n2398) );
  IV U2404 ( .A(n[123]), .Z(n3841) );
  XOR U2405 ( .A(y[123]), .B(n1674), .Z(n1675) );
  ANDN U2406 ( .B(n1675), .A(n2868), .Z(n1676) );
  XNOR U2407 ( .A(zin[122]), .B(n1676), .Z(n3840) );
  NANDN U2408 ( .A(n3841), .B(n3840), .Z(n3141) );
  XNOR U2409 ( .A(n3841), .B(n3840), .Z(n2395) );
  IV U2410 ( .A(n[122]), .Z(n3846) );
  XOR U2411 ( .A(y[122]), .B(n1677), .Z(n1678) );
  ANDN U2412 ( .B(n1678), .A(n2868), .Z(n1679) );
  XNOR U2413 ( .A(zin[121]), .B(n1679), .Z(n3845) );
  NANDN U2414 ( .A(n3846), .B(n3845), .Z(n3138) );
  XNOR U2415 ( .A(n3845), .B(n3846), .Z(n2392) );
  IV U2416 ( .A(n[121]), .Z(n3851) );
  XOR U2417 ( .A(y[121]), .B(n1680), .Z(n1681) );
  ANDN U2418 ( .B(n1681), .A(n2868), .Z(n1682) );
  XNOR U2419 ( .A(zin[120]), .B(n1682), .Z(n3850) );
  NANDN U2420 ( .A(n3851), .B(n3850), .Z(n3135) );
  XNOR U2421 ( .A(n3851), .B(n3850), .Z(n2389) );
  IV U2422 ( .A(n[120]), .Z(n3856) );
  XOR U2423 ( .A(y[120]), .B(n1683), .Z(n1684) );
  ANDN U2424 ( .B(n1684), .A(n2868), .Z(n1685) );
  XNOR U2425 ( .A(zin[119]), .B(n1685), .Z(n3855) );
  NANDN U2426 ( .A(n3856), .B(n3855), .Z(n3132) );
  XNOR U2427 ( .A(n3855), .B(n3856), .Z(n2386) );
  XOR U2428 ( .A(y[119]), .B(n1686), .Z(n1687) );
  ANDN U2429 ( .B(n1687), .A(n2868), .Z(n1688) );
  XNOR U2430 ( .A(zin[118]), .B(n1688), .Z(n3860) );
  NAND U2431 ( .A(n[119]), .B(n3860), .Z(n3129) );
  XOR U2432 ( .A(n[119]), .B(n3860), .Z(n2383) );
  IV U2433 ( .A(n[118]), .Z(n5648) );
  XOR U2434 ( .A(y[118]), .B(n1689), .Z(n1690) );
  ANDN U2435 ( .B(n1690), .A(n2868), .Z(n1691) );
  XNOR U2436 ( .A(zin[117]), .B(n1691), .Z(n3864) );
  NANDN U2437 ( .A(n5648), .B(n3864), .Z(n3126) );
  XNOR U2438 ( .A(n3864), .B(n5648), .Z(n2380) );
  IV U2439 ( .A(n[117]), .Z(n3869) );
  XOR U2440 ( .A(y[117]), .B(n1692), .Z(n1693) );
  ANDN U2441 ( .B(n1693), .A(n2868), .Z(n1694) );
  XNOR U2442 ( .A(zin[116]), .B(n1694), .Z(n3868) );
  NANDN U2443 ( .A(n3869), .B(n3868), .Z(n3123) );
  XNOR U2444 ( .A(n3869), .B(n3868), .Z(n2377) );
  IV U2445 ( .A(n[116]), .Z(n5633) );
  XOR U2446 ( .A(y[116]), .B(n1695), .Z(n1696) );
  ANDN U2447 ( .B(n1696), .A(n2868), .Z(n1697) );
  XNOR U2448 ( .A(zin[115]), .B(n1697), .Z(n3873) );
  NANDN U2449 ( .A(n5633), .B(n3873), .Z(n3120) );
  XNOR U2450 ( .A(n3873), .B(n5633), .Z(n2374) );
  IV U2451 ( .A(n[115]), .Z(n3878) );
  XOR U2452 ( .A(y[115]), .B(n1698), .Z(n1699) );
  ANDN U2453 ( .B(n1699), .A(n2868), .Z(n1700) );
  XNOR U2454 ( .A(zin[114]), .B(n1700), .Z(n3877) );
  NANDN U2455 ( .A(n3878), .B(n3877), .Z(n3117) );
  XNOR U2456 ( .A(n3878), .B(n3877), .Z(n2371) );
  IV U2457 ( .A(n[114]), .Z(n3883) );
  XOR U2458 ( .A(y[114]), .B(n1701), .Z(n1702) );
  ANDN U2459 ( .B(n1702), .A(n2868), .Z(n1703) );
  XNOR U2460 ( .A(zin[113]), .B(n1703), .Z(n3882) );
  NANDN U2461 ( .A(n3883), .B(n3882), .Z(n3114) );
  XNOR U2462 ( .A(n3882), .B(n3883), .Z(n2368) );
  IV U2463 ( .A(n[113]), .Z(n3888) );
  XOR U2464 ( .A(y[113]), .B(n1704), .Z(n1705) );
  ANDN U2465 ( .B(n1705), .A(n2868), .Z(n1706) );
  XNOR U2466 ( .A(zin[112]), .B(n1706), .Z(n3887) );
  NANDN U2467 ( .A(n3888), .B(n3887), .Z(n3111) );
  XNOR U2468 ( .A(n3888), .B(n3887), .Z(n2365) );
  IV U2469 ( .A(n[112]), .Z(n3893) );
  XOR U2470 ( .A(y[112]), .B(n1707), .Z(n1708) );
  ANDN U2471 ( .B(n1708), .A(n2868), .Z(n1709) );
  XNOR U2472 ( .A(zin[111]), .B(n1709), .Z(n3892) );
  NANDN U2473 ( .A(n3893), .B(n3892), .Z(n3108) );
  XNOR U2474 ( .A(n3892), .B(n3893), .Z(n2362) );
  IV U2475 ( .A(n[111]), .Z(n3898) );
  XOR U2476 ( .A(y[111]), .B(n1710), .Z(n1711) );
  ANDN U2477 ( .B(n1711), .A(n2868), .Z(n1712) );
  XNOR U2478 ( .A(zin[110]), .B(n1712), .Z(n3897) );
  NANDN U2479 ( .A(n3898), .B(n3897), .Z(n3105) );
  XNOR U2480 ( .A(n3898), .B(n3897), .Z(n2359) );
  IV U2481 ( .A(n[110]), .Z(n3903) );
  XOR U2482 ( .A(y[110]), .B(n1713), .Z(n1714) );
  ANDN U2483 ( .B(n1714), .A(n2868), .Z(n1715) );
  XNOR U2484 ( .A(zin[109]), .B(n1715), .Z(n3902) );
  NANDN U2485 ( .A(n3903), .B(n3902), .Z(n3102) );
  XNOR U2486 ( .A(n3902), .B(n3903), .Z(n2356) );
  XOR U2487 ( .A(y[109]), .B(n1716), .Z(n1717) );
  ANDN U2488 ( .B(n1717), .A(n2868), .Z(n1718) );
  XNOR U2489 ( .A(zin[108]), .B(n1718), .Z(n3907) );
  NAND U2490 ( .A(n[109]), .B(n3907), .Z(n3099) );
  XOR U2491 ( .A(n[109]), .B(n3907), .Z(n2353) );
  IV U2492 ( .A(n[108]), .Z(n3912) );
  XOR U2493 ( .A(y[108]), .B(n1719), .Z(n1720) );
  ANDN U2494 ( .B(n1720), .A(n2868), .Z(n1721) );
  XNOR U2495 ( .A(zin[107]), .B(n1721), .Z(n3911) );
  NANDN U2496 ( .A(n3912), .B(n3911), .Z(n3096) );
  XNOR U2497 ( .A(n3911), .B(n3912), .Z(n2350) );
  XOR U2498 ( .A(y[107]), .B(n1722), .Z(n1723) );
  ANDN U2499 ( .B(n1723), .A(n2868), .Z(n1724) );
  XNOR U2500 ( .A(zin[106]), .B(n1724), .Z(n3916) );
  NAND U2501 ( .A(n[107]), .B(n3916), .Z(n2348) );
  XOR U2502 ( .A(n3916), .B(n[107]), .Z(n2346) );
  XOR U2503 ( .A(y[106]), .B(n1725), .Z(n1726) );
  ANDN U2504 ( .B(n1726), .A(n2868), .Z(n1727) );
  XNOR U2505 ( .A(zin[105]), .B(n1727), .Z(n3920) );
  NAND U2506 ( .A(n[106]), .B(n3920), .Z(n2344) );
  XOR U2507 ( .A(n3920), .B(n[106]), .Z(n2342) );
  XOR U2508 ( .A(y[105]), .B(n1728), .Z(n1729) );
  ANDN U2509 ( .B(n1729), .A(n2868), .Z(n1730) );
  XNOR U2510 ( .A(zin[104]), .B(n1730), .Z(n3924) );
  NAND U2511 ( .A(n[105]), .B(n3924), .Z(n2340) );
  XOR U2512 ( .A(n3924), .B(n[105]), .Z(n2338) );
  XOR U2513 ( .A(y[104]), .B(n1731), .Z(n1732) );
  ANDN U2514 ( .B(n1732), .A(n2868), .Z(n1733) );
  XNOR U2515 ( .A(zin[103]), .B(n1733), .Z(n3928) );
  NAND U2516 ( .A(n[104]), .B(n3928), .Z(n2336) );
  XOR U2517 ( .A(n3928), .B(n[104]), .Z(n2334) );
  IV U2518 ( .A(n[103]), .Z(n3933) );
  XOR U2519 ( .A(y[103]), .B(n1734), .Z(n1735) );
  ANDN U2520 ( .B(n1735), .A(n2868), .Z(n1736) );
  XNOR U2521 ( .A(zin[102]), .B(n1736), .Z(n3932) );
  NANDN U2522 ( .A(n3933), .B(n3932), .Z(n3093) );
  XNOR U2523 ( .A(n3933), .B(n3932), .Z(n2331) );
  XOR U2524 ( .A(y[102]), .B(n1737), .Z(n1738) );
  ANDN U2525 ( .B(n1738), .A(n2868), .Z(n1739) );
  XNOR U2526 ( .A(zin[101]), .B(n1739), .Z(n3937) );
  NAND U2527 ( .A(n[102]), .B(n3937), .Z(n2329) );
  XOR U2528 ( .A(n3937), .B(n[102]), .Z(n2327) );
  IV U2529 ( .A(n[101]), .Z(n3942) );
  XOR U2530 ( .A(y[101]), .B(n1740), .Z(n1741) );
  ANDN U2531 ( .B(n1741), .A(n2868), .Z(n1742) );
  XNOR U2532 ( .A(zin[100]), .B(n1742), .Z(n3941) );
  NANDN U2533 ( .A(n3942), .B(n3941), .Z(n3090) );
  XNOR U2534 ( .A(n3942), .B(n3941), .Z(n2324) );
  XOR U2535 ( .A(y[100]), .B(n1743), .Z(n1744) );
  ANDN U2536 ( .B(n1744), .A(n2868), .Z(n1745) );
  XNOR U2537 ( .A(zin[99]), .B(n1745), .Z(n3946) );
  IV U2538 ( .A(n[99]), .Z(n5344) );
  XOR U2539 ( .A(y[99]), .B(n1746), .Z(n1747) );
  ANDN U2540 ( .B(n1747), .A(n2868), .Z(n1748) );
  XNOR U2541 ( .A(zin[98]), .B(n1748), .Z(n3950) );
  XOR U2542 ( .A(y[98]), .B(n1749), .Z(n1750) );
  ANDN U2543 ( .B(n1750), .A(n2868), .Z(n1751) );
  XNOR U2544 ( .A(zin[97]), .B(n1751), .Z(n3954) );
  XOR U2545 ( .A(y[97]), .B(n1752), .Z(n1753) );
  ANDN U2546 ( .B(n1753), .A(n2868), .Z(n1754) );
  XNOR U2547 ( .A(zin[96]), .B(n1754), .Z(n3958) );
  IV U2548 ( .A(n[96]), .Z(n3963) );
  XOR U2549 ( .A(y[96]), .B(n1755), .Z(n1756) );
  ANDN U2550 ( .B(n1756), .A(n2868), .Z(n1757) );
  XNOR U2551 ( .A(zin[95]), .B(n1757), .Z(n3962) );
  NANDN U2552 ( .A(n3963), .B(n3962), .Z(n3087) );
  IV U2553 ( .A(n[95]), .Z(n5529) );
  XOR U2554 ( .A(y[95]), .B(n1758), .Z(n1759) );
  ANDN U2555 ( .B(n1759), .A(n2868), .Z(n1760) );
  XNOR U2556 ( .A(zin[94]), .B(n1760), .Z(n3967) );
  NANDN U2557 ( .A(n5529), .B(n3967), .Z(n3084) );
  XNOR U2558 ( .A(n5529), .B(n3967), .Z(n2320) );
  IV U2559 ( .A(n[94]), .Z(n3969) );
  XOR U2560 ( .A(y[94]), .B(n1761), .Z(n1762) );
  ANDN U2561 ( .B(n1762), .A(n2868), .Z(n1763) );
  XNOR U2562 ( .A(zin[93]), .B(n1763), .Z(n3972) );
  NANDN U2563 ( .A(n3969), .B(n3972), .Z(n3081) );
  XNOR U2564 ( .A(n3972), .B(n3969), .Z(n2317) );
  IV U2565 ( .A(n[93]), .Z(n3974) );
  XOR U2566 ( .A(y[93]), .B(n1764), .Z(n1765) );
  ANDN U2567 ( .B(n1765), .A(n2868), .Z(n1766) );
  XNOR U2568 ( .A(zin[92]), .B(n1766), .Z(n3977) );
  NANDN U2569 ( .A(n3974), .B(n3977), .Z(n3078) );
  XNOR U2570 ( .A(n3974), .B(n3977), .Z(n2314) );
  IV U2571 ( .A(n[92]), .Z(n5353) );
  XOR U2572 ( .A(y[92]), .B(n1767), .Z(n1768) );
  ANDN U2573 ( .B(n1768), .A(n2868), .Z(n1769) );
  XNOR U2574 ( .A(zin[91]), .B(n1769), .Z(n4663) );
  NANDN U2575 ( .A(n5353), .B(n4663), .Z(n3075) );
  XNOR U2576 ( .A(n4663), .B(n5353), .Z(n2311) );
  XOR U2577 ( .A(y[91]), .B(n1770), .Z(n1771) );
  ANDN U2578 ( .B(n1771), .A(n2868), .Z(n1772) );
  XNOR U2579 ( .A(zin[90]), .B(n1772), .Z(n3981) );
  NAND U2580 ( .A(n[91]), .B(n3981), .Z(n3072) );
  XOR U2581 ( .A(n[91]), .B(n3981), .Z(n2308) );
  XOR U2582 ( .A(y[90]), .B(n1773), .Z(n1774) );
  ANDN U2583 ( .B(n1774), .A(n2868), .Z(n1775) );
  XNOR U2584 ( .A(zin[89]), .B(n1775), .Z(n3985) );
  NAND U2585 ( .A(n[90]), .B(n3985), .Z(n2306) );
  XOR U2586 ( .A(n3985), .B(n[90]), .Z(n2304) );
  XOR U2587 ( .A(y[89]), .B(n1776), .Z(n1777) );
  ANDN U2588 ( .B(n1777), .A(n2868), .Z(n1778) );
  XNOR U2589 ( .A(zin[88]), .B(n1778), .Z(n3989) );
  NAND U2590 ( .A(n[89]), .B(n3989), .Z(n3069) );
  XOR U2591 ( .A(n[89]), .B(n3989), .Z(n2301) );
  XOR U2592 ( .A(y[88]), .B(n1779), .Z(n1780) );
  ANDN U2593 ( .B(n1780), .A(n2868), .Z(n1781) );
  XNOR U2594 ( .A(zin[87]), .B(n1781), .Z(n3993) );
  NAND U2595 ( .A(n3993), .B(n[88]), .Z(n2299) );
  XOR U2596 ( .A(n[88]), .B(n3993), .Z(n2297) );
  IV U2597 ( .A(n[87]), .Z(n3998) );
  XOR U2598 ( .A(y[87]), .B(n1782), .Z(n1783) );
  ANDN U2599 ( .B(n1783), .A(n2868), .Z(n1784) );
  XNOR U2600 ( .A(zin[86]), .B(n1784), .Z(n3997) );
  NANDN U2601 ( .A(n3998), .B(n3997), .Z(n3066) );
  XNOR U2602 ( .A(n3998), .B(n3997), .Z(n2294) );
  XOR U2603 ( .A(y[86]), .B(n1785), .Z(n1786) );
  ANDN U2604 ( .B(n1786), .A(n2868), .Z(n1787) );
  XNOR U2605 ( .A(zin[85]), .B(n1787), .Z(n4002) );
  NAND U2606 ( .A(n4002), .B(n[86]), .Z(n2292) );
  XOR U2607 ( .A(n[86]), .B(n4002), .Z(n2290) );
  IV U2608 ( .A(n[85]), .Z(n5504) );
  XOR U2609 ( .A(y[85]), .B(n1788), .Z(n1789) );
  ANDN U2610 ( .B(n1789), .A(n2868), .Z(n1790) );
  XNOR U2611 ( .A(zin[84]), .B(n1790), .Z(n4006) );
  NANDN U2612 ( .A(n5504), .B(n4006), .Z(n3063) );
  XNOR U2613 ( .A(n5504), .B(n4006), .Z(n2287) );
  XOR U2614 ( .A(y[84]), .B(n1791), .Z(n1792) );
  ANDN U2615 ( .B(n1792), .A(n2868), .Z(n1793) );
  XNOR U2616 ( .A(zin[83]), .B(n1793), .Z(n4010) );
  NAND U2617 ( .A(n4010), .B(n[84]), .Z(n2285) );
  XOR U2618 ( .A(n[84]), .B(n4010), .Z(n2283) );
  XOR U2619 ( .A(y[83]), .B(n1794), .Z(n1795) );
  ANDN U2620 ( .B(n1795), .A(n2868), .Z(n1796) );
  XNOR U2621 ( .A(zin[82]), .B(n1796), .Z(n4014) );
  NAND U2622 ( .A(n[83]), .B(n4014), .Z(n2281) );
  XOR U2623 ( .A(n4014), .B(n[83]), .Z(n2279) );
  XOR U2624 ( .A(y[82]), .B(n1797), .Z(n1798) );
  ANDN U2625 ( .B(n1798), .A(n2868), .Z(n1799) );
  XNOR U2626 ( .A(zin[81]), .B(n1799), .Z(n4018) );
  NAND U2627 ( .A(n[82]), .B(n4018), .Z(n2277) );
  XOR U2628 ( .A(n4018), .B(n[82]), .Z(n2275) );
  IV U2629 ( .A(n[81]), .Z(n4023) );
  XOR U2630 ( .A(y[81]), .B(n1800), .Z(n1801) );
  ANDN U2631 ( .B(n1801), .A(n2868), .Z(n1802) );
  XNOR U2632 ( .A(zin[80]), .B(n1802), .Z(n4022) );
  NANDN U2633 ( .A(n4023), .B(n4022), .Z(n3060) );
  XNOR U2634 ( .A(n4023), .B(n4022), .Z(n2272) );
  IV U2635 ( .A(n[80]), .Z(n4028) );
  XOR U2636 ( .A(y[80]), .B(n1803), .Z(n1804) );
  ANDN U2637 ( .B(n1804), .A(n2868), .Z(n1805) );
  XNOR U2638 ( .A(zin[79]), .B(n1805), .Z(n4027) );
  NANDN U2639 ( .A(n4028), .B(n4027), .Z(n3057) );
  XNOR U2640 ( .A(n4028), .B(n4027), .Z(n2269) );
  XOR U2641 ( .A(y[79]), .B(n1806), .Z(n1807) );
  ANDN U2642 ( .B(n1807), .A(n2868), .Z(n1808) );
  XNOR U2643 ( .A(zin[78]), .B(n1808), .Z(n4032) );
  NAND U2644 ( .A(n[79]), .B(n4032), .Z(n2267) );
  XOR U2645 ( .A(n4032), .B(n[79]), .Z(n2265) );
  XOR U2646 ( .A(y[78]), .B(n1809), .Z(n1810) );
  ANDN U2647 ( .B(n1810), .A(n2868), .Z(n1811) );
  XNOR U2648 ( .A(zin[77]), .B(n1811), .Z(n4036) );
  NAND U2649 ( .A(n4036), .B(n[78]), .Z(n2263) );
  XOR U2650 ( .A(n[78]), .B(n4036), .Z(n2261) );
  IV U2651 ( .A(n[77]), .Z(n4041) );
  XOR U2652 ( .A(y[77]), .B(n1812), .Z(n1813) );
  ANDN U2653 ( .B(n1813), .A(n2868), .Z(n1814) );
  XNOR U2654 ( .A(zin[76]), .B(n1814), .Z(n4040) );
  NANDN U2655 ( .A(n4041), .B(n4040), .Z(n3054) );
  XNOR U2656 ( .A(n4041), .B(n4040), .Z(n2258) );
  XOR U2657 ( .A(y[76]), .B(n1815), .Z(n1816) );
  ANDN U2658 ( .B(n1816), .A(n2868), .Z(n1817) );
  XNOR U2659 ( .A(zin[75]), .B(n1817), .Z(n4045) );
  NAND U2660 ( .A(n4045), .B(n[76]), .Z(n2256) );
  XOR U2661 ( .A(n[76]), .B(n4045), .Z(n2254) );
  XOR U2662 ( .A(y[75]), .B(n1818), .Z(n1819) );
  ANDN U2663 ( .B(n1819), .A(n2868), .Z(n1820) );
  XNOR U2664 ( .A(zin[74]), .B(n1820), .Z(n4049) );
  NAND U2665 ( .A(n[75]), .B(n4049), .Z(n2252) );
  XOR U2666 ( .A(n4049), .B(n[75]), .Z(n2250) );
  XOR U2667 ( .A(y[74]), .B(n1821), .Z(n1822) );
  ANDN U2668 ( .B(n1822), .A(n2868), .Z(n1823) );
  XOR U2669 ( .A(zin[73]), .B(n1823), .Z(n2877) );
  NANDN U2670 ( .A(n2877), .B(n[74]), .Z(n2248) );
  XNOR U2671 ( .A(n[74]), .B(n2877), .Z(n2246) );
  XOR U2672 ( .A(y[73]), .B(n1824), .Z(n1825) );
  ANDN U2673 ( .B(n1825), .A(n2868), .Z(n1826) );
  XNOR U2674 ( .A(zin[72]), .B(n1826), .Z(n4057) );
  NAND U2675 ( .A(n[73]), .B(n4057), .Z(n2244) );
  XOR U2676 ( .A(n4057), .B(n[73]), .Z(n2242) );
  XOR U2677 ( .A(y[72]), .B(n1827), .Z(n1828) );
  ANDN U2678 ( .B(n1828), .A(n2868), .Z(n1829) );
  XOR U2679 ( .A(zin[71]), .B(n1829), .Z(n2878) );
  NANDN U2680 ( .A(n2878), .B(n[72]), .Z(n2240) );
  XNOR U2681 ( .A(n[72]), .B(n2878), .Z(n2238) );
  IV U2682 ( .A(n[71]), .Z(n5390) );
  XOR U2683 ( .A(y[71]), .B(n1830), .Z(n1831) );
  ANDN U2684 ( .B(n1831), .A(n2868), .Z(n1832) );
  XNOR U2685 ( .A(zin[70]), .B(n1832), .Z(n4065) );
  NANDN U2686 ( .A(n5390), .B(n4065), .Z(n2236) );
  XNOR U2687 ( .A(n4065), .B(n5390), .Z(n2234) );
  IV U2688 ( .A(n[70]), .Z(n5469) );
  XOR U2689 ( .A(y[70]), .B(n1833), .Z(n1834) );
  ANDN U2690 ( .B(n1834), .A(n2868), .Z(n1835) );
  XNOR U2691 ( .A(zin[69]), .B(n1835), .Z(n4069) );
  NANDN U2692 ( .A(n5469), .B(n4069), .Z(n3045) );
  XNOR U2693 ( .A(n4069), .B(n5469), .Z(n2231) );
  XOR U2694 ( .A(y[69]), .B(n1836), .Z(n1837) );
  ANDN U2695 ( .B(n1837), .A(n2868), .Z(n1838) );
  XNOR U2696 ( .A(zin[68]), .B(n1838), .Z(n4073) );
  NAND U2697 ( .A(n[69]), .B(n4073), .Z(n2229) );
  XOR U2698 ( .A(n4073), .B(n[69]), .Z(n2227) );
  XOR U2699 ( .A(y[67]), .B(n1839), .Z(n1840) );
  ANDN U2700 ( .B(n1840), .A(n2868), .Z(n1841) );
  XNOR U2701 ( .A(zin[66]), .B(n1841), .Z(n4082) );
  NAND U2702 ( .A(n[67]), .B(n4082), .Z(n1845) );
  XOR U2703 ( .A(y[68]), .B(n1842), .Z(n1843) );
  ANDN U2704 ( .B(n1843), .A(n2868), .Z(n1844) );
  XNOR U2705 ( .A(zin[67]), .B(n1844), .Z(n4077) );
  AND U2706 ( .A(n4077), .B(n[68]), .Z(n3040) );
  ANDN U2707 ( .B(n1845), .A(n3040), .Z(n2224) );
  XOR U2708 ( .A(n4082), .B(n[67]), .Z(n2222) );
  XOR U2709 ( .A(y[66]), .B(n1846), .Z(n1847) );
  ANDN U2710 ( .B(n1847), .A(n2868), .Z(n1848) );
  XNOR U2711 ( .A(zin[65]), .B(n1848), .Z(n4086) );
  NAND U2712 ( .A(n4086), .B(n[66]), .Z(n2220) );
  XOR U2713 ( .A(n[66]), .B(n4086), .Z(n2218) );
  XOR U2714 ( .A(y[65]), .B(n1849), .Z(n1850) );
  ANDN U2715 ( .B(n1850), .A(n2868), .Z(n1851) );
  XNOR U2716 ( .A(zin[64]), .B(n1851), .Z(n4090) );
  AND U2717 ( .A(n4090), .B(n[65]), .Z(n3037) );
  IV U2718 ( .A(n[65]), .Z(n4091) );
  ANDN U2719 ( .B(n4091), .A(n4090), .Z(n3038) );
  XOR U2720 ( .A(y[64]), .B(n1852), .Z(n1853) );
  ANDN U2721 ( .B(n1853), .A(n2868), .Z(n1854) );
  XOR U2722 ( .A(zin[63]), .B(n1854), .Z(n4095) );
  IV U2723 ( .A(n[64]), .Z(n5399) );
  AND U2724 ( .A(n4095), .B(n5399), .Z(n3036) );
  NOR U2725 ( .A(n3038), .B(n3036), .Z(n2215) );
  XOR U2726 ( .A(y[62]), .B(n1855), .Z(n1856) );
  ANDN U2727 ( .B(n1856), .A(n2868), .Z(n1857) );
  XOR U2728 ( .A(zin[61]), .B(n1857), .Z(n4103) );
  NANDN U2729 ( .A(n[62]), .B(n4103), .Z(n3031) );
  XOR U2730 ( .A(y[61]), .B(n1858), .Z(n1859) );
  ANDN U2731 ( .B(n1859), .A(n2868), .Z(n1860) );
  XOR U2732 ( .A(zin[60]), .B(n1860), .Z(n4107) );
  IV U2733 ( .A(n[61]), .Z(n4108) );
  AND U2734 ( .A(n4107), .B(n4108), .Z(n3030) );
  ANDN U2735 ( .B(n3031), .A(n3030), .Z(n2204) );
  XOR U2736 ( .A(y[58]), .B(n1861), .Z(n1862) );
  ANDN U2737 ( .B(n1862), .A(n2868), .Z(n1863) );
  XOR U2738 ( .A(zin[57]), .B(n1863), .Z(n4122) );
  IV U2739 ( .A(n[58]), .Z(n5411) );
  AND U2740 ( .A(n4122), .B(n5411), .Z(n3019) );
  XOR U2741 ( .A(y[59]), .B(n1864), .Z(n1865) );
  ANDN U2742 ( .B(n1865), .A(n2868), .Z(n1866) );
  XOR U2743 ( .A(zin[58]), .B(n1866), .Z(n4117) );
  IV U2744 ( .A(n[59]), .Z(n4118) );
  AND U2745 ( .A(n4117), .B(n4118), .Z(n3022) );
  NOR U2746 ( .A(n3019), .B(n3022), .Z(n2193) );
  IV U2747 ( .A(n[56]), .Z(n4131) );
  XOR U2748 ( .A(y[56]), .B(n1867), .Z(n1868) );
  ANDN U2749 ( .B(n1868), .A(n2868), .Z(n1869) );
  XNOR U2750 ( .A(zin[55]), .B(n1869), .Z(n4130) );
  ANDN U2751 ( .B(n4131), .A(n4130), .Z(n3018) );
  XOR U2752 ( .A(y[55]), .B(n1870), .Z(n1871) );
  ANDN U2753 ( .B(n1871), .A(n2868), .Z(n1872) );
  XNOR U2754 ( .A(zin[54]), .B(n1872), .Z(n4135) );
  AND U2755 ( .A(n4135), .B(n[55]), .Z(n3013) );
  XOR U2756 ( .A(y[54]), .B(n1873), .Z(n1874) );
  ANDN U2757 ( .B(n1874), .A(n2868), .Z(n1875) );
  XNOR U2758 ( .A(zin[53]), .B(n1875), .Z(n4139) );
  AND U2759 ( .A(n4139), .B(n[54]), .Z(n3010) );
  IV U2760 ( .A(n[54]), .Z(n4140) );
  ANDN U2761 ( .B(n4140), .A(n4139), .Z(n3012) );
  XOR U2762 ( .A(y[53]), .B(n1876), .Z(n1877) );
  ANDN U2763 ( .B(n1877), .A(n2868), .Z(n1878) );
  XOR U2764 ( .A(zin[52]), .B(n1878), .Z(n4144) );
  ANDN U2765 ( .B(n[53]), .A(n4144), .Z(n3009) );
  IV U2766 ( .A(n[53]), .Z(n4145) );
  AND U2767 ( .A(n4144), .B(n4145), .Z(n3007) );
  XOR U2768 ( .A(y[52]), .B(n1879), .Z(n1880) );
  ANDN U2769 ( .B(n1880), .A(n2868), .Z(n1881) );
  XNOR U2770 ( .A(zin[51]), .B(n1881), .Z(n4149) );
  AND U2771 ( .A(n4149), .B(n[52]), .Z(n3006) );
  OR U2772 ( .A(n4149), .B(n[52]), .Z(n3004) );
  XOR U2773 ( .A(y[50]), .B(n1882), .Z(n1883) );
  ANDN U2774 ( .B(n1883), .A(n2868), .Z(n1884) );
  XOR U2775 ( .A(zin[49]), .B(n1884), .Z(n4157) );
  IV U2776 ( .A(n4157), .Z(n2165) );
  NOR U2777 ( .A(n2165), .B(n[50]), .Z(n3001) );
  XOR U2778 ( .A(y[49]), .B(n1885), .Z(n1886) );
  ANDN U2779 ( .B(n1886), .A(n2868), .Z(n1887) );
  XNOR U2780 ( .A(zin[48]), .B(n1887), .Z(n4161) );
  AND U2781 ( .A(n4161), .B(n[49]), .Z(n3000) );
  XOR U2782 ( .A(y[48]), .B(n1888), .Z(n1889) );
  ANDN U2783 ( .B(n1889), .A(n2868), .Z(n1890) );
  XOR U2784 ( .A(zin[47]), .B(n1890), .Z(n4166) );
  ANDN U2785 ( .B(n[48]), .A(n4166), .Z(n2997) );
  XOR U2786 ( .A(y[47]), .B(n1891), .Z(n1892) );
  ANDN U2787 ( .B(n1892), .A(n2868), .Z(n1893) );
  XNOR U2788 ( .A(zin[46]), .B(n1893), .Z(n4170) );
  AND U2789 ( .A(n4170), .B(n[47]), .Z(n2992) );
  IV U2790 ( .A(n[47]), .Z(n6716) );
  NANDN U2791 ( .A(n4170), .B(n6716), .Z(n2994) );
  XOR U2792 ( .A(y[46]), .B(n1894), .Z(n1895) );
  ANDN U2793 ( .B(n1895), .A(n2868), .Z(n1896) );
  XOR U2794 ( .A(zin[45]), .B(n1896), .Z(n4174) );
  IV U2795 ( .A(n[46]), .Z(n6710) );
  AND U2796 ( .A(n4174), .B(n6710), .Z(n2991) );
  ANDN U2797 ( .B(n2994), .A(n2991), .Z(n2158) );
  XOR U2798 ( .A(y[44]), .B(n1897), .Z(n1898) );
  ANDN U2799 ( .B(n1898), .A(n2868), .Z(n1899) );
  XNOR U2800 ( .A(zin[43]), .B(n1899), .Z(n4470) );
  NOR U2801 ( .A(n[44]), .B(n4470), .Z(n2988) );
  XOR U2802 ( .A(y[43]), .B(n1900), .Z(n1901) );
  ANDN U2803 ( .B(n1901), .A(n2868), .Z(n1902) );
  XNOR U2804 ( .A(zin[42]), .B(n1902), .Z(n4466) );
  AND U2805 ( .A(n4466), .B(n[43]), .Z(n2985) );
  XOR U2806 ( .A(y[42]), .B(n1903), .Z(n1904) );
  ANDN U2807 ( .B(n1904), .A(n2868), .Z(n1905) );
  XOR U2808 ( .A(zin[41]), .B(n1905), .Z(n4178) );
  ANDN U2809 ( .B(n[42]), .A(n4178), .Z(n2982) );
  IV U2810 ( .A(n[42]), .Z(n4179) );
  AND U2811 ( .A(n4178), .B(n4179), .Z(n2980) );
  XOR U2812 ( .A(y[41]), .B(n1906), .Z(n1907) );
  ANDN U2813 ( .B(n1907), .A(n2868), .Z(n1908) );
  XOR U2814 ( .A(zin[40]), .B(n1908), .Z(n4183) );
  ANDN U2815 ( .B(n[41]), .A(n4183), .Z(n2979) );
  NANDN U2816 ( .A(n[41]), .B(n4183), .Z(n2977) );
  XOR U2817 ( .A(y[40]), .B(n1909), .Z(n1910) );
  ANDN U2818 ( .B(n1910), .A(n2868), .Z(n1911) );
  XOR U2819 ( .A(zin[39]), .B(n1911), .Z(n4187) );
  IV U2820 ( .A(n[40]), .Z(n4188) );
  AND U2821 ( .A(n4187), .B(n4188), .Z(n2976) );
  ANDN U2822 ( .B(n2977), .A(n2976), .Z(n2141) );
  IV U2823 ( .A(n[38]), .Z(n4197) );
  XOR U2824 ( .A(y[38]), .B(n1912), .Z(n1913) );
  ANDN U2825 ( .B(n1913), .A(n2868), .Z(n1914) );
  XNOR U2826 ( .A(zin[37]), .B(n1914), .Z(n4196) );
  ANDN U2827 ( .B(n4197), .A(n4196), .Z(n2970) );
  XOR U2828 ( .A(y[37]), .B(n1915), .Z(n1916) );
  ANDN U2829 ( .B(n1916), .A(n2868), .Z(n1917) );
  XNOR U2830 ( .A(zin[36]), .B(n1917), .Z(n4201) );
  AND U2831 ( .A(n4201), .B(n[37]), .Z(n2965) );
  XOR U2832 ( .A(y[36]), .B(n1918), .Z(n1919) );
  ANDN U2833 ( .B(n1919), .A(n2868), .Z(n1920) );
  XNOR U2834 ( .A(zin[35]), .B(n1920), .Z(n4205) );
  AND U2835 ( .A(n4205), .B(n[36]), .Z(n2962) );
  XOR U2836 ( .A(y[34]), .B(n1921), .Z(n1922) );
  ANDN U2837 ( .B(n1922), .A(n2868), .Z(n1923) );
  XNOR U2838 ( .A(zin[33]), .B(n1923), .Z(n4209) );
  NAND U2839 ( .A(n[34]), .B(n4209), .Z(n2118) );
  XOR U2840 ( .A(n4209), .B(n[34]), .Z(n2116) );
  XOR U2841 ( .A(y[33]), .B(n1924), .Z(n1925) );
  ANDN U2842 ( .B(n1925), .A(n2868), .Z(n1926) );
  XNOR U2843 ( .A(zin[32]), .B(n1926), .Z(n4213) );
  NAND U2844 ( .A(n[33]), .B(n4213), .Z(n2114) );
  XOR U2845 ( .A(n4213), .B(n[33]), .Z(n2112) );
  XOR U2846 ( .A(y[32]), .B(n1927), .Z(n1928) );
  ANDN U2847 ( .B(n1928), .A(n2868), .Z(n1929) );
  XNOR U2848 ( .A(zin[31]), .B(n1929), .Z(n4217) );
  NAND U2849 ( .A(n4217), .B(n[32]), .Z(n2110) );
  XOR U2850 ( .A(n[32]), .B(n4217), .Z(n2108) );
  IV U2851 ( .A(n[31]), .Z(n4416) );
  XOR U2852 ( .A(y[31]), .B(n1930), .Z(n1931) );
  ANDN U2853 ( .B(n1931), .A(n2868), .Z(n1932) );
  XNOR U2854 ( .A(zin[30]), .B(n1932), .Z(n4419) );
  NANDN U2855 ( .A(n4416), .B(n4419), .Z(n2961) );
  XNOR U2856 ( .A(n4416), .B(n4419), .Z(n2105) );
  IV U2857 ( .A(n[30]), .Z(n4222) );
  XOR U2858 ( .A(y[30]), .B(n1933), .Z(n1934) );
  ANDN U2859 ( .B(n1934), .A(n2868), .Z(n1935) );
  XNOR U2860 ( .A(zin[29]), .B(n1935), .Z(n4221) );
  NANDN U2861 ( .A(n4222), .B(n4221), .Z(n2958) );
  XNOR U2862 ( .A(n4221), .B(n4222), .Z(n2102) );
  IV U2863 ( .A(n[29]), .Z(n4407) );
  XOR U2864 ( .A(y[29]), .B(n1936), .Z(n1937) );
  ANDN U2865 ( .B(n1937), .A(n2868), .Z(n1938) );
  XNOR U2866 ( .A(zin[28]), .B(n1938), .Z(n4226) );
  NANDN U2867 ( .A(n4407), .B(n4226), .Z(n2955) );
  XNOR U2868 ( .A(n4407), .B(n4226), .Z(n2099) );
  XOR U2869 ( .A(y[28]), .B(n1939), .Z(n1940) );
  ANDN U2870 ( .B(n1940), .A(n2868), .Z(n1941) );
  XNOR U2871 ( .A(zin[27]), .B(n1941), .Z(n4406) );
  NAND U2872 ( .A(n[28]), .B(n4406), .Z(n2952) );
  XOR U2873 ( .A(n[28]), .B(n4406), .Z(n2096) );
  IV U2874 ( .A(n[27]), .Z(n4399) );
  XOR U2875 ( .A(y[27]), .B(n1942), .Z(n1943) );
  ANDN U2876 ( .B(n1943), .A(n2868), .Z(n1944) );
  XOR U2877 ( .A(zin[26]), .B(n1944), .Z(n4402) );
  IV U2878 ( .A(n4402), .Z(n2879) );
  NANDN U2879 ( .A(n4399), .B(n2879), .Z(n2094) );
  XNOR U2880 ( .A(n4402), .B(n[27]), .Z(n2092) );
  XOR U2881 ( .A(y[26]), .B(n1945), .Z(n1946) );
  ANDN U2882 ( .B(n1946), .A(n2868), .Z(n1947) );
  XNOR U2883 ( .A(zin[25]), .B(n1947), .Z(n4230) );
  NAND U2884 ( .A(n4230), .B(n[26]), .Z(n2090) );
  XOR U2885 ( .A(n[26]), .B(n4230), .Z(n2088) );
  XOR U2886 ( .A(y[25]), .B(n1948), .Z(n1949) );
  ANDN U2887 ( .B(n1949), .A(n2868), .Z(n1950) );
  XNOR U2888 ( .A(zin[24]), .B(n1950), .Z(n4234) );
  NAND U2889 ( .A(n[25]), .B(n4234), .Z(n2086) );
  XOR U2890 ( .A(n4234), .B(n[25]), .Z(n2084) );
  IV U2891 ( .A(n[24]), .Z(n4239) );
  XOR U2892 ( .A(y[24]), .B(n1951), .Z(n1952) );
  ANDN U2893 ( .B(n1952), .A(n2868), .Z(n1953) );
  XNOR U2894 ( .A(zin[23]), .B(n1953), .Z(n4238) );
  NANDN U2895 ( .A(n4239), .B(n4238), .Z(n2949) );
  XNOR U2896 ( .A(n4238), .B(n4239), .Z(n2081) );
  IV U2897 ( .A(n[23]), .Z(n4387) );
  XOR U2898 ( .A(y[23]), .B(n1954), .Z(n1955) );
  ANDN U2899 ( .B(n1955), .A(n2868), .Z(n1956) );
  XNOR U2900 ( .A(zin[22]), .B(n1956), .Z(n4390) );
  NANDN U2901 ( .A(n4387), .B(n4390), .Z(n2946) );
  XNOR U2902 ( .A(n4387), .B(n4390), .Z(n2078) );
  IV U2903 ( .A(n[22]), .Z(n4382) );
  XOR U2904 ( .A(y[22]), .B(n1957), .Z(n1958) );
  ANDN U2905 ( .B(n1958), .A(n2868), .Z(n1959) );
  XNOR U2906 ( .A(zin[21]), .B(n1959), .Z(n4243) );
  NANDN U2907 ( .A(n4382), .B(n4243), .Z(n2943) );
  XNOR U2908 ( .A(n4243), .B(n4382), .Z(n2075) );
  XOR U2909 ( .A(y[21]), .B(n1960), .Z(n1961) );
  ANDN U2910 ( .B(n1961), .A(n2868), .Z(n1962) );
  XNOR U2911 ( .A(zin[20]), .B(n1962), .Z(n4381) );
  NAND U2912 ( .A(n[21]), .B(n4381), .Z(n2940) );
  XOR U2913 ( .A(n[21]), .B(n4381), .Z(n2072) );
  IV U2914 ( .A(n[20]), .Z(n4248) );
  XOR U2915 ( .A(y[20]), .B(n1963), .Z(n1964) );
  ANDN U2916 ( .B(n1964), .A(n2868), .Z(n1965) );
  XNOR U2917 ( .A(zin[19]), .B(n1965), .Z(n4247) );
  NANDN U2918 ( .A(n4248), .B(n4247), .Z(n2937) );
  XNOR U2919 ( .A(n4247), .B(n4248), .Z(n2069) );
  IV U2920 ( .A(n[19]), .Z(n4370) );
  XOR U2921 ( .A(y[19]), .B(n1966), .Z(n1967) );
  ANDN U2922 ( .B(n1967), .A(n2868), .Z(n1968) );
  XNOR U2923 ( .A(zin[18]), .B(n1968), .Z(n4252) );
  NANDN U2924 ( .A(n4370), .B(n4252), .Z(n2934) );
  XNOR U2925 ( .A(n4370), .B(n4252), .Z(n2066) );
  IV U2926 ( .A(n[18]), .Z(n4257) );
  XOR U2927 ( .A(y[18]), .B(n1969), .Z(n1970) );
  ANDN U2928 ( .B(n1970), .A(n2868), .Z(n1971) );
  XNOR U2929 ( .A(zin[17]), .B(n1971), .Z(n4256) );
  NANDN U2930 ( .A(n4257), .B(n4256), .Z(n2931) );
  XNOR U2931 ( .A(n4257), .B(n4256), .Z(n2063) );
  XOR U2932 ( .A(y[17]), .B(n1972), .Z(n1973) );
  ANDN U2933 ( .B(n1973), .A(n2868), .Z(n1974) );
  XOR U2934 ( .A(zin[16]), .B(n1974), .Z(n4261) );
  ANDN U2935 ( .B(n[17]), .A(n4261), .Z(n2928) );
  XOR U2936 ( .A(y[16]), .B(n1975), .Z(n1976) );
  ANDN U2937 ( .B(n1976), .A(n2868), .Z(n1977) );
  XOR U2938 ( .A(zin[15]), .B(n1977), .Z(n4265) );
  IV U2939 ( .A(n[16]), .Z(n4266) );
  AND U2940 ( .A(n4265), .B(n4266), .Z(n2923) );
  IV U2941 ( .A(n[17]), .Z(n4362) );
  AND U2942 ( .A(n4261), .B(n4362), .Z(n2926) );
  NOR U2943 ( .A(n2923), .B(n2926), .Z(n2060) );
  ANDN U2944 ( .B(n[16]), .A(n4265), .Z(n2925) );
  XOR U2945 ( .A(y[15]), .B(n1978), .Z(n1979) );
  ANDN U2946 ( .B(n1979), .A(n2868), .Z(n1980) );
  XNOR U2947 ( .A(zin[14]), .B(n1980), .Z(n4361) );
  NOR U2948 ( .A(n[15]), .B(n4361), .Z(n2920) );
  XOR U2949 ( .A(y[13]), .B(n1981), .Z(n1982) );
  ANDN U2950 ( .B(n1982), .A(n2868), .Z(n1983) );
  XOR U2951 ( .A(zin[12]), .B(n1983), .Z(n4275) );
  ANDN U2952 ( .B(n[13]), .A(n4275), .Z(n2916) );
  XOR U2953 ( .A(y[12]), .B(n1984), .Z(n1985) );
  ANDN U2954 ( .B(n1985), .A(n2868), .Z(n1986) );
  XOR U2955 ( .A(zin[11]), .B(n1986), .Z(n4348) );
  IV U2956 ( .A(n4348), .Z(n1987) );
  AND U2957 ( .A(n[12]), .B(n1987), .Z(n2913) );
  NOR U2958 ( .A(n1987), .B(n[12]), .Z(n2911) );
  XOR U2959 ( .A(y[11]), .B(n1988), .Z(n1989) );
  ANDN U2960 ( .B(n1989), .A(n2868), .Z(n1990) );
  XOR U2961 ( .A(zin[10]), .B(n1990), .Z(n4341) );
  ANDN U2962 ( .B(n[11]), .A(n4341), .Z(n2910) );
  IV U2963 ( .A(n[11]), .Z(n4337) );
  AND U2964 ( .A(n4341), .B(n4337), .Z(n2908) );
  XOR U2965 ( .A(y[7]), .B(n1991), .Z(n1992) );
  ANDN U2966 ( .B(n1992), .A(n2868), .Z(n1993) );
  XNOR U2967 ( .A(zin[6]), .B(n1993), .Z(n4283) );
  AND U2968 ( .A(n4283), .B(n[7]), .Z(n2896) );
  OR U2969 ( .A(n4283), .B(n[7]), .Z(n2897) );
  XOR U2970 ( .A(y[6]), .B(n1994), .Z(n1995) );
  ANDN U2971 ( .B(n1995), .A(n2868), .Z(n1996) );
  XNOR U2972 ( .A(zin[5]), .B(n1996), .Z(n4287) );
  OR U2973 ( .A(n4287), .B(n[6]), .Z(n2893) );
  AND U2974 ( .A(n2897), .B(n2893), .Z(n2026) );
  XOR U2975 ( .A(y[4]), .B(n1997), .Z(n1998) );
  ANDN U2976 ( .B(n1998), .A(n2868), .Z(n1999) );
  XNOR U2977 ( .A(zin[3]), .B(n1999), .Z(n4295) );
  OR U2978 ( .A(n4295), .B(n[4]), .Z(n2887) );
  XOR U2979 ( .A(y[3]), .B(n2000), .Z(n2001) );
  ANDN U2980 ( .B(n2001), .A(n2868), .Z(n2002) );
  XNOR U2981 ( .A(zin[2]), .B(n2002), .Z(n4307) );
  OR U2982 ( .A(n4307), .B(n[3]), .Z(n2884) );
  AND U2983 ( .A(n2887), .B(n2884), .Z(n2017) );
  IV U2984 ( .A(n[2]), .Z(n6616) );
  XNOR U2985 ( .A(y[2]), .B(n2003), .Z(n2004) );
  ANDN U2986 ( .B(n2004), .A(n2868), .Z(n2005) );
  XNOR U2987 ( .A(zin[1]), .B(n2005), .Z(n4303) );
  NANDN U2988 ( .A(n6616), .B(n4303), .Z(n2014) );
  XNOR U2989 ( .A(n6616), .B(n4303), .Z(n2012) );
  NANDN U2990 ( .A(n[0]), .B(n2880), .Z(n2007) );
  NAND U2991 ( .A(n[1]), .B(n2007), .Z(n2010) );
  NANDN U2992 ( .A(n2868), .B(y[1]), .Z(n2006) );
  XNOR U2993 ( .A(zin[0]), .B(n2006), .Z(n4299) );
  XOR U2994 ( .A(n2007), .B(n[1]), .Z(n2008) );
  NANDN U2995 ( .A(n4299), .B(n2008), .Z(n2009) );
  NAND U2996 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U2997 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2998 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U2999 ( .A(n[3]), .B(n4307), .Z(n2886) );
  NANDN U3000 ( .A(n2015), .B(n2886), .Z(n2016) );
  AND U3001 ( .A(n2017), .B(n2016), .Z(n2018) );
  NAND U3002 ( .A(n[4]), .B(n4295), .Z(n2889) );
  NANDN U3003 ( .A(n2018), .B(n2889), .Z(n2022) );
  XOR U3004 ( .A(y[5]), .B(n2019), .Z(n2020) );
  ANDN U3005 ( .B(n2020), .A(n2868), .Z(n2021) );
  XOR U3006 ( .A(zin[4]), .B(n2021), .Z(n4291) );
  NANDN U3007 ( .A(n[5]), .B(n4291), .Z(n2890) );
  NAND U3008 ( .A(n2022), .B(n2890), .Z(n2023) );
  NAND U3009 ( .A(n[6]), .B(n4287), .Z(n2895) );
  NAND U3010 ( .A(n2023), .B(n2895), .Z(n2024) );
  NANDN U3011 ( .A(n4291), .B(n[5]), .Z(n2892) );
  NANDN U3012 ( .A(n2024), .B(n2892), .Z(n2025) );
  AND U3013 ( .A(n2026), .B(n2025), .Z(n2027) );
  OR U3014 ( .A(n2896), .B(n2027), .Z(n2031) );
  XOR U3015 ( .A(y[8]), .B(n2028), .Z(n2029) );
  ANDN U3016 ( .B(n2029), .A(n2868), .Z(n2030) );
  XOR U3017 ( .A(zin[7]), .B(n2030), .Z(n4279) );
  NANDN U3018 ( .A(n[8]), .B(n4279), .Z(n2900) );
  NAND U3019 ( .A(n2031), .B(n2900), .Z(n2032) );
  ANDN U3020 ( .B(n[8]), .A(n4279), .Z(n2899) );
  ANDN U3021 ( .B(n2032), .A(n2899), .Z(n2040) );
  XNOR U3022 ( .A(y[9]), .B(n2033), .Z(n2034) );
  ANDN U3023 ( .B(n2034), .A(n2868), .Z(n2035) );
  XNOR U3024 ( .A(zin[8]), .B(n2035), .Z(n4329) );
  NANDN U3025 ( .A(n2040), .B(n4329), .Z(n2039) );
  XOR U3026 ( .A(y[10]), .B(n2036), .Z(n2037) );
  ANDN U3027 ( .B(n2037), .A(n2868), .Z(n2038) );
  XNOR U3028 ( .A(zin[9]), .B(n2038), .Z(n4333) );
  AND U3029 ( .A(n4333), .B(n[10]), .Z(n2907) );
  ANDN U3030 ( .B(n2039), .A(n2907), .Z(n2043) );
  IV U3031 ( .A(n[9]), .Z(n6868) );
  XNOR U3032 ( .A(n4329), .B(n2040), .Z(n2041) );
  NANDN U3033 ( .A(n6868), .B(n2041), .Z(n2042) );
  NAND U3034 ( .A(n2043), .B(n2042), .Z(n2044) );
  NOR U3035 ( .A(n[10]), .B(n4333), .Z(n2905) );
  ANDN U3036 ( .B(n2044), .A(n2905), .Z(n2045) );
  NANDN U3037 ( .A(n2908), .B(n2045), .Z(n2046) );
  NANDN U3038 ( .A(n2910), .B(n2046), .Z(n2047) );
  NANDN U3039 ( .A(n2911), .B(n2047), .Z(n2048) );
  NANDN U3040 ( .A(n2913), .B(n2048), .Z(n2049) );
  IV U3041 ( .A(n[13]), .Z(n4349) );
  AND U3042 ( .A(n4275), .B(n4349), .Z(n2914) );
  ANDN U3043 ( .B(n2049), .A(n2914), .Z(n2053) );
  XOR U3044 ( .A(y[14]), .B(n2050), .Z(n2051) );
  ANDN U3045 ( .B(n2051), .A(n2868), .Z(n2052) );
  XOR U3046 ( .A(zin[13]), .B(n2052), .Z(n4270) );
  ANDN U3047 ( .B(n[14]), .A(n4270), .Z(n2919) );
  NOR U3048 ( .A(n2053), .B(n2919), .Z(n2054) );
  NANDN U3049 ( .A(n2916), .B(n2054), .Z(n2055) );
  IV U3050 ( .A(n[14]), .Z(n4271) );
  AND U3051 ( .A(n4270), .B(n4271), .Z(n2917) );
  ANDN U3052 ( .B(n2055), .A(n2917), .Z(n2056) );
  NANDN U3053 ( .A(n2920), .B(n2056), .Z(n2057) );
  AND U3054 ( .A(n4361), .B(n[15]), .Z(n2922) );
  ANDN U3055 ( .B(n2057), .A(n2922), .Z(n2058) );
  NANDN U3056 ( .A(n2925), .B(n2058), .Z(n2059) );
  NAND U3057 ( .A(n2060), .B(n2059), .Z(n2061) );
  NANDN U3058 ( .A(n2928), .B(n2061), .Z(n2062) );
  NAND U3059 ( .A(n2063), .B(n2062), .Z(n2064) );
  NAND U3060 ( .A(n2931), .B(n2064), .Z(n2065) );
  NAND U3061 ( .A(n2066), .B(n2065), .Z(n2067) );
  NAND U3062 ( .A(n2934), .B(n2067), .Z(n2068) );
  NAND U3063 ( .A(n2069), .B(n2068), .Z(n2070) );
  NAND U3064 ( .A(n2937), .B(n2070), .Z(n2071) );
  NAND U3065 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U3066 ( .A(n2940), .B(n2073), .Z(n2074) );
  NAND U3067 ( .A(n2075), .B(n2074), .Z(n2076) );
  NAND U3068 ( .A(n2943), .B(n2076), .Z(n2077) );
  NAND U3069 ( .A(n2078), .B(n2077), .Z(n2079) );
  NAND U3070 ( .A(n2946), .B(n2079), .Z(n2080) );
  NAND U3071 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U3072 ( .A(n2949), .B(n2082), .Z(n2083) );
  NAND U3073 ( .A(n2084), .B(n2083), .Z(n2085) );
  NAND U3074 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U3075 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U3076 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U3077 ( .A(n2092), .B(n2091), .Z(n2093) );
  NAND U3078 ( .A(n2094), .B(n2093), .Z(n2095) );
  NAND U3079 ( .A(n2096), .B(n2095), .Z(n2097) );
  NAND U3080 ( .A(n2952), .B(n2097), .Z(n2098) );
  NAND U3081 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U3082 ( .A(n2955), .B(n2100), .Z(n2101) );
  NAND U3083 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U3084 ( .A(n2958), .B(n2103), .Z(n2104) );
  NAND U3085 ( .A(n2105), .B(n2104), .Z(n2106) );
  NAND U3086 ( .A(n2961), .B(n2106), .Z(n2107) );
  NAND U3087 ( .A(n2108), .B(n2107), .Z(n2109) );
  NAND U3088 ( .A(n2110), .B(n2109), .Z(n2111) );
  NAND U3089 ( .A(n2112), .B(n2111), .Z(n2113) );
  NAND U3090 ( .A(n2114), .B(n2113), .Z(n2115) );
  NAND U3091 ( .A(n2116), .B(n2115), .Z(n2117) );
  AND U3092 ( .A(n2118), .B(n2117), .Z(n2122) );
  XOR U3093 ( .A(y[35]), .B(n2119), .Z(n2120) );
  ANDN U3094 ( .B(n2120), .A(n2868), .Z(n2121) );
  XNOR U3095 ( .A(zin[34]), .B(n2121), .Z(n4431) );
  NANDN U3096 ( .A(n2122), .B(n4431), .Z(n2125) );
  IV U3097 ( .A(n[35]), .Z(n4432) );
  XNOR U3098 ( .A(n4431), .B(n2122), .Z(n2123) );
  NANDN U3099 ( .A(n4432), .B(n2123), .Z(n2124) );
  NAND U3100 ( .A(n2125), .B(n2124), .Z(n2126) );
  IV U3101 ( .A(n[36]), .Z(n6656) );
  ANDN U3102 ( .B(n6656), .A(n4205), .Z(n2964) );
  ANDN U3103 ( .B(n2126), .A(n2964), .Z(n2127) );
  OR U3104 ( .A(n2962), .B(n2127), .Z(n2128) );
  IV U3105 ( .A(n[37]), .Z(n4438) );
  ANDN U3106 ( .B(n4438), .A(n4201), .Z(n2967) );
  ANDN U3107 ( .B(n2128), .A(n2967), .Z(n2129) );
  OR U3108 ( .A(n2965), .B(n2129), .Z(n2130) );
  NANDN U3109 ( .A(n2970), .B(n2130), .Z(n2131) );
  AND U3110 ( .A(n4196), .B(n[38]), .Z(n2968) );
  ANDN U3111 ( .B(n2131), .A(n2968), .Z(n2133) );
  IV U3112 ( .A(n[39]), .Z(n4446) );
  OR U3113 ( .A(n2133), .B(n4446), .Z(n2132) );
  ANDN U3114 ( .B(n[40]), .A(n4187), .Z(n2974) );
  ANDN U3115 ( .B(n2132), .A(n2974), .Z(n2139) );
  XOR U3116 ( .A(n4446), .B(n2133), .Z(n2137) );
  XOR U3117 ( .A(y[39]), .B(n2134), .Z(n2135) );
  ANDN U3118 ( .B(n2135), .A(n2868), .Z(n2136) );
  XNOR U3119 ( .A(zin[38]), .B(n2136), .Z(n4192) );
  NAND U3120 ( .A(n2137), .B(n4192), .Z(n2138) );
  NAND U3121 ( .A(n2139), .B(n2138), .Z(n2140) );
  NAND U3122 ( .A(n2141), .B(n2140), .Z(n2142) );
  NANDN U3123 ( .A(n2979), .B(n2142), .Z(n2143) );
  NANDN U3124 ( .A(n2980), .B(n2143), .Z(n2144) );
  NANDN U3125 ( .A(n2982), .B(n2144), .Z(n2145) );
  NOR U3126 ( .A(n[43]), .B(n4466), .Z(n2983) );
  ANDN U3127 ( .B(n2145), .A(n2983), .Z(n2146) );
  OR U3128 ( .A(n2985), .B(n2146), .Z(n2147) );
  NANDN U3129 ( .A(n2988), .B(n2147), .Z(n2148) );
  AND U3130 ( .A(n4470), .B(n[44]), .Z(n2986) );
  ANDN U3131 ( .B(n2148), .A(n2986), .Z(n2153) );
  XOR U3132 ( .A(y[45]), .B(n2149), .Z(n2150) );
  ANDN U3133 ( .B(n2150), .A(n2868), .Z(n2151) );
  XNOR U3134 ( .A(zin[44]), .B(n2151), .Z(n4474) );
  NANDN U3135 ( .A(n2153), .B(n4474), .Z(n2152) );
  ANDN U3136 ( .B(n2152), .A(n2989), .Z(n2156) );
  XNOR U3137 ( .A(n4474), .B(n2153), .Z(n2154) );
  NAND U3138 ( .A(n[45]), .B(n2154), .Z(n2155) );
  NAND U3139 ( .A(n2156), .B(n2155), .Z(n2157) );
  NAND U3140 ( .A(n2158), .B(n2157), .Z(n2159) );
  NANDN U3141 ( .A(n2992), .B(n2159), .Z(n2160) );
  NANDN U3142 ( .A(n[48]), .B(n4166), .Z(n2995) );
  NAND U3143 ( .A(n2160), .B(n2995), .Z(n2161) );
  NANDN U3144 ( .A(n2997), .B(n2161), .Z(n2162) );
  NOR U3145 ( .A(n[49]), .B(n4161), .Z(n2998) );
  ANDN U3146 ( .B(n2162), .A(n2998), .Z(n2163) );
  OR U3147 ( .A(n3000), .B(n2163), .Z(n2164) );
  NANDN U3148 ( .A(n3001), .B(n2164), .Z(n2166) );
  AND U3149 ( .A(n[50]), .B(n2165), .Z(n3003) );
  ANDN U3150 ( .B(n2166), .A(n3003), .Z(n2170) );
  XOR U3151 ( .A(y[51]), .B(n2167), .Z(n2168) );
  ANDN U3152 ( .B(n2168), .A(n2868), .Z(n2169) );
  XNOR U3153 ( .A(zin[50]), .B(n2169), .Z(n4153) );
  NANDN U3154 ( .A(n2170), .B(n4153), .Z(n2173) );
  XNOR U3155 ( .A(n4153), .B(n2170), .Z(n2171) );
  NAND U3156 ( .A(n[51]), .B(n2171), .Z(n2172) );
  NAND U3157 ( .A(n2173), .B(n2172), .Z(n2174) );
  AND U3158 ( .A(n3004), .B(n2174), .Z(n2175) );
  OR U3159 ( .A(n3006), .B(n2175), .Z(n2176) );
  NANDN U3160 ( .A(n3007), .B(n2176), .Z(n2177) );
  NANDN U3161 ( .A(n3009), .B(n2177), .Z(n2178) );
  NANDN U3162 ( .A(n3012), .B(n2178), .Z(n2179) );
  NANDN U3163 ( .A(n3010), .B(n2179), .Z(n2180) );
  NOR U3164 ( .A(n[55]), .B(n4135), .Z(n3015) );
  ANDN U3165 ( .B(n2180), .A(n3015), .Z(n2181) );
  OR U3166 ( .A(n3013), .B(n2181), .Z(n2182) );
  NANDN U3167 ( .A(n3018), .B(n2182), .Z(n2183) );
  AND U3168 ( .A(n4130), .B(n[56]), .Z(n3016) );
  ANDN U3169 ( .B(n2183), .A(n3016), .Z(n2185) );
  NANDN U3170 ( .A(n2185), .B(n[57]), .Z(n2184) );
  ANDN U3171 ( .B(n[58]), .A(n4122), .Z(n3021) );
  ANDN U3172 ( .B(n2184), .A(n3021), .Z(n2191) );
  XNOR U3173 ( .A(n[57]), .B(n2185), .Z(n2189) );
  XOR U3174 ( .A(y[57]), .B(n2186), .Z(n2187) );
  ANDN U3175 ( .B(n2187), .A(n2868), .Z(n2188) );
  XNOR U3176 ( .A(zin[56]), .B(n2188), .Z(n4126) );
  NAND U3177 ( .A(n2189), .B(n4126), .Z(n2190) );
  NAND U3178 ( .A(n2191), .B(n2190), .Z(n2192) );
  NAND U3179 ( .A(n2193), .B(n2192), .Z(n2194) );
  ANDN U3180 ( .B(n[59]), .A(n4117), .Z(n3024) );
  ANDN U3181 ( .B(n2194), .A(n3024), .Z(n2196) );
  IV U3182 ( .A(n[60]), .Z(n4113) );
  OR U3183 ( .A(n2196), .B(n4113), .Z(n2195) );
  ANDN U3184 ( .B(n[61]), .A(n4107), .Z(n3028) );
  ANDN U3185 ( .B(n2195), .A(n3028), .Z(n2202) );
  XOR U3186 ( .A(n4113), .B(n2196), .Z(n2200) );
  XOR U3187 ( .A(y[60]), .B(n2197), .Z(n2198) );
  ANDN U3188 ( .B(n2198), .A(n2868), .Z(n2199) );
  XNOR U3189 ( .A(zin[59]), .B(n2199), .Z(n4112) );
  NAND U3190 ( .A(n2200), .B(n4112), .Z(n2201) );
  NAND U3191 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U3192 ( .A(n2204), .B(n2203), .Z(n2205) );
  ANDN U3193 ( .B(n[62]), .A(n4103), .Z(n3033) );
  ANDN U3194 ( .B(n2205), .A(n3033), .Z(n2210) );
  XOR U3195 ( .A(y[63]), .B(n2206), .Z(n2207) );
  ANDN U3196 ( .B(n2207), .A(n2868), .Z(n2208) );
  XNOR U3197 ( .A(zin[62]), .B(n2208), .Z(n4099) );
  NANDN U3198 ( .A(n2210), .B(n4099), .Z(n2209) );
  ANDN U3199 ( .B(n[64]), .A(n4095), .Z(n3034) );
  ANDN U3200 ( .B(n2209), .A(n3034), .Z(n2213) );
  XNOR U3201 ( .A(n4099), .B(n2210), .Z(n2211) );
  NAND U3202 ( .A(n[63]), .B(n2211), .Z(n2212) );
  NAND U3203 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U3204 ( .A(n2215), .B(n2214), .Z(n2216) );
  NANDN U3205 ( .A(n3037), .B(n2216), .Z(n2217) );
  NAND U3206 ( .A(n2218), .B(n2217), .Z(n2219) );
  NAND U3207 ( .A(n2220), .B(n2219), .Z(n2221) );
  NAND U3208 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U3209 ( .A(n2224), .B(n2223), .Z(n2225) );
  IV U3210 ( .A(n[68]), .Z(n4078) );
  ANDN U3211 ( .B(n4078), .A(n4077), .Z(n3042) );
  ANDN U3212 ( .B(n2225), .A(n3042), .Z(n2226) );
  NAND U3213 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U3214 ( .A(n2229), .B(n2228), .Z(n2230) );
  NAND U3215 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U3216 ( .A(n3045), .B(n2232), .Z(n2233) );
  NAND U3217 ( .A(n2234), .B(n2233), .Z(n2235) );
  NAND U3218 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U3219 ( .A(n2238), .B(n2237), .Z(n2239) );
  NAND U3220 ( .A(n2240), .B(n2239), .Z(n2241) );
  NAND U3221 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U3222 ( .A(n2244), .B(n2243), .Z(n2245) );
  NAND U3223 ( .A(n2246), .B(n2245), .Z(n2247) );
  NAND U3224 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U3225 ( .A(n2250), .B(n2249), .Z(n2251) );
  NAND U3226 ( .A(n2252), .B(n2251), .Z(n2253) );
  NAND U3227 ( .A(n2254), .B(n2253), .Z(n2255) );
  NAND U3228 ( .A(n2256), .B(n2255), .Z(n2257) );
  NAND U3229 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U3230 ( .A(n3054), .B(n2259), .Z(n2260) );
  NAND U3231 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U3232 ( .A(n2263), .B(n2262), .Z(n2264) );
  NAND U3233 ( .A(n2265), .B(n2264), .Z(n2266) );
  NAND U3234 ( .A(n2267), .B(n2266), .Z(n2268) );
  NAND U3235 ( .A(n2269), .B(n2268), .Z(n2270) );
  NAND U3236 ( .A(n3057), .B(n2270), .Z(n2271) );
  NAND U3237 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U3238 ( .A(n3060), .B(n2273), .Z(n2274) );
  NAND U3239 ( .A(n2275), .B(n2274), .Z(n2276) );
  NAND U3240 ( .A(n2277), .B(n2276), .Z(n2278) );
  NAND U3241 ( .A(n2279), .B(n2278), .Z(n2280) );
  NAND U3242 ( .A(n2281), .B(n2280), .Z(n2282) );
  NAND U3243 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U3244 ( .A(n2285), .B(n2284), .Z(n2286) );
  NAND U3245 ( .A(n2287), .B(n2286), .Z(n2288) );
  NAND U3246 ( .A(n3063), .B(n2288), .Z(n2289) );
  NAND U3247 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U3248 ( .A(n2292), .B(n2291), .Z(n2293) );
  NAND U3249 ( .A(n2294), .B(n2293), .Z(n2295) );
  NAND U3250 ( .A(n3066), .B(n2295), .Z(n2296) );
  NAND U3251 ( .A(n2297), .B(n2296), .Z(n2298) );
  NAND U3252 ( .A(n2299), .B(n2298), .Z(n2300) );
  NAND U3253 ( .A(n2301), .B(n2300), .Z(n2302) );
  NAND U3254 ( .A(n3069), .B(n2302), .Z(n2303) );
  NAND U3255 ( .A(n2304), .B(n2303), .Z(n2305) );
  NAND U3256 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U3257 ( .A(n2308), .B(n2307), .Z(n2309) );
  NAND U3258 ( .A(n3072), .B(n2309), .Z(n2310) );
  NAND U3259 ( .A(n2311), .B(n2310), .Z(n2312) );
  NAND U3260 ( .A(n3075), .B(n2312), .Z(n2313) );
  NAND U3261 ( .A(n2314), .B(n2313), .Z(n2315) );
  NAND U3262 ( .A(n3078), .B(n2315), .Z(n2316) );
  NAND U3263 ( .A(n2317), .B(n2316), .Z(n2318) );
  NAND U3264 ( .A(n3081), .B(n2318), .Z(n2319) );
  NAND U3265 ( .A(n2320), .B(n2319), .Z(n2321) );
  NAND U3266 ( .A(n3084), .B(n2321), .Z(n2322) );
  NAND U3267 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U3268 ( .A(n3090), .B(n2325), .Z(n2326) );
  NAND U3269 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U3270 ( .A(n2329), .B(n2328), .Z(n2330) );
  NAND U3271 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U3272 ( .A(n3093), .B(n2332), .Z(n2333) );
  NAND U3273 ( .A(n2334), .B(n2333), .Z(n2335) );
  NAND U3274 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U3275 ( .A(n2338), .B(n2337), .Z(n2339) );
  NAND U3276 ( .A(n2340), .B(n2339), .Z(n2341) );
  NAND U3277 ( .A(n2342), .B(n2341), .Z(n2343) );
  NAND U3278 ( .A(n2344), .B(n2343), .Z(n2345) );
  NAND U3279 ( .A(n2346), .B(n2345), .Z(n2347) );
  NAND U3280 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U3281 ( .A(n2350), .B(n2349), .Z(n2351) );
  NAND U3282 ( .A(n3096), .B(n2351), .Z(n2352) );
  NAND U3283 ( .A(n2353), .B(n2352), .Z(n2354) );
  NAND U3284 ( .A(n3099), .B(n2354), .Z(n2355) );
  NAND U3285 ( .A(n2356), .B(n2355), .Z(n2357) );
  NAND U3286 ( .A(n3102), .B(n2357), .Z(n2358) );
  NAND U3287 ( .A(n2359), .B(n2358), .Z(n2360) );
  NAND U3288 ( .A(n3105), .B(n2360), .Z(n2361) );
  NAND U3289 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U3290 ( .A(n3108), .B(n2363), .Z(n2364) );
  NAND U3291 ( .A(n2365), .B(n2364), .Z(n2366) );
  NAND U3292 ( .A(n3111), .B(n2366), .Z(n2367) );
  NAND U3293 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U3294 ( .A(n3114), .B(n2369), .Z(n2370) );
  NAND U3295 ( .A(n2371), .B(n2370), .Z(n2372) );
  NAND U3296 ( .A(n3117), .B(n2372), .Z(n2373) );
  NAND U3297 ( .A(n2374), .B(n2373), .Z(n2375) );
  NAND U3298 ( .A(n3120), .B(n2375), .Z(n2376) );
  NAND U3299 ( .A(n2377), .B(n2376), .Z(n2378) );
  NAND U3300 ( .A(n3123), .B(n2378), .Z(n2379) );
  NAND U3301 ( .A(n2380), .B(n2379), .Z(n2381) );
  NAND U3302 ( .A(n3126), .B(n2381), .Z(n2382) );
  NAND U3303 ( .A(n2383), .B(n2382), .Z(n2384) );
  NAND U3304 ( .A(n3129), .B(n2384), .Z(n2385) );
  NAND U3305 ( .A(n2386), .B(n2385), .Z(n2387) );
  NAND U3306 ( .A(n3132), .B(n2387), .Z(n2388) );
  NAND U3307 ( .A(n2389), .B(n2388), .Z(n2390) );
  NAND U3308 ( .A(n3135), .B(n2390), .Z(n2391) );
  NAND U3309 ( .A(n2392), .B(n2391), .Z(n2393) );
  NAND U3310 ( .A(n3138), .B(n2393), .Z(n2394) );
  NAND U3311 ( .A(n2395), .B(n2394), .Z(n2396) );
  NAND U3312 ( .A(n3141), .B(n2396), .Z(n2397) );
  NAND U3313 ( .A(n2398), .B(n2397), .Z(n2399) );
  NAND U3314 ( .A(n2400), .B(n2399), .Z(n2401) );
  NAND U3315 ( .A(n2402), .B(n2401), .Z(n2403) );
  NAND U3316 ( .A(n3144), .B(n2403), .Z(n2404) );
  NAND U3317 ( .A(n2405), .B(n2404), .Z(n2406) );
  NAND U3318 ( .A(n2407), .B(n2406), .Z(n2408) );
  NAND U3319 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U3320 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U3321 ( .A(n2413), .B(n2412), .Z(n2414) );
  NAND U3322 ( .A(n3147), .B(n2414), .Z(n2415) );
  NAND U3323 ( .A(n2416), .B(n2415), .Z(n2417) );
  NAND U3324 ( .A(n2418), .B(n2417), .Z(n2419) );
  NAND U3325 ( .A(n2420), .B(n2419), .Z(n2421) );
  NAND U3326 ( .A(n3150), .B(n2421), .Z(n2422) );
  NAND U3327 ( .A(n2423), .B(n2422), .Z(n2424) );
  NAND U3328 ( .A(n3153), .B(n2424), .Z(n2425) );
  NAND U3329 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U3330 ( .A(n2428), .B(n2427), .Z(n2429) );
  NAND U3331 ( .A(n2430), .B(n2429), .Z(n2431) );
  NAND U3332 ( .A(n3156), .B(n2431), .Z(n2432) );
  NAND U3333 ( .A(n2433), .B(n2432), .Z(n2434) );
  NAND U3334 ( .A(n2435), .B(n2434), .Z(n2436) );
  NAND U3335 ( .A(n2437), .B(n2436), .Z(n2438) );
  NAND U3336 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U3337 ( .A(n2441), .B(n2440), .Z(n2442) );
  NAND U3338 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U3339 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U3340 ( .A(n2447), .B(n2446), .Z(n2448) );
  NAND U3341 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U3342 ( .A(n2451), .B(n2450), .Z(n2452) );
  NAND U3343 ( .A(n2453), .B(n2452), .Z(n2454) );
  NAND U3344 ( .A(n2455), .B(n2454), .Z(n2456) );
  NAND U3345 ( .A(n2457), .B(n2456), .Z(n2458) );
  NAND U3346 ( .A(n3159), .B(n2458), .Z(n2459) );
  NAND U3347 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U3348 ( .A(n2462), .B(n2461), .Z(n2463) );
  NAND U3349 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U3350 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U3351 ( .A(n2468), .B(n2467), .Z(n2469) );
  NAND U3352 ( .A(n2470), .B(n2469), .Z(n2471) );
  NAND U3353 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U3354 ( .A(n3165), .B(n2473), .Z(n2474) );
  NAND U3355 ( .A(n2475), .B(n2474), .Z(n2476) );
  NAND U3356 ( .A(n3168), .B(n2476), .Z(n2477) );
  NAND U3357 ( .A(n2478), .B(n2477), .Z(n2479) );
  NAND U3358 ( .A(n2480), .B(n2479), .Z(n2481) );
  NAND U3359 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U3360 ( .A(n3171), .B(n2483), .Z(n2484) );
  NAND U3361 ( .A(n2485), .B(n2484), .Z(n2486) );
  NAND U3362 ( .A(n2487), .B(n2486), .Z(n2488) );
  NAND U3363 ( .A(n2489), .B(n2488), .Z(n2490) );
  NAND U3364 ( .A(n2491), .B(n2490), .Z(n2492) );
  NAND U3365 ( .A(n2493), .B(n2492), .Z(n2494) );
  NAND U3366 ( .A(n2495), .B(n2494), .Z(n2496) );
  NAND U3367 ( .A(n2497), .B(n2496), .Z(n2498) );
  NAND U3368 ( .A(n3174), .B(n2498), .Z(n2499) );
  NAND U3369 ( .A(n2500), .B(n2499), .Z(n2501) );
  NAND U3370 ( .A(n2502), .B(n2501), .Z(n2503) );
  NAND U3371 ( .A(n2504), .B(n2503), .Z(n2505) );
  NAND U3372 ( .A(n3177), .B(n2505), .Z(n2506) );
  NAND U3373 ( .A(n2507), .B(n2506), .Z(n2508) );
  NAND U3374 ( .A(n3180), .B(n2508), .Z(n2509) );
  NAND U3375 ( .A(n2510), .B(n2509), .Z(n2511) );
  NAND U3376 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U3377 ( .A(n2514), .B(n2513), .Z(n2515) );
  NAND U3378 ( .A(n3183), .B(n2515), .Z(n2516) );
  NAND U3379 ( .A(n2517), .B(n2516), .Z(n2518) );
  NAND U3380 ( .A(n3186), .B(n2518), .Z(n2519) );
  NAND U3381 ( .A(n2520), .B(n2519), .Z(n2521) );
  NAND U3382 ( .A(n3189), .B(n2521), .Z(n2522) );
  NAND U3383 ( .A(n2523), .B(n2522), .Z(n2524) );
  NAND U3384 ( .A(n2525), .B(n2524), .Z(n2526) );
  NAND U3385 ( .A(n2527), .B(n2526), .Z(n2528) );
  NAND U3386 ( .A(n3192), .B(n2528), .Z(n2529) );
  NAND U3387 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U3388 ( .A(n2532), .B(n2531), .Z(n2533) );
  NAND U3389 ( .A(n2534), .B(n2533), .Z(n2535) );
  NAND U3390 ( .A(n2536), .B(n2535), .Z(n2537) );
  NAND U3391 ( .A(n2538), .B(n2537), .Z(n2539) );
  NAND U3392 ( .A(n2540), .B(n2539), .Z(n2541) );
  NAND U3393 ( .A(n2542), .B(n2541), .Z(n2543) );
  NAND U3394 ( .A(n3195), .B(n2543), .Z(n2544) );
  NAND U3395 ( .A(n2545), .B(n2544), .Z(n2546) );
  NAND U3396 ( .A(n3198), .B(n2546), .Z(n2547) );
  NAND U3397 ( .A(n2548), .B(n2547), .Z(n2549) );
  NAND U3398 ( .A(n3201), .B(n2549), .Z(n2550) );
  NAND U3399 ( .A(n2551), .B(n2550), .Z(n2552) );
  NAND U3400 ( .A(n3204), .B(n2552), .Z(n2553) );
  NAND U3401 ( .A(n2554), .B(n2553), .Z(n2555) );
  NAND U3402 ( .A(n3207), .B(n2555), .Z(n2556) );
  NAND U3403 ( .A(n2557), .B(n2556), .Z(n2558) );
  NAND U3404 ( .A(n2559), .B(n2558), .Z(n2560) );
  NAND U3405 ( .A(n2561), .B(n2560), .Z(n2562) );
  NAND U3406 ( .A(n3210), .B(n2562), .Z(n2563) );
  NAND U3407 ( .A(n2564), .B(n2563), .Z(n2565) );
  NAND U3408 ( .A(n3213), .B(n2565), .Z(n2566) );
  NAND U3409 ( .A(n2567), .B(n2566), .Z(n2568) );
  NAND U3410 ( .A(n3216), .B(n2568), .Z(n2569) );
  NAND U3411 ( .A(n2570), .B(n2569), .Z(n2571) );
  NAND U3412 ( .A(n3219), .B(n2571), .Z(n2572) );
  NAND U3413 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U3414 ( .A(n2575), .B(n2574), .Z(n2576) );
  NAND U3415 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U3416 ( .A(n3222), .B(n2578), .Z(n2579) );
  NAND U3417 ( .A(n2580), .B(n2579), .Z(n2581) );
  NAND U3418 ( .A(n2582), .B(n2581), .Z(n2583) );
  NAND U3419 ( .A(n2584), .B(n2583), .Z(n2585) );
  NAND U3420 ( .A(n3225), .B(n2585), .Z(n2586) );
  NAND U3421 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U3422 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U3423 ( .A(n2591), .B(n2590), .Z(n2592) );
  NAND U3424 ( .A(n2593), .B(n2592), .Z(n2594) );
  NAND U3425 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U3426 ( .A(n2597), .B(n2596), .Z(n2598) );
  NAND U3427 ( .A(n2599), .B(n2598), .Z(n2600) );
  NAND U3428 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U3429 ( .A(n2603), .B(n2602), .Z(n2604) );
  NAND U3430 ( .A(n2605), .B(n2604), .Z(n2606) );
  NAND U3431 ( .A(n2607), .B(n2606), .Z(n2608) );
  NAND U3432 ( .A(n3228), .B(n2608), .Z(n2609) );
  NAND U3433 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U3434 ( .A(n3231), .B(n2611), .Z(n2612) );
  NAND U3435 ( .A(n2613), .B(n2612), .Z(n2614) );
  NAND U3436 ( .A(n2615), .B(n2614), .Z(n2616) );
  NAND U3437 ( .A(n2617), .B(n2616), .Z(n2618) );
  NAND U3438 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U3439 ( .A(n2621), .B(n2620), .Z(n2622) );
  NAND U3440 ( .A(n3234), .B(n2622), .Z(n2623) );
  NAND U3441 ( .A(n2624), .B(n2623), .Z(n2625) );
  NAND U3442 ( .A(n3237), .B(n2625), .Z(n2626) );
  NAND U3443 ( .A(n2627), .B(n2626), .Z(n2628) );
  NAND U3444 ( .A(n2629), .B(n2628), .Z(n2630) );
  NAND U3445 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U3446 ( .A(n3240), .B(n2632), .Z(n2633) );
  NAND U3447 ( .A(n2634), .B(n2633), .Z(n2635) );
  NAND U3448 ( .A(n3243), .B(n2635), .Z(n2636) );
  NAND U3449 ( .A(n2637), .B(n2636), .Z(n2638) );
  NAND U3450 ( .A(n2639), .B(n2638), .Z(n2640) );
  NAND U3451 ( .A(n2641), .B(n2640), .Z(n2642) );
  NAND U3452 ( .A(n2643), .B(n2642), .Z(n2644) );
  NAND U3453 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U3454 ( .A(n2647), .B(n2646), .Z(n2648) );
  NAND U3455 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U3456 ( .A(n3246), .B(n2650), .Z(n2651) );
  NAND U3457 ( .A(n2652), .B(n2651), .Z(n2653) );
  NAND U3458 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U3459 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U3460 ( .A(n2658), .B(n2657), .Z(n2659) );
  NAND U3461 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U3462 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U3463 ( .A(n2664), .B(n2663), .Z(n2665) );
  NAND U3464 ( .A(n2666), .B(n2665), .Z(n2667) );
  NAND U3465 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U3466 ( .A(n3249), .B(n2669), .Z(n2670) );
  NAND U3467 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND U3468 ( .A(n3252), .B(n2672), .Z(n2673) );
  NAND U3469 ( .A(n2674), .B(n2673), .Z(n2675) );
  NAND U3470 ( .A(n2676), .B(n2675), .Z(n2677) );
  NAND U3471 ( .A(n2678), .B(n2677), .Z(n2679) );
  NAND U3472 ( .A(n3255), .B(n2679), .Z(n2680) );
  NAND U3473 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U3474 ( .A(n2683), .B(n2682), .Z(n2684) );
  NAND U3475 ( .A(n2685), .B(n2684), .Z(n2686) );
  NAND U3476 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U3477 ( .A(n2689), .B(n2688), .Z(n2690) );
  NAND U3478 ( .A(n3258), .B(n2690), .Z(n2691) );
  NAND U3479 ( .A(n2692), .B(n2691), .Z(n2693) );
  NAND U3480 ( .A(n2694), .B(n2693), .Z(n2695) );
  NAND U3481 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U3482 ( .A(n3261), .B(n2697), .Z(n2698) );
  NAND U3483 ( .A(n2699), .B(n2698), .Z(n2700) );
  NAND U3484 ( .A(n2701), .B(n2700), .Z(n2702) );
  NAND U3485 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U3486 ( .A(n2705), .B(n2704), .Z(n2706) );
  NAND U3487 ( .A(n2707), .B(n2706), .Z(n2708) );
  NAND U3488 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U3489 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U3490 ( .A(n2713), .B(n2712), .Z(n2714) );
  NAND U3491 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U3492 ( .A(n3264), .B(n2716), .Z(n2717) );
  NAND U3493 ( .A(n2718), .B(n2717), .Z(n2719) );
  NAND U3494 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U3495 ( .A(n2722), .B(n2721), .Z(n2723) );
  NAND U3496 ( .A(n2724), .B(n2723), .Z(n2725) );
  NAND U3497 ( .A(n2726), .B(n2725), .Z(n2727) );
  NAND U3498 ( .A(n2728), .B(n2727), .Z(n2729) );
  NAND U3499 ( .A(n2730), .B(n2729), .Z(n2731) );
  NAND U3500 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U3501 ( .A(n2734), .B(n2733), .Z(n2735) );
  NAND U3502 ( .A(n3267), .B(n2735), .Z(n2736) );
  NAND U3503 ( .A(n2737), .B(n2736), .Z(n2738) );
  NAND U3504 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND U3505 ( .A(n2741), .B(n2740), .Z(n2742) );
  NAND U3506 ( .A(n2743), .B(n2742), .Z(n2744) );
  NAND U3507 ( .A(n2745), .B(n2744), .Z(n2746) );
  NAND U3508 ( .A(n2747), .B(n2746), .Z(n2748) );
  NAND U3509 ( .A(n2749), .B(n2748), .Z(n2750) );
  NAND U3510 ( .A(n3270), .B(n2750), .Z(n2751) );
  NAND U3511 ( .A(n2752), .B(n2751), .Z(n2753) );
  NAND U3512 ( .A(n2754), .B(n2753), .Z(n2755) );
  NAND U3513 ( .A(n2756), .B(n2755), .Z(n2757) );
  NAND U3514 ( .A(n2758), .B(n2757), .Z(n2759) );
  NAND U3515 ( .A(n2760), .B(n2759), .Z(n2761) );
  NAND U3516 ( .A(n3273), .B(n2761), .Z(n2762) );
  NAND U3517 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U3518 ( .A(n2765), .B(n2764), .Z(n2766) );
  NAND U3519 ( .A(n2767), .B(n2766), .Z(n2768) );
  NAND U3520 ( .A(n2769), .B(n2768), .Z(n2770) );
  NAND U3521 ( .A(n2771), .B(n2770), .Z(n2772) );
  NAND U3522 ( .A(n2773), .B(n2772), .Z(n2774) );
  NAND U3523 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3524 ( .A(n2777), .B(n2776), .Z(n2778) );
  NAND U3525 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U3526 ( .A(n2781), .B(n2780), .Z(n2782) );
  NAND U3527 ( .A(n2783), .B(n2782), .Z(n2784) );
  NAND U3528 ( .A(n3279), .B(n2784), .Z(n2785) );
  NAND U3529 ( .A(n2786), .B(n2785), .Z(n2787) );
  NAND U3530 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U3531 ( .A(n2790), .B(n2789), .Z(n2791) );
  NAND U3532 ( .A(n2792), .B(n2791), .Z(n2793) );
  NAND U3533 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U3534 ( .A(n2796), .B(n2795), .Z(n2797) );
  NAND U3535 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U3536 ( .A(n2800), .B(n2799), .Z(n2801) );
  NAND U3537 ( .A(n2802), .B(n2801), .Z(n2803) );
  NAND U3538 ( .A(n2804), .B(n2803), .Z(n2805) );
  NAND U3539 ( .A(n2806), .B(n2805), .Z(n2807) );
  NAND U3540 ( .A(n2808), .B(n2807), .Z(n2809) );
  NAND U3541 ( .A(n2810), .B(n2809), .Z(n2811) );
  NAND U3542 ( .A(n2812), .B(n2811), .Z(n2813) );
  NAND U3543 ( .A(n2814), .B(n2813), .Z(n2815) );
  NAND U3544 ( .A(n3282), .B(n2815), .Z(n2816) );
  NAND U3545 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U3546 ( .A(n2819), .B(n2818), .Z(n2820) );
  NAND U3547 ( .A(n2821), .B(n2820), .Z(n2822) );
  NAND U3548 ( .A(n2823), .B(n2822), .Z(n2824) );
  NAND U3549 ( .A(n2825), .B(n2824), .Z(n2826) );
  NAND U3550 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U3551 ( .A(n2829), .B(n2828), .Z(n2830) );
  NAND U3552 ( .A(n2831), .B(n2830), .Z(n2832) );
  NAND U3553 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U3554 ( .A(n3285), .B(n2834), .Z(n2835) );
  NAND U3555 ( .A(n2836), .B(n2835), .Z(n2837) );
  NAND U3556 ( .A(n3288), .B(n2837), .Z(n2838) );
  NAND U3557 ( .A(n2839), .B(n2838), .Z(n2840) );
  NAND U3558 ( .A(n3291), .B(n2840), .Z(n2841) );
  NAND U3559 ( .A(n2842), .B(n2841), .Z(n2843) );
  NAND U3560 ( .A(n3294), .B(n2843), .Z(n2844) );
  NAND U3561 ( .A(n2845), .B(n2844), .Z(n2846) );
  NAND U3562 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U3563 ( .A(n2849), .B(n2848), .Z(n2850) );
  NAND U3564 ( .A(n3297), .B(n2850), .Z(n2851) );
  NAND U3565 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3566 ( .A(n2854), .B(n2853), .Z(n2855) );
  NAND U3567 ( .A(y[254]), .B(zin[253]), .Z(n2860) );
  XOR U3568 ( .A(zin[253]), .B(y[254]), .Z(n2858) );
  NAND U3569 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U3570 ( .A(n2860), .B(n2859), .Z(n2864) );
  XOR U3571 ( .A(y[255]), .B(n2864), .Z(n2861) );
  ANDN U3572 ( .B(n2861), .A(n2868), .Z(n2862) );
  XNOR U3573 ( .A(zin[254]), .B(n2862), .Z(n3308) );
  AND U3574 ( .A(y[255]), .B(zin[254]), .Z(n2866) );
  XOR U3575 ( .A(zin[254]), .B(y[255]), .Z(n2863) );
  AND U3576 ( .A(n2864), .B(n2863), .Z(n2865) );
  OR U3577 ( .A(n2866), .B(n2865), .Z(n2867) );
  NANDN U3578 ( .A(n2868), .B(n2867), .Z(n2870) );
  ANDN U3579 ( .B(zin[255]), .A(n2870), .Z(n2869) );
  XOR U3580 ( .A(n2869), .B(zin[256]), .Z(n3313) );
  XNOR U3581 ( .A(n2870), .B(zin[255]), .Z(n3312) );
  NANDN U3582 ( .A(n524), .B(n[0]), .Z(n2871) );
  XNOR U3583 ( .A(n2880), .B(n2871), .Z(n5342) );
  NOR U3584 ( .A(n[254]), .B(n3318), .Z(n3301) );
  NOR U3585 ( .A(n[252]), .B(n3326), .Z(n3298) );
  NOR U3586 ( .A(n[249]), .B(n3339), .Z(n3295) );
  NOR U3587 ( .A(n[247]), .B(n3347), .Z(n3292) );
  NOR U3588 ( .A(n[246]), .B(n3352), .Z(n3289) );
  NOR U3589 ( .A(n[245]), .B(n3356), .Z(n3286) );
  NOR U3590 ( .A(n[244]), .B(n3360), .Z(n3283) );
  NOR U3591 ( .A(n[239]), .B(n3381), .Z(n3280) );
  NOR U3592 ( .A(n[231]), .B(n3411), .Z(n3277) );
  IV U3593 ( .A(n2873), .Z(n3419) );
  OR U3594 ( .A(n[228]), .B(n3419), .Z(n3276) );
  ANDN U3595 ( .B(n[228]), .A(n2873), .Z(n3274) );
  NOR U3596 ( .A(n[225]), .B(n3431), .Z(n3271) );
  NOR U3597 ( .A(n[222]), .B(n3443), .Z(n3268) );
  NOR U3598 ( .A(n[218]), .B(n3459), .Z(n3265) );
  NOR U3599 ( .A(n[213]), .B(n3475), .Z(n3262) );
  NOR U3600 ( .A(n[208]), .B(n3498), .Z(n3259) );
  NOR U3601 ( .A(n[206]), .B(n3507), .Z(n3256) );
  NOR U3602 ( .A(n[203]), .B(n3520), .Z(n3253) );
  NOR U3603 ( .A(n[201]), .B(n3528), .Z(n3250) );
  NOR U3604 ( .A(n[200]), .B(n3533), .Z(n3247) );
  NOR U3605 ( .A(n[195]), .B(n3554), .Z(n3244) );
  NOR U3606 ( .A(n[191]), .B(n3572), .Z(n3241) );
  NOR U3607 ( .A(n[190]), .B(n3576), .Z(n3238) );
  NOR U3608 ( .A(n[188]), .B(n3585), .Z(n3235) );
  NOR U3609 ( .A(n[187]), .B(n3590), .Z(n3232) );
  NOR U3610 ( .A(n[184]), .B(n3598), .Z(n3229) );
  NOR U3611 ( .A(n[183]), .B(n3602), .Z(n3226) );
  NOR U3612 ( .A(n[177]), .B(n3623), .Z(n3223) );
  NOR U3613 ( .A(n[175]), .B(n3632), .Z(n3220) );
  NOR U3614 ( .A(n[173]), .B(n3640), .Z(n3217) );
  NOR U3615 ( .A(n[172]), .B(n3645), .Z(n3214) );
  NOR U3616 ( .A(n[171]), .B(n3650), .Z(n3211) );
  NOR U3617 ( .A(n[170]), .B(n3654), .Z(n3208) );
  NOR U3618 ( .A(n[168]), .B(n3663), .Z(n3205) );
  NOR U3619 ( .A(n[167]), .B(n3668), .Z(n3202) );
  NOR U3620 ( .A(n[166]), .B(n3672), .Z(n3199) );
  NOR U3621 ( .A(n[165]), .B(n3677), .Z(n3196) );
  NOR U3622 ( .A(n[164]), .B(n3681), .Z(n3193) );
  NOR U3623 ( .A(n[160]), .B(n3697), .Z(n3190) );
  NOR U3624 ( .A(n[158]), .B(n3706), .Z(n3187) );
  NOR U3625 ( .A(n[157]), .B(n4937), .Z(n3184) );
  NOR U3626 ( .A(n[156]), .B(n3710), .Z(n3181) );
  NOR U3627 ( .A(n[154]), .B(n3714), .Z(n3178) );
  NOR U3628 ( .A(n[153]), .B(n4913), .Z(n3175) );
  NOR U3629 ( .A(n[151]), .B(n3722), .Z(n3172) );
  NOR U3630 ( .A(n[147]), .B(n3738), .Z(n3169) );
  NOR U3631 ( .A(n[145]), .B(n3747), .Z(n3166) );
  NOR U3632 ( .A(n[144]), .B(n3751), .Z(n3163) );
  IV U3633 ( .A(n2876), .Z(n3760) );
  OR U3634 ( .A(n[142]), .B(n3760), .Z(n3162) );
  ANDN U3635 ( .B(n[142]), .A(n2876), .Z(n3160) );
  NOR U3636 ( .A(n[140]), .B(n3768), .Z(n3157) );
  NOR U3637 ( .A(n[133]), .B(n3797), .Z(n3154) );
  NOR U3638 ( .A(n[131]), .B(n3806), .Z(n3151) );
  NOR U3639 ( .A(n[130]), .B(n3810), .Z(n3148) );
  NOR U3640 ( .A(n[128]), .B(n3819), .Z(n3145) );
  NOR U3641 ( .A(n[125]), .B(n3831), .Z(n3142) );
  NOR U3642 ( .A(n[123]), .B(n3840), .Z(n3139) );
  NOR U3643 ( .A(n[122]), .B(n3845), .Z(n3136) );
  NOR U3644 ( .A(n[121]), .B(n3850), .Z(n3133) );
  NOR U3645 ( .A(n[120]), .B(n3855), .Z(n3130) );
  NOR U3646 ( .A(n[119]), .B(n3860), .Z(n3127) );
  NOR U3647 ( .A(n[118]), .B(n3864), .Z(n3124) );
  NOR U3648 ( .A(n[117]), .B(n3868), .Z(n3121) );
  NOR U3649 ( .A(n[116]), .B(n3873), .Z(n3118) );
  NOR U3650 ( .A(n[115]), .B(n3877), .Z(n3115) );
  NOR U3651 ( .A(n[114]), .B(n3882), .Z(n3112) );
  NOR U3652 ( .A(n[113]), .B(n3887), .Z(n3109) );
  NOR U3653 ( .A(n[112]), .B(n3892), .Z(n3106) );
  NOR U3654 ( .A(n[111]), .B(n3897), .Z(n3103) );
  NOR U3655 ( .A(n[110]), .B(n3902), .Z(n3100) );
  NOR U3656 ( .A(n[109]), .B(n3907), .Z(n3097) );
  NOR U3657 ( .A(n[108]), .B(n3911), .Z(n3094) );
  NOR U3658 ( .A(n[103]), .B(n3932), .Z(n3091) );
  NOR U3659 ( .A(n[101]), .B(n3941), .Z(n3088) );
  NOR U3660 ( .A(n[96]), .B(n3962), .Z(n3085) );
  NOR U3661 ( .A(n[95]), .B(n3967), .Z(n3082) );
  NOR U3662 ( .A(n[94]), .B(n3972), .Z(n3079) );
  NOR U3663 ( .A(n[93]), .B(n3977), .Z(n3076) );
  NOR U3664 ( .A(n[92]), .B(n4663), .Z(n3073) );
  NOR U3665 ( .A(n[91]), .B(n3981), .Z(n3070) );
  NOR U3666 ( .A(n[89]), .B(n3989), .Z(n3067) );
  NOR U3667 ( .A(n[87]), .B(n3997), .Z(n3064) );
  NOR U3668 ( .A(n[85]), .B(n4006), .Z(n3061) );
  NOR U3669 ( .A(n[81]), .B(n4022), .Z(n3058) );
  NOR U3670 ( .A(n[80]), .B(n4027), .Z(n3055) );
  NOR U3671 ( .A(n[77]), .B(n4040), .Z(n3052) );
  IV U3672 ( .A(n2877), .Z(n4053) );
  OR U3673 ( .A(n[74]), .B(n4053), .Z(n3051) );
  ANDN U3674 ( .B(n[74]), .A(n2877), .Z(n3049) );
  IV U3675 ( .A(n2878), .Z(n4061) );
  OR U3676 ( .A(n[72]), .B(n4061), .Z(n3048) );
  ANDN U3677 ( .B(n[72]), .A(n2878), .Z(n3046) );
  NOR U3678 ( .A(n[70]), .B(n4069), .Z(n3043) );
  NANDN U3679 ( .A(n4113), .B(n4112), .Z(n3027) );
  NOR U3680 ( .A(n[60]), .B(n4112), .Z(n3025) );
  NANDN U3681 ( .A(n4446), .B(n4192), .Z(n2973) );
  NOR U3682 ( .A(n[39]), .B(n4192), .Z(n2971) );
  NOR U3683 ( .A(n[31]), .B(n4419), .Z(n2959) );
  NOR U3684 ( .A(n[30]), .B(n4221), .Z(n2956) );
  NOR U3685 ( .A(n[29]), .B(n4226), .Z(n2953) );
  NOR U3686 ( .A(n[28]), .B(n4406), .Z(n2950) );
  NOR U3687 ( .A(n[24]), .B(n4238), .Z(n2947) );
  NOR U3688 ( .A(n[23]), .B(n4390), .Z(n2944) );
  NOR U3689 ( .A(n[22]), .B(n4243), .Z(n2941) );
  NOR U3690 ( .A(n[21]), .B(n4381), .Z(n2938) );
  NOR U3691 ( .A(n[20]), .B(n4247), .Z(n2935) );
  NOR U3692 ( .A(n[19]), .B(n4252), .Z(n2932) );
  NOR U3693 ( .A(n[18]), .B(n4256), .Z(n2929) );
  NANDN U3694 ( .A(n6868), .B(n4329), .Z(n2904) );
  ANDN U3695 ( .B(n[0]), .A(n2880), .Z(n4296) );
  NANDN U3696 ( .A(n6616), .B(n4300), .Z(n2883) );
  NOR U3697 ( .A(n[2]), .B(n4300), .Z(n2881) );
  NANDN U3698 ( .A(n2881), .B(n4303), .Z(n2882) );
  NAND U3699 ( .A(n2883), .B(n2882), .Z(n4304) );
  NAND U3700 ( .A(n4304), .B(n2884), .Z(n2885) );
  NAND U3701 ( .A(n2886), .B(n2885), .Z(n4292) );
  NAND U3702 ( .A(n4292), .B(n2887), .Z(n2888) );
  NAND U3703 ( .A(n2889), .B(n2888), .Z(n4288) );
  NAND U3704 ( .A(n4288), .B(n2890), .Z(n2891) );
  NAND U3705 ( .A(n2892), .B(n2891), .Z(n4284) );
  NAND U3706 ( .A(n4284), .B(n2893), .Z(n2894) );
  NAND U3707 ( .A(n2895), .B(n2894), .Z(n4280) );
  OR U3708 ( .A(n2896), .B(n4280), .Z(n2898) );
  AND U3709 ( .A(n2898), .B(n2897), .Z(n4276) );
  OR U3710 ( .A(n4276), .B(n2899), .Z(n2901) );
  NAND U3711 ( .A(n2901), .B(n2900), .Z(n4326) );
  NOR U3712 ( .A(n[9]), .B(n4329), .Z(n2902) );
  OR U3713 ( .A(n4326), .B(n2902), .Z(n2903) );
  NAND U3714 ( .A(n2904), .B(n2903), .Z(n4330) );
  NANDN U3715 ( .A(n2905), .B(n4330), .Z(n2906) );
  NANDN U3716 ( .A(n2907), .B(n2906), .Z(n4338) );
  NANDN U3717 ( .A(n2908), .B(n4338), .Z(n2909) );
  NANDN U3718 ( .A(n2910), .B(n2909), .Z(n4345) );
  NANDN U3719 ( .A(n2911), .B(n4345), .Z(n2912) );
  NANDN U3720 ( .A(n2913), .B(n2912), .Z(n4272) );
  NANDN U3721 ( .A(n2914), .B(n4272), .Z(n2915) );
  NANDN U3722 ( .A(n2916), .B(n2915), .Z(n4267) );
  NANDN U3723 ( .A(n2917), .B(n4267), .Z(n2918) );
  NANDN U3724 ( .A(n2919), .B(n2918), .Z(n4357) );
  NANDN U3725 ( .A(n2920), .B(n4357), .Z(n2921) );
  NANDN U3726 ( .A(n2922), .B(n2921), .Z(n4262) );
  NANDN U3727 ( .A(n2923), .B(n4262), .Z(n2924) );
  NANDN U3728 ( .A(n2925), .B(n2924), .Z(n4258) );
  NANDN U3729 ( .A(n2926), .B(n4258), .Z(n2927) );
  NANDN U3730 ( .A(n2928), .B(n2927), .Z(n4253) );
  NANDN U3731 ( .A(n2929), .B(n4253), .Z(n2930) );
  NAND U3732 ( .A(n2931), .B(n2930), .Z(n4249) );
  NANDN U3733 ( .A(n2932), .B(n4249), .Z(n2933) );
  NAND U3734 ( .A(n2934), .B(n2933), .Z(n4244) );
  NANDN U3735 ( .A(n2935), .B(n4244), .Z(n2936) );
  NAND U3736 ( .A(n2937), .B(n2936), .Z(n4378) );
  NANDN U3737 ( .A(n2938), .B(n4378), .Z(n2939) );
  NAND U3738 ( .A(n2940), .B(n2939), .Z(n4240) );
  NANDN U3739 ( .A(n2941), .B(n4240), .Z(n2942) );
  NAND U3740 ( .A(n2943), .B(n2942), .Z(n4386) );
  NANDN U3741 ( .A(n2944), .B(n4386), .Z(n2945) );
  NAND U3742 ( .A(n2946), .B(n2945), .Z(n4235) );
  NANDN U3743 ( .A(n2947), .B(n4235), .Z(n2948) );
  NAND U3744 ( .A(n2949), .B(n2948), .Z(n4231) );
  OR U3745 ( .A(n2950), .B(n4403), .Z(n2951) );
  NAND U3746 ( .A(n2952), .B(n2951), .Z(n4223) );
  NANDN U3747 ( .A(n2953), .B(n4223), .Z(n2954) );
  NAND U3748 ( .A(n2955), .B(n2954), .Z(n4218) );
  NANDN U3749 ( .A(n2956), .B(n4218), .Z(n2957) );
  NAND U3750 ( .A(n2958), .B(n2957), .Z(n4415) );
  NANDN U3751 ( .A(n2959), .B(n4415), .Z(n2960) );
  NAND U3752 ( .A(n2961), .B(n2960), .Z(n4214) );
  NANDN U3753 ( .A(n2962), .B(n4202), .Z(n2963) );
  NANDN U3754 ( .A(n2964), .B(n2963), .Z(n4198) );
  NANDN U3755 ( .A(n2965), .B(n4198), .Z(n2966) );
  NANDN U3756 ( .A(n2967), .B(n2966), .Z(n4193) );
  NANDN U3757 ( .A(n2968), .B(n4193), .Z(n2969) );
  NANDN U3758 ( .A(n2970), .B(n2969), .Z(n4189) );
  OR U3759 ( .A(n2971), .B(n4189), .Z(n2972) );
  NAND U3760 ( .A(n2973), .B(n2972), .Z(n4184) );
  OR U3761 ( .A(n2974), .B(n4184), .Z(n2975) );
  NANDN U3762 ( .A(n2976), .B(n2975), .Z(n4180) );
  NANDN U3763 ( .A(n4180), .B(n2977), .Z(n2978) );
  NANDN U3764 ( .A(n2979), .B(n2978), .Z(n4175) );
  NANDN U3765 ( .A(n2980), .B(n4175), .Z(n2981) );
  NANDN U3766 ( .A(n2982), .B(n2981), .Z(n4462) );
  NANDN U3767 ( .A(n2983), .B(n4462), .Z(n2984) );
  NANDN U3768 ( .A(n2985), .B(n2984), .Z(n4467) );
  OR U3769 ( .A(n2986), .B(n4467), .Z(n2987) );
  NANDN U3770 ( .A(n2988), .B(n2987), .Z(n4471) );
  NANDN U3771 ( .A(n2989), .B(n4171), .Z(n2990) );
  NANDN U3772 ( .A(n2991), .B(n2990), .Z(n4167) );
  NANDN U3773 ( .A(n2992), .B(n4167), .Z(n2993) );
  NAND U3774 ( .A(n2994), .B(n2993), .Z(n4163) );
  NANDN U3775 ( .A(n4163), .B(n2995), .Z(n2996) );
  NANDN U3776 ( .A(n2997), .B(n2996), .Z(n4158) );
  NANDN U3777 ( .A(n2998), .B(n4158), .Z(n2999) );
  NANDN U3778 ( .A(n3000), .B(n2999), .Z(n4154) );
  NANDN U3779 ( .A(n3001), .B(n4154), .Z(n3002) );
  NANDN U3780 ( .A(n3003), .B(n3002), .Z(n4150) );
  NANDN U3781 ( .A(n4146), .B(n3004), .Z(n3005) );
  NANDN U3782 ( .A(n3006), .B(n3005), .Z(n4141) );
  NANDN U3783 ( .A(n3007), .B(n4141), .Z(n3008) );
  NANDN U3784 ( .A(n3009), .B(n3008), .Z(n4136) );
  OR U3785 ( .A(n3010), .B(n4136), .Z(n3011) );
  NANDN U3786 ( .A(n3012), .B(n3011), .Z(n4132) );
  NANDN U3787 ( .A(n3013), .B(n4132), .Z(n3014) );
  NANDN U3788 ( .A(n3015), .B(n3014), .Z(n4127) );
  NANDN U3789 ( .A(n3016), .B(n4127), .Z(n3017) );
  NANDN U3790 ( .A(n3018), .B(n3017), .Z(n4123) );
  NANDN U3791 ( .A(n3019), .B(n4119), .Z(n3020) );
  NANDN U3792 ( .A(n3021), .B(n3020), .Z(n4114) );
  NANDN U3793 ( .A(n3022), .B(n4114), .Z(n3023) );
  NANDN U3794 ( .A(n3024), .B(n3023), .Z(n4109) );
  NANDN U3795 ( .A(n3025), .B(n4109), .Z(n3026) );
  NAND U3796 ( .A(n3027), .B(n3026), .Z(n4104) );
  OR U3797 ( .A(n3028), .B(n4104), .Z(n3029) );
  NANDN U3798 ( .A(n3030), .B(n3029), .Z(n4100) );
  NANDN U3799 ( .A(n4100), .B(n3031), .Z(n3032) );
  NANDN U3800 ( .A(n3033), .B(n3032), .Z(n4096) );
  NANDN U3801 ( .A(n3034), .B(n4092), .Z(n3035) );
  NANDN U3802 ( .A(n3036), .B(n3035), .Z(n4087) );
  NANDN U3803 ( .A(n3037), .B(n4087), .Z(n3039) );
  ANDN U3804 ( .B(n3039), .A(n3038), .Z(n4083) );
  NANDN U3805 ( .A(n3040), .B(n4074), .Z(n3041) );
  NANDN U3806 ( .A(n3042), .B(n3041), .Z(n4070) );
  OR U3807 ( .A(n3043), .B(n4066), .Z(n3044) );
  NAND U3808 ( .A(n3045), .B(n3044), .Z(n4062) );
  NANDN U3809 ( .A(n3046), .B(n4058), .Z(n3047) );
  NAND U3810 ( .A(n3048), .B(n3047), .Z(n4054) );
  NANDN U3811 ( .A(n3049), .B(n4050), .Z(n3050) );
  NAND U3812 ( .A(n3051), .B(n3050), .Z(n4046) );
  OR U3813 ( .A(n3052), .B(n4037), .Z(n3053) );
  NAND U3814 ( .A(n3054), .B(n3053), .Z(n4033) );
  OR U3815 ( .A(n3055), .B(n4024), .Z(n3056) );
  NAND U3816 ( .A(n3057), .B(n3056), .Z(n4019) );
  NANDN U3817 ( .A(n3058), .B(n4019), .Z(n3059) );
  NAND U3818 ( .A(n3060), .B(n3059), .Z(n4015) );
  OR U3819 ( .A(n3061), .B(n4003), .Z(n3062) );
  NAND U3820 ( .A(n3063), .B(n3062), .Z(n3999) );
  OR U3821 ( .A(n3064), .B(n3994), .Z(n3065) );
  NAND U3822 ( .A(n3066), .B(n3065), .Z(n3990) );
  OR U3823 ( .A(n3067), .B(n3986), .Z(n3068) );
  NAND U3824 ( .A(n3069), .B(n3068), .Z(n3982) );
  OR U3825 ( .A(n3070), .B(n3978), .Z(n3071) );
  NAND U3826 ( .A(n3072), .B(n3071), .Z(n4660) );
  NANDN U3827 ( .A(n3073), .B(n4660), .Z(n3074) );
  NAND U3828 ( .A(n3075), .B(n3074), .Z(n3973) );
  NANDN U3829 ( .A(n3076), .B(n3973), .Z(n3077) );
  NAND U3830 ( .A(n3078), .B(n3077), .Z(n3968) );
  NANDN U3831 ( .A(n3079), .B(n3968), .Z(n3080) );
  NAND U3832 ( .A(n3081), .B(n3080), .Z(n3964) );
  NANDN U3833 ( .A(n3082), .B(n3964), .Z(n3083) );
  NAND U3834 ( .A(n3084), .B(n3083), .Z(n3959) );
  NANDN U3835 ( .A(n3085), .B(n3959), .Z(n3086) );
  NAND U3836 ( .A(n3087), .B(n3086), .Z(n3955) );
  OR U3837 ( .A(n3088), .B(n3938), .Z(n3089) );
  NAND U3838 ( .A(n3090), .B(n3089), .Z(n3934) );
  OR U3839 ( .A(n3091), .B(n3929), .Z(n3092) );
  NAND U3840 ( .A(n3093), .B(n3092), .Z(n3925) );
  OR U3841 ( .A(n3094), .B(n3908), .Z(n3095) );
  NAND U3842 ( .A(n3096), .B(n3095), .Z(n3904) );
  NANDN U3843 ( .A(n3097), .B(n3904), .Z(n3098) );
  NAND U3844 ( .A(n3099), .B(n3098), .Z(n3899) );
  NANDN U3845 ( .A(n3100), .B(n3899), .Z(n3101) );
  NAND U3846 ( .A(n3102), .B(n3101), .Z(n3894) );
  NANDN U3847 ( .A(n3103), .B(n3894), .Z(n3104) );
  NAND U3848 ( .A(n3105), .B(n3104), .Z(n3889) );
  NANDN U3849 ( .A(n3106), .B(n3889), .Z(n3107) );
  NAND U3850 ( .A(n3108), .B(n3107), .Z(n3884) );
  NANDN U3851 ( .A(n3109), .B(n3884), .Z(n3110) );
  NAND U3852 ( .A(n3111), .B(n3110), .Z(n3879) );
  NANDN U3853 ( .A(n3112), .B(n3879), .Z(n3113) );
  NAND U3854 ( .A(n3114), .B(n3113), .Z(n3874) );
  NANDN U3855 ( .A(n3115), .B(n3874), .Z(n3116) );
  NAND U3856 ( .A(n3117), .B(n3116), .Z(n3870) );
  NANDN U3857 ( .A(n3118), .B(n3870), .Z(n3119) );
  NAND U3858 ( .A(n3120), .B(n3119), .Z(n3865) );
  NANDN U3859 ( .A(n3121), .B(n3865), .Z(n3122) );
  NAND U3860 ( .A(n3123), .B(n3122), .Z(n3861) );
  NANDN U3861 ( .A(n3124), .B(n3861), .Z(n3125) );
  NAND U3862 ( .A(n3126), .B(n3125), .Z(n3857) );
  NANDN U3863 ( .A(n3127), .B(n3857), .Z(n3128) );
  NAND U3864 ( .A(n3129), .B(n3128), .Z(n3852) );
  NANDN U3865 ( .A(n3130), .B(n3852), .Z(n3131) );
  NAND U3866 ( .A(n3132), .B(n3131), .Z(n3847) );
  NANDN U3867 ( .A(n3133), .B(n3847), .Z(n3134) );
  NAND U3868 ( .A(n3135), .B(n3134), .Z(n3842) );
  NANDN U3869 ( .A(n3136), .B(n3842), .Z(n3137) );
  NAND U3870 ( .A(n3138), .B(n3137), .Z(n3837) );
  NANDN U3871 ( .A(n3139), .B(n3837), .Z(n3140) );
  NAND U3872 ( .A(n3141), .B(n3140), .Z(n3833) );
  OR U3873 ( .A(n3142), .B(n3828), .Z(n3143) );
  NAND U3874 ( .A(n3144), .B(n3143), .Z(n3824) );
  OR U3875 ( .A(n3145), .B(n3816), .Z(n3146) );
  NAND U3876 ( .A(n3147), .B(n3146), .Z(n3812) );
  OR U3877 ( .A(n3148), .B(n3807), .Z(n3149) );
  NAND U3878 ( .A(n3150), .B(n3149), .Z(n3803) );
  NANDN U3879 ( .A(n3151), .B(n3803), .Z(n3152) );
  NAND U3880 ( .A(n3153), .B(n3152), .Z(n3799) );
  OR U3881 ( .A(n3154), .B(n3794), .Z(n3155) );
  NAND U3882 ( .A(n3156), .B(n3155), .Z(n3790) );
  OR U3883 ( .A(n3157), .B(n3765), .Z(n3158) );
  NAND U3884 ( .A(n3159), .B(n3158), .Z(n3761) );
  NANDN U3885 ( .A(n3160), .B(n3757), .Z(n3161) );
  NAND U3886 ( .A(n3162), .B(n3161), .Z(n3753) );
  OR U3887 ( .A(n3163), .B(n3748), .Z(n3164) );
  NAND U3888 ( .A(n3165), .B(n3164), .Z(n3744) );
  NANDN U3889 ( .A(n3166), .B(n3744), .Z(n3167) );
  NAND U3890 ( .A(n3168), .B(n3167), .Z(n3740) );
  OR U3891 ( .A(n3169), .B(n3735), .Z(n3170) );
  NAND U3892 ( .A(n3171), .B(n3170), .Z(n3731) );
  OR U3893 ( .A(n3172), .B(n3719), .Z(n3173) );
  NAND U3894 ( .A(n3174), .B(n3173), .Z(n3715) );
  OR U3895 ( .A(n3175), .B(n4909), .Z(n3176) );
  NAND U3896 ( .A(n3177), .B(n3176), .Z(n3711) );
  NANDN U3897 ( .A(n3178), .B(n3711), .Z(n3179) );
  NAND U3898 ( .A(n3180), .B(n3179), .Z(n4923) );
  OR U3899 ( .A(n3181), .B(n3707), .Z(n3182) );
  NAND U3900 ( .A(n3183), .B(n3182), .Z(n4934) );
  NANDN U3901 ( .A(n3184), .B(n4934), .Z(n3185) );
  NAND U3902 ( .A(n3186), .B(n3185), .Z(n3703) );
  NANDN U3903 ( .A(n3187), .B(n3703), .Z(n3188) );
  NAND U3904 ( .A(n3189), .B(n3188), .Z(n3699) );
  OR U3905 ( .A(n3190), .B(n3694), .Z(n3191) );
  NAND U3906 ( .A(n3192), .B(n3191), .Z(n3690) );
  OR U3907 ( .A(n3193), .B(n3678), .Z(n3194) );
  NAND U3908 ( .A(n3195), .B(n3194), .Z(n3674) );
  NANDN U3909 ( .A(n3196), .B(n3674), .Z(n3197) );
  NAND U3910 ( .A(n3198), .B(n3197), .Z(n3669) );
  NANDN U3911 ( .A(n3199), .B(n3669), .Z(n3200) );
  NAND U3912 ( .A(n3201), .B(n3200), .Z(n3665) );
  NANDN U3913 ( .A(n3202), .B(n3665), .Z(n3203) );
  NAND U3914 ( .A(n3204), .B(n3203), .Z(n3660) );
  NANDN U3915 ( .A(n3205), .B(n3660), .Z(n3206) );
  NAND U3916 ( .A(n3207), .B(n3206), .Z(n3656) );
  OR U3917 ( .A(n3208), .B(n3651), .Z(n3209) );
  NAND U3918 ( .A(n3210), .B(n3209), .Z(n3647) );
  NANDN U3919 ( .A(n3211), .B(n3647), .Z(n3212) );
  NAND U3920 ( .A(n3213), .B(n3212), .Z(n3642) );
  NANDN U3921 ( .A(n3214), .B(n3642), .Z(n3215) );
  NAND U3922 ( .A(n3216), .B(n3215), .Z(n3637) );
  NANDN U3923 ( .A(n3217), .B(n3637), .Z(n3218) );
  NAND U3924 ( .A(n3219), .B(n3218), .Z(n3633) );
  OR U3925 ( .A(n3220), .B(n3629), .Z(n3221) );
  NAND U3926 ( .A(n3222), .B(n3221), .Z(n3625) );
  OR U3927 ( .A(n3223), .B(n3620), .Z(n3224) );
  NAND U3928 ( .A(n3225), .B(n3224), .Z(n3616) );
  OR U3929 ( .A(n3226), .B(n3599), .Z(n3227) );
  NAND U3930 ( .A(n3228), .B(n3227), .Z(n3595) );
  NANDN U3931 ( .A(n3229), .B(n3595), .Z(n3230) );
  NAND U3932 ( .A(n3231), .B(n3230), .Z(n5051) );
  OR U3933 ( .A(n3232), .B(n3587), .Z(n3233) );
  NAND U3934 ( .A(n3234), .B(n3233), .Z(n3582) );
  NANDN U3935 ( .A(n3235), .B(n3582), .Z(n3236) );
  NAND U3936 ( .A(n3237), .B(n3236), .Z(n3577) );
  OR U3937 ( .A(n3238), .B(n3573), .Z(n3239) );
  NAND U3938 ( .A(n3240), .B(n3239), .Z(n3569) );
  NANDN U3939 ( .A(n3241), .B(n3569), .Z(n3242) );
  NAND U3940 ( .A(n3243), .B(n3242), .Z(n3565) );
  OR U3941 ( .A(n3244), .B(n3551), .Z(n3245) );
  NAND U3942 ( .A(n3246), .B(n3245), .Z(n3547) );
  OR U3943 ( .A(n3247), .B(n3530), .Z(n3248) );
  NAND U3944 ( .A(n3249), .B(n3248), .Z(n3525) );
  NANDN U3945 ( .A(n3250), .B(n3525), .Z(n3251) );
  NAND U3946 ( .A(n3252), .B(n3251), .Z(n3521) );
  OR U3947 ( .A(n3253), .B(n3517), .Z(n3254) );
  NAND U3948 ( .A(n3255), .B(n3254), .Z(n3513) );
  OR U3949 ( .A(n3256), .B(n3504), .Z(n3257) );
  NAND U3950 ( .A(n3258), .B(n3257), .Z(n3500) );
  OR U3951 ( .A(n3259), .B(n3495), .Z(n3260) );
  NAND U3952 ( .A(n3261), .B(n3260), .Z(n3489) );
  OR U3953 ( .A(n3262), .B(n3472), .Z(n3263) );
  NAND U3954 ( .A(n3264), .B(n3263), .Z(n3468) );
  OR U3955 ( .A(n3265), .B(n3456), .Z(n3266) );
  NAND U3956 ( .A(n3267), .B(n3266), .Z(n3452) );
  OR U3957 ( .A(n3268), .B(n3440), .Z(n3269) );
  NAND U3958 ( .A(n3270), .B(n3269), .Z(n3436) );
  OR U3959 ( .A(n3271), .B(n3428), .Z(n3272) );
  NAND U3960 ( .A(n3273), .B(n3272), .Z(n3424) );
  NANDN U3961 ( .A(n3274), .B(n3416), .Z(n3275) );
  NAND U3962 ( .A(n3276), .B(n3275), .Z(n3412) );
  OR U3963 ( .A(n3277), .B(n3408), .Z(n3278) );
  NAND U3964 ( .A(n3279), .B(n3278), .Z(n3404) );
  OR U3965 ( .A(n3280), .B(n3378), .Z(n3281) );
  NAND U3966 ( .A(n3282), .B(n3281), .Z(n3374) );
  OR U3967 ( .A(n3283), .B(n3357), .Z(n3284) );
  NAND U3968 ( .A(n3285), .B(n3284), .Z(n3353) );
  NANDN U3969 ( .A(n3286), .B(n3353), .Z(n3287) );
  NAND U3970 ( .A(n3288), .B(n3287), .Z(n3349) );
  NANDN U3971 ( .A(n3289), .B(n3349), .Z(n3290) );
  NAND U3972 ( .A(n3291), .B(n3290), .Z(n3344) );
  NANDN U3973 ( .A(n3292), .B(n3344), .Z(n3293) );
  NAND U3974 ( .A(n3294), .B(n3293), .Z(n3340) );
  OR U3975 ( .A(n3295), .B(n3336), .Z(n3296) );
  NAND U3976 ( .A(n3297), .B(n3296), .Z(n3332) );
  OR U3977 ( .A(n3298), .B(n3323), .Z(n3299) );
  NAND U3978 ( .A(n3300), .B(n3299), .Z(n3319) );
  OR U3979 ( .A(n3301), .B(n3315), .Z(n3302) );
  NAND U3980 ( .A(n3303), .B(n3302), .Z(n3305) );
  XOR U3981 ( .A(n[255]), .B(n3305), .Z(n3304) );
  AND U3982 ( .A(n3304), .B(n523), .Z(n3307) );
  XOR U3983 ( .A(n3308), .B(n3307), .Z(n6580) );
  OR U3984 ( .A(n6580), .B(n[255]), .Z(n3314) );
  NAND U3985 ( .A(n[255]), .B(n3305), .Z(n3306) );
  OR U3986 ( .A(n3306), .B(n524), .Z(n3310) );
  NAND U3987 ( .A(n3308), .B(n3307), .Z(n3309) );
  NAND U3988 ( .A(n3310), .B(n3309), .Z(n3311) );
  XNOR U3989 ( .A(n3312), .B(n3311), .Z(n6594) );
  NANDN U3990 ( .A(n3313), .B(n6594), .Z(n6577) );
  ANDN U3991 ( .B(n3314), .A(n6577), .Z(n5340) );
  XOR U3992 ( .A(n6582), .B(n3315), .Z(n3316) );
  NANDN U3993 ( .A(n524), .B(n3316), .Z(n3317) );
  XNOR U3994 ( .A(n3318), .B(n3317), .Z(n6583) );
  NANDN U3995 ( .A(n6582), .B(n6583), .Z(n5336) );
  XNOR U3996 ( .A(n6582), .B(n6583), .Z(n5334) );
  XOR U3997 ( .A(n[253]), .B(n3319), .Z(n3320) );
  NANDN U3998 ( .A(n524), .B(n3320), .Z(n3321) );
  XNOR U3999 ( .A(n3322), .B(n3321), .Z(n6571) );
  NAND U4000 ( .A(n[253]), .B(n6571), .Z(n5332) );
  XOR U4001 ( .A(n6571), .B(n[253]), .Z(n5330) );
  XOR U4002 ( .A(n3327), .B(n3323), .Z(n3324) );
  NANDN U4003 ( .A(n524), .B(n3324), .Z(n3325) );
  XNOR U4004 ( .A(n3326), .B(n3325), .Z(n6564) );
  NANDN U4005 ( .A(n3327), .B(n6564), .Z(n5328) );
  XNOR U4006 ( .A(n3327), .B(n6564), .Z(n5326) );
  XNOR U4007 ( .A(n[251]), .B(n3328), .Z(n3329) );
  NANDN U4008 ( .A(n524), .B(n3329), .Z(n3330) );
  XNOR U4009 ( .A(n3331), .B(n3330), .Z(n6558) );
  NAND U4010 ( .A(n[251]), .B(n6558), .Z(n5324) );
  XOR U4011 ( .A(n6558), .B(n[251]), .Z(n5322) );
  XOR U4012 ( .A(n[250]), .B(n3332), .Z(n3333) );
  NANDN U4013 ( .A(n524), .B(n3333), .Z(n3334) );
  XNOR U4014 ( .A(n3335), .B(n3334), .Z(n6552) );
  NAND U4015 ( .A(n[250]), .B(n6552), .Z(n5320) );
  XOR U4016 ( .A(n[250]), .B(n6552), .Z(n5318) );
  XOR U4017 ( .A(n6534), .B(n3336), .Z(n3337) );
  NANDN U4018 ( .A(n524), .B(n3337), .Z(n3338) );
  XNOR U4019 ( .A(n3339), .B(n3338), .Z(n6546) );
  NANDN U4020 ( .A(n6534), .B(n6546), .Z(n5316) );
  XNOR U4021 ( .A(n6546), .B(n6534), .Z(n5314) );
  XOR U4022 ( .A(n[248]), .B(n3340), .Z(n3341) );
  NANDN U4023 ( .A(n524), .B(n3341), .Z(n3342) );
  XNOR U4024 ( .A(n3343), .B(n3342), .Z(n6528) );
  NAND U4025 ( .A(n[248]), .B(n6528), .Z(n5312) );
  XOR U4026 ( .A(n[248]), .B(n6528), .Z(n5310) );
  XNOR U4027 ( .A(n3348), .B(n3344), .Z(n3345) );
  NANDN U4028 ( .A(n524), .B(n3345), .Z(n3346) );
  XNOR U4029 ( .A(n3347), .B(n3346), .Z(n6522) );
  NANDN U4030 ( .A(n3348), .B(n6522), .Z(n5308) );
  XNOR U4031 ( .A(n6522), .B(n3348), .Z(n5306) );
  XNOR U4032 ( .A(n6514), .B(n3349), .Z(n3350) );
  NANDN U4033 ( .A(n524), .B(n3350), .Z(n3351) );
  XNOR U4034 ( .A(n3352), .B(n3351), .Z(n6515) );
  NANDN U4035 ( .A(n6514), .B(n6515), .Z(n5304) );
  XNOR U4036 ( .A(n6514), .B(n6515), .Z(n5302) );
  XOR U4037 ( .A(n[245]), .B(n3353), .Z(n3354) );
  NANDN U4038 ( .A(n524), .B(n3354), .Z(n3355) );
  XNOR U4039 ( .A(n3356), .B(n3355), .Z(n6508) );
  NAND U4040 ( .A(n[245]), .B(n6508), .Z(n5300) );
  XOR U4041 ( .A(n6508), .B(n[245]), .Z(n5298) );
  XOR U4042 ( .A(n3361), .B(n3357), .Z(n3358) );
  NANDN U4043 ( .A(n524), .B(n3358), .Z(n3359) );
  XNOR U4044 ( .A(n3360), .B(n3359), .Z(n6503) );
  NANDN U4045 ( .A(n3361), .B(n6503), .Z(n5296) );
  XNOR U4046 ( .A(n3361), .B(n6503), .Z(n5294) );
  XNOR U4047 ( .A(n[243]), .B(n3362), .Z(n3363) );
  NANDN U4048 ( .A(n524), .B(n3363), .Z(n3364) );
  XNOR U4049 ( .A(n3365), .B(n3364), .Z(n6496) );
  NAND U4050 ( .A(n[243]), .B(n6496), .Z(n5292) );
  XOR U4051 ( .A(n6496), .B(n[243]), .Z(n5290) );
  XNOR U4052 ( .A(n[242]), .B(n3366), .Z(n3367) );
  NANDN U4053 ( .A(n524), .B(n3367), .Z(n3368) );
  XNOR U4054 ( .A(n3369), .B(n3368), .Z(n6490) );
  NAND U4055 ( .A(n[242]), .B(n6490), .Z(n5288) );
  XOR U4056 ( .A(n[242]), .B(n6490), .Z(n5286) );
  XNOR U4057 ( .A(n[241]), .B(n3370), .Z(n3371) );
  NANDN U4058 ( .A(n524), .B(n3371), .Z(n3372) );
  XNOR U4059 ( .A(n3373), .B(n3372), .Z(n6483) );
  NAND U4060 ( .A(n[241]), .B(n6483), .Z(n5284) );
  XOR U4061 ( .A(n6483), .B(n[241]), .Z(n5282) );
  XOR U4062 ( .A(n[240]), .B(n3374), .Z(n3375) );
  NANDN U4063 ( .A(n524), .B(n3375), .Z(n3376) );
  XNOR U4064 ( .A(n3377), .B(n3376), .Z(n6477) );
  NAND U4065 ( .A(n[240]), .B(n6477), .Z(n5280) );
  XOR U4066 ( .A(n[240]), .B(n6477), .Z(n5278) );
  XOR U4067 ( .A(n3382), .B(n3378), .Z(n3379) );
  NANDN U4068 ( .A(n524), .B(n3379), .Z(n3380) );
  XNOR U4069 ( .A(n3381), .B(n3380), .Z(n6474) );
  NANDN U4070 ( .A(n3382), .B(n6474), .Z(n5276) );
  XNOR U4071 ( .A(n6474), .B(n3382), .Z(n5274) );
  XNOR U4072 ( .A(n[238]), .B(n3383), .Z(n3384) );
  NANDN U4073 ( .A(n524), .B(n3384), .Z(n3385) );
  XNOR U4074 ( .A(n3386), .B(n3385), .Z(n6466) );
  NAND U4075 ( .A(n[238]), .B(n6466), .Z(n5272) );
  XOR U4076 ( .A(n[238]), .B(n6466), .Z(n5270) );
  XOR U4077 ( .A(n6449), .B(n3387), .Z(n3388) );
  NANDN U4078 ( .A(n524), .B(n3388), .Z(n3389) );
  XOR U4079 ( .A(n3390), .B(n3389), .Z(n5263) );
  IV U4080 ( .A(n5263), .Z(n6450) );
  XNOR U4081 ( .A(n[235]), .B(n3391), .Z(n3392) );
  NANDN U4082 ( .A(n524), .B(n3392), .Z(n3393) );
  XNOR U4083 ( .A(n3394), .B(n3393), .Z(n6443) );
  NAND U4084 ( .A(n[235]), .B(n6443), .Z(n5256) );
  XOR U4085 ( .A(n6443), .B(n[235]), .Z(n5254) );
  XOR U4086 ( .A(n3399), .B(n3395), .Z(n3396) );
  NANDN U4087 ( .A(n524), .B(n3396), .Z(n3397) );
  XOR U4088 ( .A(n3398), .B(n3397), .Z(n6439) );
  NANDN U4089 ( .A(n3399), .B(n6439), .Z(n5252) );
  XNOR U4090 ( .A(n3399), .B(n6439), .Z(n5250) );
  XNOR U4091 ( .A(n[233]), .B(n3400), .Z(n3401) );
  NANDN U4092 ( .A(n524), .B(n3401), .Z(n3402) );
  XNOR U4093 ( .A(n3403), .B(n3402), .Z(n6434) );
  NAND U4094 ( .A(n[233]), .B(n6434), .Z(n5248) );
  XOR U4095 ( .A(n6434), .B(n[233]), .Z(n5246) );
  XOR U4096 ( .A(n[232]), .B(n3404), .Z(n3405) );
  NANDN U4097 ( .A(n524), .B(n3405), .Z(n3406) );
  XNOR U4098 ( .A(n3407), .B(n3406), .Z(n6427) );
  NAND U4099 ( .A(n[232]), .B(n6427), .Z(n5244) );
  XOR U4100 ( .A(n[232]), .B(n6427), .Z(n5242) );
  XOR U4101 ( .A(n6413), .B(n3408), .Z(n3409) );
  NANDN U4102 ( .A(n524), .B(n3409), .Z(n3410) );
  XNOR U4103 ( .A(n3411), .B(n3410), .Z(n6415) );
  OR U4104 ( .A(n6415), .B(n[231]), .Z(n5239) );
  XNOR U4105 ( .A(n[229]), .B(n3412), .Z(n3413) );
  NANDN U4106 ( .A(n524), .B(n3413), .Z(n3414) );
  XNOR U4107 ( .A(n3415), .B(n3414), .Z(n6407) );
  NAND U4108 ( .A(n[229]), .B(n6407), .Z(n5229) );
  XOR U4109 ( .A(n6407), .B(n[229]), .Z(n5227) );
  XNOR U4110 ( .A(n[228]), .B(n3416), .Z(n3417) );
  NANDN U4111 ( .A(n524), .B(n3417), .Z(n3418) );
  XNOR U4112 ( .A(n3419), .B(n3418), .Z(n6397) );
  NAND U4113 ( .A(n[228]), .B(n6397), .Z(n5225) );
  XOR U4114 ( .A(n6397), .B(n[228]), .Z(n5223) );
  XNOR U4115 ( .A(n[227]), .B(n3420), .Z(n3421) );
  NANDN U4116 ( .A(n524), .B(n3421), .Z(n3422) );
  XNOR U4117 ( .A(n3423), .B(n3422), .Z(n6390) );
  NAND U4118 ( .A(n[227]), .B(n6390), .Z(n5221) );
  XOR U4119 ( .A(n[227]), .B(n6390), .Z(n5219) );
  XOR U4120 ( .A(n[226]), .B(n3424), .Z(n3425) );
  NANDN U4121 ( .A(n524), .B(n3425), .Z(n3426) );
  XNOR U4122 ( .A(n3427), .B(n3426), .Z(n6383) );
  NAND U4123 ( .A(n[226]), .B(n6383), .Z(n5217) );
  XOR U4124 ( .A(n6383), .B(n[226]), .Z(n5215) );
  XOR U4125 ( .A(n6376), .B(n3428), .Z(n3429) );
  NANDN U4126 ( .A(n524), .B(n3429), .Z(n3430) );
  XNOR U4127 ( .A(n3431), .B(n3430), .Z(n6377) );
  NANDN U4128 ( .A(n6376), .B(n6377), .Z(n5213) );
  XNOR U4129 ( .A(n6376), .B(n6377), .Z(n5211) );
  XNOR U4130 ( .A(n[224]), .B(n3432), .Z(n3433) );
  NANDN U4131 ( .A(n524), .B(n3433), .Z(n3434) );
  XNOR U4132 ( .A(n3435), .B(n3434), .Z(n6371) );
  NAND U4133 ( .A(n[224]), .B(n6371), .Z(n5209) );
  XOR U4134 ( .A(n6371), .B(n[224]), .Z(n5207) );
  XOR U4135 ( .A(n[223]), .B(n3436), .Z(n3437) );
  NANDN U4136 ( .A(n524), .B(n3437), .Z(n3438) );
  XNOR U4137 ( .A(n3439), .B(n3438), .Z(n6365) );
  NAND U4138 ( .A(n[223]), .B(n6365), .Z(n5205) );
  XOR U4139 ( .A(n[223]), .B(n6365), .Z(n5203) );
  XOR U4140 ( .A(n6357), .B(n3440), .Z(n3441) );
  NANDN U4141 ( .A(n524), .B(n3441), .Z(n3442) );
  XNOR U4142 ( .A(n3443), .B(n3442), .Z(n6358) );
  NANDN U4143 ( .A(n6357), .B(n6358), .Z(n5201) );
  XNOR U4144 ( .A(n6358), .B(n6357), .Z(n5199) );
  XNOR U4145 ( .A(n[221]), .B(n3444), .Z(n3445) );
  NANDN U4146 ( .A(n524), .B(n3445), .Z(n3446) );
  XNOR U4147 ( .A(n3447), .B(n3446), .Z(n6351) );
  NAND U4148 ( .A(n[221]), .B(n6351), .Z(n5197) );
  XOR U4149 ( .A(n6351), .B(n[221]), .Z(n5195) );
  XNOR U4150 ( .A(n[220]), .B(n3448), .Z(n3449) );
  NANDN U4151 ( .A(n524), .B(n3449), .Z(n3450) );
  XNOR U4152 ( .A(n3451), .B(n3450), .Z(n6342) );
  NAND U4153 ( .A(n[220]), .B(n6342), .Z(n5193) );
  XOR U4154 ( .A(n[220]), .B(n6342), .Z(n5191) );
  XOR U4155 ( .A(n[219]), .B(n3452), .Z(n3453) );
  NANDN U4156 ( .A(n524), .B(n3453), .Z(n3454) );
  XNOR U4157 ( .A(n3455), .B(n3454), .Z(n6335) );
  NAND U4158 ( .A(n[219]), .B(n6335), .Z(n5189) );
  XOR U4159 ( .A(n6335), .B(n[219]), .Z(n5187) );
  XOR U4160 ( .A(n6317), .B(n3456), .Z(n3457) );
  NANDN U4161 ( .A(n524), .B(n3457), .Z(n3458) );
  XNOR U4162 ( .A(n3459), .B(n3458), .Z(n6319) );
  NANDN U4163 ( .A(n6317), .B(n6319), .Z(n6326) );
  XNOR U4164 ( .A(n[216]), .B(n3460), .Z(n3461) );
  NANDN U4165 ( .A(n524), .B(n3461), .Z(n3462) );
  XNOR U4166 ( .A(n3463), .B(n3462), .Z(n6311) );
  NAND U4167 ( .A(n[216]), .B(n6311), .Z(n5174) );
  XOR U4168 ( .A(n6311), .B(n[216]), .Z(n5172) );
  XNOR U4169 ( .A(n[215]), .B(n3464), .Z(n3465) );
  NANDN U4170 ( .A(n524), .B(n3465), .Z(n3466) );
  XNOR U4171 ( .A(n3467), .B(n3466), .Z(n6305) );
  NAND U4172 ( .A(n[215]), .B(n6305), .Z(n5170) );
  XOR U4173 ( .A(n[215]), .B(n6305), .Z(n5168) );
  XOR U4174 ( .A(n[214]), .B(n3468), .Z(n3469) );
  NANDN U4175 ( .A(n524), .B(n3469), .Z(n3470) );
  XOR U4176 ( .A(n3471), .B(n3470), .Z(n6302) );
  NANDN U4177 ( .A(n6302), .B(n[214]), .Z(n5166) );
  XNOR U4178 ( .A(n6302), .B(n[214]), .Z(n5164) );
  XOR U4179 ( .A(n3476), .B(n3472), .Z(n3473) );
  NANDN U4180 ( .A(n524), .B(n3473), .Z(n3474) );
  XNOR U4181 ( .A(n3475), .B(n3474), .Z(n6295) );
  NANDN U4182 ( .A(n3476), .B(n6295), .Z(n5162) );
  XNOR U4183 ( .A(n3476), .B(n6295), .Z(n5160) );
  XNOR U4184 ( .A(n[212]), .B(n3477), .Z(n3478) );
  NANDN U4185 ( .A(n524), .B(n3478), .Z(n3479) );
  XNOR U4186 ( .A(n3480), .B(n3479), .Z(n6289) );
  NAND U4187 ( .A(n[212]), .B(n6289), .Z(n5158) );
  XOR U4188 ( .A(n6289), .B(n[212]), .Z(n5156) );
  XNOR U4189 ( .A(n[211]), .B(n3481), .Z(n3482) );
  NANDN U4190 ( .A(n524), .B(n3482), .Z(n3483) );
  XNOR U4191 ( .A(n3484), .B(n3483), .Z(n6283) );
  NAND U4192 ( .A(n[211]), .B(n6283), .Z(n5154) );
  XOR U4193 ( .A(n[211]), .B(n6283), .Z(n5152) );
  XOR U4194 ( .A(n6268), .B(n3485), .Z(n3486) );
  NANDN U4195 ( .A(n524), .B(n3486), .Z(n3487) );
  XOR U4196 ( .A(n3488), .B(n3487), .Z(n6270) );
  ANDN U4197 ( .B(n6270), .A(n6268), .Z(n6278) );
  XNOR U4198 ( .A(n6256), .B(n3489), .Z(n3490) );
  NANDN U4199 ( .A(n524), .B(n3490), .Z(n3491) );
  XOR U4200 ( .A(n3492), .B(n3491), .Z(n6271) );
  NANDN U4201 ( .A(n[209]), .B(n6271), .Z(n3494) );
  NOR U4202 ( .A(n[210]), .B(n6270), .Z(n3493) );
  ANDN U4203 ( .B(n3494), .A(n3493), .Z(n5149) );
  XOR U4204 ( .A(n3499), .B(n3495), .Z(n3496) );
  NANDN U4205 ( .A(n524), .B(n3496), .Z(n3497) );
  XNOR U4206 ( .A(n3498), .B(n3497), .Z(n6254) );
  NANDN U4207 ( .A(n3499), .B(n6254), .Z(n5145) );
  XNOR U4208 ( .A(n3499), .B(n6254), .Z(n5143) );
  XOR U4209 ( .A(n[207]), .B(n3500), .Z(n3501) );
  NANDN U4210 ( .A(n524), .B(n3501), .Z(n3502) );
  XNOR U4211 ( .A(n3503), .B(n3502), .Z(n6249) );
  NAND U4212 ( .A(n[207]), .B(n6249), .Z(n5141) );
  XOR U4213 ( .A(n6249), .B(n[207]), .Z(n5139) );
  XOR U4214 ( .A(n3508), .B(n3504), .Z(n3505) );
  NANDN U4215 ( .A(n524), .B(n3505), .Z(n3506) );
  XNOR U4216 ( .A(n3507), .B(n3506), .Z(n6242) );
  NANDN U4217 ( .A(n3508), .B(n6242), .Z(n5137) );
  XNOR U4218 ( .A(n3508), .B(n6242), .Z(n5135) );
  XNOR U4219 ( .A(n[205]), .B(n3509), .Z(n3510) );
  NANDN U4220 ( .A(n524), .B(n3510), .Z(n3511) );
  XNOR U4221 ( .A(n3512), .B(n3511), .Z(n6239) );
  NAND U4222 ( .A(n[205]), .B(n6239), .Z(n5133) );
  XOR U4223 ( .A(n6239), .B(n[205]), .Z(n5131) );
  XOR U4224 ( .A(n[204]), .B(n3513), .Z(n3514) );
  NANDN U4225 ( .A(n524), .B(n3514), .Z(n3515) );
  XNOR U4226 ( .A(n3516), .B(n3515), .Z(n6232) );
  NAND U4227 ( .A(n[204]), .B(n6232), .Z(n5129) );
  XOR U4228 ( .A(n[204]), .B(n6232), .Z(n5127) );
  XOR U4229 ( .A(n6225), .B(n3517), .Z(n3518) );
  NANDN U4230 ( .A(n524), .B(n3518), .Z(n3519) );
  XNOR U4231 ( .A(n3520), .B(n3519), .Z(n6226) );
  NANDN U4232 ( .A(n6225), .B(n6226), .Z(n5125) );
  XNOR U4233 ( .A(n6226), .B(n6225), .Z(n5123) );
  XOR U4234 ( .A(n[202]), .B(n3521), .Z(n3522) );
  NANDN U4235 ( .A(n524), .B(n3522), .Z(n3523) );
  XNOR U4236 ( .A(n3524), .B(n3523), .Z(n6219) );
  NAND U4237 ( .A(n[202]), .B(n6219), .Z(n5121) );
  XOR U4238 ( .A(n[202]), .B(n6219), .Z(n5119) );
  XNOR U4239 ( .A(n3529), .B(n3525), .Z(n3526) );
  NANDN U4240 ( .A(n524), .B(n3526), .Z(n3527) );
  XNOR U4241 ( .A(n3528), .B(n3527), .Z(n6213) );
  NANDN U4242 ( .A(n3529), .B(n6213), .Z(n5117) );
  XNOR U4243 ( .A(n6213), .B(n3529), .Z(n5115) );
  XOR U4244 ( .A(n6199), .B(n3530), .Z(n3531) );
  NANDN U4245 ( .A(n524), .B(n3531), .Z(n3532) );
  XNOR U4246 ( .A(n3533), .B(n3532), .Z(n6201) );
  NANDN U4247 ( .A(n6199), .B(n6201), .Z(n6208) );
  XNOR U4248 ( .A(n[199]), .B(n3534), .Z(n3535) );
  NANDN U4249 ( .A(n524), .B(n3535), .Z(n3536) );
  XNOR U4250 ( .A(n3537), .B(n3536), .Z(n6202) );
  NAND U4251 ( .A(n[199]), .B(n6202), .Z(n3538) );
  AND U4252 ( .A(n6208), .B(n3538), .Z(n5111) );
  XOR U4253 ( .A(n6202), .B(n[199]), .Z(n5109) );
  XNOR U4254 ( .A(n[198]), .B(n3539), .Z(n3540) );
  NANDN U4255 ( .A(n524), .B(n3540), .Z(n3541) );
  XNOR U4256 ( .A(n3542), .B(n3541), .Z(n6188) );
  NAND U4257 ( .A(n[198]), .B(n6188), .Z(n5107) );
  XOR U4258 ( .A(n[198]), .B(n6188), .Z(n5105) );
  XNOR U4259 ( .A(n[197]), .B(n3543), .Z(n3544) );
  NANDN U4260 ( .A(n524), .B(n3544), .Z(n3545) );
  XNOR U4261 ( .A(n3546), .B(n3545), .Z(n6181) );
  NAND U4262 ( .A(n[197]), .B(n6181), .Z(n5103) );
  XOR U4263 ( .A(n6181), .B(n[197]), .Z(n5101) );
  XNOR U4264 ( .A(n6166), .B(n3547), .Z(n3548) );
  NANDN U4265 ( .A(n524), .B(n3548), .Z(n3549) );
  XNOR U4266 ( .A(n3550), .B(n3549), .Z(n6168) );
  NANDN U4267 ( .A(n6166), .B(n6168), .Z(n6175) );
  XOR U4268 ( .A(n3556), .B(n3551), .Z(n3552) );
  NANDN U4269 ( .A(n524), .B(n3552), .Z(n3553) );
  XNOR U4270 ( .A(n3554), .B(n3553), .Z(n6169) );
  NANDN U4271 ( .A(n3556), .B(n6169), .Z(n3555) );
  AND U4272 ( .A(n6175), .B(n3555), .Z(n5097) );
  XNOR U4273 ( .A(n6169), .B(n3556), .Z(n5095) );
  XNOR U4274 ( .A(n[194]), .B(n3557), .Z(n3558) );
  NANDN U4275 ( .A(n524), .B(n3558), .Z(n3559) );
  XNOR U4276 ( .A(n3560), .B(n3559), .Z(n6160) );
  NAND U4277 ( .A(n[194]), .B(n6160), .Z(n5093) );
  XOR U4278 ( .A(n[194]), .B(n6160), .Z(n5091) );
  XNOR U4279 ( .A(n[193]), .B(n3561), .Z(n3562) );
  NANDN U4280 ( .A(n524), .B(n3562), .Z(n3563) );
  XNOR U4281 ( .A(n3564), .B(n3563), .Z(n6154) );
  NAND U4282 ( .A(n[193]), .B(n6154), .Z(n5089) );
  XOR U4283 ( .A(n6154), .B(n[193]), .Z(n5087) );
  XOR U4284 ( .A(n[192]), .B(n3565), .Z(n3566) );
  NANDN U4285 ( .A(n524), .B(n3566), .Z(n3567) );
  XNOR U4286 ( .A(n3568), .B(n3567), .Z(n6148) );
  NAND U4287 ( .A(n[192]), .B(n6148), .Z(n5085) );
  XOR U4288 ( .A(n[192]), .B(n6148), .Z(n5083) );
  XOR U4289 ( .A(n[191]), .B(n3569), .Z(n3570) );
  NANDN U4290 ( .A(n524), .B(n3570), .Z(n3571) );
  XNOR U4291 ( .A(n3572), .B(n3571), .Z(n6142) );
  NAND U4292 ( .A(n[191]), .B(n6142), .Z(n5081) );
  XOR U4293 ( .A(n6142), .B(n[191]), .Z(n5079) );
  XOR U4294 ( .A(n6135), .B(n3573), .Z(n3574) );
  NANDN U4295 ( .A(n524), .B(n3574), .Z(n3575) );
  XNOR U4296 ( .A(n3576), .B(n3575), .Z(n6136) );
  NANDN U4297 ( .A(n6135), .B(n6136), .Z(n5077) );
  XNOR U4298 ( .A(n6136), .B(n6135), .Z(n5075) );
  XNOR U4299 ( .A(n3581), .B(n3577), .Z(n3578) );
  NANDN U4300 ( .A(n524), .B(n3578), .Z(n3579) );
  XOR U4301 ( .A(n3580), .B(n3579), .Z(n6130) );
  NANDN U4302 ( .A(n3581), .B(n6130), .Z(n5073) );
  XNOR U4303 ( .A(n3581), .B(n6130), .Z(n5071) );
  XNOR U4304 ( .A(n3586), .B(n3582), .Z(n3583) );
  NANDN U4305 ( .A(n524), .B(n3583), .Z(n3584) );
  XNOR U4306 ( .A(n3585), .B(n3584), .Z(n6113) );
  NANDN U4307 ( .A(n3586), .B(n6113), .Z(n5069) );
  XNOR U4308 ( .A(n6113), .B(n3586), .Z(n5067) );
  XOR U4309 ( .A(n6106), .B(n3587), .Z(n3588) );
  NANDN U4310 ( .A(n524), .B(n3588), .Z(n3589) );
  XNOR U4311 ( .A(n3590), .B(n3589), .Z(n6107) );
  NANDN U4312 ( .A(n6106), .B(n6107), .Z(n5065) );
  XNOR U4313 ( .A(n6106), .B(n6107), .Z(n5063) );
  XNOR U4314 ( .A(n[186]), .B(n3591), .Z(n3592) );
  NANDN U4315 ( .A(n524), .B(n3592), .Z(n3593) );
  XNOR U4316 ( .A(n3594), .B(n3593), .Z(n6100) );
  NAND U4317 ( .A(n[186]), .B(n6100), .Z(n5061) );
  XOR U4318 ( .A(n6100), .B(n[186]), .Z(n5059) );
  XNOR U4319 ( .A(n6086), .B(n3595), .Z(n3596) );
  NANDN U4320 ( .A(n524), .B(n3596), .Z(n3597) );
  XNOR U4321 ( .A(n3598), .B(n3597), .Z(n6087) );
  NANDN U4322 ( .A(n6086), .B(n6087), .Z(n5049) );
  XNOR U4323 ( .A(n6086), .B(n6087), .Z(n5047) );
  XOR U4324 ( .A(n3603), .B(n3599), .Z(n3600) );
  NANDN U4325 ( .A(n524), .B(n3600), .Z(n3601) );
  XNOR U4326 ( .A(n3602), .B(n3601), .Z(n6080) );
  NANDN U4327 ( .A(n3603), .B(n6080), .Z(n5045) );
  XNOR U4328 ( .A(n6080), .B(n3603), .Z(n5043) );
  XNOR U4329 ( .A(n[182]), .B(n3604), .Z(n3605) );
  NANDN U4330 ( .A(n524), .B(n3605), .Z(n3606) );
  XNOR U4331 ( .A(n3607), .B(n3606), .Z(n6073) );
  NAND U4332 ( .A(n[182]), .B(n6073), .Z(n5041) );
  XOR U4333 ( .A(n6073), .B(n[182]), .Z(n5039) );
  XNOR U4334 ( .A(n[181]), .B(n3608), .Z(n3609) );
  NANDN U4335 ( .A(n524), .B(n3609), .Z(n3610) );
  XNOR U4336 ( .A(n3611), .B(n3610), .Z(n6067) );
  NAND U4337 ( .A(n[181]), .B(n6067), .Z(n5037) );
  XOR U4338 ( .A(n[181]), .B(n6067), .Z(n5035) );
  XNOR U4339 ( .A(n[180]), .B(n3612), .Z(n3613) );
  NANDN U4340 ( .A(n524), .B(n3613), .Z(n3614) );
  XNOR U4341 ( .A(n3615), .B(n3614), .Z(n6061) );
  NAND U4342 ( .A(n[180]), .B(n6061), .Z(n5033) );
  XOR U4343 ( .A(n6061), .B(n[180]), .Z(n5031) );
  XNOR U4344 ( .A(n6039), .B(n3616), .Z(n3617) );
  NANDN U4345 ( .A(n524), .B(n3617), .Z(n3618) );
  XOR U4346 ( .A(n3619), .B(n3618), .Z(n6041) );
  NANDN U4347 ( .A(n[178]), .B(n6041), .Z(n5021) );
  NANDN U4348 ( .A(n6041), .B(n[178]), .Z(n6049) );
  XOR U4349 ( .A(n6042), .B(n3620), .Z(n3621) );
  NANDN U4350 ( .A(n524), .B(n3621), .Z(n3622) );
  XNOR U4351 ( .A(n3623), .B(n3622), .Z(n6043) );
  NANDN U4352 ( .A(n6042), .B(n6043), .Z(n3624) );
  AND U4353 ( .A(n6049), .B(n3624), .Z(n5019) );
  XNOR U4354 ( .A(n6043), .B(n6042), .Z(n5017) );
  XNOR U4355 ( .A(n6025), .B(n3625), .Z(n3626) );
  NANDN U4356 ( .A(n524), .B(n3626), .Z(n3627) );
  XOR U4357 ( .A(n3628), .B(n3627), .Z(n6033) );
  NANDN U4358 ( .A(n6033), .B(n[176]), .Z(n5015) );
  XNOR U4359 ( .A(n[176]), .B(n6033), .Z(n5013) );
  XOR U4360 ( .A(n6024), .B(n3629), .Z(n3630) );
  NANDN U4361 ( .A(n524), .B(n3630), .Z(n3631) );
  XNOR U4362 ( .A(n3632), .B(n3631), .Z(n6026) );
  NANDN U4363 ( .A(n6024), .B(n6026), .Z(n5011) );
  XNOR U4364 ( .A(n6026), .B(n6024), .Z(n5009) );
  XOR U4365 ( .A(n[174]), .B(n3633), .Z(n3634) );
  NANDN U4366 ( .A(n524), .B(n3634), .Z(n3635) );
  XNOR U4367 ( .A(n3636), .B(n3635), .Z(n6018) );
  NAND U4368 ( .A(n[174]), .B(n6018), .Z(n5007) );
  XOR U4369 ( .A(n[174]), .B(n6018), .Z(n5005) );
  XNOR U4370 ( .A(n3641), .B(n3637), .Z(n3638) );
  NANDN U4371 ( .A(n524), .B(n3638), .Z(n3639) );
  XNOR U4372 ( .A(n3640), .B(n3639), .Z(n6012) );
  NANDN U4373 ( .A(n3641), .B(n6012), .Z(n5003) );
  XNOR U4374 ( .A(n6012), .B(n3641), .Z(n5001) );
  XNOR U4375 ( .A(n3646), .B(n3642), .Z(n3643) );
  NANDN U4376 ( .A(n524), .B(n3643), .Z(n3644) );
  XNOR U4377 ( .A(n3645), .B(n3644), .Z(n6005) );
  NANDN U4378 ( .A(n3646), .B(n6005), .Z(n4999) );
  XNOR U4379 ( .A(n6005), .B(n3646), .Z(n4997) );
  XNOR U4380 ( .A(n5998), .B(n3647), .Z(n3648) );
  NANDN U4381 ( .A(n524), .B(n3648), .Z(n3649) );
  XNOR U4382 ( .A(n3650), .B(n3649), .Z(n5999) );
  NANDN U4383 ( .A(n5998), .B(n5999), .Z(n4995) );
  XNOR U4384 ( .A(n5998), .B(n5999), .Z(n4993) );
  XOR U4385 ( .A(n3655), .B(n3651), .Z(n3652) );
  NANDN U4386 ( .A(n524), .B(n3652), .Z(n3653) );
  XOR U4387 ( .A(n3654), .B(n3653), .Z(n5993) );
  IV U4388 ( .A(n5993), .Z(n5994) );
  NANDN U4389 ( .A(n3655), .B(n5994), .Z(n4991) );
  XNOR U4390 ( .A(n5993), .B(n[170]), .Z(n4989) );
  XOR U4391 ( .A(n[169]), .B(n3656), .Z(n3657) );
  NANDN U4392 ( .A(n524), .B(n3657), .Z(n3658) );
  XNOR U4393 ( .A(n3659), .B(n3658), .Z(n5986) );
  NAND U4394 ( .A(n[169]), .B(n5986), .Z(n4987) );
  XOR U4395 ( .A(n5986), .B(n[169]), .Z(n4985) );
  XNOR U4396 ( .A(n3664), .B(n3660), .Z(n3661) );
  NANDN U4397 ( .A(n524), .B(n3661), .Z(n3662) );
  XNOR U4398 ( .A(n3663), .B(n3662), .Z(n5970) );
  NANDN U4399 ( .A(n3664), .B(n5970), .Z(n4983) );
  XNOR U4400 ( .A(n3664), .B(n5970), .Z(n4981) );
  XOR U4401 ( .A(n[167]), .B(n3665), .Z(n3666) );
  NANDN U4402 ( .A(n524), .B(n3666), .Z(n3667) );
  XNOR U4403 ( .A(n3668), .B(n3667), .Z(n5964) );
  NAND U4404 ( .A(n[167]), .B(n5964), .Z(n4979) );
  XOR U4405 ( .A(n5964), .B(n[167]), .Z(n4977) );
  XNOR U4406 ( .A(n3673), .B(n3669), .Z(n3670) );
  NANDN U4407 ( .A(n524), .B(n3670), .Z(n3671) );
  XNOR U4408 ( .A(n3672), .B(n3671), .Z(n5958) );
  NANDN U4409 ( .A(n3673), .B(n5958), .Z(n4975) );
  XNOR U4410 ( .A(n3673), .B(n5958), .Z(n4973) );
  XOR U4411 ( .A(n[165]), .B(n3674), .Z(n3675) );
  NANDN U4412 ( .A(n524), .B(n3675), .Z(n3676) );
  XNOR U4413 ( .A(n3677), .B(n3676), .Z(n5951) );
  NAND U4414 ( .A(n[165]), .B(n5951), .Z(n4971) );
  XOR U4415 ( .A(n5951), .B(n[165]), .Z(n4969) );
  XOR U4416 ( .A(n5943), .B(n3678), .Z(n3679) );
  NANDN U4417 ( .A(n524), .B(n3679), .Z(n3680) );
  XNOR U4418 ( .A(n3681), .B(n3680), .Z(n5945) );
  NANDN U4419 ( .A(n5943), .B(n5945), .Z(n4967) );
  XNOR U4420 ( .A(n5943), .B(n5945), .Z(n4965) );
  XNOR U4421 ( .A(n[163]), .B(n3682), .Z(n3683) );
  NANDN U4422 ( .A(n524), .B(n3683), .Z(n3684) );
  XNOR U4423 ( .A(n3685), .B(n3684), .Z(n5937) );
  NAND U4424 ( .A(n[163]), .B(n5937), .Z(n4963) );
  XOR U4425 ( .A(n5937), .B(n[163]), .Z(n4961) );
  XNOR U4426 ( .A(n[162]), .B(n3686), .Z(n3687) );
  NANDN U4427 ( .A(n524), .B(n3687), .Z(n3688) );
  XNOR U4428 ( .A(n3689), .B(n3688), .Z(n5931) );
  NAND U4429 ( .A(n[162]), .B(n5931), .Z(n4959) );
  XOR U4430 ( .A(n[162]), .B(n5931), .Z(n4957) );
  XOR U4431 ( .A(n[161]), .B(n3690), .Z(n3691) );
  NANDN U4432 ( .A(n524), .B(n3691), .Z(n3692) );
  XNOR U4433 ( .A(n3693), .B(n3692), .Z(n5928) );
  NAND U4434 ( .A(n[161]), .B(n5928), .Z(n4955) );
  XOR U4435 ( .A(n5928), .B(n[161]), .Z(n4953) );
  XOR U4436 ( .A(n3698), .B(n3694), .Z(n3695) );
  NANDN U4437 ( .A(n524), .B(n3695), .Z(n3696) );
  XNOR U4438 ( .A(n3697), .B(n3696), .Z(n5924) );
  NANDN U4439 ( .A(n3698), .B(n5924), .Z(n4951) );
  XNOR U4440 ( .A(n3698), .B(n5924), .Z(n4949) );
  XOR U4441 ( .A(n[159]), .B(n3699), .Z(n3700) );
  NANDN U4442 ( .A(n524), .B(n3700), .Z(n3701) );
  XNOR U4443 ( .A(n3702), .B(n3701), .Z(n5919) );
  NAND U4444 ( .A(n[159]), .B(n5919), .Z(n4947) );
  XOR U4445 ( .A(n5919), .B(n[159]), .Z(n4945) );
  XNOR U4446 ( .A(n5903), .B(n3703), .Z(n3704) );
  NANDN U4447 ( .A(n524), .B(n3704), .Z(n3705) );
  XNOR U4448 ( .A(n3706), .B(n3705), .Z(n5905) );
  ANDN U4449 ( .B(n5905), .A(n5903), .Z(n5912) );
  XOR U4450 ( .A(n5889), .B(n3707), .Z(n3708) );
  NANDN U4451 ( .A(n524), .B(n3708), .Z(n3709) );
  XOR U4452 ( .A(n3710), .B(n3709), .Z(n5891) );
  NANDN U4453 ( .A(n[156]), .B(n5891), .Z(n4931) );
  NANDN U4454 ( .A(n5891), .B(n[156]), .Z(n5898) );
  XOR U4455 ( .A(n[154]), .B(n3711), .Z(n3712) );
  NANDN U4456 ( .A(n524), .B(n3712), .Z(n3713) );
  XNOR U4457 ( .A(n3714), .B(n3713), .Z(n5883) );
  NAND U4458 ( .A(n[154]), .B(n5883), .Z(n4920) );
  XOR U4459 ( .A(n5883), .B(n[154]), .Z(n4918) );
  XOR U4460 ( .A(n[152]), .B(n3715), .Z(n3716) );
  NANDN U4461 ( .A(n524), .B(n3716), .Z(n3717) );
  XNOR U4462 ( .A(n3718), .B(n3717), .Z(n5872) );
  NAND U4463 ( .A(n[152]), .B(n5872), .Z(n4907) );
  XOR U4464 ( .A(n[152]), .B(n5872), .Z(n4905) );
  XNOR U4465 ( .A(n[151]), .B(n3719), .Z(n3720) );
  NANDN U4466 ( .A(n524), .B(n3720), .Z(n3721) );
  XNOR U4467 ( .A(n3722), .B(n3721), .Z(n5866) );
  NAND U4468 ( .A(n[151]), .B(n5866), .Z(n4903) );
  XOR U4469 ( .A(n5866), .B(n[151]), .Z(n4901) );
  XNOR U4470 ( .A(n[150]), .B(n3723), .Z(n3724) );
  NANDN U4471 ( .A(n524), .B(n3724), .Z(n3725) );
  XNOR U4472 ( .A(n3726), .B(n3725), .Z(n5861) );
  NAND U4473 ( .A(n[150]), .B(n5861), .Z(n4899) );
  XOR U4474 ( .A(n5861), .B(n[150]), .Z(n4897) );
  XNOR U4475 ( .A(n[149]), .B(n3727), .Z(n3728) );
  NANDN U4476 ( .A(n524), .B(n3728), .Z(n3729) );
  XNOR U4477 ( .A(n3730), .B(n3729), .Z(n5854) );
  NAND U4478 ( .A(n[149]), .B(n5854), .Z(n4895) );
  XOR U4479 ( .A(n[149]), .B(n5854), .Z(n4893) );
  XOR U4480 ( .A(n[148]), .B(n3731), .Z(n3732) );
  NANDN U4481 ( .A(n524), .B(n3732), .Z(n3733) );
  XNOR U4482 ( .A(n3734), .B(n3733), .Z(n5838) );
  NAND U4483 ( .A(n[148]), .B(n5838), .Z(n4891) );
  XOR U4484 ( .A(n5838), .B(n[148]), .Z(n4889) );
  XOR U4485 ( .A(n3739), .B(n3735), .Z(n3736) );
  NANDN U4486 ( .A(n524), .B(n3736), .Z(n3737) );
  XNOR U4487 ( .A(n3738), .B(n3737), .Z(n5832) );
  NANDN U4488 ( .A(n3739), .B(n5832), .Z(n4887) );
  XNOR U4489 ( .A(n5832), .B(n3739), .Z(n4885) );
  XOR U4490 ( .A(n[146]), .B(n3740), .Z(n3741) );
  NANDN U4491 ( .A(n524), .B(n3741), .Z(n3742) );
  XNOR U4492 ( .A(n3743), .B(n3742), .Z(n5826) );
  NAND U4493 ( .A(n[146]), .B(n5826), .Z(n4883) );
  XOR U4494 ( .A(n[146]), .B(n5826), .Z(n4881) );
  XOR U4495 ( .A(n[145]), .B(n3744), .Z(n3745) );
  NANDN U4496 ( .A(n524), .B(n3745), .Z(n3746) );
  XNOR U4497 ( .A(n3747), .B(n3746), .Z(n5820) );
  NAND U4498 ( .A(n[145]), .B(n5820), .Z(n4879) );
  XOR U4499 ( .A(n5820), .B(n[145]), .Z(n4877) );
  XOR U4500 ( .A(n3752), .B(n3748), .Z(n3749) );
  NANDN U4501 ( .A(n524), .B(n3749), .Z(n3750) );
  XNOR U4502 ( .A(n3751), .B(n3750), .Z(n5813) );
  NANDN U4503 ( .A(n3752), .B(n5813), .Z(n4875) );
  XNOR U4504 ( .A(n5813), .B(n3752), .Z(n4873) );
  XNOR U4505 ( .A(n[143]), .B(n3753), .Z(n3754) );
  NANDN U4506 ( .A(n524), .B(n3754), .Z(n3755) );
  XNOR U4507 ( .A(n3756), .B(n3755), .Z(n5806) );
  NAND U4508 ( .A(n[143]), .B(n5806), .Z(n4871) );
  XOR U4509 ( .A(n[143]), .B(n5806), .Z(n4869) );
  XNOR U4510 ( .A(n[142]), .B(n3757), .Z(n3758) );
  NANDN U4511 ( .A(n524), .B(n3758), .Z(n3759) );
  XNOR U4512 ( .A(n3760), .B(n3759), .Z(n5800) );
  NAND U4513 ( .A(n[142]), .B(n5800), .Z(n4867) );
  XOR U4514 ( .A(n5800), .B(n[142]), .Z(n4865) );
  XOR U4515 ( .A(n[141]), .B(n3761), .Z(n3762) );
  NANDN U4516 ( .A(n524), .B(n3762), .Z(n3763) );
  XOR U4517 ( .A(n3764), .B(n3763), .Z(n5796) );
  NANDN U4518 ( .A(n5796), .B(n[141]), .Z(n4863) );
  XNOR U4519 ( .A(n[141]), .B(n5796), .Z(n4861) );
  XOR U4520 ( .A(n3769), .B(n3765), .Z(n3766) );
  NANDN U4521 ( .A(n524), .B(n3766), .Z(n3767) );
  XNOR U4522 ( .A(n3768), .B(n3767), .Z(n5789) );
  NANDN U4523 ( .A(n3769), .B(n5789), .Z(n4859) );
  XNOR U4524 ( .A(n5789), .B(n3769), .Z(n4857) );
  XNOR U4525 ( .A(n[139]), .B(n3770), .Z(n3771) );
  NANDN U4526 ( .A(n524), .B(n3771), .Z(n3772) );
  XNOR U4527 ( .A(n3773), .B(n3772), .Z(n5783) );
  NAND U4528 ( .A(n[139]), .B(n5783), .Z(n4855) );
  XOR U4529 ( .A(n5783), .B(n[139]), .Z(n4853) );
  XNOR U4530 ( .A(n[138]), .B(n3774), .Z(n3775) );
  NANDN U4531 ( .A(n524), .B(n3775), .Z(n3776) );
  XNOR U4532 ( .A(n3777), .B(n3776), .Z(n5776) );
  NAND U4533 ( .A(n[138]), .B(n5776), .Z(n4851) );
  XOR U4534 ( .A(n[138]), .B(n5776), .Z(n4849) );
  XNOR U4535 ( .A(n[137]), .B(n3778), .Z(n3779) );
  NANDN U4536 ( .A(n524), .B(n3779), .Z(n3780) );
  XNOR U4537 ( .A(n3781), .B(n3780), .Z(n5770) );
  NAND U4538 ( .A(n[137]), .B(n5770), .Z(n4847) );
  XOR U4539 ( .A(n5770), .B(n[137]), .Z(n4845) );
  XNOR U4540 ( .A(n[136]), .B(n3782), .Z(n3783) );
  NANDN U4541 ( .A(n524), .B(n3783), .Z(n3784) );
  XNOR U4542 ( .A(n3785), .B(n3784), .Z(n5764) );
  NAND U4543 ( .A(n[136]), .B(n5764), .Z(n4843) );
  XOR U4544 ( .A(n[136]), .B(n5764), .Z(n4841) );
  XNOR U4545 ( .A(n[135]), .B(n3786), .Z(n3787) );
  NANDN U4546 ( .A(n524), .B(n3787), .Z(n3788) );
  XNOR U4547 ( .A(n3789), .B(n3788), .Z(n5758) );
  NAND U4548 ( .A(n[135]), .B(n5758), .Z(n4839) );
  XOR U4549 ( .A(n5758), .B(n[135]), .Z(n4837) );
  XOR U4550 ( .A(n[134]), .B(n3790), .Z(n3791) );
  NANDN U4551 ( .A(n524), .B(n3791), .Z(n3792) );
  XNOR U4552 ( .A(n3793), .B(n3792), .Z(n5752) );
  NAND U4553 ( .A(n[134]), .B(n5752), .Z(n4835) );
  XOR U4554 ( .A(n[134]), .B(n5752), .Z(n4833) );
  XOR U4555 ( .A(n3798), .B(n3794), .Z(n3795) );
  NANDN U4556 ( .A(n524), .B(n3795), .Z(n3796) );
  XNOR U4557 ( .A(n3797), .B(n3796), .Z(n5746) );
  NANDN U4558 ( .A(n3798), .B(n5746), .Z(n4831) );
  XNOR U4559 ( .A(n5746), .B(n3798), .Z(n4829) );
  XOR U4560 ( .A(n[132]), .B(n3799), .Z(n3800) );
  NANDN U4561 ( .A(n524), .B(n3800), .Z(n3801) );
  XNOR U4562 ( .A(n3802), .B(n3801), .Z(n5739) );
  NAND U4563 ( .A(n[132]), .B(n5739), .Z(n4827) );
  XOR U4564 ( .A(n[132]), .B(n5739), .Z(n4825) );
  XOR U4565 ( .A(n[131]), .B(n3803), .Z(n3804) );
  NANDN U4566 ( .A(n524), .B(n3804), .Z(n3805) );
  XNOR U4567 ( .A(n3806), .B(n3805), .Z(n5733) );
  NAND U4568 ( .A(n[131]), .B(n5733), .Z(n4823) );
  XOR U4569 ( .A(n5733), .B(n[131]), .Z(n4821) );
  XOR U4570 ( .A(n3811), .B(n3807), .Z(n3808) );
  NANDN U4571 ( .A(n524), .B(n3808), .Z(n3809) );
  XNOR U4572 ( .A(n3810), .B(n3809), .Z(n5727) );
  NANDN U4573 ( .A(n3811), .B(n5727), .Z(n4819) );
  XNOR U4574 ( .A(n3811), .B(n5727), .Z(n4817) );
  XOR U4575 ( .A(n[129]), .B(n3812), .Z(n3813) );
  NANDN U4576 ( .A(n524), .B(n3813), .Z(n3814) );
  XNOR U4577 ( .A(n3815), .B(n3814), .Z(n5720) );
  NAND U4578 ( .A(n[129]), .B(n5720), .Z(n4815) );
  XOR U4579 ( .A(n5720), .B(n[129]), .Z(n4813) );
  XNOR U4580 ( .A(n[128]), .B(n3816), .Z(n3817) );
  NANDN U4581 ( .A(n524), .B(n3817), .Z(n3818) );
  XNOR U4582 ( .A(n3819), .B(n3818), .Z(n5710) );
  NAND U4583 ( .A(n[128]), .B(n5710), .Z(n4811) );
  XOR U4584 ( .A(n5710), .B(n[128]), .Z(n4809) );
  XNOR U4585 ( .A(n[127]), .B(n3820), .Z(n3821) );
  NANDN U4586 ( .A(n524), .B(n3821), .Z(n3822) );
  XNOR U4587 ( .A(n3823), .B(n3822), .Z(n5704) );
  NAND U4588 ( .A(n[127]), .B(n5704), .Z(n4807) );
  XOR U4589 ( .A(n[127]), .B(n5704), .Z(n4805) );
  XOR U4590 ( .A(n[126]), .B(n3824), .Z(n3825) );
  NANDN U4591 ( .A(n524), .B(n3825), .Z(n3826) );
  XNOR U4592 ( .A(n3827), .B(n3826), .Z(n5697) );
  NAND U4593 ( .A(n[126]), .B(n5697), .Z(n4803) );
  XOR U4594 ( .A(n5697), .B(n[126]), .Z(n4801) );
  XOR U4595 ( .A(n3832), .B(n3828), .Z(n3829) );
  NANDN U4596 ( .A(n524), .B(n3829), .Z(n3830) );
  XNOR U4597 ( .A(n3831), .B(n3830), .Z(n5694) );
  NANDN U4598 ( .A(n3832), .B(n5694), .Z(n4799) );
  XNOR U4599 ( .A(n3832), .B(n5694), .Z(n4797) );
  XOR U4600 ( .A(n[124]), .B(n3833), .Z(n3834) );
  NANDN U4601 ( .A(n524), .B(n3834), .Z(n3835) );
  XNOR U4602 ( .A(n3836), .B(n3835), .Z(n5687) );
  NAND U4603 ( .A(n[124]), .B(n5687), .Z(n4795) );
  XOR U4604 ( .A(n5687), .B(n[124]), .Z(n4793) );
  XNOR U4605 ( .A(n3841), .B(n3837), .Z(n3838) );
  NANDN U4606 ( .A(n524), .B(n3838), .Z(n3839) );
  XNOR U4607 ( .A(n3840), .B(n3839), .Z(n5681) );
  NANDN U4608 ( .A(n3841), .B(n5681), .Z(n4791) );
  XNOR U4609 ( .A(n3841), .B(n5681), .Z(n4789) );
  XNOR U4610 ( .A(n3846), .B(n3842), .Z(n3843) );
  NANDN U4611 ( .A(n524), .B(n3843), .Z(n3844) );
  XNOR U4612 ( .A(n3845), .B(n3844), .Z(n5675) );
  NANDN U4613 ( .A(n3846), .B(n5675), .Z(n4787) );
  XNOR U4614 ( .A(n5675), .B(n3846), .Z(n4785) );
  XNOR U4615 ( .A(n3851), .B(n3847), .Z(n3848) );
  NANDN U4616 ( .A(n524), .B(n3848), .Z(n3849) );
  XNOR U4617 ( .A(n3850), .B(n3849), .Z(n5669) );
  NANDN U4618 ( .A(n3851), .B(n5669), .Z(n4783) );
  XNOR U4619 ( .A(n3851), .B(n5669), .Z(n4781) );
  XNOR U4620 ( .A(n3856), .B(n3852), .Z(n3853) );
  NANDN U4621 ( .A(n524), .B(n3853), .Z(n3854) );
  XNOR U4622 ( .A(n3855), .B(n3854), .Z(n5666) );
  NANDN U4623 ( .A(n3856), .B(n5666), .Z(n4779) );
  XNOR U4624 ( .A(n5666), .B(n3856), .Z(n4777) );
  XOR U4625 ( .A(n[119]), .B(n3857), .Z(n3858) );
  NANDN U4626 ( .A(n524), .B(n3858), .Z(n3859) );
  XNOR U4627 ( .A(n3860), .B(n3859), .Z(n5659) );
  NAND U4628 ( .A(n[119]), .B(n5659), .Z(n4775) );
  XOR U4629 ( .A(n5659), .B(n[119]), .Z(n4773) );
  XNOR U4630 ( .A(n5648), .B(n3861), .Z(n3862) );
  NANDN U4631 ( .A(n524), .B(n3862), .Z(n3863) );
  XNOR U4632 ( .A(n3864), .B(n3863), .Z(n5649) );
  NANDN U4633 ( .A(n5648), .B(n5649), .Z(n4771) );
  XNOR U4634 ( .A(n5648), .B(n5649), .Z(n4769) );
  XNOR U4635 ( .A(n3869), .B(n3865), .Z(n3866) );
  NANDN U4636 ( .A(n524), .B(n3866), .Z(n3867) );
  XNOR U4637 ( .A(n3868), .B(n3867), .Z(n5641) );
  NANDN U4638 ( .A(n3869), .B(n5641), .Z(n4767) );
  XNOR U4639 ( .A(n5641), .B(n3869), .Z(n4765) );
  XNOR U4640 ( .A(n5633), .B(n3870), .Z(n3871) );
  NANDN U4641 ( .A(n524), .B(n3871), .Z(n3872) );
  XNOR U4642 ( .A(n3873), .B(n3872), .Z(n5634) );
  NANDN U4643 ( .A(n5633), .B(n5634), .Z(n4763) );
  XNOR U4644 ( .A(n5633), .B(n5634), .Z(n4761) );
  XNOR U4645 ( .A(n3878), .B(n3874), .Z(n3875) );
  NANDN U4646 ( .A(n524), .B(n3875), .Z(n3876) );
  XNOR U4647 ( .A(n3877), .B(n3876), .Z(n5627) );
  NANDN U4648 ( .A(n3878), .B(n5627), .Z(n4759) );
  XNOR U4649 ( .A(n5627), .B(n3878), .Z(n4757) );
  XNOR U4650 ( .A(n3883), .B(n3879), .Z(n3880) );
  NANDN U4651 ( .A(n524), .B(n3880), .Z(n3881) );
  XNOR U4652 ( .A(n3882), .B(n3881), .Z(n5625) );
  NANDN U4653 ( .A(n3883), .B(n5625), .Z(n4755) );
  XNOR U4654 ( .A(n3883), .B(n5625), .Z(n4753) );
  XNOR U4655 ( .A(n3888), .B(n3884), .Z(n3885) );
  NANDN U4656 ( .A(n524), .B(n3885), .Z(n3886) );
  XNOR U4657 ( .A(n3887), .B(n3886), .Z(n5621) );
  NANDN U4658 ( .A(n3888), .B(n5621), .Z(n4751) );
  XNOR U4659 ( .A(n5621), .B(n3888), .Z(n4749) );
  XNOR U4660 ( .A(n3893), .B(n3889), .Z(n3890) );
  NANDN U4661 ( .A(n524), .B(n3890), .Z(n3891) );
  XNOR U4662 ( .A(n3892), .B(n3891), .Z(n5616) );
  NANDN U4663 ( .A(n3893), .B(n5616), .Z(n4747) );
  XNOR U4664 ( .A(n5616), .B(n3893), .Z(n4745) );
  XNOR U4665 ( .A(n3898), .B(n3894), .Z(n3895) );
  NANDN U4666 ( .A(n524), .B(n3895), .Z(n3896) );
  XNOR U4667 ( .A(n3897), .B(n3896), .Z(n5612) );
  NANDN U4668 ( .A(n3898), .B(n5612), .Z(n4743) );
  XNOR U4669 ( .A(n5612), .B(n3898), .Z(n4741) );
  XNOR U4670 ( .A(n3903), .B(n3899), .Z(n3900) );
  NANDN U4671 ( .A(n524), .B(n3900), .Z(n3901) );
  XNOR U4672 ( .A(n3902), .B(n3901), .Z(n5605) );
  NANDN U4673 ( .A(n3903), .B(n5605), .Z(n4739) );
  XNOR U4674 ( .A(n3903), .B(n5605), .Z(n4737) );
  XOR U4675 ( .A(n[109]), .B(n3904), .Z(n3905) );
  NANDN U4676 ( .A(n524), .B(n3905), .Z(n3906) );
  XNOR U4677 ( .A(n3907), .B(n3906), .Z(n5599) );
  NAND U4678 ( .A(n[109]), .B(n5599), .Z(n4735) );
  XOR U4679 ( .A(n5599), .B(n[109]), .Z(n4733) );
  XOR U4680 ( .A(n3912), .B(n3908), .Z(n3909) );
  NANDN U4681 ( .A(n524), .B(n3909), .Z(n3910) );
  XNOR U4682 ( .A(n3911), .B(n3910), .Z(n5589) );
  NANDN U4683 ( .A(n3912), .B(n5589), .Z(n4731) );
  XNOR U4684 ( .A(n3912), .B(n5589), .Z(n4729) );
  XNOR U4685 ( .A(n[107]), .B(n3913), .Z(n3914) );
  NANDN U4686 ( .A(n524), .B(n3914), .Z(n3915) );
  XNOR U4687 ( .A(n3916), .B(n3915), .Z(n5582) );
  NAND U4688 ( .A(n[107]), .B(n5582), .Z(n4727) );
  XOR U4689 ( .A(n5582), .B(n[107]), .Z(n4725) );
  XNOR U4690 ( .A(n[106]), .B(n3917), .Z(n3918) );
  NANDN U4691 ( .A(n524), .B(n3918), .Z(n3919) );
  XNOR U4692 ( .A(n3920), .B(n3919), .Z(n5577) );
  NAND U4693 ( .A(n[106]), .B(n5577), .Z(n4723) );
  XOR U4694 ( .A(n5577), .B(n[106]), .Z(n4721) );
  XNOR U4695 ( .A(n[105]), .B(n3921), .Z(n3922) );
  NANDN U4696 ( .A(n524), .B(n3922), .Z(n3923) );
  XNOR U4697 ( .A(n3924), .B(n3923), .Z(n5570) );
  NAND U4698 ( .A(n[105]), .B(n5570), .Z(n4719) );
  XOR U4699 ( .A(n[105]), .B(n5570), .Z(n4717) );
  XOR U4700 ( .A(n[104]), .B(n3925), .Z(n3926) );
  NANDN U4701 ( .A(n524), .B(n3926), .Z(n3927) );
  XNOR U4702 ( .A(n3928), .B(n3927), .Z(n5567) );
  NAND U4703 ( .A(n[104]), .B(n5567), .Z(n4715) );
  XOR U4704 ( .A(n5567), .B(n[104]), .Z(n4713) );
  XOR U4705 ( .A(n3933), .B(n3929), .Z(n3930) );
  NANDN U4706 ( .A(n524), .B(n3930), .Z(n3931) );
  XNOR U4707 ( .A(n3932), .B(n3931), .Z(n5561) );
  NANDN U4708 ( .A(n3933), .B(n5561), .Z(n4711) );
  XNOR U4709 ( .A(n5561), .B(n3933), .Z(n4709) );
  XOR U4710 ( .A(n[102]), .B(n3934), .Z(n3935) );
  NANDN U4711 ( .A(n524), .B(n3935), .Z(n3936) );
  XNOR U4712 ( .A(n3937), .B(n3936), .Z(n5554) );
  NAND U4713 ( .A(n[102]), .B(n5554), .Z(n4707) );
  XOR U4714 ( .A(n[102]), .B(n5554), .Z(n4705) );
  XOR U4715 ( .A(n3942), .B(n3938), .Z(n3939) );
  NANDN U4716 ( .A(n524), .B(n3939), .Z(n3940) );
  XNOR U4717 ( .A(n3941), .B(n3940), .Z(n5551) );
  NANDN U4718 ( .A(n3942), .B(n5551), .Z(n4703) );
  XNOR U4719 ( .A(n5551), .B(n3942), .Z(n4701) );
  XNOR U4720 ( .A(n[100]), .B(n3943), .Z(n3944) );
  NANDN U4721 ( .A(n524), .B(n3944), .Z(n3945) );
  XNOR U4722 ( .A(n3946), .B(n3945), .Z(n5544) );
  NAND U4723 ( .A(n[100]), .B(n5544), .Z(n4699) );
  XOR U4724 ( .A(n[100]), .B(n5544), .Z(n4697) );
  XOR U4725 ( .A(n5344), .B(n3947), .Z(n3948) );
  NANDN U4726 ( .A(n524), .B(n3948), .Z(n3949) );
  XNOR U4727 ( .A(n3950), .B(n3949), .Z(n6866) );
  NANDN U4728 ( .A(n5344), .B(n6866), .Z(n4695) );
  XNOR U4729 ( .A(n6866), .B(n5344), .Z(n4693) );
  XNOR U4730 ( .A(n[98]), .B(n3951), .Z(n3952) );
  NANDN U4731 ( .A(n524), .B(n3952), .Z(n3953) );
  XNOR U4732 ( .A(n3954), .B(n3953), .Z(n5347) );
  NAND U4733 ( .A(n[98]), .B(n5347), .Z(n4691) );
  XOR U4734 ( .A(n[98]), .B(n5347), .Z(n4689) );
  XOR U4735 ( .A(n[97]), .B(n3955), .Z(n3956) );
  NANDN U4736 ( .A(n524), .B(n3956), .Z(n3957) );
  XNOR U4737 ( .A(n3958), .B(n3957), .Z(n6860) );
  NAND U4738 ( .A(n[97]), .B(n6860), .Z(n4687) );
  XOR U4739 ( .A(n6860), .B(n[97]), .Z(n4685) );
  XNOR U4740 ( .A(n3963), .B(n3959), .Z(n3960) );
  NANDN U4741 ( .A(n524), .B(n3960), .Z(n3961) );
  XNOR U4742 ( .A(n3962), .B(n3961), .Z(n5535) );
  NANDN U4743 ( .A(n3963), .B(n5535), .Z(n4683) );
  XNOR U4744 ( .A(n3963), .B(n5535), .Z(n4681) );
  XNOR U4745 ( .A(n5529), .B(n3964), .Z(n3965) );
  NANDN U4746 ( .A(n524), .B(n3965), .Z(n3966) );
  XNOR U4747 ( .A(n3967), .B(n3966), .Z(n5531) );
  XOR U4748 ( .A(n[95]), .B(n5531), .Z(n4677) );
  XNOR U4749 ( .A(n3969), .B(n3968), .Z(n3970) );
  NANDN U4750 ( .A(n524), .B(n3970), .Z(n3971) );
  XNOR U4751 ( .A(n3972), .B(n3971), .Z(n5350) );
  XNOR U4752 ( .A(n3974), .B(n3973), .Z(n3975) );
  NANDN U4753 ( .A(n524), .B(n3975), .Z(n3976) );
  XNOR U4754 ( .A(n3977), .B(n3976), .Z(n5352) );
  OR U4755 ( .A(n5352), .B(n[93]), .Z(n4671) );
  XOR U4756 ( .A(n5352), .B(n[93]), .Z(n4669) );
  XNOR U4757 ( .A(n[91]), .B(n3978), .Z(n3979) );
  NANDN U4758 ( .A(n524), .B(n3979), .Z(n3980) );
  XNOR U4759 ( .A(n3981), .B(n3980), .Z(n5359) );
  NAND U4760 ( .A(n[91]), .B(n5359), .Z(n4659) );
  XOR U4761 ( .A(n5359), .B(n[91]), .Z(n4657) );
  XOR U4762 ( .A(n[90]), .B(n3982), .Z(n3983) );
  NANDN U4763 ( .A(n524), .B(n3983), .Z(n3984) );
  XNOR U4764 ( .A(n3985), .B(n3984), .Z(n5361) );
  NAND U4765 ( .A(n[90]), .B(n5361), .Z(n4655) );
  XOR U4766 ( .A(n[90]), .B(n5361), .Z(n4653) );
  XNOR U4767 ( .A(n[89]), .B(n3986), .Z(n3987) );
  NANDN U4768 ( .A(n524), .B(n3987), .Z(n3988) );
  XNOR U4769 ( .A(n3989), .B(n3988), .Z(n5364) );
  NAND U4770 ( .A(n[89]), .B(n5364), .Z(n4651) );
  XOR U4771 ( .A(n5364), .B(n[89]), .Z(n4649) );
  XOR U4772 ( .A(n[88]), .B(n3990), .Z(n3991) );
  NANDN U4773 ( .A(n524), .B(n3991), .Z(n3992) );
  XNOR U4774 ( .A(n3993), .B(n3992), .Z(n5514) );
  NAND U4775 ( .A(n[88]), .B(n5514), .Z(n4647) );
  XOR U4776 ( .A(n[88]), .B(n5514), .Z(n4645) );
  XOR U4777 ( .A(n3998), .B(n3994), .Z(n3995) );
  NANDN U4778 ( .A(n524), .B(n3995), .Z(n3996) );
  XNOR U4779 ( .A(n3997), .B(n3996), .Z(n5366) );
  NANDN U4780 ( .A(n3998), .B(n5366), .Z(n4643) );
  XNOR U4781 ( .A(n5366), .B(n3998), .Z(n4641) );
  XOR U4782 ( .A(n[86]), .B(n3999), .Z(n4000) );
  NANDN U4783 ( .A(n524), .B(n4000), .Z(n4001) );
  XNOR U4784 ( .A(n4002), .B(n4001), .Z(n5368) );
  NAND U4785 ( .A(n[86]), .B(n5368), .Z(n4639) );
  XOR U4786 ( .A(n[86]), .B(n5368), .Z(n4637) );
  XOR U4787 ( .A(n5504), .B(n4003), .Z(n4004) );
  NANDN U4788 ( .A(n524), .B(n4004), .Z(n4005) );
  XNOR U4789 ( .A(n4006), .B(n4005), .Z(n5506) );
  NANDN U4790 ( .A(n5504), .B(n5506), .Z(n4635) );
  XNOR U4791 ( .A(n5506), .B(n5504), .Z(n4633) );
  XNOR U4792 ( .A(n[84]), .B(n4007), .Z(n4008) );
  NANDN U4793 ( .A(n524), .B(n4008), .Z(n4009) );
  XNOR U4794 ( .A(n4010), .B(n4009), .Z(n5370) );
  NAND U4795 ( .A(n[84]), .B(n5370), .Z(n4631) );
  XOR U4796 ( .A(n[84]), .B(n5370), .Z(n4629) );
  XNOR U4797 ( .A(n[83]), .B(n4011), .Z(n4012) );
  NANDN U4798 ( .A(n524), .B(n4012), .Z(n4013) );
  XNOR U4799 ( .A(n4014), .B(n4013), .Z(n5372) );
  NAND U4800 ( .A(n[83]), .B(n5372), .Z(n4627) );
  XOR U4801 ( .A(n5372), .B(n[83]), .Z(n4625) );
  XOR U4802 ( .A(n[82]), .B(n4015), .Z(n4016) );
  NANDN U4803 ( .A(n524), .B(n4016), .Z(n4017) );
  XNOR U4804 ( .A(n4018), .B(n4017), .Z(n5375) );
  NAND U4805 ( .A(n[82]), .B(n5375), .Z(n4623) );
  XOR U4806 ( .A(n5375), .B(n[82]), .Z(n4621) );
  XNOR U4807 ( .A(n4023), .B(n4019), .Z(n4020) );
  NANDN U4808 ( .A(n524), .B(n4020), .Z(n4021) );
  XNOR U4809 ( .A(n4022), .B(n4021), .Z(n5377) );
  NANDN U4810 ( .A(n4023), .B(n5377), .Z(n4619) );
  XNOR U4811 ( .A(n4023), .B(n5377), .Z(n4617) );
  XOR U4812 ( .A(n4028), .B(n4024), .Z(n4025) );
  NANDN U4813 ( .A(n524), .B(n4025), .Z(n4026) );
  XNOR U4814 ( .A(n4027), .B(n4026), .Z(n5379) );
  NANDN U4815 ( .A(n4028), .B(n5379), .Z(n4615) );
  XNOR U4816 ( .A(n5379), .B(n4028), .Z(n4613) );
  XNOR U4817 ( .A(n[79]), .B(n4029), .Z(n4030) );
  NANDN U4818 ( .A(n524), .B(n4030), .Z(n4031) );
  XNOR U4819 ( .A(n4032), .B(n4031), .Z(n6810) );
  NAND U4820 ( .A(n[79]), .B(n6810), .Z(n4611) );
  XOR U4821 ( .A(n6810), .B(n[79]), .Z(n4609) );
  XOR U4822 ( .A(n[78]), .B(n4033), .Z(n4034) );
  NANDN U4823 ( .A(n524), .B(n4034), .Z(n4035) );
  XNOR U4824 ( .A(n4036), .B(n4035), .Z(n5381) );
  NAND U4825 ( .A(n[78]), .B(n5381), .Z(n4607) );
  XOR U4826 ( .A(n[78]), .B(n5381), .Z(n4605) );
  XOR U4827 ( .A(n4041), .B(n4037), .Z(n4038) );
  NANDN U4828 ( .A(n524), .B(n4038), .Z(n4039) );
  XNOR U4829 ( .A(n4040), .B(n4039), .Z(n6804) );
  NANDN U4830 ( .A(n4041), .B(n6804), .Z(n4603) );
  XNOR U4831 ( .A(n6804), .B(n4041), .Z(n4601) );
  XNOR U4832 ( .A(n[76]), .B(n4042), .Z(n4043) );
  NANDN U4833 ( .A(n524), .B(n4043), .Z(n4044) );
  XNOR U4834 ( .A(n4045), .B(n4044), .Z(n5383) );
  NAND U4835 ( .A(n[76]), .B(n5383), .Z(n4599) );
  XOR U4836 ( .A(n5383), .B(n[76]), .Z(n4597) );
  XNOR U4837 ( .A(n[75]), .B(n4046), .Z(n4047) );
  NANDN U4838 ( .A(n524), .B(n4047), .Z(n4048) );
  XNOR U4839 ( .A(n4049), .B(n4048), .Z(n5487) );
  NAND U4840 ( .A(n[75]), .B(n5487), .Z(n4595) );
  XOR U4841 ( .A(n[75]), .B(n5487), .Z(n4593) );
  XNOR U4842 ( .A(n[74]), .B(n4050), .Z(n4051) );
  NANDN U4843 ( .A(n524), .B(n4051), .Z(n4052) );
  XNOR U4844 ( .A(n4053), .B(n4052), .Z(n5386) );
  NAND U4845 ( .A(n[74]), .B(n5386), .Z(n4591) );
  XOR U4846 ( .A(n5386), .B(n[74]), .Z(n4589) );
  XNOR U4847 ( .A(n[73]), .B(n4054), .Z(n4055) );
  NANDN U4848 ( .A(n524), .B(n4055), .Z(n4056) );
  XNOR U4849 ( .A(n4057), .B(n4056), .Z(n5388) );
  NAND U4850 ( .A(n[73]), .B(n5388), .Z(n4587) );
  XOR U4851 ( .A(n[73]), .B(n5388), .Z(n4585) );
  XNOR U4852 ( .A(n[72]), .B(n4058), .Z(n4059) );
  NANDN U4853 ( .A(n524), .B(n4059), .Z(n4060) );
  XNOR U4854 ( .A(n4061), .B(n4060), .Z(n5479) );
  NAND U4855 ( .A(n[72]), .B(n5479), .Z(n4583) );
  XOR U4856 ( .A(n5479), .B(n[72]), .Z(n4581) );
  XNOR U4857 ( .A(n5390), .B(n4062), .Z(n4063) );
  NANDN U4858 ( .A(n524), .B(n4063), .Z(n4064) );
  XOR U4859 ( .A(n4065), .B(n4064), .Z(n5475) );
  NANDN U4860 ( .A(n5475), .B(n[71]), .Z(n4579) );
  XOR U4861 ( .A(n5469), .B(n4066), .Z(n4067) );
  NANDN U4862 ( .A(n524), .B(n4067), .Z(n4068) );
  XOR U4863 ( .A(n4069), .B(n4068), .Z(n4573) );
  IV U4864 ( .A(n4573), .Z(n5471) );
  XNOR U4865 ( .A(n[69]), .B(n4070), .Z(n4071) );
  NANDN U4866 ( .A(n524), .B(n4071), .Z(n4072) );
  XNOR U4867 ( .A(n4073), .B(n4072), .Z(n5393) );
  NAND U4868 ( .A(n[69]), .B(n5393), .Z(n4570) );
  XOR U4869 ( .A(n5393), .B(n[69]), .Z(n4568) );
  XOR U4870 ( .A(n4078), .B(n4074), .Z(n4075) );
  NANDN U4871 ( .A(n524), .B(n4075), .Z(n4076) );
  XNOR U4872 ( .A(n4077), .B(n4076), .Z(n6774) );
  NANDN U4873 ( .A(n4078), .B(n6774), .Z(n4566) );
  XNOR U4874 ( .A(n4078), .B(n6774), .Z(n4564) );
  XNOR U4875 ( .A(n[67]), .B(n4079), .Z(n4080) );
  NANDN U4876 ( .A(n524), .B(n4080), .Z(n4081) );
  XNOR U4877 ( .A(n4082), .B(n4081), .Z(n5396) );
  NAND U4878 ( .A(n[67]), .B(n5396), .Z(n4562) );
  XOR U4879 ( .A(n5396), .B(n[67]), .Z(n4560) );
  XOR U4880 ( .A(n[66]), .B(n4083), .Z(n4084) );
  NANDN U4881 ( .A(n524), .B(n4084), .Z(n4085) );
  XNOR U4882 ( .A(n4086), .B(n4085), .Z(n6768) );
  NAND U4883 ( .A(n[66]), .B(n6768), .Z(n4558) );
  XOR U4884 ( .A(n6768), .B(n[66]), .Z(n4556) );
  XOR U4885 ( .A(n4091), .B(n4087), .Z(n4088) );
  NANDN U4886 ( .A(n524), .B(n4088), .Z(n4089) );
  XNOR U4887 ( .A(n4090), .B(n4089), .Z(n5398) );
  NANDN U4888 ( .A(n4091), .B(n5398), .Z(n4554) );
  XNOR U4889 ( .A(n4091), .B(n5398), .Z(n4552) );
  XOR U4890 ( .A(n5399), .B(n4092), .Z(n4093) );
  NANDN U4891 ( .A(n524), .B(n4093), .Z(n4094) );
  XOR U4892 ( .A(n4095), .B(n4094), .Z(n5402) );
  NANDN U4893 ( .A(n5399), .B(n5402), .Z(n4550) );
  XNOR U4894 ( .A(n5402), .B(n5399), .Z(n4548) );
  XOR U4895 ( .A(n[63]), .B(n4096), .Z(n4097) );
  NANDN U4896 ( .A(n524), .B(n4097), .Z(n4098) );
  XNOR U4897 ( .A(n4099), .B(n4098), .Z(n5458) );
  NAND U4898 ( .A(n[63]), .B(n5458), .Z(n4546) );
  XOR U4899 ( .A(n[63]), .B(n5458), .Z(n4544) );
  XNOR U4900 ( .A(n[62]), .B(n4100), .Z(n4101) );
  NANDN U4901 ( .A(n524), .B(n4101), .Z(n4102) );
  XOR U4902 ( .A(n4103), .B(n4102), .Z(n5404) );
  NAND U4903 ( .A(n[62]), .B(n5404), .Z(n4542) );
  XOR U4904 ( .A(n5404), .B(n[62]), .Z(n4540) );
  XNOR U4905 ( .A(n4108), .B(n4104), .Z(n4105) );
  NANDN U4906 ( .A(n524), .B(n4105), .Z(n4106) );
  XOR U4907 ( .A(n4107), .B(n4106), .Z(n5406) );
  NANDN U4908 ( .A(n4108), .B(n5406), .Z(n4538) );
  XNOR U4909 ( .A(n4108), .B(n5406), .Z(n4536) );
  XNOR U4910 ( .A(n4113), .B(n4109), .Z(n4110) );
  NANDN U4911 ( .A(n524), .B(n4110), .Z(n4111) );
  XNOR U4912 ( .A(n4112), .B(n4111), .Z(n5408) );
  NANDN U4913 ( .A(n4113), .B(n5408), .Z(n4534) );
  XNOR U4914 ( .A(n5408), .B(n4113), .Z(n4532) );
  XNOR U4915 ( .A(n4118), .B(n4114), .Z(n4115) );
  NANDN U4916 ( .A(n524), .B(n4115), .Z(n4116) );
  XOR U4917 ( .A(n4117), .B(n4116), .Z(n5410) );
  NANDN U4918 ( .A(n4118), .B(n5410), .Z(n4530) );
  XNOR U4919 ( .A(n4118), .B(n5410), .Z(n4528) );
  XNOR U4920 ( .A(n5411), .B(n4119), .Z(n4120) );
  NANDN U4921 ( .A(n524), .B(n4120), .Z(n4121) );
  XOR U4922 ( .A(n4122), .B(n4121), .Z(n5414) );
  NANDN U4923 ( .A(n5411), .B(n5414), .Z(n4526) );
  XNOR U4924 ( .A(n5414), .B(n5411), .Z(n4524) );
  XNOR U4925 ( .A(n[57]), .B(n4123), .Z(n4124) );
  NANDN U4926 ( .A(n524), .B(n4124), .Z(n4125) );
  XNOR U4927 ( .A(n4126), .B(n4125), .Z(n5417) );
  NAND U4928 ( .A(n[57]), .B(n5417), .Z(n4522) );
  XOR U4929 ( .A(n5417), .B(n[57]), .Z(n4520) );
  XOR U4930 ( .A(n4131), .B(n4127), .Z(n4128) );
  NANDN U4931 ( .A(n524), .B(n4128), .Z(n4129) );
  XNOR U4932 ( .A(n4130), .B(n4129), .Z(n5419) );
  NANDN U4933 ( .A(n4131), .B(n5419), .Z(n4518) );
  XNOR U4934 ( .A(n4131), .B(n5419), .Z(n4516) );
  XNOR U4935 ( .A(n[55]), .B(n4132), .Z(n4133) );
  NANDN U4936 ( .A(n524), .B(n4133), .Z(n4134) );
  XNOR U4937 ( .A(n4135), .B(n4134), .Z(n5421) );
  NAND U4938 ( .A(n[55]), .B(n5421), .Z(n4514) );
  XOR U4939 ( .A(n5421), .B(n[55]), .Z(n4512) );
  XNOR U4940 ( .A(n4140), .B(n4136), .Z(n4137) );
  NANDN U4941 ( .A(n524), .B(n4137), .Z(n4138) );
  XNOR U4942 ( .A(n4139), .B(n4138), .Z(n5423) );
  NANDN U4943 ( .A(n4140), .B(n5423), .Z(n4510) );
  XNOR U4944 ( .A(n4140), .B(n5423), .Z(n4508) );
  XNOR U4945 ( .A(n4145), .B(n4141), .Z(n4142) );
  NANDN U4946 ( .A(n524), .B(n4142), .Z(n4143) );
  XOR U4947 ( .A(n4144), .B(n4143), .Z(n6739) );
  NANDN U4948 ( .A(n4145), .B(n6739), .Z(n4506) );
  XNOR U4949 ( .A(n6739), .B(n4145), .Z(n4504) );
  XNOR U4950 ( .A(n[52]), .B(n4146), .Z(n4147) );
  NANDN U4951 ( .A(n524), .B(n4147), .Z(n4148) );
  XNOR U4952 ( .A(n4149), .B(n4148), .Z(n5426) );
  NAND U4953 ( .A(n5426), .B(n[52]), .Z(n4502) );
  XOR U4954 ( .A(n[52]), .B(n5426), .Z(n4500) );
  XOR U4955 ( .A(n[51]), .B(n4150), .Z(n4151) );
  NANDN U4956 ( .A(n524), .B(n4151), .Z(n4152) );
  XNOR U4957 ( .A(n4153), .B(n4152), .Z(n5428) );
  NAND U4958 ( .A(n[51]), .B(n5428), .Z(n4498) );
  XOR U4959 ( .A(n5428), .B(n[51]), .Z(n4496) );
  XOR U4960 ( .A(n[50]), .B(n4154), .Z(n4155) );
  NANDN U4961 ( .A(n524), .B(n4155), .Z(n4156) );
  XOR U4962 ( .A(n4157), .B(n4156), .Z(n6731) );
  NAND U4963 ( .A(n[50]), .B(n6731), .Z(n4494) );
  XOR U4964 ( .A(n[50]), .B(n6731), .Z(n4492) );
  IV U4965 ( .A(n[49]), .Z(n4162) );
  XNOR U4966 ( .A(n4162), .B(n4158), .Z(n4159) );
  NANDN U4967 ( .A(n524), .B(n4159), .Z(n4160) );
  XNOR U4968 ( .A(n4161), .B(n4160), .Z(n6723) );
  NANDN U4969 ( .A(n4162), .B(n6723), .Z(n4490) );
  XNOR U4970 ( .A(n6723), .B(n4162), .Z(n4488) );
  XNOR U4971 ( .A(n[48]), .B(n4163), .Z(n4164) );
  NANDN U4972 ( .A(n524), .B(n4164), .Z(n4165) );
  XOR U4973 ( .A(n4166), .B(n4165), .Z(n5432) );
  NAND U4974 ( .A(n[48]), .B(n5432), .Z(n4486) );
  XOR U4975 ( .A(n6716), .B(n4167), .Z(n4168) );
  NANDN U4976 ( .A(n524), .B(n4168), .Z(n4169) );
  XNOR U4977 ( .A(n4170), .B(n4169), .Z(n6719) );
  NANDN U4978 ( .A(n6716), .B(n6719), .Z(n4483) );
  XNOR U4979 ( .A(n6716), .B(n6719), .Z(n4481) );
  XOR U4980 ( .A(n6710), .B(n4171), .Z(n4172) );
  NANDN U4981 ( .A(n524), .B(n4172), .Z(n4173) );
  XOR U4982 ( .A(n4174), .B(n4173), .Z(n6714) );
  NANDN U4983 ( .A(n6710), .B(n6714), .Z(n4480) );
  NOR U4984 ( .A(n[46]), .B(n6714), .Z(n4478) );
  XNOR U4985 ( .A(n4179), .B(n4175), .Z(n4176) );
  NANDN U4986 ( .A(n524), .B(n4176), .Z(n4177) );
  XOR U4987 ( .A(n4178), .B(n4177), .Z(n6697) );
  NANDN U4988 ( .A(n4179), .B(n6697), .Z(n4461) );
  XNOR U4989 ( .A(n4179), .B(n6697), .Z(n4459) );
  IV U4990 ( .A(n[41]), .Z(n4454) );
  XOR U4991 ( .A(n4454), .B(n4180), .Z(n4181) );
  NANDN U4992 ( .A(n524), .B(n4181), .Z(n4182) );
  XOR U4993 ( .A(n4183), .B(n4182), .Z(n6690) );
  NANDN U4994 ( .A(n4454), .B(n6690), .Z(n4457) );
  XNOR U4995 ( .A(n4188), .B(n4184), .Z(n4185) );
  NANDN U4996 ( .A(n524), .B(n4185), .Z(n4186) );
  XOR U4997 ( .A(n4187), .B(n4186), .Z(n6686) );
  NANDN U4998 ( .A(n4188), .B(n6686), .Z(n4453) );
  XNOR U4999 ( .A(n4188), .B(n6686), .Z(n4451) );
  XOR U5000 ( .A(n4446), .B(n4189), .Z(n4190) );
  NANDN U5001 ( .A(n524), .B(n4190), .Z(n4191) );
  XNOR U5002 ( .A(n4192), .B(n4191), .Z(n6679) );
  NANDN U5003 ( .A(n4446), .B(n6679), .Z(n4449) );
  XOR U5004 ( .A(n4197), .B(n4193), .Z(n4194) );
  NANDN U5005 ( .A(n524), .B(n4194), .Z(n4195) );
  XNOR U5006 ( .A(n4196), .B(n4195), .Z(n6671) );
  NANDN U5007 ( .A(n4197), .B(n6671), .Z(n4445) );
  XNOR U5008 ( .A(n4197), .B(n6671), .Z(n4443) );
  XOR U5009 ( .A(n4438), .B(n4198), .Z(n4199) );
  NANDN U5010 ( .A(n524), .B(n4199), .Z(n4200) );
  XNOR U5011 ( .A(n4201), .B(n4200), .Z(n6664) );
  NANDN U5012 ( .A(n4438), .B(n6664), .Z(n4441) );
  XOR U5013 ( .A(n6656), .B(n4202), .Z(n4203) );
  NANDN U5014 ( .A(n524), .B(n4203), .Z(n4204) );
  XNOR U5015 ( .A(n4205), .B(n4204), .Z(n6658) );
  NANDN U5016 ( .A(n6656), .B(n6658), .Z(n4437) );
  XNOR U5017 ( .A(n[34]), .B(n4206), .Z(n4207) );
  NANDN U5018 ( .A(n524), .B(n4207), .Z(n4208) );
  XNOR U5019 ( .A(n4209), .B(n4208), .Z(n6648) );
  NAND U5020 ( .A(n[34]), .B(n6648), .Z(n4425) );
  XNOR U5021 ( .A(n[33]), .B(n4210), .Z(n4211) );
  NANDN U5022 ( .A(n524), .B(n4211), .Z(n4212) );
  XNOR U5023 ( .A(n4213), .B(n4212), .Z(n6644) );
  NAND U5024 ( .A(n[33]), .B(n6644), .Z(n4422) );
  XOR U5025 ( .A(n[32]), .B(n4214), .Z(n4215) );
  NANDN U5026 ( .A(n524), .B(n4215), .Z(n4216) );
  XNOR U5027 ( .A(n4217), .B(n4216), .Z(n6640) );
  XNOR U5028 ( .A(n4222), .B(n4218), .Z(n4219) );
  NANDN U5029 ( .A(n524), .B(n4219), .Z(n4220) );
  XNOR U5030 ( .A(n4221), .B(n4220), .Z(n6629) );
  NANDN U5031 ( .A(n4222), .B(n6629), .Z(n4414) );
  XNOR U5032 ( .A(n4222), .B(n6629), .Z(n4412) );
  XNOR U5033 ( .A(n4407), .B(n4223), .Z(n4224) );
  NANDN U5034 ( .A(n524), .B(n4224), .Z(n4225) );
  XNOR U5035 ( .A(n4226), .B(n4225), .Z(n6622) );
  NANDN U5036 ( .A(n4407), .B(n6622), .Z(n4410) );
  XNOR U5037 ( .A(n[26]), .B(n4227), .Z(n4228) );
  NANDN U5038 ( .A(n524), .B(n4228), .Z(n4229) );
  XNOR U5039 ( .A(n4230), .B(n4229), .Z(n6605) );
  NAND U5040 ( .A(n[26]), .B(n6605), .Z(n4397) );
  XOR U5041 ( .A(n[26]), .B(n6605), .Z(n4395) );
  XOR U5042 ( .A(n[25]), .B(n4231), .Z(n4232) );
  NANDN U5043 ( .A(n524), .B(n4232), .Z(n4233) );
  XNOR U5044 ( .A(n4234), .B(n4233), .Z(n6598) );
  NAND U5045 ( .A(n[25]), .B(n6598), .Z(n4393) );
  XNOR U5046 ( .A(n4239), .B(n4235), .Z(n4236) );
  NANDN U5047 ( .A(n524), .B(n4236), .Z(n4237) );
  XNOR U5048 ( .A(n4238), .B(n4237), .Z(n6544) );
  XNOR U5049 ( .A(n4382), .B(n4240), .Z(n4241) );
  NANDN U5050 ( .A(n524), .B(n4241), .Z(n4242) );
  XNOR U5051 ( .A(n4243), .B(n4242), .Z(n6406) );
  NANDN U5052 ( .A(n4382), .B(n6406), .Z(n4385) );
  XNOR U5053 ( .A(n4248), .B(n4244), .Z(n4245) );
  NANDN U5054 ( .A(n524), .B(n4245), .Z(n4246) );
  XNOR U5055 ( .A(n4247), .B(n4246), .Z(n6267) );
  NANDN U5056 ( .A(n4248), .B(n6267), .Z(n4377) );
  XNOR U5057 ( .A(n4248), .B(n6267), .Z(n4375) );
  XNOR U5058 ( .A(n4370), .B(n4249), .Z(n4250) );
  NANDN U5059 ( .A(n524), .B(n4250), .Z(n4251) );
  XNOR U5060 ( .A(n4252), .B(n4251), .Z(n6260) );
  NANDN U5061 ( .A(n4370), .B(n6260), .Z(n4373) );
  XNOR U5062 ( .A(n4257), .B(n4253), .Z(n4254) );
  NANDN U5063 ( .A(n524), .B(n4254), .Z(n4255) );
  XNOR U5064 ( .A(n4256), .B(n4255), .Z(n6129) );
  NANDN U5065 ( .A(n4257), .B(n6129), .Z(n4369) );
  XNOR U5066 ( .A(n4257), .B(n6129), .Z(n4367) );
  XNOR U5067 ( .A(n4362), .B(n4258), .Z(n4259) );
  NANDN U5068 ( .A(n524), .B(n4259), .Z(n4260) );
  XOR U5069 ( .A(n4261), .B(n4260), .Z(n6122) );
  NANDN U5070 ( .A(n4362), .B(n6122), .Z(n4365) );
  XNOR U5071 ( .A(n4266), .B(n4262), .Z(n4263) );
  NANDN U5072 ( .A(n524), .B(n4263), .Z(n4264) );
  XOR U5073 ( .A(n4265), .B(n4264), .Z(n5985) );
  IV U5074 ( .A(n[15]), .Z(n4358) );
  XNOR U5075 ( .A(n4271), .B(n4267), .Z(n4268) );
  NANDN U5076 ( .A(n524), .B(n4268), .Z(n4269) );
  XOR U5077 ( .A(n4270), .B(n4269), .Z(n5853) );
  NANDN U5078 ( .A(n4271), .B(n5853), .Z(n4356) );
  XNOR U5079 ( .A(n4271), .B(n5853), .Z(n4354) );
  XNOR U5080 ( .A(n4349), .B(n4272), .Z(n4273) );
  NANDN U5081 ( .A(n524), .B(n4273), .Z(n4274) );
  XOR U5082 ( .A(n4275), .B(n4274), .Z(n5846) );
  NANDN U5083 ( .A(n4349), .B(n5846), .Z(n4352) );
  XOR U5084 ( .A(n4276), .B(n[8]), .Z(n4277) );
  ANDN U5085 ( .B(n4277), .A(n524), .Z(n4278) );
  XNOR U5086 ( .A(n4279), .B(n4278), .Z(n6844) );
  NAND U5087 ( .A(n6844), .B(n[8]), .Z(n4325) );
  XOR U5088 ( .A(n[8]), .B(n6844), .Z(n4323) );
  IV U5089 ( .A(n[7]), .Z(n4318) );
  XNOR U5090 ( .A(n4318), .B(n4280), .Z(n4281) );
  ANDN U5091 ( .B(n4281), .A(n524), .Z(n4282) );
  XOR U5092 ( .A(n4283), .B(n4282), .Z(n6837) );
  NANDN U5093 ( .A(n4318), .B(n6837), .Z(n4321) );
  XOR U5094 ( .A(n[6]), .B(n4284), .Z(n4285) );
  NANDN U5095 ( .A(n524), .B(n4285), .Z(n4286) );
  XNOR U5096 ( .A(n4287), .B(n4286), .Z(n6788) );
  NAND U5097 ( .A(n[6]), .B(n6788), .Z(n4317) );
  XOR U5098 ( .A(n[6]), .B(n6788), .Z(n4315) );
  XOR U5099 ( .A(n4288), .B(n[5]), .Z(n4289) );
  ANDN U5100 ( .B(n4289), .A(n524), .Z(n4290) );
  XNOR U5101 ( .A(n4291), .B(n4290), .Z(n6781) );
  NAND U5102 ( .A(n[5]), .B(n6781), .Z(n4313) );
  XOR U5103 ( .A(n[4]), .B(n4292), .Z(n4293) );
  NANDN U5104 ( .A(n524), .B(n4293), .Z(n4294) );
  XNOR U5105 ( .A(n4295), .B(n4294), .Z(n6729) );
  NAND U5106 ( .A(n[4]), .B(n6729), .Z(n4310) );
  ANDN U5107 ( .B(n[0]), .A(n5342), .Z(n6195) );
  XOR U5108 ( .A(n[1]), .B(n4296), .Z(n4297) );
  NANDN U5109 ( .A(n524), .B(n4297), .Z(n4298) );
  XNOR U5110 ( .A(n4299), .B(n4298), .Z(n6198) );
  XNOR U5111 ( .A(n4300), .B(n6616), .Z(n4301) );
  ANDN U5112 ( .B(n4301), .A(n524), .Z(n4302) );
  XOR U5113 ( .A(n4303), .B(n4302), .Z(n6619) );
  XOR U5114 ( .A(n[3]), .B(n4304), .Z(n4305) );
  NANDN U5115 ( .A(n524), .B(n4305), .Z(n4306) );
  XNOR U5116 ( .A(n4307), .B(n4306), .Z(n6676) );
  XOR U5117 ( .A(n6729), .B(n[4]), .Z(n4308) );
  NANDN U5118 ( .A(n6726), .B(n4308), .Z(n4309) );
  AND U5119 ( .A(n4310), .B(n4309), .Z(n6754) );
  XOR U5120 ( .A(n6781), .B(n[5]), .Z(n4311) );
  NANDN U5121 ( .A(n6754), .B(n4311), .Z(n4312) );
  NAND U5122 ( .A(n4313), .B(n4312), .Z(n4314) );
  NAND U5123 ( .A(n4315), .B(n4314), .Z(n4316) );
  AND U5124 ( .A(n4317), .B(n4316), .Z(n6813) );
  XNOR U5125 ( .A(n6837), .B(n4318), .Z(n4319) );
  NANDN U5126 ( .A(n6813), .B(n4319), .Z(n4320) );
  NAND U5127 ( .A(n4321), .B(n4320), .Z(n4322) );
  NAND U5128 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U5129 ( .A(n4325), .B(n4324), .Z(n6867) );
  XOR U5130 ( .A(n6868), .B(n4326), .Z(n4327) );
  NANDN U5131 ( .A(n524), .B(n4327), .Z(n4328) );
  XNOR U5132 ( .A(n4329), .B(n4328), .Z(n6871) );
  XOR U5133 ( .A(n[10]), .B(n4330), .Z(n4331) );
  NANDN U5134 ( .A(n524), .B(n4331), .Z(n4332) );
  XNOR U5135 ( .A(n4333), .B(n4332), .Z(n5598) );
  XOR U5136 ( .A(n[10]), .B(n5598), .Z(n4334) );
  NANDN U5137 ( .A(n5595), .B(n4334), .Z(n4336) );
  NAND U5138 ( .A(n5598), .B(n[10]), .Z(n4335) );
  NAND U5139 ( .A(n4336), .B(n4335), .Z(n5655) );
  ANDN U5140 ( .B(n5655), .A(n4337), .Z(n4342) );
  XNOR U5141 ( .A(n4338), .B(n4337), .Z(n4339) );
  ANDN U5142 ( .B(n4339), .A(n524), .Z(n4340) );
  XNOR U5143 ( .A(n4341), .B(n4340), .Z(n5658) );
  OR U5144 ( .A(n4342), .B(n5658), .Z(n4344) );
  NOR U5145 ( .A(n[11]), .B(n5655), .Z(n4343) );
  ANDN U5146 ( .B(n4344), .A(n4343), .Z(n5716) );
  XOR U5147 ( .A(n[12]), .B(n4345), .Z(n4346) );
  NANDN U5148 ( .A(n524), .B(n4346), .Z(n4347) );
  XOR U5149 ( .A(n4348), .B(n4347), .Z(n5719) );
  XNOR U5150 ( .A(n5846), .B(n4349), .Z(n4350) );
  NANDN U5151 ( .A(n5782), .B(n4350), .Z(n4351) );
  NAND U5152 ( .A(n4352), .B(n4351), .Z(n4353) );
  NAND U5153 ( .A(n4354), .B(n4353), .Z(n4355) );
  NAND U5154 ( .A(n4356), .B(n4355), .Z(n5918) );
  XNOR U5155 ( .A(n4358), .B(n4357), .Z(n4359) );
  NANDN U5156 ( .A(n524), .B(n4359), .Z(n4360) );
  XNOR U5157 ( .A(n4361), .B(n4360), .Z(n5978) );
  XNOR U5158 ( .A(n6122), .B(n4362), .Z(n4363) );
  NANDN U5159 ( .A(n6054), .B(n4363), .Z(n4364) );
  NAND U5160 ( .A(n4365), .B(n4364), .Z(n4366) );
  NAND U5161 ( .A(n4367), .B(n4366), .Z(n4368) );
  AND U5162 ( .A(n4369), .B(n4368), .Z(n6194) );
  XNOR U5163 ( .A(n6260), .B(n4370), .Z(n4371) );
  NANDN U5164 ( .A(n6194), .B(n4371), .Z(n4372) );
  NAND U5165 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U5166 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U5167 ( .A(n4377), .B(n4376), .Z(n6331) );
  XOR U5168 ( .A(n[21]), .B(n4378), .Z(n4379) );
  NANDN U5169 ( .A(n524), .B(n4379), .Z(n4380) );
  XNOR U5170 ( .A(n4381), .B(n4380), .Z(n6334) );
  XNOR U5171 ( .A(n6406), .B(n4382), .Z(n4383) );
  NANDN U5172 ( .A(n6403), .B(n4383), .Z(n4384) );
  NAND U5173 ( .A(n4385), .B(n4384), .Z(n6473) );
  XNOR U5174 ( .A(n4387), .B(n4386), .Z(n4388) );
  NANDN U5175 ( .A(n524), .B(n4388), .Z(n4389) );
  XNOR U5176 ( .A(n4390), .B(n4389), .Z(n6537) );
  XOR U5177 ( .A(n6598), .B(n[25]), .Z(n4391) );
  NANDN U5178 ( .A(n6595), .B(n4391), .Z(n4392) );
  NAND U5179 ( .A(n4393), .B(n4392), .Z(n4394) );
  NAND U5180 ( .A(n4395), .B(n4394), .Z(n4396) );
  NAND U5181 ( .A(n4397), .B(n4396), .Z(n6606) );
  XOR U5182 ( .A(n4399), .B(n4398), .Z(n4400) );
  NANDN U5183 ( .A(n524), .B(n4400), .Z(n4401) );
  XOR U5184 ( .A(n4402), .B(n4401), .Z(n6609) );
  XNOR U5185 ( .A(n[28]), .B(n4403), .Z(n4404) );
  NANDN U5186 ( .A(n524), .B(n4404), .Z(n4405) );
  XNOR U5187 ( .A(n4406), .B(n4405), .Z(n6613) );
  XNOR U5188 ( .A(n6622), .B(n4407), .Z(n4408) );
  NANDN U5189 ( .A(n6614), .B(n4408), .Z(n4409) );
  NAND U5190 ( .A(n4410), .B(n4409), .Z(n4411) );
  NAND U5191 ( .A(n4412), .B(n4411), .Z(n4413) );
  NAND U5192 ( .A(n4414), .B(n4413), .Z(n6630) );
  XNOR U5193 ( .A(n4416), .B(n4415), .Z(n4417) );
  NANDN U5194 ( .A(n524), .B(n4417), .Z(n4418) );
  XNOR U5195 ( .A(n4419), .B(n4418), .Z(n6633) );
  XOR U5196 ( .A(n6644), .B(n[33]), .Z(n4420) );
  NANDN U5197 ( .A(n6641), .B(n4420), .Z(n4421) );
  AND U5198 ( .A(n4422), .B(n4421), .Z(n6645) );
  XOR U5199 ( .A(n[34]), .B(n6648), .Z(n4423) );
  NANDN U5200 ( .A(n6645), .B(n4423), .Z(n4424) );
  AND U5201 ( .A(n4425), .B(n4424), .Z(n6649) );
  NANDN U5202 ( .A(n[35]), .B(n6649), .Z(n4427) );
  NOR U5203 ( .A(n[36]), .B(n6658), .Z(n4426) );
  ANDN U5204 ( .B(n4427), .A(n4426), .Z(n4435) );
  XOR U5205 ( .A(n4432), .B(n4428), .Z(n4429) );
  NANDN U5206 ( .A(n524), .B(n4429), .Z(n4430) );
  XNOR U5207 ( .A(n4431), .B(n4430), .Z(n6650) );
  XOR U5208 ( .A(n4432), .B(n6649), .Z(n4433) );
  NANDN U5209 ( .A(n6650), .B(n4433), .Z(n4434) );
  NAND U5210 ( .A(n4435), .B(n4434), .Z(n4436) );
  AND U5211 ( .A(n4437), .B(n4436), .Z(n6661) );
  XNOR U5212 ( .A(n6664), .B(n4438), .Z(n4439) );
  NANDN U5213 ( .A(n6661), .B(n4439), .Z(n4440) );
  NAND U5214 ( .A(n4441), .B(n4440), .Z(n4442) );
  NAND U5215 ( .A(n4443), .B(n4442), .Z(n4444) );
  AND U5216 ( .A(n4445), .B(n4444), .Z(n6672) );
  XNOR U5217 ( .A(n6679), .B(n4446), .Z(n4447) );
  NANDN U5218 ( .A(n6672), .B(n4447), .Z(n4448) );
  NAND U5219 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U5220 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U5221 ( .A(n4453), .B(n4452), .Z(n6687) );
  XNOR U5222 ( .A(n6690), .B(n4454), .Z(n4455) );
  NANDN U5223 ( .A(n6687), .B(n4455), .Z(n4456) );
  NAND U5224 ( .A(n4457), .B(n4456), .Z(n4458) );
  NAND U5225 ( .A(n4459), .B(n4458), .Z(n4460) );
  NAND U5226 ( .A(n4461), .B(n4460), .Z(n6698) );
  IV U5227 ( .A(n[43]), .Z(n4463) );
  XNOR U5228 ( .A(n4463), .B(n4462), .Z(n4464) );
  NANDN U5229 ( .A(n524), .B(n4464), .Z(n4465) );
  XNOR U5230 ( .A(n4466), .B(n4465), .Z(n6701) );
  XOR U5231 ( .A(n[44]), .B(n4467), .Z(n4468) );
  NANDN U5232 ( .A(n524), .B(n4468), .Z(n4469) );
  XNOR U5233 ( .A(n4470), .B(n4469), .Z(n6705) );
  XNOR U5234 ( .A(n[45]), .B(n4471), .Z(n4472) );
  NANDN U5235 ( .A(n524), .B(n4472), .Z(n4473) );
  XNOR U5236 ( .A(n4474), .B(n4473), .Z(n6709) );
  XOR U5237 ( .A(n[45]), .B(n6709), .Z(n4475) );
  NANDN U5238 ( .A(n6706), .B(n4475), .Z(n4477) );
  NAND U5239 ( .A(n[45]), .B(n6709), .Z(n4476) );
  NAND U5240 ( .A(n4477), .B(n4476), .Z(n6711) );
  NANDN U5241 ( .A(n4478), .B(n6711), .Z(n4479) );
  NAND U5242 ( .A(n4480), .B(n4479), .Z(n6715) );
  NAND U5243 ( .A(n4481), .B(n6715), .Z(n4482) );
  AND U5244 ( .A(n4483), .B(n4482), .Z(n5430) );
  XOR U5245 ( .A(n5432), .B(n[48]), .Z(n4484) );
  NANDN U5246 ( .A(n5430), .B(n4484), .Z(n4485) );
  NAND U5247 ( .A(n4486), .B(n4485), .Z(n4487) );
  NAND U5248 ( .A(n4488), .B(n4487), .Z(n4489) );
  NAND U5249 ( .A(n4490), .B(n4489), .Z(n4491) );
  NAND U5250 ( .A(n4492), .B(n4491), .Z(n4493) );
  NAND U5251 ( .A(n4494), .B(n4493), .Z(n4495) );
  NAND U5252 ( .A(n4496), .B(n4495), .Z(n4497) );
  NAND U5253 ( .A(n4498), .B(n4497), .Z(n4499) );
  NAND U5254 ( .A(n4500), .B(n4499), .Z(n4501) );
  NAND U5255 ( .A(n4502), .B(n4501), .Z(n4503) );
  NAND U5256 ( .A(n4504), .B(n4503), .Z(n4505) );
  NAND U5257 ( .A(n4506), .B(n4505), .Z(n4507) );
  NAND U5258 ( .A(n4508), .B(n4507), .Z(n4509) );
  NAND U5259 ( .A(n4510), .B(n4509), .Z(n4511) );
  NAND U5260 ( .A(n4512), .B(n4511), .Z(n4513) );
  NAND U5261 ( .A(n4514), .B(n4513), .Z(n4515) );
  NAND U5262 ( .A(n4516), .B(n4515), .Z(n4517) );
  NAND U5263 ( .A(n4518), .B(n4517), .Z(n4519) );
  NAND U5264 ( .A(n4520), .B(n4519), .Z(n4521) );
  NAND U5265 ( .A(n4522), .B(n4521), .Z(n4523) );
  NAND U5266 ( .A(n4524), .B(n4523), .Z(n4525) );
  NAND U5267 ( .A(n4526), .B(n4525), .Z(n4527) );
  NAND U5268 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U5269 ( .A(n4530), .B(n4529), .Z(n4531) );
  NAND U5270 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U5271 ( .A(n4534), .B(n4533), .Z(n4535) );
  NAND U5272 ( .A(n4536), .B(n4535), .Z(n4537) );
  NAND U5273 ( .A(n4538), .B(n4537), .Z(n4539) );
  NAND U5274 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U5275 ( .A(n4542), .B(n4541), .Z(n4543) );
  NAND U5276 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U5277 ( .A(n4546), .B(n4545), .Z(n4547) );
  NAND U5278 ( .A(n4548), .B(n4547), .Z(n4549) );
  NAND U5279 ( .A(n4550), .B(n4549), .Z(n4551) );
  NAND U5280 ( .A(n4552), .B(n4551), .Z(n4553) );
  NAND U5281 ( .A(n4554), .B(n4553), .Z(n4555) );
  NAND U5282 ( .A(n4556), .B(n4555), .Z(n4557) );
  NAND U5283 ( .A(n4558), .B(n4557), .Z(n4559) );
  NAND U5284 ( .A(n4560), .B(n4559), .Z(n4561) );
  NAND U5285 ( .A(n4562), .B(n4561), .Z(n4563) );
  NAND U5286 ( .A(n4564), .B(n4563), .Z(n4565) );
  NAND U5287 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U5288 ( .A(n4568), .B(n4567), .Z(n4569) );
  AND U5289 ( .A(n4570), .B(n4569), .Z(n4574) );
  NANDN U5290 ( .A(n5471), .B(n4574), .Z(n4572) );
  ANDN U5291 ( .B(n5475), .A(n[71]), .Z(n4571) );
  ANDN U5292 ( .B(n4572), .A(n4571), .Z(n4577) );
  XOR U5293 ( .A(n4574), .B(n4573), .Z(n4575) );
  NANDN U5294 ( .A(n[70]), .B(n4575), .Z(n4576) );
  NAND U5295 ( .A(n4577), .B(n4576), .Z(n4578) );
  NAND U5296 ( .A(n4579), .B(n4578), .Z(n4580) );
  NAND U5297 ( .A(n4581), .B(n4580), .Z(n4582) );
  NAND U5298 ( .A(n4583), .B(n4582), .Z(n4584) );
  NAND U5299 ( .A(n4585), .B(n4584), .Z(n4586) );
  NAND U5300 ( .A(n4587), .B(n4586), .Z(n4588) );
  NAND U5301 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U5302 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U5303 ( .A(n4593), .B(n4592), .Z(n4594) );
  NAND U5304 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U5305 ( .A(n4597), .B(n4596), .Z(n4598) );
  NAND U5306 ( .A(n4599), .B(n4598), .Z(n4600) );
  NAND U5307 ( .A(n4601), .B(n4600), .Z(n4602) );
  NAND U5308 ( .A(n4603), .B(n4602), .Z(n4604) );
  NAND U5309 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U5310 ( .A(n4607), .B(n4606), .Z(n4608) );
  NAND U5311 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U5312 ( .A(n4611), .B(n4610), .Z(n4612) );
  NAND U5313 ( .A(n4613), .B(n4612), .Z(n4614) );
  NAND U5314 ( .A(n4615), .B(n4614), .Z(n4616) );
  NAND U5315 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U5316 ( .A(n4619), .B(n4618), .Z(n4620) );
  NAND U5317 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U5318 ( .A(n4623), .B(n4622), .Z(n4624) );
  NAND U5319 ( .A(n4625), .B(n4624), .Z(n4626) );
  NAND U5320 ( .A(n4627), .B(n4626), .Z(n4628) );
  NAND U5321 ( .A(n4629), .B(n4628), .Z(n4630) );
  NAND U5322 ( .A(n4631), .B(n4630), .Z(n4632) );
  NAND U5323 ( .A(n4633), .B(n4632), .Z(n4634) );
  NAND U5324 ( .A(n4635), .B(n4634), .Z(n4636) );
  NAND U5325 ( .A(n4637), .B(n4636), .Z(n4638) );
  NAND U5326 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U5327 ( .A(n4641), .B(n4640), .Z(n4642) );
  NAND U5328 ( .A(n4643), .B(n4642), .Z(n4644) );
  NAND U5329 ( .A(n4645), .B(n4644), .Z(n4646) );
  NAND U5330 ( .A(n4647), .B(n4646), .Z(n4648) );
  NAND U5331 ( .A(n4649), .B(n4648), .Z(n4650) );
  NAND U5332 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U5333 ( .A(n4653), .B(n4652), .Z(n4654) );
  NAND U5334 ( .A(n4655), .B(n4654), .Z(n4656) );
  NAND U5335 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U5336 ( .A(n4659), .B(n4658), .Z(n4665) );
  XNOR U5337 ( .A(n5353), .B(n4660), .Z(n4661) );
  NANDN U5338 ( .A(n524), .B(n4661), .Z(n4662) );
  XNOR U5339 ( .A(n4663), .B(n4662), .Z(n5356) );
  XNOR U5340 ( .A(n4665), .B(n5356), .Z(n4664) );
  NANDN U5341 ( .A(n5353), .B(n4664), .Z(n4667) );
  NANDN U5342 ( .A(n4665), .B(n5356), .Z(n4666) );
  AND U5343 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U5344 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U5345 ( .A(n4671), .B(n4670), .Z(n4672) );
  OR U5346 ( .A(n5350), .B(n4672), .Z(n4675) );
  XOR U5347 ( .A(n5350), .B(n4672), .Z(n4673) );
  NANDN U5348 ( .A(n[94]), .B(n4673), .Z(n4674) );
  NAND U5349 ( .A(n4675), .B(n4674), .Z(n4676) );
  NAND U5350 ( .A(n4677), .B(n4676), .Z(n4679) );
  NANDN U5351 ( .A(n5531), .B(n5529), .Z(n4678) );
  AND U5352 ( .A(n4679), .B(n4678), .Z(n4680) );
  NAND U5353 ( .A(n4681), .B(n4680), .Z(n4682) );
  NAND U5354 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U5355 ( .A(n4685), .B(n4684), .Z(n4686) );
  NAND U5356 ( .A(n4687), .B(n4686), .Z(n4688) );
  NAND U5357 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U5358 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U5359 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U5360 ( .A(n4695), .B(n4694), .Z(n4696) );
  NAND U5361 ( .A(n4697), .B(n4696), .Z(n4698) );
  NAND U5362 ( .A(n4699), .B(n4698), .Z(n4700) );
  NAND U5363 ( .A(n4701), .B(n4700), .Z(n4702) );
  NAND U5364 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U5365 ( .A(n4705), .B(n4704), .Z(n4706) );
  NAND U5366 ( .A(n4707), .B(n4706), .Z(n4708) );
  NAND U5367 ( .A(n4709), .B(n4708), .Z(n4710) );
  NAND U5368 ( .A(n4711), .B(n4710), .Z(n4712) );
  NAND U5369 ( .A(n4713), .B(n4712), .Z(n4714) );
  NAND U5370 ( .A(n4715), .B(n4714), .Z(n4716) );
  NAND U5371 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U5372 ( .A(n4719), .B(n4718), .Z(n4720) );
  NAND U5373 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U5374 ( .A(n4723), .B(n4722), .Z(n4724) );
  NAND U5375 ( .A(n4725), .B(n4724), .Z(n4726) );
  NAND U5376 ( .A(n4727), .B(n4726), .Z(n4728) );
  NAND U5377 ( .A(n4729), .B(n4728), .Z(n4730) );
  NAND U5378 ( .A(n4731), .B(n4730), .Z(n4732) );
  NAND U5379 ( .A(n4733), .B(n4732), .Z(n4734) );
  NAND U5380 ( .A(n4735), .B(n4734), .Z(n4736) );
  NAND U5381 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U5382 ( .A(n4739), .B(n4738), .Z(n4740) );
  NAND U5383 ( .A(n4741), .B(n4740), .Z(n4742) );
  NAND U5384 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U5385 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U5386 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U5387 ( .A(n4749), .B(n4748), .Z(n4750) );
  NAND U5388 ( .A(n4751), .B(n4750), .Z(n4752) );
  NAND U5389 ( .A(n4753), .B(n4752), .Z(n4754) );
  NAND U5390 ( .A(n4755), .B(n4754), .Z(n4756) );
  NAND U5391 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5392 ( .A(n4759), .B(n4758), .Z(n4760) );
  NAND U5393 ( .A(n4761), .B(n4760), .Z(n4762) );
  NAND U5394 ( .A(n4763), .B(n4762), .Z(n4764) );
  NAND U5395 ( .A(n4765), .B(n4764), .Z(n4766) );
  NAND U5396 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U5397 ( .A(n4769), .B(n4768), .Z(n4770) );
  NAND U5398 ( .A(n4771), .B(n4770), .Z(n4772) );
  NAND U5399 ( .A(n4773), .B(n4772), .Z(n4774) );
  NAND U5400 ( .A(n4775), .B(n4774), .Z(n4776) );
  NAND U5401 ( .A(n4777), .B(n4776), .Z(n4778) );
  NAND U5402 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U5403 ( .A(n4781), .B(n4780), .Z(n4782) );
  NAND U5404 ( .A(n4783), .B(n4782), .Z(n4784) );
  NAND U5405 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U5406 ( .A(n4787), .B(n4786), .Z(n4788) );
  NAND U5407 ( .A(n4789), .B(n4788), .Z(n4790) );
  NAND U5408 ( .A(n4791), .B(n4790), .Z(n4792) );
  NAND U5409 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U5410 ( .A(n4795), .B(n4794), .Z(n4796) );
  NAND U5411 ( .A(n4797), .B(n4796), .Z(n4798) );
  NAND U5412 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U5413 ( .A(n4801), .B(n4800), .Z(n4802) );
  NAND U5414 ( .A(n4803), .B(n4802), .Z(n4804) );
  NAND U5415 ( .A(n4805), .B(n4804), .Z(n4806) );
  NAND U5416 ( .A(n4807), .B(n4806), .Z(n4808) );
  NAND U5417 ( .A(n4809), .B(n4808), .Z(n4810) );
  NAND U5418 ( .A(n4811), .B(n4810), .Z(n4812) );
  NAND U5419 ( .A(n4813), .B(n4812), .Z(n4814) );
  NAND U5420 ( .A(n4815), .B(n4814), .Z(n4816) );
  NAND U5421 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U5422 ( .A(n4819), .B(n4818), .Z(n4820) );
  NAND U5423 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U5424 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U5425 ( .A(n4825), .B(n4824), .Z(n4826) );
  NAND U5426 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5427 ( .A(n4829), .B(n4828), .Z(n4830) );
  NAND U5428 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U5429 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U5430 ( .A(n4835), .B(n4834), .Z(n4836) );
  NAND U5431 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U5432 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U5433 ( .A(n4841), .B(n4840), .Z(n4842) );
  NAND U5434 ( .A(n4843), .B(n4842), .Z(n4844) );
  NAND U5435 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5436 ( .A(n4847), .B(n4846), .Z(n4848) );
  NAND U5437 ( .A(n4849), .B(n4848), .Z(n4850) );
  NAND U5438 ( .A(n4851), .B(n4850), .Z(n4852) );
  NAND U5439 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U5440 ( .A(n4855), .B(n4854), .Z(n4856) );
  NAND U5441 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U5442 ( .A(n4859), .B(n4858), .Z(n4860) );
  NAND U5443 ( .A(n4861), .B(n4860), .Z(n4862) );
  NAND U5444 ( .A(n4863), .B(n4862), .Z(n4864) );
  NAND U5445 ( .A(n4865), .B(n4864), .Z(n4866) );
  NAND U5446 ( .A(n4867), .B(n4866), .Z(n4868) );
  NAND U5447 ( .A(n4869), .B(n4868), .Z(n4870) );
  NAND U5448 ( .A(n4871), .B(n4870), .Z(n4872) );
  NAND U5449 ( .A(n4873), .B(n4872), .Z(n4874) );
  NAND U5450 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U5451 ( .A(n4877), .B(n4876), .Z(n4878) );
  NAND U5452 ( .A(n4879), .B(n4878), .Z(n4880) );
  NAND U5453 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U5454 ( .A(n4883), .B(n4882), .Z(n4884) );
  NAND U5455 ( .A(n4885), .B(n4884), .Z(n4886) );
  NAND U5456 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U5457 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U5458 ( .A(n4891), .B(n4890), .Z(n4892) );
  NAND U5459 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U5460 ( .A(n4895), .B(n4894), .Z(n4896) );
  NAND U5461 ( .A(n4897), .B(n4896), .Z(n4898) );
  NAND U5462 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U5463 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U5464 ( .A(n4903), .B(n4902), .Z(n4904) );
  NAND U5465 ( .A(n4905), .B(n4904), .Z(n4906) );
  AND U5466 ( .A(n4907), .B(n4906), .Z(n4908) );
  OR U5467 ( .A(n4908), .B(n4910), .Z(n4916) );
  XOR U5468 ( .A(n4908), .B(n4910), .Z(n4914) );
  XOR U5469 ( .A(n4910), .B(n4909), .Z(n4911) );
  NANDN U5470 ( .A(n524), .B(n4911), .Z(n4912) );
  XNOR U5471 ( .A(n4913), .B(n4912), .Z(n5879) );
  NAND U5472 ( .A(n4914), .B(n5879), .Z(n4915) );
  NAND U5473 ( .A(n4916), .B(n4915), .Z(n4917) );
  NAND U5474 ( .A(n4918), .B(n4917), .Z(n4919) );
  AND U5475 ( .A(n4920), .B(n4919), .Z(n4922) );
  NANDN U5476 ( .A(n4922), .B(n[155]), .Z(n4921) );
  AND U5477 ( .A(n5898), .B(n4921), .Z(n4929) );
  XNOR U5478 ( .A(n[155]), .B(n4922), .Z(n4927) );
  XOR U5479 ( .A(n[155]), .B(n4923), .Z(n4924) );
  NANDN U5480 ( .A(n524), .B(n4924), .Z(n4925) );
  XNOR U5481 ( .A(n4926), .B(n4925), .Z(n5892) );
  NAND U5482 ( .A(n4927), .B(n5892), .Z(n4928) );
  NAND U5483 ( .A(n4929), .B(n4928), .Z(n4930) );
  NAND U5484 ( .A(n4931), .B(n4930), .Z(n4938) );
  NANDN U5485 ( .A(n[157]), .B(n4938), .Z(n4933) );
  NOR U5486 ( .A(n[158]), .B(n5905), .Z(n4932) );
  ANDN U5487 ( .B(n4933), .A(n4932), .Z(n4942) );
  XNOR U5488 ( .A(n4939), .B(n4934), .Z(n4935) );
  NANDN U5489 ( .A(n524), .B(n4935), .Z(n4936) );
  XNOR U5490 ( .A(n4937), .B(n4936), .Z(n5906) );
  XOR U5491 ( .A(n4939), .B(n4938), .Z(n4940) );
  NANDN U5492 ( .A(n5906), .B(n4940), .Z(n4941) );
  NAND U5493 ( .A(n4942), .B(n4941), .Z(n4943) );
  NANDN U5494 ( .A(n5912), .B(n4943), .Z(n4944) );
  NAND U5495 ( .A(n4945), .B(n4944), .Z(n4946) );
  NAND U5496 ( .A(n4947), .B(n4946), .Z(n4948) );
  NAND U5497 ( .A(n4949), .B(n4948), .Z(n4950) );
  NAND U5498 ( .A(n4951), .B(n4950), .Z(n4952) );
  NAND U5499 ( .A(n4953), .B(n4952), .Z(n4954) );
  NAND U5500 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U5501 ( .A(n4957), .B(n4956), .Z(n4958) );
  NAND U5502 ( .A(n4959), .B(n4958), .Z(n4960) );
  NAND U5503 ( .A(n4961), .B(n4960), .Z(n4962) );
  NAND U5504 ( .A(n4963), .B(n4962), .Z(n4964) );
  NAND U5505 ( .A(n4965), .B(n4964), .Z(n4966) );
  NAND U5506 ( .A(n4967), .B(n4966), .Z(n4968) );
  NAND U5507 ( .A(n4969), .B(n4968), .Z(n4970) );
  NAND U5508 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U5509 ( .A(n4973), .B(n4972), .Z(n4974) );
  NAND U5510 ( .A(n4975), .B(n4974), .Z(n4976) );
  NAND U5511 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5512 ( .A(n4979), .B(n4978), .Z(n4980) );
  NAND U5513 ( .A(n4981), .B(n4980), .Z(n4982) );
  NAND U5514 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5515 ( .A(n4985), .B(n4984), .Z(n4986) );
  NAND U5516 ( .A(n4987), .B(n4986), .Z(n4988) );
  NAND U5517 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U5518 ( .A(n4991), .B(n4990), .Z(n4992) );
  NAND U5519 ( .A(n4993), .B(n4992), .Z(n4994) );
  NAND U5520 ( .A(n4995), .B(n4994), .Z(n4996) );
  NAND U5521 ( .A(n4997), .B(n4996), .Z(n4998) );
  NAND U5522 ( .A(n4999), .B(n4998), .Z(n5000) );
  NAND U5523 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U5524 ( .A(n5003), .B(n5002), .Z(n5004) );
  NAND U5525 ( .A(n5005), .B(n5004), .Z(n5006) );
  NAND U5526 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U5527 ( .A(n5009), .B(n5008), .Z(n5010) );
  NAND U5528 ( .A(n5011), .B(n5010), .Z(n5012) );
  NAND U5529 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U5530 ( .A(n5015), .B(n5014), .Z(n5016) );
  NAND U5531 ( .A(n5017), .B(n5016), .Z(n5018) );
  NAND U5532 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U5533 ( .A(n5021), .B(n5020), .Z(n5022) );
  NANDN U5534 ( .A(n5022), .B(n[179]), .Z(n5029) );
  XNOR U5535 ( .A(n5022), .B(n[179]), .Z(n5027) );
  XNOR U5536 ( .A(n[179]), .B(n5023), .Z(n5024) );
  NANDN U5537 ( .A(n524), .B(n5024), .Z(n5025) );
  XNOR U5538 ( .A(n5026), .B(n5025), .Z(n6055) );
  NAND U5539 ( .A(n5027), .B(n6055), .Z(n5028) );
  NAND U5540 ( .A(n5029), .B(n5028), .Z(n5030) );
  NAND U5541 ( .A(n5031), .B(n5030), .Z(n5032) );
  NAND U5542 ( .A(n5033), .B(n5032), .Z(n5034) );
  NAND U5543 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U5544 ( .A(n5037), .B(n5036), .Z(n5038) );
  NAND U5545 ( .A(n5039), .B(n5038), .Z(n5040) );
  NAND U5546 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U5547 ( .A(n5043), .B(n5042), .Z(n5044) );
  NAND U5548 ( .A(n5045), .B(n5044), .Z(n5046) );
  NAND U5549 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U5550 ( .A(n5049), .B(n5048), .Z(n5050) );
  NANDN U5551 ( .A(n5050), .B(n[185]), .Z(n5057) );
  XNOR U5552 ( .A(n5050), .B(n[185]), .Z(n5055) );
  XOR U5553 ( .A(n[185]), .B(n5051), .Z(n5052) );
  NANDN U5554 ( .A(n524), .B(n5052), .Z(n5053) );
  XNOR U5555 ( .A(n5054), .B(n5053), .Z(n6093) );
  NAND U5556 ( .A(n5055), .B(n6093), .Z(n5056) );
  NAND U5557 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U5558 ( .A(n5059), .B(n5058), .Z(n5060) );
  NAND U5559 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U5560 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U5561 ( .A(n5065), .B(n5064), .Z(n5066) );
  NAND U5562 ( .A(n5067), .B(n5066), .Z(n5068) );
  NAND U5563 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND U5564 ( .A(n5071), .B(n5070), .Z(n5072) );
  NAND U5565 ( .A(n5073), .B(n5072), .Z(n5074) );
  NAND U5566 ( .A(n5075), .B(n5074), .Z(n5076) );
  NAND U5567 ( .A(n5077), .B(n5076), .Z(n5078) );
  NAND U5568 ( .A(n5079), .B(n5078), .Z(n5080) );
  NAND U5569 ( .A(n5081), .B(n5080), .Z(n5082) );
  NAND U5570 ( .A(n5083), .B(n5082), .Z(n5084) );
  NAND U5571 ( .A(n5085), .B(n5084), .Z(n5086) );
  NAND U5572 ( .A(n5087), .B(n5086), .Z(n5088) );
  NAND U5573 ( .A(n5089), .B(n5088), .Z(n5090) );
  NAND U5574 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U5575 ( .A(n5093), .B(n5092), .Z(n5094) );
  NAND U5576 ( .A(n5095), .B(n5094), .Z(n5096) );
  NAND U5577 ( .A(n5097), .B(n5096), .Z(n5099) );
  OR U5578 ( .A(n6168), .B(n[196]), .Z(n5098) );
  AND U5579 ( .A(n5099), .B(n5098), .Z(n5100) );
  NAND U5580 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U5581 ( .A(n5103), .B(n5102), .Z(n5104) );
  NAND U5582 ( .A(n5105), .B(n5104), .Z(n5106) );
  NAND U5583 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U5584 ( .A(n5109), .B(n5108), .Z(n5110) );
  NAND U5585 ( .A(n5111), .B(n5110), .Z(n5113) );
  OR U5586 ( .A(n6201), .B(n[200]), .Z(n5112) );
  AND U5587 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5588 ( .A(n5115), .B(n5114), .Z(n5116) );
  NAND U5589 ( .A(n5117), .B(n5116), .Z(n5118) );
  NAND U5590 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U5591 ( .A(n5121), .B(n5120), .Z(n5122) );
  NAND U5592 ( .A(n5123), .B(n5122), .Z(n5124) );
  NAND U5593 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U5594 ( .A(n5127), .B(n5126), .Z(n5128) );
  NAND U5595 ( .A(n5129), .B(n5128), .Z(n5130) );
  NAND U5596 ( .A(n5131), .B(n5130), .Z(n5132) );
  NAND U5597 ( .A(n5133), .B(n5132), .Z(n5134) );
  NAND U5598 ( .A(n5135), .B(n5134), .Z(n5136) );
  NAND U5599 ( .A(n5137), .B(n5136), .Z(n5138) );
  NAND U5600 ( .A(n5139), .B(n5138), .Z(n5140) );
  NAND U5601 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5602 ( .A(n5143), .B(n5142), .Z(n5144) );
  NAND U5603 ( .A(n5145), .B(n5144), .Z(n5147) );
  XNOR U5604 ( .A(n6271), .B(n[209]), .Z(n5146) );
  NANDN U5605 ( .A(n5147), .B(n5146), .Z(n5148) );
  NAND U5606 ( .A(n5149), .B(n5148), .Z(n5150) );
  NANDN U5607 ( .A(n6278), .B(n5150), .Z(n5151) );
  NAND U5608 ( .A(n5152), .B(n5151), .Z(n5153) );
  NAND U5609 ( .A(n5154), .B(n5153), .Z(n5155) );
  NAND U5610 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U5611 ( .A(n5158), .B(n5157), .Z(n5159) );
  NAND U5612 ( .A(n5160), .B(n5159), .Z(n5161) );
  NAND U5613 ( .A(n5162), .B(n5161), .Z(n5163) );
  NAND U5614 ( .A(n5164), .B(n5163), .Z(n5165) );
  NAND U5615 ( .A(n5166), .B(n5165), .Z(n5167) );
  NAND U5616 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U5617 ( .A(n5170), .B(n5169), .Z(n5171) );
  NAND U5618 ( .A(n5172), .B(n5171), .Z(n5173) );
  AND U5619 ( .A(n5174), .B(n5173), .Z(n5180) );
  XNOR U5620 ( .A(n[217]), .B(n5175), .Z(n5176) );
  NANDN U5621 ( .A(n524), .B(n5176), .Z(n5177) );
  XNOR U5622 ( .A(n5178), .B(n5177), .Z(n6320) );
  NANDN U5623 ( .A(n5180), .B(n6320), .Z(n5179) );
  AND U5624 ( .A(n6326), .B(n5179), .Z(n5183) );
  XNOR U5625 ( .A(n6320), .B(n5180), .Z(n5181) );
  NAND U5626 ( .A(n[217]), .B(n5181), .Z(n5182) );
  NAND U5627 ( .A(n5183), .B(n5182), .Z(n5185) );
  OR U5628 ( .A(n6319), .B(n[218]), .Z(n5184) );
  AND U5629 ( .A(n5185), .B(n5184), .Z(n5186) );
  NAND U5630 ( .A(n5187), .B(n5186), .Z(n5188) );
  NAND U5631 ( .A(n5189), .B(n5188), .Z(n5190) );
  NAND U5632 ( .A(n5191), .B(n5190), .Z(n5192) );
  NAND U5633 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U5634 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U5635 ( .A(n5197), .B(n5196), .Z(n5198) );
  NAND U5636 ( .A(n5199), .B(n5198), .Z(n5200) );
  NAND U5637 ( .A(n5201), .B(n5200), .Z(n5202) );
  NAND U5638 ( .A(n5203), .B(n5202), .Z(n5204) );
  NAND U5639 ( .A(n5205), .B(n5204), .Z(n5206) );
  NAND U5640 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U5641 ( .A(n5209), .B(n5208), .Z(n5210) );
  NAND U5642 ( .A(n5211), .B(n5210), .Z(n5212) );
  NAND U5643 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5644 ( .A(n5215), .B(n5214), .Z(n5216) );
  NAND U5645 ( .A(n5217), .B(n5216), .Z(n5218) );
  NAND U5646 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U5647 ( .A(n5221), .B(n5220), .Z(n5222) );
  NAND U5648 ( .A(n5223), .B(n5222), .Z(n5224) );
  NAND U5649 ( .A(n5225), .B(n5224), .Z(n5226) );
  NAND U5650 ( .A(n5227), .B(n5226), .Z(n5228) );
  AND U5651 ( .A(n5229), .B(n5228), .Z(n5234) );
  XNOR U5652 ( .A(n[230]), .B(n5230), .Z(n5231) );
  NANDN U5653 ( .A(n524), .B(n5231), .Z(n5232) );
  XNOR U5654 ( .A(n5233), .B(n5232), .Z(n6416) );
  NANDN U5655 ( .A(n5234), .B(n6416), .Z(n5237) );
  XNOR U5656 ( .A(n6416), .B(n5234), .Z(n5235) );
  NAND U5657 ( .A(n[230]), .B(n5235), .Z(n5236) );
  NAND U5658 ( .A(n5237), .B(n5236), .Z(n5238) );
  AND U5659 ( .A(n5239), .B(n5238), .Z(n5240) );
  ANDN U5660 ( .B(n6415), .A(n6413), .Z(n6422) );
  OR U5661 ( .A(n5240), .B(n6422), .Z(n5241) );
  NAND U5662 ( .A(n5242), .B(n5241), .Z(n5243) );
  NAND U5663 ( .A(n5244), .B(n5243), .Z(n5245) );
  NAND U5664 ( .A(n5246), .B(n5245), .Z(n5247) );
  NAND U5665 ( .A(n5248), .B(n5247), .Z(n5249) );
  NAND U5666 ( .A(n5250), .B(n5249), .Z(n5251) );
  NAND U5667 ( .A(n5252), .B(n5251), .Z(n5253) );
  NAND U5668 ( .A(n5254), .B(n5253), .Z(n5255) );
  AND U5669 ( .A(n5256), .B(n5255), .Z(n5264) );
  NANDN U5670 ( .A(n6450), .B(n5264), .Z(n5262) );
  XOR U5671 ( .A(n6456), .B(n5257), .Z(n5258) );
  NANDN U5672 ( .A(n524), .B(n5258), .Z(n5259) );
  XOR U5673 ( .A(n5260), .B(n5259), .Z(n6457) );
  ANDN U5674 ( .B(n6457), .A(n[237]), .Z(n5261) );
  ANDN U5675 ( .B(n5262), .A(n5261), .Z(n5267) );
  XOR U5676 ( .A(n5264), .B(n5263), .Z(n5265) );
  NANDN U5677 ( .A(n[236]), .B(n5265), .Z(n5266) );
  NAND U5678 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U5679 ( .A(n5268), .B(n6459), .Z(n5269) );
  NAND U5680 ( .A(n5270), .B(n5269), .Z(n5271) );
  NAND U5681 ( .A(n5272), .B(n5271), .Z(n5273) );
  NAND U5682 ( .A(n5274), .B(n5273), .Z(n5275) );
  NAND U5683 ( .A(n5276), .B(n5275), .Z(n5277) );
  NAND U5684 ( .A(n5278), .B(n5277), .Z(n5279) );
  NAND U5685 ( .A(n5280), .B(n5279), .Z(n5281) );
  NAND U5686 ( .A(n5282), .B(n5281), .Z(n5283) );
  NAND U5687 ( .A(n5284), .B(n5283), .Z(n5285) );
  NAND U5688 ( .A(n5286), .B(n5285), .Z(n5287) );
  NAND U5689 ( .A(n5288), .B(n5287), .Z(n5289) );
  NAND U5690 ( .A(n5290), .B(n5289), .Z(n5291) );
  NAND U5691 ( .A(n5292), .B(n5291), .Z(n5293) );
  NAND U5692 ( .A(n5294), .B(n5293), .Z(n5295) );
  NAND U5693 ( .A(n5296), .B(n5295), .Z(n5297) );
  NAND U5694 ( .A(n5298), .B(n5297), .Z(n5299) );
  NAND U5695 ( .A(n5300), .B(n5299), .Z(n5301) );
  NAND U5696 ( .A(n5302), .B(n5301), .Z(n5303) );
  NAND U5697 ( .A(n5304), .B(n5303), .Z(n5305) );
  NAND U5698 ( .A(n5306), .B(n5305), .Z(n5307) );
  NAND U5699 ( .A(n5308), .B(n5307), .Z(n5309) );
  NAND U5700 ( .A(n5310), .B(n5309), .Z(n5311) );
  NAND U5701 ( .A(n5312), .B(n5311), .Z(n5313) );
  NAND U5702 ( .A(n5314), .B(n5313), .Z(n5315) );
  NAND U5703 ( .A(n5316), .B(n5315), .Z(n5317) );
  NAND U5704 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U5705 ( .A(n5320), .B(n5319), .Z(n5321) );
  NAND U5706 ( .A(n5322), .B(n5321), .Z(n5323) );
  NAND U5707 ( .A(n5324), .B(n5323), .Z(n5325) );
  NAND U5708 ( .A(n5326), .B(n5325), .Z(n5327) );
  NAND U5709 ( .A(n5328), .B(n5327), .Z(n5329) );
  NAND U5710 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5711 ( .A(n5332), .B(n5331), .Z(n5333) );
  NAND U5712 ( .A(n5334), .B(n5333), .Z(n5335) );
  NAND U5713 ( .A(n5336), .B(n5335), .Z(n5338) );
  XOR U5714 ( .A(n[255]), .B(n6580), .Z(n5337) );
  NANDN U5715 ( .A(n5338), .B(n5337), .Z(n5339) );
  NAND U5716 ( .A(n5340), .B(n5339), .Z(n6814) );
  ANDN U5717 ( .B(n[0]), .A(n525), .Z(n5341) );
  XOR U5718 ( .A(n5342), .B(n5341), .Z(zout[0]) );
  NANDN U5719 ( .A(n525), .B(n[100]), .Z(n5343) );
  XOR U5720 ( .A(n5544), .B(n5343), .Z(n5547) );
  NANDN U5721 ( .A(n5344), .B(n6814), .Z(n5541) );
  AND U5722 ( .A(n5347), .B(n[98]), .Z(n5345) );
  NANDN U5723 ( .A(n525), .B(n5345), .Z(n5539) );
  NANDN U5724 ( .A(n525), .B(n[98]), .Z(n5346) );
  XOR U5725 ( .A(n5347), .B(n5346), .Z(n6863) );
  AND U5726 ( .A(n6814), .B(n[96]), .Z(n5534) );
  OR U5727 ( .A(n5534), .B(n5535), .Z(n5537) );
  ANDN U5728 ( .B(n5531), .A(n5529), .Z(n5348) );
  NANDN U5729 ( .A(n525), .B(n5348), .Z(n5533) );
  NANDN U5730 ( .A(n525), .B(n[94]), .Z(n5349) );
  NANDN U5731 ( .A(n5349), .B(n5350), .Z(n5528) );
  XOR U5732 ( .A(n5350), .B(n5349), .Z(n6854) );
  NANDN U5733 ( .A(n525), .B(n[93]), .Z(n5351) );
  NANDN U5734 ( .A(n5351), .B(n5352), .Z(n5526) );
  XOR U5735 ( .A(n5352), .B(n5351), .Z(n6852) );
  ANDN U5736 ( .B(n5356), .A(n5353), .Z(n5354) );
  NANDN U5737 ( .A(n525), .B(n5354), .Z(n5524) );
  NANDN U5738 ( .A(n525), .B(n[92]), .Z(n5355) );
  XOR U5739 ( .A(n5356), .B(n5355), .Z(n6850) );
  AND U5740 ( .A(n5359), .B(n[91]), .Z(n5357) );
  NANDN U5741 ( .A(n525), .B(n5357), .Z(n5522) );
  NANDN U5742 ( .A(n525), .B(n[91]), .Z(n5358) );
  XOR U5743 ( .A(n5359), .B(n5358), .Z(n6848) );
  NANDN U5744 ( .A(n525), .B(n[90]), .Z(n5360) );
  NANDN U5745 ( .A(n5360), .B(n5361), .Z(n5520) );
  XOR U5746 ( .A(n5361), .B(n5360), .Z(n6846) );
  AND U5747 ( .A(n5364), .B(n[89]), .Z(n5362) );
  NANDN U5748 ( .A(n525), .B(n5362), .Z(n5518) );
  NANDN U5749 ( .A(n525), .B(n[89]), .Z(n5363) );
  XOR U5750 ( .A(n5364), .B(n5363), .Z(n6834) );
  NANDN U5751 ( .A(n525), .B(n[87]), .Z(n5365) );
  NANDN U5752 ( .A(n5365), .B(n5366), .Z(n5512) );
  XOR U5753 ( .A(n5366), .B(n5365), .Z(n6830) );
  NANDN U5754 ( .A(n525), .B(n[86]), .Z(n5367) );
  NANDN U5755 ( .A(n5367), .B(n5368), .Z(n5510) );
  XOR U5756 ( .A(n5368), .B(n5367), .Z(n6828) );
  NANDN U5757 ( .A(n525), .B(n[84]), .Z(n5369) );
  NANDN U5758 ( .A(n5369), .B(n5370), .Z(n5503) );
  XOR U5759 ( .A(n5370), .B(n5369), .Z(n6824) );
  NANDN U5760 ( .A(n525), .B(n[83]), .Z(n5371) );
  NANDN U5761 ( .A(n5371), .B(n5372), .Z(n5501) );
  XOR U5762 ( .A(n5372), .B(n5371), .Z(n6822) );
  AND U5763 ( .A(n5375), .B(n[82]), .Z(n5373) );
  NANDN U5764 ( .A(n525), .B(n5373), .Z(n5499) );
  NANDN U5765 ( .A(n525), .B(n[82]), .Z(n5374) );
  XOR U5766 ( .A(n5375), .B(n5374), .Z(n6820) );
  NANDN U5767 ( .A(n525), .B(n[81]), .Z(n5376) );
  NANDN U5768 ( .A(n5376), .B(n5377), .Z(n5497) );
  XOR U5769 ( .A(n5377), .B(n5376), .Z(n6818) );
  NANDN U5770 ( .A(n525), .B(n[80]), .Z(n5378) );
  NANDN U5771 ( .A(n5378), .B(n5379), .Z(n5495) );
  XOR U5772 ( .A(n5379), .B(n5378), .Z(n6815) );
  NANDN U5773 ( .A(n525), .B(n[78]), .Z(n5380) );
  NANDN U5774 ( .A(n5380), .B(n5381), .Z(n5493) );
  XOR U5775 ( .A(n5381), .B(n5380), .Z(n6808) );
  NANDN U5776 ( .A(n525), .B(n[76]), .Z(n5382) );
  NANDN U5777 ( .A(n5382), .B(n5383), .Z(n5491) );
  XOR U5778 ( .A(n5383), .B(n5382), .Z(n6802) );
  AND U5779 ( .A(n5386), .B(n[74]), .Z(n5384) );
  NANDN U5780 ( .A(n525), .B(n5384), .Z(n5485) );
  NANDN U5781 ( .A(n525), .B(n[74]), .Z(n5385) );
  XOR U5782 ( .A(n5386), .B(n5385), .Z(n6798) );
  NANDN U5783 ( .A(n525), .B(n[73]), .Z(n5387) );
  NANDN U5784 ( .A(n5387), .B(n5388), .Z(n5483) );
  XOR U5785 ( .A(n5388), .B(n5387), .Z(n6796) );
  AND U5786 ( .A(n5479), .B(n[72]), .Z(n5389) );
  NANDN U5787 ( .A(n525), .B(n5389), .Z(n5481) );
  NANDN U5788 ( .A(n5390), .B(n6814), .Z(n5474) );
  AND U5789 ( .A(n5475), .B(n5474), .Z(n5477) );
  ANDN U5790 ( .B(n5471), .A(n5469), .Z(n5391) );
  NANDN U5791 ( .A(n525), .B(n5391), .Z(n5473) );
  NANDN U5792 ( .A(n525), .B(n[69]), .Z(n5392) );
  NANDN U5793 ( .A(n5392), .B(n5393), .Z(n5468) );
  XOR U5794 ( .A(n5393), .B(n5392), .Z(n6777) );
  AND U5795 ( .A(n5396), .B(n[67]), .Z(n5394) );
  NANDN U5796 ( .A(n525), .B(n5394), .Z(n5466) );
  NANDN U5797 ( .A(n525), .B(n[67]), .Z(n5395) );
  XOR U5798 ( .A(n5396), .B(n5395), .Z(n6771) );
  NANDN U5799 ( .A(n525), .B(n[65]), .Z(n5397) );
  NANDN U5800 ( .A(n5397), .B(n5398), .Z(n5464) );
  XOR U5801 ( .A(n5398), .B(n5397), .Z(n6766) );
  ANDN U5802 ( .B(n5402), .A(n5399), .Z(n5400) );
  NANDN U5803 ( .A(n525), .B(n5400), .Z(n5462) );
  NANDN U5804 ( .A(n525), .B(n[64]), .Z(n5401) );
  XOR U5805 ( .A(n5402), .B(n5401), .Z(n6764) );
  NANDN U5806 ( .A(n525), .B(n[62]), .Z(n5403) );
  NANDN U5807 ( .A(n5403), .B(n5404), .Z(n5456) );
  XOR U5808 ( .A(n5404), .B(n5403), .Z(n6760) );
  NANDN U5809 ( .A(n525), .B(n[61]), .Z(n5405) );
  NANDN U5810 ( .A(n5405), .B(n5406), .Z(n5454) );
  XOR U5811 ( .A(n5406), .B(n5405), .Z(n6758) );
  NANDN U5812 ( .A(n525), .B(n[60]), .Z(n5407) );
  NANDN U5813 ( .A(n5407), .B(n5408), .Z(n5452) );
  XOR U5814 ( .A(n5408), .B(n5407), .Z(n6756) );
  NANDN U5815 ( .A(n525), .B(n[59]), .Z(n5409) );
  NANDN U5816 ( .A(n5409), .B(n5410), .Z(n5450) );
  XOR U5817 ( .A(n5410), .B(n5409), .Z(n6753) );
  ANDN U5818 ( .B(n5414), .A(n5411), .Z(n5412) );
  NANDN U5819 ( .A(n525), .B(n5412), .Z(n5448) );
  NANDN U5820 ( .A(n525), .B(n[58]), .Z(n5413) );
  XOR U5821 ( .A(n5414), .B(n5413), .Z(n6751) );
  AND U5822 ( .A(n5417), .B(n[57]), .Z(n5415) );
  NANDN U5823 ( .A(n525), .B(n5415), .Z(n5446) );
  NANDN U5824 ( .A(n525), .B(n[57]), .Z(n5416) );
  XOR U5825 ( .A(n5417), .B(n5416), .Z(n6749) );
  NANDN U5826 ( .A(n525), .B(n[56]), .Z(n5418) );
  NANDN U5827 ( .A(n5418), .B(n5419), .Z(n5444) );
  XOR U5828 ( .A(n5419), .B(n5418), .Z(n6747) );
  NANDN U5829 ( .A(n525), .B(n[55]), .Z(n5420) );
  NANDN U5830 ( .A(n5420), .B(n5421), .Z(n5442) );
  XOR U5831 ( .A(n5421), .B(n5420), .Z(n6745) );
  NANDN U5832 ( .A(n525), .B(n[54]), .Z(n5422) );
  NANDN U5833 ( .A(n5422), .B(n5423), .Z(n5440) );
  XOR U5834 ( .A(n5423), .B(n5422), .Z(n6742) );
  AND U5835 ( .A(n5426), .B(n[52]), .Z(n5424) );
  NANDN U5836 ( .A(n525), .B(n5424), .Z(n5438) );
  NANDN U5837 ( .A(n525), .B(n[52]), .Z(n5425) );
  XOR U5838 ( .A(n5426), .B(n5425), .Z(n6737) );
  NANDN U5839 ( .A(n525), .B(n[51]), .Z(n5427) );
  NANDN U5840 ( .A(n5427), .B(n5428), .Z(n5436) );
  XOR U5841 ( .A(n5428), .B(n5427), .Z(n6734) );
  AND U5842 ( .A(n5432), .B(n[48]), .Z(n5429) );
  NANDN U5843 ( .A(n525), .B(n5429), .Z(n5434) );
  OR U5844 ( .A(n5430), .B(n525), .Z(n6721) );
  NANDN U5845 ( .A(n525), .B(n[48]), .Z(n5431) );
  XOR U5846 ( .A(n5432), .B(n5431), .Z(n6720) );
  OR U5847 ( .A(n6721), .B(n6720), .Z(n5433) );
  NAND U5848 ( .A(n5434), .B(n5433), .Z(n6725) );
  AND U5849 ( .A(n6814), .B(n[49]), .Z(n6722) );
  AND U5850 ( .A(n[50]), .B(n6814), .Z(n6733) );
  OR U5851 ( .A(n6734), .B(n6735), .Z(n5435) );
  AND U5852 ( .A(n5436), .B(n5435), .Z(n6736) );
  OR U5853 ( .A(n6737), .B(n6736), .Z(n5437) );
  AND U5854 ( .A(n5438), .B(n5437), .Z(n6738) );
  NANDN U5855 ( .A(n525), .B(n[53]), .Z(n6741) );
  NANDN U5856 ( .A(n6742), .B(n6743), .Z(n5439) );
  AND U5857 ( .A(n5440), .B(n5439), .Z(n6744) );
  OR U5858 ( .A(n6745), .B(n6744), .Z(n5441) );
  AND U5859 ( .A(n5442), .B(n5441), .Z(n6746) );
  OR U5860 ( .A(n6747), .B(n6746), .Z(n5443) );
  AND U5861 ( .A(n5444), .B(n5443), .Z(n6748) );
  OR U5862 ( .A(n6749), .B(n6748), .Z(n5445) );
  AND U5863 ( .A(n5446), .B(n5445), .Z(n6750) );
  OR U5864 ( .A(n6751), .B(n6750), .Z(n5447) );
  AND U5865 ( .A(n5448), .B(n5447), .Z(n6752) );
  OR U5866 ( .A(n6753), .B(n6752), .Z(n5449) );
  AND U5867 ( .A(n5450), .B(n5449), .Z(n6755) );
  OR U5868 ( .A(n6756), .B(n6755), .Z(n5451) );
  AND U5869 ( .A(n5452), .B(n5451), .Z(n6757) );
  OR U5870 ( .A(n6758), .B(n6757), .Z(n5453) );
  AND U5871 ( .A(n5454), .B(n5453), .Z(n6759) );
  OR U5872 ( .A(n6760), .B(n6759), .Z(n5455) );
  NAND U5873 ( .A(n5456), .B(n5455), .Z(n5457) );
  NAND U5874 ( .A(n5457), .B(n5458), .Z(n5460) );
  NANDN U5875 ( .A(n525), .B(n[63]), .Z(n6761) );
  XOR U5876 ( .A(n5458), .B(n5457), .Z(n6762) );
  NANDN U5877 ( .A(n6761), .B(n6762), .Z(n5459) );
  AND U5878 ( .A(n5460), .B(n5459), .Z(n6763) );
  OR U5879 ( .A(n6764), .B(n6763), .Z(n5461) );
  AND U5880 ( .A(n5462), .B(n5461), .Z(n6765) );
  OR U5881 ( .A(n6766), .B(n6765), .Z(n5463) );
  AND U5882 ( .A(n5464), .B(n5463), .Z(n6767) );
  NANDN U5883 ( .A(n525), .B(n[66]), .Z(n6770) );
  NANDN U5884 ( .A(n6771), .B(n6772), .Z(n5465) );
  AND U5885 ( .A(n5466), .B(n5465), .Z(n6773) );
  NANDN U5886 ( .A(n525), .B(n[68]), .Z(n6776) );
  NANDN U5887 ( .A(n6777), .B(n6778), .Z(n5467) );
  AND U5888 ( .A(n5468), .B(n5467), .Z(n6789) );
  NANDN U5889 ( .A(n5469), .B(n6814), .Z(n5470) );
  XNOR U5890 ( .A(n5471), .B(n5470), .Z(n6790) );
  NANDN U5891 ( .A(n6789), .B(n6790), .Z(n5472) );
  NAND U5892 ( .A(n5473), .B(n5472), .Z(n6791) );
  XOR U5893 ( .A(n5475), .B(n5474), .Z(n6792) );
  NANDN U5894 ( .A(n6791), .B(n6792), .Z(n5476) );
  NANDN U5895 ( .A(n5477), .B(n5476), .Z(n6794) );
  NANDN U5896 ( .A(n525), .B(n[72]), .Z(n5478) );
  XOR U5897 ( .A(n5479), .B(n5478), .Z(n6793) );
  OR U5898 ( .A(n6794), .B(n6793), .Z(n5480) );
  AND U5899 ( .A(n5481), .B(n5480), .Z(n6795) );
  OR U5900 ( .A(n6796), .B(n6795), .Z(n5482) );
  AND U5901 ( .A(n5483), .B(n5482), .Z(n6797) );
  OR U5902 ( .A(n6798), .B(n6797), .Z(n5484) );
  NAND U5903 ( .A(n5485), .B(n5484), .Z(n5486) );
  NAND U5904 ( .A(n5486), .B(n5487), .Z(n5489) );
  NANDN U5905 ( .A(n525), .B(n[75]), .Z(n6799) );
  XOR U5906 ( .A(n5487), .B(n5486), .Z(n6800) );
  NANDN U5907 ( .A(n6799), .B(n6800), .Z(n5488) );
  AND U5908 ( .A(n5489), .B(n5488), .Z(n6801) );
  OR U5909 ( .A(n6802), .B(n6801), .Z(n5490) );
  NAND U5910 ( .A(n5491), .B(n5490), .Z(n6806) );
  AND U5911 ( .A(n6814), .B(n[77]), .Z(n6803) );
  OR U5912 ( .A(n6808), .B(n6807), .Z(n5492) );
  NAND U5913 ( .A(n5493), .B(n5492), .Z(n6812) );
  AND U5914 ( .A(n[79]), .B(n6814), .Z(n6809) );
  OR U5915 ( .A(n6815), .B(n6816), .Z(n5494) );
  AND U5916 ( .A(n5495), .B(n5494), .Z(n6817) );
  OR U5917 ( .A(n6818), .B(n6817), .Z(n5496) );
  AND U5918 ( .A(n5497), .B(n5496), .Z(n6819) );
  OR U5919 ( .A(n6820), .B(n6819), .Z(n5498) );
  AND U5920 ( .A(n5499), .B(n5498), .Z(n6821) );
  OR U5921 ( .A(n6822), .B(n6821), .Z(n5500) );
  AND U5922 ( .A(n5501), .B(n5500), .Z(n6823) );
  OR U5923 ( .A(n6824), .B(n6823), .Z(n5502) );
  NAND U5924 ( .A(n5503), .B(n5502), .Z(n5505) );
  NAND U5925 ( .A(n5505), .B(n5506), .Z(n5508) );
  NANDN U5926 ( .A(n5504), .B(n6814), .Z(n6825) );
  XOR U5927 ( .A(n5506), .B(n5505), .Z(n6826) );
  NANDN U5928 ( .A(n6825), .B(n6826), .Z(n5507) );
  AND U5929 ( .A(n5508), .B(n5507), .Z(n6827) );
  OR U5930 ( .A(n6828), .B(n6827), .Z(n5509) );
  AND U5931 ( .A(n5510), .B(n5509), .Z(n6829) );
  OR U5932 ( .A(n6830), .B(n6829), .Z(n5511) );
  NAND U5933 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U5934 ( .A(n5513), .B(n5514), .Z(n5516) );
  NANDN U5935 ( .A(n525), .B(n[88]), .Z(n6831) );
  XOR U5936 ( .A(n5514), .B(n5513), .Z(n6832) );
  NANDN U5937 ( .A(n6831), .B(n6832), .Z(n5515) );
  AND U5938 ( .A(n5516), .B(n5515), .Z(n6833) );
  OR U5939 ( .A(n6834), .B(n6833), .Z(n5517) );
  AND U5940 ( .A(n5518), .B(n5517), .Z(n6845) );
  OR U5941 ( .A(n6846), .B(n6845), .Z(n5519) );
  AND U5942 ( .A(n5520), .B(n5519), .Z(n6847) );
  OR U5943 ( .A(n6848), .B(n6847), .Z(n5521) );
  AND U5944 ( .A(n5522), .B(n5521), .Z(n6849) );
  OR U5945 ( .A(n6850), .B(n6849), .Z(n5523) );
  AND U5946 ( .A(n5524), .B(n5523), .Z(n6851) );
  OR U5947 ( .A(n6852), .B(n6851), .Z(n5525) );
  AND U5948 ( .A(n5526), .B(n5525), .Z(n6853) );
  OR U5949 ( .A(n6854), .B(n6853), .Z(n5527) );
  AND U5950 ( .A(n5528), .B(n5527), .Z(n6855) );
  NANDN U5951 ( .A(n5529), .B(n6814), .Z(n5530) );
  XNOR U5952 ( .A(n5531), .B(n5530), .Z(n6856) );
  NANDN U5953 ( .A(n6855), .B(n6856), .Z(n5532) );
  NAND U5954 ( .A(n5533), .B(n5532), .Z(n6858) );
  XOR U5955 ( .A(n5535), .B(n5534), .Z(n6857) );
  NANDN U5956 ( .A(n6858), .B(n6857), .Z(n5536) );
  NAND U5957 ( .A(n5537), .B(n5536), .Z(n6859) );
  NANDN U5958 ( .A(n525), .B(n[97]), .Z(n6862) );
  NANDN U5959 ( .A(n6863), .B(n6864), .Z(n5538) );
  AND U5960 ( .A(n5539), .B(n5538), .Z(n5540) );
  OR U5961 ( .A(n5541), .B(n5540), .Z(n5543) );
  XNOR U5962 ( .A(n5541), .B(n5540), .Z(n6865) );
  NANDN U5963 ( .A(n6865), .B(n6866), .Z(n5542) );
  AND U5964 ( .A(n5543), .B(n5542), .Z(n5546) );
  XNOR U5965 ( .A(n5547), .B(n5546), .Z(zout[100]) );
  AND U5966 ( .A(n5544), .B(n[100]), .Z(n5545) );
  NANDN U5967 ( .A(n525), .B(n5545), .Z(n5549) );
  OR U5968 ( .A(n5547), .B(n5546), .Z(n5548) );
  NAND U5969 ( .A(n5549), .B(n5548), .Z(n5552) );
  AND U5970 ( .A(n6814), .B(n[101]), .Z(n5553) );
  XOR U5971 ( .A(n5551), .B(n5553), .Z(n5550) );
  XNOR U5972 ( .A(n5552), .B(n5550), .Z(zout[101]) );
  NANDN U5973 ( .A(n525), .B(n[102]), .Z(n5555) );
  XOR U5974 ( .A(n5554), .B(n5555), .Z(n5557) );
  XNOR U5975 ( .A(n5556), .B(n5557), .Z(zout[102]) );
  NANDN U5976 ( .A(n5555), .B(n5554), .Z(n5559) );
  OR U5977 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U5978 ( .A(n5559), .B(n5558), .Z(n5560) );
  XOR U5979 ( .A(n5561), .B(n5560), .Z(n5562) );
  AND U5980 ( .A(n6814), .B(n[103]), .Z(n5563) );
  XNOR U5981 ( .A(n5562), .B(n5563), .Z(zout[103]) );
  NANDN U5982 ( .A(n525), .B(n[104]), .Z(n5569) );
  OR U5983 ( .A(n5561), .B(n5560), .Z(n5565) );
  NANDN U5984 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U5985 ( .A(n5565), .B(n5564), .Z(n5568) );
  XOR U5986 ( .A(n5567), .B(n5568), .Z(n5566) );
  XNOR U5987 ( .A(n5569), .B(n5566), .Z(zout[104]) );
  NANDN U5988 ( .A(n525), .B(n[105]), .Z(n5571) );
  XOR U5989 ( .A(n5570), .B(n5571), .Z(n5573) );
  XOR U5990 ( .A(n5572), .B(n5573), .Z(zout[105]) );
  NANDN U5991 ( .A(n5571), .B(n5570), .Z(n5575) );
  NANDN U5992 ( .A(n5573), .B(n5572), .Z(n5574) );
  NAND U5993 ( .A(n5575), .B(n5574), .Z(n5576) );
  XOR U5994 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U5995 ( .A(n[106]), .B(n6814), .Z(n5579) );
  XNOR U5996 ( .A(n5578), .B(n5579), .Z(zout[106]) );
  OR U5997 ( .A(n5577), .B(n5576), .Z(n5581) );
  NANDN U5998 ( .A(n5579), .B(n5578), .Z(n5580) );
  AND U5999 ( .A(n5581), .B(n5580), .Z(n5583) );
  XOR U6000 ( .A(n5582), .B(n5583), .Z(n5584) );
  NANDN U6001 ( .A(n525), .B(n[107]), .Z(n5585) );
  XOR U6002 ( .A(n5584), .B(n5585), .Z(zout[107]) );
  NANDN U6003 ( .A(n525), .B(n[108]), .Z(n5590) );
  XOR U6004 ( .A(n5589), .B(n5590), .Z(n5592) );
  NAND U6005 ( .A(n5583), .B(n5582), .Z(n5587) );
  NANDN U6006 ( .A(n5585), .B(n5584), .Z(n5586) );
  AND U6007 ( .A(n5587), .B(n5586), .Z(n5591) );
  XNOR U6008 ( .A(n5592), .B(n5591), .Z(zout[108]) );
  NANDN U6009 ( .A(n525), .B(n[109]), .Z(n5588) );
  XOR U6010 ( .A(n5599), .B(n5588), .Z(n5602) );
  NANDN U6011 ( .A(n5590), .B(n5589), .Z(n5594) );
  OR U6012 ( .A(n5592), .B(n5591), .Z(n5593) );
  AND U6013 ( .A(n5594), .B(n5593), .Z(n5601) );
  XNOR U6014 ( .A(n5602), .B(n5601), .Z(zout[109]) );
  XNOR U6015 ( .A(n[10]), .B(n5595), .Z(n5596) );
  NANDN U6016 ( .A(n525), .B(n5596), .Z(n5597) );
  XOR U6017 ( .A(n5598), .B(n5597), .Z(zout[10]) );
  NANDN U6018 ( .A(n525), .B(n[110]), .Z(n5606) );
  XOR U6019 ( .A(n5605), .B(n5606), .Z(n5608) );
  AND U6020 ( .A(n5599), .B(n[109]), .Z(n5600) );
  NANDN U6021 ( .A(n525), .B(n5600), .Z(n5604) );
  OR U6022 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U6023 ( .A(n5604), .B(n5603), .Z(n5607) );
  XNOR U6024 ( .A(n5608), .B(n5607), .Z(zout[110]) );
  NANDN U6025 ( .A(n5606), .B(n5605), .Z(n5610) );
  OR U6026 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U6027 ( .A(n5610), .B(n5609), .Z(n5613) );
  AND U6028 ( .A(n6814), .B(n[111]), .Z(n5614) );
  XOR U6029 ( .A(n5612), .B(n5614), .Z(n5611) );
  XNOR U6030 ( .A(n5613), .B(n5611), .Z(zout[111]) );
  NANDN U6031 ( .A(n525), .B(n[112]), .Z(n5618) );
  XNOR U6032 ( .A(n5616), .B(n5617), .Z(n5615) );
  XNOR U6033 ( .A(n5618), .B(n5615), .Z(zout[112]) );
  NANDN U6034 ( .A(n525), .B(n[113]), .Z(n5622) );
  XNOR U6035 ( .A(n5621), .B(n5620), .Z(n5619) );
  XNOR U6036 ( .A(n5622), .B(n5619), .Z(zout[113]) );
  NANDN U6037 ( .A(n525), .B(n[114]), .Z(n5626) );
  XNOR U6038 ( .A(n5625), .B(n5624), .Z(n5623) );
  XNOR U6039 ( .A(n5626), .B(n5623), .Z(zout[114]) );
  NANDN U6040 ( .A(n525), .B(n[115]), .Z(n5628) );
  XOR U6041 ( .A(n5627), .B(n5628), .Z(n5630) );
  XOR U6042 ( .A(n5629), .B(n5630), .Z(zout[115]) );
  NANDN U6043 ( .A(n5628), .B(n5627), .Z(n5632) );
  NANDN U6044 ( .A(n5630), .B(n5629), .Z(n5631) );
  NAND U6045 ( .A(n5632), .B(n5631), .Z(n5635) );
  XOR U6046 ( .A(n5634), .B(n5635), .Z(n5636) );
  NANDN U6047 ( .A(n5633), .B(n6814), .Z(n5637) );
  XOR U6048 ( .A(n5636), .B(n5637), .Z(zout[116]) );
  NANDN U6049 ( .A(n525), .B(n[117]), .Z(n5642) );
  XOR U6050 ( .A(n5641), .B(n5642), .Z(n5644) );
  NAND U6051 ( .A(n5635), .B(n5634), .Z(n5639) );
  NANDN U6052 ( .A(n5637), .B(n5636), .Z(n5638) );
  AND U6053 ( .A(n5639), .B(n5638), .Z(n5643) );
  XNOR U6054 ( .A(n5644), .B(n5643), .Z(zout[117]) );
  NANDN U6055 ( .A(n5648), .B(n6814), .Z(n5640) );
  XOR U6056 ( .A(n5649), .B(n5640), .Z(n5652) );
  NANDN U6057 ( .A(n5642), .B(n5641), .Z(n5646) );
  OR U6058 ( .A(n5644), .B(n5643), .Z(n5645) );
  AND U6059 ( .A(n5646), .B(n5645), .Z(n5651) );
  XNOR U6060 ( .A(n5652), .B(n5651), .Z(zout[118]) );
  NANDN U6061 ( .A(n525), .B(n[119]), .Z(n5647) );
  XOR U6062 ( .A(n5659), .B(n5647), .Z(n5662) );
  ANDN U6063 ( .B(n5649), .A(n5648), .Z(n5650) );
  NANDN U6064 ( .A(n525), .B(n5650), .Z(n5654) );
  OR U6065 ( .A(n5652), .B(n5651), .Z(n5653) );
  AND U6066 ( .A(n5654), .B(n5653), .Z(n5661) );
  XNOR U6067 ( .A(n5662), .B(n5661), .Z(zout[119]) );
  XOR U6068 ( .A(n[11]), .B(n5655), .Z(n5656) );
  ANDN U6069 ( .B(n5656), .A(n525), .Z(n5657) );
  XNOR U6070 ( .A(n5658), .B(n5657), .Z(zout[11]) );
  AND U6071 ( .A(n5659), .B(n[119]), .Z(n5660) );
  NANDN U6072 ( .A(n525), .B(n5660), .Z(n5664) );
  OR U6073 ( .A(n5662), .B(n5661), .Z(n5663) );
  NAND U6074 ( .A(n5664), .B(n5663), .Z(n5667) );
  AND U6075 ( .A(n6814), .B(n[120]), .Z(n5668) );
  XOR U6076 ( .A(n5666), .B(n5668), .Z(n5665) );
  XNOR U6077 ( .A(n5667), .B(n5665), .Z(zout[120]) );
  NANDN U6078 ( .A(n525), .B(n[121]), .Z(n5670) );
  XOR U6079 ( .A(n5669), .B(n5670), .Z(n5672) );
  XNOR U6080 ( .A(n5671), .B(n5672), .Z(zout[121]) );
  NANDN U6081 ( .A(n525), .B(n[122]), .Z(n5676) );
  XOR U6082 ( .A(n5675), .B(n5676), .Z(n5678) );
  NANDN U6083 ( .A(n5670), .B(n5669), .Z(n5674) );
  OR U6084 ( .A(n5672), .B(n5671), .Z(n5673) );
  AND U6085 ( .A(n5674), .B(n5673), .Z(n5677) );
  XNOR U6086 ( .A(n5678), .B(n5677), .Z(zout[122]) );
  NANDN U6087 ( .A(n525), .B(n[123]), .Z(n5682) );
  XOR U6088 ( .A(n5681), .B(n5682), .Z(n5684) );
  NANDN U6089 ( .A(n5676), .B(n5675), .Z(n5680) );
  OR U6090 ( .A(n5678), .B(n5677), .Z(n5679) );
  AND U6091 ( .A(n5680), .B(n5679), .Z(n5683) );
  XNOR U6092 ( .A(n5684), .B(n5683), .Z(zout[123]) );
  NANDN U6093 ( .A(n525), .B(n[124]), .Z(n5688) );
  XOR U6094 ( .A(n5687), .B(n5688), .Z(n5690) );
  NANDN U6095 ( .A(n5682), .B(n5681), .Z(n5686) );
  OR U6096 ( .A(n5684), .B(n5683), .Z(n5685) );
  AND U6097 ( .A(n5686), .B(n5685), .Z(n5689) );
  XNOR U6098 ( .A(n5690), .B(n5689), .Z(zout[124]) );
  NANDN U6099 ( .A(n525), .B(n[125]), .Z(n5696) );
  NANDN U6100 ( .A(n5688), .B(n5687), .Z(n5692) );
  OR U6101 ( .A(n5690), .B(n5689), .Z(n5691) );
  AND U6102 ( .A(n5692), .B(n5691), .Z(n5695) );
  XOR U6103 ( .A(n5694), .B(n5695), .Z(n5693) );
  XNOR U6104 ( .A(n5696), .B(n5693), .Z(zout[125]) );
  NANDN U6105 ( .A(n525), .B(n[126]), .Z(n5698) );
  XOR U6106 ( .A(n5697), .B(n5698), .Z(n5700) );
  XOR U6107 ( .A(n5699), .B(n5700), .Z(zout[126]) );
  NANDN U6108 ( .A(n525), .B(n[127]), .Z(n5705) );
  XOR U6109 ( .A(n5704), .B(n5705), .Z(n5707) );
  NANDN U6110 ( .A(n5698), .B(n5697), .Z(n5702) );
  NANDN U6111 ( .A(n5700), .B(n5699), .Z(n5701) );
  AND U6112 ( .A(n5702), .B(n5701), .Z(n5706) );
  XNOR U6113 ( .A(n5707), .B(n5706), .Z(zout[127]) );
  NANDN U6114 ( .A(n525), .B(n[128]), .Z(n5703) );
  XOR U6115 ( .A(n5710), .B(n5703), .Z(n5713) );
  NANDN U6116 ( .A(n5705), .B(n5704), .Z(n5709) );
  OR U6117 ( .A(n5707), .B(n5706), .Z(n5708) );
  AND U6118 ( .A(n5709), .B(n5708), .Z(n5712) );
  XNOR U6119 ( .A(n5713), .B(n5712), .Z(zout[128]) );
  NANDN U6120 ( .A(n525), .B(n[129]), .Z(n5721) );
  XOR U6121 ( .A(n5720), .B(n5721), .Z(n5723) );
  AND U6122 ( .A(n5710), .B(n[128]), .Z(n5711) );
  NANDN U6123 ( .A(n525), .B(n5711), .Z(n5715) );
  OR U6124 ( .A(n5713), .B(n5712), .Z(n5714) );
  AND U6125 ( .A(n5715), .B(n5714), .Z(n5722) );
  XNOR U6126 ( .A(n5723), .B(n5722), .Z(zout[129]) );
  XOR U6127 ( .A(n[12]), .B(n5716), .Z(n5717) );
  NANDN U6128 ( .A(n525), .B(n5717), .Z(n5718) );
  XOR U6129 ( .A(n5719), .B(n5718), .Z(zout[12]) );
  NANDN U6130 ( .A(n525), .B(n[130]), .Z(n5728) );
  XOR U6131 ( .A(n5727), .B(n5728), .Z(n5730) );
  NANDN U6132 ( .A(n5721), .B(n5720), .Z(n5725) );
  OR U6133 ( .A(n5723), .B(n5722), .Z(n5724) );
  AND U6134 ( .A(n5725), .B(n5724), .Z(n5729) );
  XNOR U6135 ( .A(n5730), .B(n5729), .Z(zout[130]) );
  NANDN U6136 ( .A(n525), .B(n[131]), .Z(n5726) );
  XOR U6137 ( .A(n5733), .B(n5726), .Z(n5736) );
  NANDN U6138 ( .A(n5728), .B(n5727), .Z(n5732) );
  OR U6139 ( .A(n5730), .B(n5729), .Z(n5731) );
  AND U6140 ( .A(n5732), .B(n5731), .Z(n5735) );
  XNOR U6141 ( .A(n5736), .B(n5735), .Z(zout[131]) );
  NANDN U6142 ( .A(n525), .B(n[132]), .Z(n5740) );
  XOR U6143 ( .A(n5739), .B(n5740), .Z(n5742) );
  AND U6144 ( .A(n5733), .B(n[131]), .Z(n5734) );
  NANDN U6145 ( .A(n525), .B(n5734), .Z(n5738) );
  OR U6146 ( .A(n5736), .B(n5735), .Z(n5737) );
  AND U6147 ( .A(n5738), .B(n5737), .Z(n5741) );
  XNOR U6148 ( .A(n5742), .B(n5741), .Z(zout[132]) );
  NANDN U6149 ( .A(n525), .B(n[133]), .Z(n5747) );
  XOR U6150 ( .A(n5746), .B(n5747), .Z(n5749) );
  NANDN U6151 ( .A(n5740), .B(n5739), .Z(n5744) );
  OR U6152 ( .A(n5742), .B(n5741), .Z(n5743) );
  AND U6153 ( .A(n5744), .B(n5743), .Z(n5748) );
  XNOR U6154 ( .A(n5749), .B(n5748), .Z(zout[133]) );
  NANDN U6155 ( .A(n525), .B(n[134]), .Z(n5745) );
  XOR U6156 ( .A(n5752), .B(n5745), .Z(n5755) );
  NANDN U6157 ( .A(n5747), .B(n5746), .Z(n5751) );
  OR U6158 ( .A(n5749), .B(n5748), .Z(n5750) );
  AND U6159 ( .A(n5751), .B(n5750), .Z(n5754) );
  XNOR U6160 ( .A(n5755), .B(n5754), .Z(zout[134]) );
  NANDN U6161 ( .A(n525), .B(n[135]), .Z(n5759) );
  XOR U6162 ( .A(n5758), .B(n5759), .Z(n5761) );
  AND U6163 ( .A(n5752), .B(n[134]), .Z(n5753) );
  NANDN U6164 ( .A(n525), .B(n5753), .Z(n5757) );
  OR U6165 ( .A(n5755), .B(n5754), .Z(n5756) );
  AND U6166 ( .A(n5757), .B(n5756), .Z(n5760) );
  XNOR U6167 ( .A(n5761), .B(n5760), .Z(zout[135]) );
  NANDN U6168 ( .A(n525), .B(n[136]), .Z(n5765) );
  XOR U6169 ( .A(n5764), .B(n5765), .Z(n5767) );
  NANDN U6170 ( .A(n5759), .B(n5758), .Z(n5763) );
  OR U6171 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U6172 ( .A(n5763), .B(n5762), .Z(n5766) );
  XNOR U6173 ( .A(n5767), .B(n5766), .Z(zout[136]) );
  NANDN U6174 ( .A(n525), .B(n[137]), .Z(n5771) );
  XOR U6175 ( .A(n5770), .B(n5771), .Z(n5773) );
  NANDN U6176 ( .A(n5765), .B(n5764), .Z(n5769) );
  OR U6177 ( .A(n5767), .B(n5766), .Z(n5768) );
  AND U6178 ( .A(n5769), .B(n5768), .Z(n5772) );
  XNOR U6179 ( .A(n5773), .B(n5772), .Z(zout[137]) );
  NANDN U6180 ( .A(n5771), .B(n5770), .Z(n5775) );
  OR U6181 ( .A(n5773), .B(n5772), .Z(n5774) );
  NAND U6182 ( .A(n5775), .B(n5774), .Z(n5777) );
  XOR U6183 ( .A(n5776), .B(n5777), .Z(n5778) );
  NANDN U6184 ( .A(n525), .B(n[138]), .Z(n5779) );
  XOR U6185 ( .A(n5778), .B(n5779), .Z(zout[138]) );
  NAND U6186 ( .A(n5777), .B(n5776), .Z(n5781) );
  NANDN U6187 ( .A(n5779), .B(n5778), .Z(n5780) );
  NAND U6188 ( .A(n5781), .B(n5780), .Z(n5784) );
  XOR U6189 ( .A(n5783), .B(n5784), .Z(n5785) );
  NANDN U6190 ( .A(n525), .B(n[139]), .Z(n5786) );
  XOR U6191 ( .A(n5785), .B(n5786), .Z(zout[139]) );
  AND U6192 ( .A(n6814), .B(n[13]), .Z(n5847) );
  XNOR U6193 ( .A(n5846), .B(n5847), .Z(n5844) );
  NOR U6194 ( .A(n525), .B(n5782), .Z(n5845) );
  XOR U6195 ( .A(n5844), .B(n5845), .Z(zout[13]) );
  NANDN U6196 ( .A(n525), .B(n[140]), .Z(n5790) );
  XOR U6197 ( .A(n5789), .B(n5790), .Z(n5792) );
  NAND U6198 ( .A(n5784), .B(n5783), .Z(n5788) );
  NANDN U6199 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U6200 ( .A(n5788), .B(n5787), .Z(n5791) );
  XNOR U6201 ( .A(n5792), .B(n5791), .Z(zout[140]) );
  AND U6202 ( .A(n[141]), .B(n6814), .Z(n5798) );
  NANDN U6203 ( .A(n5790), .B(n5789), .Z(n5794) );
  OR U6204 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6205 ( .A(n5794), .B(n5793), .Z(n5797) );
  XNOR U6206 ( .A(n5796), .B(n5797), .Z(n5795) );
  XOR U6207 ( .A(n5798), .B(n5795), .Z(zout[141]) );
  NANDN U6208 ( .A(n525), .B(n[142]), .Z(n5799) );
  XOR U6209 ( .A(n5800), .B(n5799), .Z(n5802) );
  XNOR U6210 ( .A(n5803), .B(n5802), .Z(zout[142]) );
  AND U6211 ( .A(n5800), .B(n[142]), .Z(n5801) );
  NANDN U6212 ( .A(n525), .B(n5801), .Z(n5805) );
  OR U6213 ( .A(n5803), .B(n5802), .Z(n5804) );
  NAND U6214 ( .A(n5805), .B(n5804), .Z(n5807) );
  XOR U6215 ( .A(n5806), .B(n5807), .Z(n5808) );
  NANDN U6216 ( .A(n525), .B(n[143]), .Z(n5809) );
  XOR U6217 ( .A(n5808), .B(n5809), .Z(zout[143]) );
  NANDN U6218 ( .A(n525), .B(n[144]), .Z(n5814) );
  XOR U6219 ( .A(n5813), .B(n5814), .Z(n5816) );
  NAND U6220 ( .A(n5807), .B(n5806), .Z(n5811) );
  NANDN U6221 ( .A(n5809), .B(n5808), .Z(n5810) );
  AND U6222 ( .A(n5811), .B(n5810), .Z(n5815) );
  XNOR U6223 ( .A(n5816), .B(n5815), .Z(zout[144]) );
  NANDN U6224 ( .A(n525), .B(n[145]), .Z(n5812) );
  XOR U6225 ( .A(n5820), .B(n5812), .Z(n5823) );
  NANDN U6226 ( .A(n5814), .B(n5813), .Z(n5818) );
  OR U6227 ( .A(n5816), .B(n5815), .Z(n5817) );
  AND U6228 ( .A(n5818), .B(n5817), .Z(n5822) );
  XNOR U6229 ( .A(n5823), .B(n5822), .Z(zout[145]) );
  NANDN U6230 ( .A(n525), .B(n[146]), .Z(n5819) );
  XOR U6231 ( .A(n5826), .B(n5819), .Z(n5829) );
  AND U6232 ( .A(n5820), .B(n[145]), .Z(n5821) );
  NANDN U6233 ( .A(n525), .B(n5821), .Z(n5825) );
  OR U6234 ( .A(n5823), .B(n5822), .Z(n5824) );
  AND U6235 ( .A(n5825), .B(n5824), .Z(n5828) );
  XNOR U6236 ( .A(n5829), .B(n5828), .Z(zout[146]) );
  NANDN U6237 ( .A(n525), .B(n[147]), .Z(n5833) );
  XOR U6238 ( .A(n5832), .B(n5833), .Z(n5835) );
  AND U6239 ( .A(n5826), .B(n[146]), .Z(n5827) );
  NANDN U6240 ( .A(n525), .B(n5827), .Z(n5831) );
  OR U6241 ( .A(n5829), .B(n5828), .Z(n5830) );
  AND U6242 ( .A(n5831), .B(n5830), .Z(n5834) );
  XNOR U6243 ( .A(n5835), .B(n5834), .Z(zout[147]) );
  NANDN U6244 ( .A(n525), .B(n[148]), .Z(n5839) );
  XOR U6245 ( .A(n5838), .B(n5839), .Z(n5841) );
  NANDN U6246 ( .A(n5833), .B(n5832), .Z(n5837) );
  OR U6247 ( .A(n5835), .B(n5834), .Z(n5836) );
  AND U6248 ( .A(n5837), .B(n5836), .Z(n5840) );
  XNOR U6249 ( .A(n5841), .B(n5840), .Z(zout[148]) );
  NANDN U6250 ( .A(n525), .B(n[149]), .Z(n5855) );
  XOR U6251 ( .A(n5854), .B(n5855), .Z(n5857) );
  NANDN U6252 ( .A(n5839), .B(n5838), .Z(n5843) );
  OR U6253 ( .A(n5841), .B(n5840), .Z(n5842) );
  AND U6254 ( .A(n5843), .B(n5842), .Z(n5856) );
  XNOR U6255 ( .A(n5857), .B(n5856), .Z(zout[149]) );
  OR U6256 ( .A(n5845), .B(n5844), .Z(n5849) );
  OR U6257 ( .A(n5847), .B(n5846), .Z(n5848) );
  AND U6258 ( .A(n5849), .B(n5848), .Z(n5851) );
  NANDN U6259 ( .A(n525), .B(n[14]), .Z(n5850) );
  XNOR U6260 ( .A(n5851), .B(n5850), .Z(n5852) );
  XNOR U6261 ( .A(n5853), .B(n5852), .Z(zout[14]) );
  NANDN U6262 ( .A(n525), .B(n[150]), .Z(n5863) );
  NANDN U6263 ( .A(n5855), .B(n5854), .Z(n5859) );
  OR U6264 ( .A(n5857), .B(n5856), .Z(n5858) );
  AND U6265 ( .A(n5859), .B(n5858), .Z(n5862) );
  XOR U6266 ( .A(n5861), .B(n5862), .Z(n5860) );
  XNOR U6267 ( .A(n5863), .B(n5860), .Z(zout[150]) );
  NANDN U6268 ( .A(n525), .B(n[151]), .Z(n5864) );
  XOR U6269 ( .A(n5866), .B(n5864), .Z(n5869) );
  XOR U6270 ( .A(n5868), .B(n5869), .Z(zout[151]) );
  NANDN U6271 ( .A(n525), .B(n[152]), .Z(n5865) );
  XOR U6272 ( .A(n5872), .B(n5865), .Z(n5875) );
  AND U6273 ( .A(n5866), .B(n[151]), .Z(n5867) );
  NANDN U6274 ( .A(n525), .B(n5867), .Z(n5871) );
  NANDN U6275 ( .A(n5869), .B(n5868), .Z(n5870) );
  AND U6276 ( .A(n5871), .B(n5870), .Z(n5874) );
  XNOR U6277 ( .A(n5875), .B(n5874), .Z(zout[152]) );
  NANDN U6278 ( .A(n525), .B(n[153]), .Z(n5881) );
  AND U6279 ( .A(n5872), .B(n[152]), .Z(n5873) );
  NANDN U6280 ( .A(n525), .B(n5873), .Z(n5877) );
  OR U6281 ( .A(n5875), .B(n5874), .Z(n5876) );
  AND U6282 ( .A(n5877), .B(n5876), .Z(n5880) );
  XOR U6283 ( .A(n5879), .B(n5880), .Z(n5878) );
  XNOR U6284 ( .A(n5881), .B(n5878), .Z(zout[153]) );
  NANDN U6285 ( .A(n525), .B(n[154]), .Z(n5882) );
  XOR U6286 ( .A(n5883), .B(n5882), .Z(n5886) );
  XOR U6287 ( .A(n5885), .B(n5886), .Z(zout[154]) );
  NANDN U6288 ( .A(n525), .B(n[155]), .Z(n5893) );
  XOR U6289 ( .A(n5892), .B(n5893), .Z(n5895) );
  AND U6290 ( .A(n5883), .B(n[154]), .Z(n5884) );
  NANDN U6291 ( .A(n525), .B(n5884), .Z(n5888) );
  NANDN U6292 ( .A(n5886), .B(n5885), .Z(n5887) );
  AND U6293 ( .A(n5888), .B(n5887), .Z(n5894) );
  XNOR U6294 ( .A(n5895), .B(n5894), .Z(zout[155]) );
  NANDN U6295 ( .A(n5889), .B(n6814), .Z(n5890) );
  XOR U6296 ( .A(n5891), .B(n5890), .Z(n5899) );
  NANDN U6297 ( .A(n5893), .B(n5892), .Z(n5897) );
  OR U6298 ( .A(n5895), .B(n5894), .Z(n5896) );
  AND U6299 ( .A(n5897), .B(n5896), .Z(n5900) );
  XOR U6300 ( .A(n5899), .B(n5900), .Z(zout[156]) );
  NANDN U6301 ( .A(n525), .B(n[157]), .Z(n5907) );
  XOR U6302 ( .A(n5906), .B(n5907), .Z(n5909) );
  OR U6303 ( .A(n5898), .B(n525), .Z(n5902) );
  NANDN U6304 ( .A(n5900), .B(n5899), .Z(n5901) );
  AND U6305 ( .A(n5902), .B(n5901), .Z(n5908) );
  XNOR U6306 ( .A(n5909), .B(n5908), .Z(zout[157]) );
  NANDN U6307 ( .A(n5903), .B(n6814), .Z(n5904) );
  XNOR U6308 ( .A(n5905), .B(n5904), .Z(n5913) );
  NANDN U6309 ( .A(n5907), .B(n5906), .Z(n5911) );
  OR U6310 ( .A(n5909), .B(n5908), .Z(n5910) );
  AND U6311 ( .A(n5911), .B(n5910), .Z(n5914) );
  XOR U6312 ( .A(n5913), .B(n5914), .Z(zout[158]) );
  NANDN U6313 ( .A(n525), .B(n5912), .Z(n5916) );
  NANDN U6314 ( .A(n5914), .B(n5913), .Z(n5915) );
  NAND U6315 ( .A(n5916), .B(n5915), .Z(n5920) );
  AND U6316 ( .A(n[159]), .B(n6814), .Z(n5921) );
  XOR U6317 ( .A(n5919), .B(n5921), .Z(n5917) );
  XNOR U6318 ( .A(n5920), .B(n5917), .Z(zout[159]) );
  AND U6319 ( .A(n6814), .B(n[15]), .Z(n5979) );
  XNOR U6320 ( .A(n5978), .B(n5979), .Z(n5976) );
  AND U6321 ( .A(n6814), .B(n5918), .Z(n5977) );
  XOR U6322 ( .A(n5976), .B(n5977), .Z(zout[15]) );
  NANDN U6323 ( .A(n525), .B(n[160]), .Z(n5923) );
  XNOR U6324 ( .A(n5924), .B(n5925), .Z(n5922) );
  XNOR U6325 ( .A(n5923), .B(n5922), .Z(zout[160]) );
  AND U6326 ( .A(n[161]), .B(n6814), .Z(n5929) );
  XNOR U6327 ( .A(n5928), .B(n5927), .Z(n5926) );
  XNOR U6328 ( .A(n5929), .B(n5926), .Z(zout[161]) );
  NANDN U6329 ( .A(n525), .B(n[162]), .Z(n5932) );
  XOR U6330 ( .A(n5931), .B(n5932), .Z(n5934) );
  XNOR U6331 ( .A(n5933), .B(n5934), .Z(zout[162]) );
  NANDN U6332 ( .A(n525), .B(n[163]), .Z(n5930) );
  XOR U6333 ( .A(n5937), .B(n5930), .Z(n5940) );
  NANDN U6334 ( .A(n5932), .B(n5931), .Z(n5936) );
  OR U6335 ( .A(n5934), .B(n5933), .Z(n5935) );
  AND U6336 ( .A(n5936), .B(n5935), .Z(n5939) );
  XNOR U6337 ( .A(n5940), .B(n5939), .Z(zout[163]) );
  AND U6338 ( .A(n5937), .B(n[163]), .Z(n5938) );
  NANDN U6339 ( .A(n525), .B(n5938), .Z(n5942) );
  OR U6340 ( .A(n5940), .B(n5939), .Z(n5941) );
  NAND U6341 ( .A(n5942), .B(n5941), .Z(n5946) );
  XOR U6342 ( .A(n5945), .B(n5946), .Z(n5947) );
  NANDN U6343 ( .A(n5943), .B(n6814), .Z(n5948) );
  XOR U6344 ( .A(n5947), .B(n5948), .Z(zout[164]) );
  NANDN U6345 ( .A(n525), .B(n[165]), .Z(n5944) );
  XOR U6346 ( .A(n5951), .B(n5944), .Z(n5954) );
  NAND U6347 ( .A(n5946), .B(n5945), .Z(n5950) );
  NANDN U6348 ( .A(n5948), .B(n5947), .Z(n5949) );
  AND U6349 ( .A(n5950), .B(n5949), .Z(n5953) );
  XNOR U6350 ( .A(n5954), .B(n5953), .Z(zout[165]) );
  NANDN U6351 ( .A(n525), .B(n[166]), .Z(n5959) );
  XOR U6352 ( .A(n5958), .B(n5959), .Z(n5961) );
  AND U6353 ( .A(n5951), .B(n[165]), .Z(n5952) );
  NANDN U6354 ( .A(n525), .B(n5952), .Z(n5956) );
  OR U6355 ( .A(n5954), .B(n5953), .Z(n5955) );
  AND U6356 ( .A(n5956), .B(n5955), .Z(n5960) );
  XNOR U6357 ( .A(n5961), .B(n5960), .Z(zout[166]) );
  NANDN U6358 ( .A(n525), .B(n[167]), .Z(n5957) );
  XOR U6359 ( .A(n5964), .B(n5957), .Z(n5967) );
  NANDN U6360 ( .A(n5959), .B(n5958), .Z(n5963) );
  OR U6361 ( .A(n5961), .B(n5960), .Z(n5962) );
  AND U6362 ( .A(n5963), .B(n5962), .Z(n5966) );
  XNOR U6363 ( .A(n5967), .B(n5966), .Z(zout[167]) );
  NANDN U6364 ( .A(n525), .B(n[168]), .Z(n5971) );
  XOR U6365 ( .A(n5970), .B(n5971), .Z(n5973) );
  AND U6366 ( .A(n5964), .B(n[167]), .Z(n5965) );
  NANDN U6367 ( .A(n525), .B(n5965), .Z(n5969) );
  OR U6368 ( .A(n5967), .B(n5966), .Z(n5968) );
  AND U6369 ( .A(n5969), .B(n5968), .Z(n5972) );
  XNOR U6370 ( .A(n5973), .B(n5972), .Z(zout[168]) );
  NANDN U6371 ( .A(n5971), .B(n5970), .Z(n5975) );
  OR U6372 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U6373 ( .A(n5975), .B(n5974), .Z(n5987) );
  XOR U6374 ( .A(n5986), .B(n5987), .Z(n5988) );
  NANDN U6375 ( .A(n525), .B(n[169]), .Z(n5989) );
  XOR U6376 ( .A(n5988), .B(n5989), .Z(zout[169]) );
  OR U6377 ( .A(n5977), .B(n5976), .Z(n5981) );
  OR U6378 ( .A(n5979), .B(n5978), .Z(n5980) );
  AND U6379 ( .A(n5981), .B(n5980), .Z(n5983) );
  NANDN U6380 ( .A(n525), .B(n[16]), .Z(n5982) );
  XNOR U6381 ( .A(n5983), .B(n5982), .Z(n5984) );
  XNOR U6382 ( .A(n5985), .B(n5984), .Z(zout[16]) );
  AND U6383 ( .A(n6814), .B(n[170]), .Z(n5996) );
  NAND U6384 ( .A(n5987), .B(n5986), .Z(n5991) );
  NANDN U6385 ( .A(n5989), .B(n5988), .Z(n5990) );
  AND U6386 ( .A(n5991), .B(n5990), .Z(n5995) );
  XNOR U6387 ( .A(n5993), .B(n5995), .Z(n5992) );
  XOR U6388 ( .A(n5996), .B(n5992), .Z(zout[170]) );
  NANDN U6389 ( .A(n5998), .B(n6814), .Z(n5997) );
  XOR U6390 ( .A(n5999), .B(n5997), .Z(n6001) );
  XNOR U6391 ( .A(n6002), .B(n6001), .Z(zout[171]) );
  NANDN U6392 ( .A(n525), .B(n[172]), .Z(n6006) );
  XOR U6393 ( .A(n6005), .B(n6006), .Z(n6008) );
  ANDN U6394 ( .B(n5999), .A(n5998), .Z(n6000) );
  NANDN U6395 ( .A(n525), .B(n6000), .Z(n6004) );
  OR U6396 ( .A(n6002), .B(n6001), .Z(n6003) );
  AND U6397 ( .A(n6004), .B(n6003), .Z(n6007) );
  XNOR U6398 ( .A(n6008), .B(n6007), .Z(zout[172]) );
  NANDN U6399 ( .A(n525), .B(n[173]), .Z(n6013) );
  XOR U6400 ( .A(n6012), .B(n6013), .Z(n6015) );
  NANDN U6401 ( .A(n6006), .B(n6005), .Z(n6010) );
  OR U6402 ( .A(n6008), .B(n6007), .Z(n6009) );
  AND U6403 ( .A(n6010), .B(n6009), .Z(n6014) );
  XNOR U6404 ( .A(n6015), .B(n6014), .Z(zout[173]) );
  NANDN U6405 ( .A(n525), .B(n[174]), .Z(n6011) );
  XOR U6406 ( .A(n6018), .B(n6011), .Z(n6021) );
  NANDN U6407 ( .A(n6013), .B(n6012), .Z(n6017) );
  OR U6408 ( .A(n6015), .B(n6014), .Z(n6016) );
  AND U6409 ( .A(n6017), .B(n6016), .Z(n6020) );
  XNOR U6410 ( .A(n6021), .B(n6020), .Z(zout[174]) );
  AND U6411 ( .A(n6018), .B(n[174]), .Z(n6019) );
  NANDN U6412 ( .A(n525), .B(n6019), .Z(n6023) );
  OR U6413 ( .A(n6021), .B(n6020), .Z(n6022) );
  NAND U6414 ( .A(n6023), .B(n6022), .Z(n6027) );
  XOR U6415 ( .A(n6026), .B(n6027), .Z(n6028) );
  NANDN U6416 ( .A(n6024), .B(n6814), .Z(n6029) );
  XOR U6417 ( .A(n6028), .B(n6029), .Z(zout[175]) );
  NANDN U6418 ( .A(n6025), .B(n6814), .Z(n6032) );
  XOR U6419 ( .A(n6033), .B(n6032), .Z(n6034) );
  NAND U6420 ( .A(n6027), .B(n6026), .Z(n6031) );
  NANDN U6421 ( .A(n6029), .B(n6028), .Z(n6030) );
  NAND U6422 ( .A(n6031), .B(n6030), .Z(n6035) );
  XNOR U6423 ( .A(n6034), .B(n6035), .Z(zout[176]) );
  AND U6424 ( .A(n6033), .B(n6032), .Z(n6037) );
  NANDN U6425 ( .A(n6035), .B(n6034), .Z(n6036) );
  NANDN U6426 ( .A(n6037), .B(n6036), .Z(n6046) );
  NANDN U6427 ( .A(n525), .B(n[177]), .Z(n6038) );
  XOR U6428 ( .A(n6043), .B(n6038), .Z(n6045) );
  XNOR U6429 ( .A(n6046), .B(n6045), .Z(zout[177]) );
  NANDN U6430 ( .A(n6039), .B(n6814), .Z(n6040) );
  XOR U6431 ( .A(n6041), .B(n6040), .Z(n6050) );
  ANDN U6432 ( .B(n6043), .A(n6042), .Z(n6044) );
  NANDN U6433 ( .A(n525), .B(n6044), .Z(n6048) );
  OR U6434 ( .A(n6046), .B(n6045), .Z(n6047) );
  AND U6435 ( .A(n6048), .B(n6047), .Z(n6051) );
  XOR U6436 ( .A(n6050), .B(n6051), .Z(zout[178]) );
  NANDN U6437 ( .A(n525), .B(n[179]), .Z(n6056) );
  XOR U6438 ( .A(n6055), .B(n6056), .Z(n6058) );
  OR U6439 ( .A(n6049), .B(n525), .Z(n6053) );
  NANDN U6440 ( .A(n6051), .B(n6050), .Z(n6052) );
  AND U6441 ( .A(n6053), .B(n6052), .Z(n6057) );
  XNOR U6442 ( .A(n6058), .B(n6057), .Z(zout[179]) );
  NOR U6443 ( .A(n525), .B(n6054), .Z(n6123) );
  XNOR U6444 ( .A(n6122), .B(n6123), .Z(n6120) );
  AND U6445 ( .A(n6814), .B(n[17]), .Z(n6121) );
  XOR U6446 ( .A(n6120), .B(n6121), .Z(zout[17]) );
  NANDN U6447 ( .A(n6056), .B(n6055), .Z(n6060) );
  OR U6448 ( .A(n6058), .B(n6057), .Z(n6059) );
  NAND U6449 ( .A(n6060), .B(n6059), .Z(n6062) );
  XOR U6450 ( .A(n6061), .B(n6062), .Z(n6063) );
  NANDN U6451 ( .A(n525), .B(n[180]), .Z(n6064) );
  XOR U6452 ( .A(n6063), .B(n6064), .Z(zout[180]) );
  NANDN U6453 ( .A(n525), .B(n[181]), .Z(n6068) );
  XOR U6454 ( .A(n6067), .B(n6068), .Z(n6070) );
  NAND U6455 ( .A(n6062), .B(n6061), .Z(n6066) );
  NANDN U6456 ( .A(n6064), .B(n6063), .Z(n6065) );
  AND U6457 ( .A(n6066), .B(n6065), .Z(n6069) );
  XNOR U6458 ( .A(n6070), .B(n6069), .Z(zout[181]) );
  NANDN U6459 ( .A(n525), .B(n[182]), .Z(n6074) );
  XOR U6460 ( .A(n6073), .B(n6074), .Z(n6076) );
  NANDN U6461 ( .A(n6068), .B(n6067), .Z(n6072) );
  OR U6462 ( .A(n6070), .B(n6069), .Z(n6071) );
  AND U6463 ( .A(n6072), .B(n6071), .Z(n6075) );
  XNOR U6464 ( .A(n6076), .B(n6075), .Z(zout[182]) );
  NANDN U6465 ( .A(n525), .B(n[183]), .Z(n6081) );
  XOR U6466 ( .A(n6080), .B(n6081), .Z(n6083) );
  NANDN U6467 ( .A(n6074), .B(n6073), .Z(n6078) );
  OR U6468 ( .A(n6076), .B(n6075), .Z(n6077) );
  AND U6469 ( .A(n6078), .B(n6077), .Z(n6082) );
  XNOR U6470 ( .A(n6083), .B(n6082), .Z(zout[183]) );
  NANDN U6471 ( .A(n6086), .B(n6814), .Z(n6079) );
  XOR U6472 ( .A(n6087), .B(n6079), .Z(n6090) );
  NANDN U6473 ( .A(n6081), .B(n6080), .Z(n6085) );
  OR U6474 ( .A(n6083), .B(n6082), .Z(n6084) );
  AND U6475 ( .A(n6085), .B(n6084), .Z(n6089) );
  XNOR U6476 ( .A(n6090), .B(n6089), .Z(zout[184]) );
  ANDN U6477 ( .B(n6087), .A(n6086), .Z(n6088) );
  NANDN U6478 ( .A(n525), .B(n6088), .Z(n6092) );
  OR U6479 ( .A(n6090), .B(n6089), .Z(n6091) );
  NAND U6480 ( .A(n6092), .B(n6091), .Z(n6094) );
  XOR U6481 ( .A(n6093), .B(n6094), .Z(n6095) );
  NANDN U6482 ( .A(n525), .B(n[185]), .Z(n6096) );
  XOR U6483 ( .A(n6095), .B(n6096), .Z(zout[185]) );
  NANDN U6484 ( .A(n525), .B(n[186]), .Z(n6101) );
  XOR U6485 ( .A(n6100), .B(n6101), .Z(n6103) );
  NAND U6486 ( .A(n6094), .B(n6093), .Z(n6098) );
  NANDN U6487 ( .A(n6096), .B(n6095), .Z(n6097) );
  AND U6488 ( .A(n6098), .B(n6097), .Z(n6102) );
  XNOR U6489 ( .A(n6103), .B(n6102), .Z(zout[186]) );
  NANDN U6490 ( .A(n6106), .B(n6814), .Z(n6099) );
  XOR U6491 ( .A(n6107), .B(n6099), .Z(n6110) );
  NANDN U6492 ( .A(n6101), .B(n6100), .Z(n6105) );
  OR U6493 ( .A(n6103), .B(n6102), .Z(n6104) );
  AND U6494 ( .A(n6105), .B(n6104), .Z(n6109) );
  XNOR U6495 ( .A(n6110), .B(n6109), .Z(zout[187]) );
  NANDN U6496 ( .A(n525), .B(n[188]), .Z(n6114) );
  XOR U6497 ( .A(n6113), .B(n6114), .Z(n6116) );
  ANDN U6498 ( .B(n6107), .A(n6106), .Z(n6108) );
  NANDN U6499 ( .A(n525), .B(n6108), .Z(n6112) );
  OR U6500 ( .A(n6110), .B(n6109), .Z(n6111) );
  AND U6501 ( .A(n6112), .B(n6111), .Z(n6115) );
  XNOR U6502 ( .A(n6116), .B(n6115), .Z(zout[188]) );
  NANDN U6503 ( .A(n6114), .B(n6113), .Z(n6118) );
  OR U6504 ( .A(n6116), .B(n6115), .Z(n6117) );
  NAND U6505 ( .A(n6118), .B(n6117), .Z(n6131) );
  AND U6506 ( .A(n6814), .B(n[189]), .Z(n6132) );
  XOR U6507 ( .A(n6130), .B(n6132), .Z(n6119) );
  XNOR U6508 ( .A(n6131), .B(n6119), .Z(zout[189]) );
  OR U6509 ( .A(n6121), .B(n6120), .Z(n6125) );
  OR U6510 ( .A(n6123), .B(n6122), .Z(n6124) );
  AND U6511 ( .A(n6125), .B(n6124), .Z(n6127) );
  NANDN U6512 ( .A(n525), .B(n[18]), .Z(n6126) );
  XNOR U6513 ( .A(n6127), .B(n6126), .Z(n6128) );
  XNOR U6514 ( .A(n6129), .B(n6128), .Z(zout[18]) );
  NANDN U6515 ( .A(n525), .B(n[190]), .Z(n6133) );
  XOR U6516 ( .A(n6136), .B(n6133), .Z(n6138) );
  XNOR U6517 ( .A(n6139), .B(n6138), .Z(zout[190]) );
  NANDN U6518 ( .A(n525), .B(n[191]), .Z(n6134) );
  XOR U6519 ( .A(n6142), .B(n6134), .Z(n6145) );
  ANDN U6520 ( .B(n6136), .A(n6135), .Z(n6137) );
  NANDN U6521 ( .A(n525), .B(n6137), .Z(n6141) );
  OR U6522 ( .A(n6139), .B(n6138), .Z(n6140) );
  AND U6523 ( .A(n6141), .B(n6140), .Z(n6144) );
  XNOR U6524 ( .A(n6145), .B(n6144), .Z(zout[191]) );
  NANDN U6525 ( .A(n525), .B(n[192]), .Z(n6149) );
  XOR U6526 ( .A(n6148), .B(n6149), .Z(n6151) );
  AND U6527 ( .A(n6142), .B(n[191]), .Z(n6143) );
  NANDN U6528 ( .A(n525), .B(n6143), .Z(n6147) );
  OR U6529 ( .A(n6145), .B(n6144), .Z(n6146) );
  AND U6530 ( .A(n6147), .B(n6146), .Z(n6150) );
  XNOR U6531 ( .A(n6151), .B(n6150), .Z(zout[192]) );
  NANDN U6532 ( .A(n525), .B(n[193]), .Z(n6155) );
  XOR U6533 ( .A(n6154), .B(n6155), .Z(n6157) );
  NANDN U6534 ( .A(n6149), .B(n6148), .Z(n6153) );
  OR U6535 ( .A(n6151), .B(n6150), .Z(n6152) );
  AND U6536 ( .A(n6153), .B(n6152), .Z(n6156) );
  XNOR U6537 ( .A(n6157), .B(n6156), .Z(zout[193]) );
  NANDN U6538 ( .A(n525), .B(n[194]), .Z(n6161) );
  XOR U6539 ( .A(n6160), .B(n6161), .Z(n6163) );
  NANDN U6540 ( .A(n6155), .B(n6154), .Z(n6159) );
  OR U6541 ( .A(n6157), .B(n6156), .Z(n6158) );
  AND U6542 ( .A(n6159), .B(n6158), .Z(n6162) );
  XNOR U6543 ( .A(n6163), .B(n6162), .Z(zout[194]) );
  NANDN U6544 ( .A(n525), .B(n[195]), .Z(n6170) );
  XOR U6545 ( .A(n6169), .B(n6170), .Z(n6172) );
  NANDN U6546 ( .A(n6161), .B(n6160), .Z(n6165) );
  OR U6547 ( .A(n6163), .B(n6162), .Z(n6164) );
  AND U6548 ( .A(n6165), .B(n6164), .Z(n6171) );
  XNOR U6549 ( .A(n6172), .B(n6171), .Z(zout[195]) );
  NANDN U6550 ( .A(n6166), .B(n6814), .Z(n6167) );
  XNOR U6551 ( .A(n6168), .B(n6167), .Z(n6176) );
  NANDN U6552 ( .A(n6170), .B(n6169), .Z(n6174) );
  OR U6553 ( .A(n6172), .B(n6171), .Z(n6173) );
  AND U6554 ( .A(n6174), .B(n6173), .Z(n6177) );
  XOR U6555 ( .A(n6176), .B(n6177), .Z(zout[196]) );
  NANDN U6556 ( .A(n525), .B(n[197]), .Z(n6182) );
  XOR U6557 ( .A(n6181), .B(n6182), .Z(n6184) );
  OR U6558 ( .A(n6175), .B(n525), .Z(n6179) );
  NANDN U6559 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U6560 ( .A(n6179), .B(n6178), .Z(n6183) );
  XNOR U6561 ( .A(n6184), .B(n6183), .Z(zout[197]) );
  NANDN U6562 ( .A(n525), .B(n[198]), .Z(n6180) );
  XOR U6563 ( .A(n6188), .B(n6180), .Z(n6191) );
  NANDN U6564 ( .A(n6182), .B(n6181), .Z(n6186) );
  OR U6565 ( .A(n6184), .B(n6183), .Z(n6185) );
  AND U6566 ( .A(n6186), .B(n6185), .Z(n6190) );
  XNOR U6567 ( .A(n6191), .B(n6190), .Z(zout[198]) );
  NANDN U6568 ( .A(n525), .B(n[199]), .Z(n6187) );
  XOR U6569 ( .A(n6202), .B(n6187), .Z(n6205) );
  AND U6570 ( .A(n6188), .B(n[198]), .Z(n6189) );
  NANDN U6571 ( .A(n525), .B(n6189), .Z(n6193) );
  OR U6572 ( .A(n6191), .B(n6190), .Z(n6192) );
  AND U6573 ( .A(n6193), .B(n6192), .Z(n6204) );
  XNOR U6574 ( .A(n6205), .B(n6204), .Z(zout[199]) );
  AND U6575 ( .A(n6814), .B(n[19]), .Z(n6261) );
  XNOR U6576 ( .A(n6260), .B(n6261), .Z(n6258) );
  NOR U6577 ( .A(n525), .B(n6194), .Z(n6259) );
  XOR U6578 ( .A(n6258), .B(n6259), .Z(zout[19]) );
  XOR U6579 ( .A(n[1]), .B(n6195), .Z(n6196) );
  NANDN U6580 ( .A(n525), .B(n6196), .Z(n6197) );
  XNOR U6581 ( .A(n6198), .B(n6197), .Z(zout[1]) );
  NANDN U6582 ( .A(n6199), .B(n6814), .Z(n6200) );
  XNOR U6583 ( .A(n6201), .B(n6200), .Z(n6209) );
  AND U6584 ( .A(n6202), .B(n[199]), .Z(n6203) );
  NANDN U6585 ( .A(n525), .B(n6203), .Z(n6207) );
  OR U6586 ( .A(n6205), .B(n6204), .Z(n6206) );
  AND U6587 ( .A(n6207), .B(n6206), .Z(n6210) );
  XOR U6588 ( .A(n6209), .B(n6210), .Z(zout[200]) );
  NANDN U6589 ( .A(n525), .B(n[201]), .Z(n6214) );
  XOR U6590 ( .A(n6213), .B(n6214), .Z(n6216) );
  OR U6591 ( .A(n6208), .B(n525), .Z(n6212) );
  NANDN U6592 ( .A(n6210), .B(n6209), .Z(n6211) );
  AND U6593 ( .A(n6212), .B(n6211), .Z(n6215) );
  XNOR U6594 ( .A(n6216), .B(n6215), .Z(zout[201]) );
  NANDN U6595 ( .A(n6214), .B(n6213), .Z(n6218) );
  OR U6596 ( .A(n6216), .B(n6215), .Z(n6217) );
  NAND U6597 ( .A(n6218), .B(n6217), .Z(n6220) );
  XOR U6598 ( .A(n6219), .B(n6220), .Z(n6221) );
  NANDN U6599 ( .A(n525), .B(n[202]), .Z(n6222) );
  XOR U6600 ( .A(n6221), .B(n6222), .Z(zout[202]) );
  NAND U6601 ( .A(n6220), .B(n6219), .Z(n6224) );
  NANDN U6602 ( .A(n6222), .B(n6221), .Z(n6223) );
  NAND U6603 ( .A(n6224), .B(n6223), .Z(n6227) );
  XOR U6604 ( .A(n6226), .B(n6227), .Z(n6228) );
  NANDN U6605 ( .A(n6225), .B(n6814), .Z(n6229) );
  XOR U6606 ( .A(n6228), .B(n6229), .Z(zout[203]) );
  NANDN U6607 ( .A(n525), .B(n[204]), .Z(n6233) );
  XOR U6608 ( .A(n6232), .B(n6233), .Z(n6235) );
  NAND U6609 ( .A(n6227), .B(n6226), .Z(n6231) );
  NANDN U6610 ( .A(n6229), .B(n6228), .Z(n6230) );
  AND U6611 ( .A(n6231), .B(n6230), .Z(n6234) );
  XNOR U6612 ( .A(n6235), .B(n6234), .Z(zout[204]) );
  NANDN U6613 ( .A(n6233), .B(n6232), .Z(n6237) );
  OR U6614 ( .A(n6235), .B(n6234), .Z(n6236) );
  NAND U6615 ( .A(n6237), .B(n6236), .Z(n6240) );
  AND U6616 ( .A(n[205]), .B(n6814), .Z(n6241) );
  XOR U6617 ( .A(n6239), .B(n6241), .Z(n6238) );
  XNOR U6618 ( .A(n6240), .B(n6238), .Z(zout[205]) );
  NANDN U6619 ( .A(n525), .B(n[206]), .Z(n6243) );
  XOR U6620 ( .A(n6242), .B(n6243), .Z(n6245) );
  XNOR U6621 ( .A(n6244), .B(n6245), .Z(zout[206]) );
  NANDN U6622 ( .A(n525), .B(n[207]), .Z(n6251) );
  NANDN U6623 ( .A(n6243), .B(n6242), .Z(n6247) );
  OR U6624 ( .A(n6245), .B(n6244), .Z(n6246) );
  AND U6625 ( .A(n6247), .B(n6246), .Z(n6250) );
  XOR U6626 ( .A(n6249), .B(n6250), .Z(n6248) );
  XNOR U6627 ( .A(n6251), .B(n6248), .Z(zout[207]) );
  AND U6628 ( .A(n6814), .B(n[208]), .Z(n6255) );
  XNOR U6629 ( .A(n6254), .B(n6253), .Z(n6252) );
  XNOR U6630 ( .A(n6255), .B(n6252), .Z(zout[208]) );
  NANDN U6631 ( .A(n6256), .B(n6814), .Z(n6257) );
  XOR U6632 ( .A(n6271), .B(n6257), .Z(n6273) );
  XOR U6633 ( .A(n6274), .B(n6273), .Z(zout[209]) );
  OR U6634 ( .A(n6259), .B(n6258), .Z(n6263) );
  OR U6635 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U6636 ( .A(n6263), .B(n6262), .Z(n6265) );
  NANDN U6637 ( .A(n525), .B(n[20]), .Z(n6264) );
  XNOR U6638 ( .A(n6265), .B(n6264), .Z(n6266) );
  XNOR U6639 ( .A(n6267), .B(n6266), .Z(zout[20]) );
  NANDN U6640 ( .A(n6268), .B(n6814), .Z(n6269) );
  XNOR U6641 ( .A(n6270), .B(n6269), .Z(n6279) );
  ANDN U6642 ( .B(n[209]), .A(n6271), .Z(n6272) );
  NANDN U6643 ( .A(n525), .B(n6272), .Z(n6276) );
  NANDN U6644 ( .A(n6274), .B(n6273), .Z(n6275) );
  AND U6645 ( .A(n6276), .B(n6275), .Z(n6280) );
  XOR U6646 ( .A(n6279), .B(n6280), .Z(zout[210]) );
  NANDN U6647 ( .A(n525), .B(n[211]), .Z(n6277) );
  XOR U6648 ( .A(n6283), .B(n6277), .Z(n6286) );
  NANDN U6649 ( .A(n525), .B(n6278), .Z(n6282) );
  NANDN U6650 ( .A(n6280), .B(n6279), .Z(n6281) );
  AND U6651 ( .A(n6282), .B(n6281), .Z(n6285) );
  XNOR U6652 ( .A(n6286), .B(n6285), .Z(zout[211]) );
  NANDN U6653 ( .A(n525), .B(n[212]), .Z(n6290) );
  XOR U6654 ( .A(n6289), .B(n6290), .Z(n6292) );
  AND U6655 ( .A(n6283), .B(n[211]), .Z(n6284) );
  NANDN U6656 ( .A(n525), .B(n6284), .Z(n6288) );
  OR U6657 ( .A(n6286), .B(n6285), .Z(n6287) );
  AND U6658 ( .A(n6288), .B(n6287), .Z(n6291) );
  XNOR U6659 ( .A(n6292), .B(n6291), .Z(zout[212]) );
  NANDN U6660 ( .A(n525), .B(n[213]), .Z(n6296) );
  XOR U6661 ( .A(n6295), .B(n6296), .Z(n6298) );
  NANDN U6662 ( .A(n6290), .B(n6289), .Z(n6294) );
  OR U6663 ( .A(n6292), .B(n6291), .Z(n6293) );
  AND U6664 ( .A(n6294), .B(n6293), .Z(n6297) );
  XNOR U6665 ( .A(n6298), .B(n6297), .Z(zout[213]) );
  AND U6666 ( .A(n[214]), .B(n6814), .Z(n6304) );
  NANDN U6667 ( .A(n6296), .B(n6295), .Z(n6300) );
  OR U6668 ( .A(n6298), .B(n6297), .Z(n6299) );
  AND U6669 ( .A(n6300), .B(n6299), .Z(n6303) );
  XNOR U6670 ( .A(n6302), .B(n6303), .Z(n6301) );
  XOR U6671 ( .A(n6304), .B(n6301), .Z(zout[214]) );
  NANDN U6672 ( .A(n525), .B(n[215]), .Z(n6306) );
  XOR U6673 ( .A(n6305), .B(n6306), .Z(n6308) );
  XNOR U6674 ( .A(n6307), .B(n6308), .Z(zout[215]) );
  NANDN U6675 ( .A(n525), .B(n[216]), .Z(n6312) );
  XOR U6676 ( .A(n6311), .B(n6312), .Z(n6314) );
  NANDN U6677 ( .A(n6306), .B(n6305), .Z(n6310) );
  OR U6678 ( .A(n6308), .B(n6307), .Z(n6309) );
  AND U6679 ( .A(n6310), .B(n6309), .Z(n6313) );
  XNOR U6680 ( .A(n6314), .B(n6313), .Z(zout[216]) );
  NANDN U6681 ( .A(n6312), .B(n6311), .Z(n6316) );
  OR U6682 ( .A(n6314), .B(n6313), .Z(n6315) );
  NAND U6683 ( .A(n6316), .B(n6315), .Z(n6321) );
  XOR U6684 ( .A(n6320), .B(n6321), .Z(n6322) );
  NANDN U6685 ( .A(n525), .B(n[217]), .Z(n6323) );
  XOR U6686 ( .A(n6322), .B(n6323), .Z(zout[217]) );
  NANDN U6687 ( .A(n6317), .B(n6814), .Z(n6318) );
  XNOR U6688 ( .A(n6319), .B(n6318), .Z(n6327) );
  NAND U6689 ( .A(n6321), .B(n6320), .Z(n6325) );
  NANDN U6690 ( .A(n6323), .B(n6322), .Z(n6324) );
  AND U6691 ( .A(n6325), .B(n6324), .Z(n6328) );
  XOR U6692 ( .A(n6327), .B(n6328), .Z(zout[218]) );
  NANDN U6693 ( .A(n525), .B(n[219]), .Z(n6336) );
  XOR U6694 ( .A(n6335), .B(n6336), .Z(n6338) );
  OR U6695 ( .A(n6326), .B(n525), .Z(n6330) );
  NANDN U6696 ( .A(n6328), .B(n6327), .Z(n6329) );
  AND U6697 ( .A(n6330), .B(n6329), .Z(n6337) );
  XNOR U6698 ( .A(n6338), .B(n6337), .Z(zout[219]) );
  XOR U6699 ( .A(n[21]), .B(n6331), .Z(n6332) );
  NANDN U6700 ( .A(n525), .B(n6332), .Z(n6333) );
  XOR U6701 ( .A(n6334), .B(n6333), .Z(zout[21]) );
  NANDN U6702 ( .A(n6336), .B(n6335), .Z(n6340) );
  OR U6703 ( .A(n6338), .B(n6337), .Z(n6339) );
  AND U6704 ( .A(n6340), .B(n6339), .Z(n6347) );
  AND U6705 ( .A(n6342), .B(n[220]), .Z(n6341) );
  NAND U6706 ( .A(n6814), .B(n6341), .Z(n6346) );
  NANDN U6707 ( .A(n525), .B(n[220]), .Z(n6343) );
  ANDN U6708 ( .B(n6343), .A(n6342), .Z(n6349) );
  ANDN U6709 ( .B(n6346), .A(n6349), .Z(n6344) );
  XOR U6710 ( .A(n6347), .B(n6344), .Z(zout[220]) );
  NANDN U6711 ( .A(n525), .B(n[221]), .Z(n6345) );
  XOR U6712 ( .A(n6351), .B(n6345), .Z(n6354) );
  NAND U6713 ( .A(n6347), .B(n6346), .Z(n6348) );
  NANDN U6714 ( .A(n6349), .B(n6348), .Z(n6353) );
  XNOR U6715 ( .A(n6354), .B(n6353), .Z(zout[221]) );
  NANDN U6716 ( .A(n525), .B(n[222]), .Z(n6350) );
  XOR U6717 ( .A(n6358), .B(n6350), .Z(n6361) );
  AND U6718 ( .A(n6351), .B(n[221]), .Z(n6352) );
  NANDN U6719 ( .A(n525), .B(n6352), .Z(n6356) );
  OR U6720 ( .A(n6354), .B(n6353), .Z(n6355) );
  AND U6721 ( .A(n6356), .B(n6355), .Z(n6360) );
  XNOR U6722 ( .A(n6361), .B(n6360), .Z(zout[222]) );
  ANDN U6723 ( .B(n6358), .A(n6357), .Z(n6359) );
  NANDN U6724 ( .A(n525), .B(n6359), .Z(n6363) );
  OR U6725 ( .A(n6361), .B(n6360), .Z(n6362) );
  NAND U6726 ( .A(n6363), .B(n6362), .Z(n6364) );
  XOR U6727 ( .A(n6365), .B(n6364), .Z(n6366) );
  AND U6728 ( .A(n[223]), .B(n6814), .Z(n6367) );
  XNOR U6729 ( .A(n6366), .B(n6367), .Z(zout[223]) );
  OR U6730 ( .A(n6365), .B(n6364), .Z(n6369) );
  NANDN U6731 ( .A(n6367), .B(n6366), .Z(n6368) );
  AND U6732 ( .A(n6369), .B(n6368), .Z(n6370) );
  XOR U6733 ( .A(n6371), .B(n6370), .Z(n6372) );
  AND U6734 ( .A(n[224]), .B(n6814), .Z(n6373) );
  XNOR U6735 ( .A(n6372), .B(n6373), .Z(zout[224]) );
  OR U6736 ( .A(n6371), .B(n6370), .Z(n6375) );
  NANDN U6737 ( .A(n6373), .B(n6372), .Z(n6374) );
  AND U6738 ( .A(n6375), .B(n6374), .Z(n6378) );
  XOR U6739 ( .A(n6377), .B(n6378), .Z(n6379) );
  NANDN U6740 ( .A(n6376), .B(n6814), .Z(n6380) );
  XOR U6741 ( .A(n6379), .B(n6380), .Z(zout[225]) );
  NANDN U6742 ( .A(n525), .B(n[226]), .Z(n6384) );
  XOR U6743 ( .A(n6383), .B(n6384), .Z(n6386) );
  NAND U6744 ( .A(n6378), .B(n6377), .Z(n6382) );
  NANDN U6745 ( .A(n6380), .B(n6379), .Z(n6381) );
  AND U6746 ( .A(n6382), .B(n6381), .Z(n6385) );
  XNOR U6747 ( .A(n6386), .B(n6385), .Z(zout[226]) );
  NANDN U6748 ( .A(n525), .B(n[227]), .Z(n6391) );
  XOR U6749 ( .A(n6390), .B(n6391), .Z(n6393) );
  NANDN U6750 ( .A(n6384), .B(n6383), .Z(n6388) );
  OR U6751 ( .A(n6386), .B(n6385), .Z(n6387) );
  AND U6752 ( .A(n6388), .B(n6387), .Z(n6392) );
  XNOR U6753 ( .A(n6393), .B(n6392), .Z(zout[227]) );
  NANDN U6754 ( .A(n525), .B(n[228]), .Z(n6389) );
  XOR U6755 ( .A(n6397), .B(n6389), .Z(n6400) );
  NANDN U6756 ( .A(n6391), .B(n6390), .Z(n6395) );
  OR U6757 ( .A(n6393), .B(n6392), .Z(n6394) );
  AND U6758 ( .A(n6395), .B(n6394), .Z(n6399) );
  XNOR U6759 ( .A(n6400), .B(n6399), .Z(zout[228]) );
  NANDN U6760 ( .A(n525), .B(n[229]), .Z(n6396) );
  XOR U6761 ( .A(n6407), .B(n6396), .Z(n6410) );
  AND U6762 ( .A(n6397), .B(n[228]), .Z(n6398) );
  NANDN U6763 ( .A(n525), .B(n6398), .Z(n6402) );
  OR U6764 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U6765 ( .A(n6402), .B(n6401), .Z(n6409) );
  XNOR U6766 ( .A(n6410), .B(n6409), .Z(zout[229]) );
  XNOR U6767 ( .A(n[22]), .B(n6403), .Z(n6404) );
  NANDN U6768 ( .A(n525), .B(n6404), .Z(n6405) );
  XOR U6769 ( .A(n6406), .B(n6405), .Z(zout[22]) );
  NANDN U6770 ( .A(n525), .B(n[230]), .Z(n6417) );
  XOR U6771 ( .A(n6416), .B(n6417), .Z(n6419) );
  AND U6772 ( .A(n6407), .B(n[229]), .Z(n6408) );
  NANDN U6773 ( .A(n525), .B(n6408), .Z(n6412) );
  OR U6774 ( .A(n6410), .B(n6409), .Z(n6411) );
  AND U6775 ( .A(n6412), .B(n6411), .Z(n6418) );
  XNOR U6776 ( .A(n6419), .B(n6418), .Z(zout[230]) );
  NANDN U6777 ( .A(n6413), .B(n6814), .Z(n6414) );
  XNOR U6778 ( .A(n6415), .B(n6414), .Z(n6423) );
  NANDN U6779 ( .A(n6417), .B(n6416), .Z(n6421) );
  OR U6780 ( .A(n6419), .B(n6418), .Z(n6420) );
  AND U6781 ( .A(n6421), .B(n6420), .Z(n6424) );
  XOR U6782 ( .A(n6423), .B(n6424), .Z(zout[231]) );
  NANDN U6783 ( .A(n525), .B(n[232]), .Z(n6428) );
  XOR U6784 ( .A(n6427), .B(n6428), .Z(n6430) );
  NANDN U6785 ( .A(n525), .B(n6422), .Z(n6426) );
  NANDN U6786 ( .A(n6424), .B(n6423), .Z(n6425) );
  AND U6787 ( .A(n6426), .B(n6425), .Z(n6429) );
  XNOR U6788 ( .A(n6430), .B(n6429), .Z(zout[232]) );
  NANDN U6789 ( .A(n525), .B(n[233]), .Z(n6436) );
  NANDN U6790 ( .A(n6428), .B(n6427), .Z(n6432) );
  OR U6791 ( .A(n6430), .B(n6429), .Z(n6431) );
  AND U6792 ( .A(n6432), .B(n6431), .Z(n6435) );
  XOR U6793 ( .A(n6434), .B(n6435), .Z(n6433) );
  XNOR U6794 ( .A(n6436), .B(n6433), .Z(zout[233]) );
  NANDN U6795 ( .A(n525), .B(n[234]), .Z(n6440) );
  XNOR U6796 ( .A(n6439), .B(n6438), .Z(n6437) );
  XNOR U6797 ( .A(n6440), .B(n6437), .Z(zout[234]) );
  NANDN U6798 ( .A(n525), .B(n[235]), .Z(n6441) );
  XOR U6799 ( .A(n6443), .B(n6441), .Z(n6446) );
  XOR U6800 ( .A(n6445), .B(n6446), .Z(zout[235]) );
  NANDN U6801 ( .A(n6449), .B(n6814), .Z(n6442) );
  XNOR U6802 ( .A(n6450), .B(n6442), .Z(n6452) );
  AND U6803 ( .A(n6443), .B(n[235]), .Z(n6444) );
  NANDN U6804 ( .A(n525), .B(n6444), .Z(n6448) );
  NANDN U6805 ( .A(n6446), .B(n6445), .Z(n6447) );
  AND U6806 ( .A(n6448), .B(n6447), .Z(n6453) );
  XOR U6807 ( .A(n6452), .B(n6453), .Z(zout[236]) );
  ANDN U6808 ( .B(n6450), .A(n6449), .Z(n6451) );
  NANDN U6809 ( .A(n525), .B(n6451), .Z(n6455) );
  NANDN U6810 ( .A(n6453), .B(n6452), .Z(n6454) );
  NAND U6811 ( .A(n6455), .B(n6454), .Z(n6461) );
  NANDN U6812 ( .A(n6456), .B(n6814), .Z(n6458) );
  AND U6813 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U6814 ( .A(n6459), .B(n6814), .Z(n6463) );
  NANDN U6815 ( .A(n6462), .B(n6463), .Z(n6460) );
  XOR U6816 ( .A(n6461), .B(n6460), .Z(zout[237]) );
  NANDN U6817 ( .A(n6462), .B(n6461), .Z(n6464) );
  AND U6818 ( .A(n6464), .B(n6463), .Z(n6469) );
  NANDN U6819 ( .A(n525), .B(n[238]), .Z(n6465) );
  XOR U6820 ( .A(n6466), .B(n6465), .Z(n6468) );
  XNOR U6821 ( .A(n6469), .B(n6468), .Z(zout[238]) );
  AND U6822 ( .A(n6466), .B(n[238]), .Z(n6467) );
  NANDN U6823 ( .A(n525), .B(n6467), .Z(n6471) );
  OR U6824 ( .A(n6469), .B(n6468), .Z(n6470) );
  NAND U6825 ( .A(n6471), .B(n6470), .Z(n6475) );
  AND U6826 ( .A(n6814), .B(n[239]), .Z(n6476) );
  XOR U6827 ( .A(n6474), .B(n6476), .Z(n6472) );
  XNOR U6828 ( .A(n6475), .B(n6472), .Z(zout[239]) );
  AND U6829 ( .A(n6814), .B(n[23]), .Z(n6538) );
  XNOR U6830 ( .A(n6537), .B(n6538), .Z(n6535) );
  AND U6831 ( .A(n6814), .B(n6473), .Z(n6536) );
  XOR U6832 ( .A(n6535), .B(n6536), .Z(zout[23]) );
  NANDN U6833 ( .A(n525), .B(n[240]), .Z(n6478) );
  XOR U6834 ( .A(n6477), .B(n6478), .Z(n6480) );
  XNOR U6835 ( .A(n6480), .B(n6479), .Z(zout[240]) );
  NANDN U6836 ( .A(n525), .B(n[241]), .Z(n6484) );
  XOR U6837 ( .A(n6483), .B(n6484), .Z(n6486) );
  NANDN U6838 ( .A(n6478), .B(n6477), .Z(n6482) );
  OR U6839 ( .A(n6480), .B(n6479), .Z(n6481) );
  AND U6840 ( .A(n6482), .B(n6481), .Z(n6485) );
  XNOR U6841 ( .A(n6486), .B(n6485), .Z(zout[241]) );
  NANDN U6842 ( .A(n525), .B(n[242]), .Z(n6491) );
  XOR U6843 ( .A(n6490), .B(n6491), .Z(n6493) );
  NANDN U6844 ( .A(n6484), .B(n6483), .Z(n6488) );
  OR U6845 ( .A(n6486), .B(n6485), .Z(n6487) );
  AND U6846 ( .A(n6488), .B(n6487), .Z(n6492) );
  XNOR U6847 ( .A(n6493), .B(n6492), .Z(zout[242]) );
  NANDN U6848 ( .A(n525), .B(n[243]), .Z(n6489) );
  XOR U6849 ( .A(n6496), .B(n6489), .Z(n6499) );
  NANDN U6850 ( .A(n6491), .B(n6490), .Z(n6495) );
  OR U6851 ( .A(n6493), .B(n6492), .Z(n6494) );
  AND U6852 ( .A(n6495), .B(n6494), .Z(n6498) );
  XNOR U6853 ( .A(n6499), .B(n6498), .Z(zout[243]) );
  NANDN U6854 ( .A(n525), .B(n[244]), .Z(n6505) );
  AND U6855 ( .A(n6496), .B(n[243]), .Z(n6497) );
  NANDN U6856 ( .A(n525), .B(n6497), .Z(n6501) );
  OR U6857 ( .A(n6499), .B(n6498), .Z(n6500) );
  AND U6858 ( .A(n6501), .B(n6500), .Z(n6504) );
  XOR U6859 ( .A(n6503), .B(n6504), .Z(n6502) );
  XNOR U6860 ( .A(n6505), .B(n6502), .Z(zout[244]) );
  NANDN U6861 ( .A(n525), .B(n[245]), .Z(n6506) );
  XOR U6862 ( .A(n6508), .B(n6506), .Z(n6511) );
  XOR U6863 ( .A(n6510), .B(n6511), .Z(zout[245]) );
  NANDN U6864 ( .A(n6514), .B(n6814), .Z(n6507) );
  XOR U6865 ( .A(n6515), .B(n6507), .Z(n6518) );
  AND U6866 ( .A(n6508), .B(n[245]), .Z(n6509) );
  NANDN U6867 ( .A(n525), .B(n6509), .Z(n6513) );
  NANDN U6868 ( .A(n6511), .B(n6510), .Z(n6512) );
  AND U6869 ( .A(n6513), .B(n6512), .Z(n6517) );
  XNOR U6870 ( .A(n6518), .B(n6517), .Z(zout[246]) );
  NANDN U6871 ( .A(n525), .B(n[247]), .Z(n6523) );
  XOR U6872 ( .A(n6522), .B(n6523), .Z(n6525) );
  ANDN U6873 ( .B(n6515), .A(n6514), .Z(n6516) );
  NANDN U6874 ( .A(n525), .B(n6516), .Z(n6520) );
  OR U6875 ( .A(n6518), .B(n6517), .Z(n6519) );
  AND U6876 ( .A(n6520), .B(n6519), .Z(n6524) );
  XNOR U6877 ( .A(n6525), .B(n6524), .Z(zout[247]) );
  NANDN U6878 ( .A(n525), .B(n[248]), .Z(n6521) );
  XOR U6879 ( .A(n6528), .B(n6521), .Z(n6531) );
  NANDN U6880 ( .A(n6523), .B(n6522), .Z(n6527) );
  OR U6881 ( .A(n6525), .B(n6524), .Z(n6526) );
  AND U6882 ( .A(n6527), .B(n6526), .Z(n6530) );
  XNOR U6883 ( .A(n6531), .B(n6530), .Z(zout[248]) );
  AND U6884 ( .A(n6528), .B(n[248]), .Z(n6529) );
  NANDN U6885 ( .A(n525), .B(n6529), .Z(n6533) );
  OR U6886 ( .A(n6531), .B(n6530), .Z(n6532) );
  NAND U6887 ( .A(n6533), .B(n6532), .Z(n6547) );
  XOR U6888 ( .A(n6546), .B(n6547), .Z(n6548) );
  NANDN U6889 ( .A(n6534), .B(n6814), .Z(n6549) );
  XOR U6890 ( .A(n6548), .B(n6549), .Z(zout[249]) );
  OR U6891 ( .A(n6536), .B(n6535), .Z(n6540) );
  OR U6892 ( .A(n6538), .B(n6537), .Z(n6539) );
  AND U6893 ( .A(n6540), .B(n6539), .Z(n6542) );
  NANDN U6894 ( .A(n525), .B(n[24]), .Z(n6541) );
  XNOR U6895 ( .A(n6542), .B(n6541), .Z(n6543) );
  XNOR U6896 ( .A(n6544), .B(n6543), .Z(zout[24]) );
  NANDN U6897 ( .A(n525), .B(n[250]), .Z(n6545) );
  XOR U6898 ( .A(n6552), .B(n6545), .Z(n6555) );
  NAND U6899 ( .A(n6547), .B(n6546), .Z(n6551) );
  NANDN U6900 ( .A(n6549), .B(n6548), .Z(n6550) );
  AND U6901 ( .A(n6551), .B(n6550), .Z(n6554) );
  XNOR U6902 ( .A(n6555), .B(n6554), .Z(zout[250]) );
  NANDN U6903 ( .A(n525), .B(n[251]), .Z(n6559) );
  XOR U6904 ( .A(n6558), .B(n6559), .Z(n6561) );
  AND U6905 ( .A(n6552), .B(n[250]), .Z(n6553) );
  NANDN U6906 ( .A(n525), .B(n6553), .Z(n6557) );
  OR U6907 ( .A(n6555), .B(n6554), .Z(n6556) );
  AND U6908 ( .A(n6557), .B(n6556), .Z(n6560) );
  XNOR U6909 ( .A(n6561), .B(n6560), .Z(zout[251]) );
  NANDN U6910 ( .A(n525), .B(n[252]), .Z(n6565) );
  XOR U6911 ( .A(n6564), .B(n6565), .Z(n6567) );
  NANDN U6912 ( .A(n6559), .B(n6558), .Z(n6563) );
  OR U6913 ( .A(n6561), .B(n6560), .Z(n6562) );
  AND U6914 ( .A(n6563), .B(n6562), .Z(n6566) );
  XNOR U6915 ( .A(n6567), .B(n6566), .Z(zout[252]) );
  NANDN U6916 ( .A(n6565), .B(n6564), .Z(n6569) );
  OR U6917 ( .A(n6567), .B(n6566), .Z(n6568) );
  NAND U6918 ( .A(n6569), .B(n6568), .Z(n6572) );
  XOR U6919 ( .A(n6571), .B(n6572), .Z(n6573) );
  NANDN U6920 ( .A(n525), .B(n[253]), .Z(n6574) );
  XOR U6921 ( .A(n6573), .B(n6574), .Z(zout[253]) );
  NANDN U6922 ( .A(n6582), .B(n6814), .Z(n6570) );
  XOR U6923 ( .A(n6583), .B(n6570), .Z(n6586) );
  NAND U6924 ( .A(n6572), .B(n6571), .Z(n6576) );
  NANDN U6925 ( .A(n6574), .B(n6573), .Z(n6575) );
  AND U6926 ( .A(n6576), .B(n6575), .Z(n6585) );
  XNOR U6927 ( .A(n6586), .B(n6585), .Z(zout[254]) );
  AND U6928 ( .A(n6580), .B(n[255]), .Z(n6578) );
  NAND U6929 ( .A(n6578), .B(n6577), .Z(n6592) );
  NANDN U6930 ( .A(n525), .B(n[255]), .Z(n6579) );
  NANDN U6931 ( .A(n6580), .B(n6579), .Z(n6581) );
  NAND U6932 ( .A(n6592), .B(n6581), .Z(n6590) );
  ANDN U6933 ( .B(n6583), .A(n6582), .Z(n6584) );
  NANDN U6934 ( .A(n525), .B(n6584), .Z(n6588) );
  OR U6935 ( .A(n6586), .B(n6585), .Z(n6587) );
  AND U6936 ( .A(n6588), .B(n6587), .Z(n6589) );
  XNOR U6937 ( .A(n6590), .B(n6589), .Z(zout[255]) );
  NOR U6938 ( .A(n6590), .B(n6589), .Z(n6591) );
  ANDN U6939 ( .B(n6592), .A(n6591), .Z(n6593) );
  XOR U6940 ( .A(n6594), .B(n6593), .Z(zout[256]) );
  NOR U6941 ( .A(n525), .B(n6595), .Z(n6599) );
  XNOR U6942 ( .A(n6598), .B(n6599), .Z(n6596) );
  AND U6943 ( .A(n[25]), .B(n6814), .Z(n6597) );
  XOR U6944 ( .A(n6596), .B(n6597), .Z(zout[25]) );
  OR U6945 ( .A(n6597), .B(n6596), .Z(n6601) );
  OR U6946 ( .A(n6599), .B(n6598), .Z(n6600) );
  AND U6947 ( .A(n6601), .B(n6600), .Z(n6603) );
  NANDN U6948 ( .A(n525), .B(n[26]), .Z(n6602) );
  XNOR U6949 ( .A(n6603), .B(n6602), .Z(n6604) );
  XNOR U6950 ( .A(n6605), .B(n6604), .Z(zout[26]) );
  XOR U6951 ( .A(n[27]), .B(n6606), .Z(n6607) );
  NANDN U6952 ( .A(n525), .B(n6607), .Z(n6608) );
  XOR U6953 ( .A(n6609), .B(n6608), .Z(zout[27]) );
  XOR U6954 ( .A(n[28]), .B(n6610), .Z(n6611) );
  NANDN U6955 ( .A(n525), .B(n6611), .Z(n6612) );
  XOR U6956 ( .A(n6613), .B(n6612), .Z(zout[28]) );
  AND U6957 ( .A(n6814), .B(n[29]), .Z(n6623) );
  XNOR U6958 ( .A(n6622), .B(n6623), .Z(n6620) );
  NOR U6959 ( .A(n525), .B(n6614), .Z(n6621) );
  XOR U6960 ( .A(n6620), .B(n6621), .Z(zout[29]) );
  XNOR U6961 ( .A(n6616), .B(n6615), .Z(n6617) );
  NANDN U6962 ( .A(n525), .B(n6617), .Z(n6618) );
  XOR U6963 ( .A(n6619), .B(n6618), .Z(zout[2]) );
  OR U6964 ( .A(n6621), .B(n6620), .Z(n6625) );
  OR U6965 ( .A(n6623), .B(n6622), .Z(n6624) );
  AND U6966 ( .A(n6625), .B(n6624), .Z(n6627) );
  NANDN U6967 ( .A(n525), .B(n[30]), .Z(n6626) );
  XNOR U6968 ( .A(n6627), .B(n6626), .Z(n6628) );
  XNOR U6969 ( .A(n6629), .B(n6628), .Z(zout[30]) );
  AND U6970 ( .A(n6814), .B(n[31]), .Z(n6634) );
  XNOR U6971 ( .A(n6633), .B(n6634), .Z(n6631) );
  AND U6972 ( .A(n6814), .B(n6630), .Z(n6632) );
  XOR U6973 ( .A(n6631), .B(n6632), .Z(zout[31]) );
  OR U6974 ( .A(n6632), .B(n6631), .Z(n6636) );
  OR U6975 ( .A(n6634), .B(n6633), .Z(n6635) );
  AND U6976 ( .A(n6636), .B(n6635), .Z(n6638) );
  NANDN U6977 ( .A(n525), .B(n[32]), .Z(n6637) );
  XNOR U6978 ( .A(n6638), .B(n6637), .Z(n6639) );
  XNOR U6979 ( .A(n6640), .B(n6639), .Z(zout[32]) );
  XNOR U6980 ( .A(n[33]), .B(n6641), .Z(n6642) );
  ANDN U6981 ( .B(n6642), .A(n525), .Z(n6643) );
  XNOR U6982 ( .A(n6644), .B(n6643), .Z(zout[33]) );
  XNOR U6983 ( .A(n[34]), .B(n6645), .Z(n6646) );
  ANDN U6984 ( .B(n6646), .A(n525), .Z(n6647) );
  XNOR U6985 ( .A(n6648), .B(n6647), .Z(zout[34]) );
  ANDN U6986 ( .B(n6814), .A(n6649), .Z(n6651) );
  XOR U6987 ( .A(n6650), .B(n6651), .Z(n6652) );
  AND U6988 ( .A(n6814), .B(n[35]), .Z(n6653) );
  XNOR U6989 ( .A(n6652), .B(n6653), .Z(zout[35]) );
  OR U6990 ( .A(n6651), .B(n6650), .Z(n6655) );
  NANDN U6991 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U6992 ( .A(n6655), .B(n6654), .Z(n6660) );
  NANDN U6993 ( .A(n6656), .B(n6814), .Z(n6657) );
  XNOR U6994 ( .A(n6658), .B(n6657), .Z(n6659) );
  XNOR U6995 ( .A(n6660), .B(n6659), .Z(zout[36]) );
  NOR U6996 ( .A(n525), .B(n6661), .Z(n6665) );
  XNOR U6997 ( .A(n6664), .B(n6665), .Z(n6662) );
  AND U6998 ( .A(n6814), .B(n[37]), .Z(n6663) );
  XOR U6999 ( .A(n6662), .B(n6663), .Z(zout[37]) );
  OR U7000 ( .A(n6663), .B(n6662), .Z(n6667) );
  OR U7001 ( .A(n6665), .B(n6664), .Z(n6666) );
  AND U7002 ( .A(n6667), .B(n6666), .Z(n6669) );
  NANDN U7003 ( .A(n525), .B(n[38]), .Z(n6668) );
  XNOR U7004 ( .A(n6669), .B(n6668), .Z(n6670) );
  XNOR U7005 ( .A(n6671), .B(n6670), .Z(zout[38]) );
  AND U7006 ( .A(n6814), .B(n[39]), .Z(n6680) );
  XNOR U7007 ( .A(n6679), .B(n6680), .Z(n6677) );
  NOR U7008 ( .A(n525), .B(n6672), .Z(n6678) );
  XOR U7009 ( .A(n6677), .B(n6678), .Z(zout[39]) );
  XOR U7010 ( .A(n[3]), .B(n6673), .Z(n6674) );
  NANDN U7011 ( .A(n525), .B(n6674), .Z(n6675) );
  XOR U7012 ( .A(n6676), .B(n6675), .Z(zout[3]) );
  OR U7013 ( .A(n6678), .B(n6677), .Z(n6682) );
  OR U7014 ( .A(n6680), .B(n6679), .Z(n6681) );
  AND U7015 ( .A(n6682), .B(n6681), .Z(n6684) );
  NANDN U7016 ( .A(n525), .B(n[40]), .Z(n6683) );
  XNOR U7017 ( .A(n6684), .B(n6683), .Z(n6685) );
  XNOR U7018 ( .A(n6686), .B(n6685), .Z(zout[40]) );
  AND U7019 ( .A(n6814), .B(n[41]), .Z(n6691) );
  XNOR U7020 ( .A(n6690), .B(n6691), .Z(n6688) );
  NOR U7021 ( .A(n525), .B(n6687), .Z(n6689) );
  XOR U7022 ( .A(n6688), .B(n6689), .Z(zout[41]) );
  OR U7023 ( .A(n6689), .B(n6688), .Z(n6693) );
  OR U7024 ( .A(n6691), .B(n6690), .Z(n6692) );
  AND U7025 ( .A(n6693), .B(n6692), .Z(n6695) );
  NANDN U7026 ( .A(n525), .B(n[42]), .Z(n6694) );
  XNOR U7027 ( .A(n6695), .B(n6694), .Z(n6696) );
  XNOR U7028 ( .A(n6697), .B(n6696), .Z(zout[42]) );
  XOR U7029 ( .A(n[43]), .B(n6698), .Z(n6699) );
  NANDN U7030 ( .A(n525), .B(n6699), .Z(n6700) );
  XOR U7031 ( .A(n6701), .B(n6700), .Z(zout[43]) );
  XOR U7032 ( .A(n[44]), .B(n6702), .Z(n6703) );
  NANDN U7033 ( .A(n525), .B(n6703), .Z(n6704) );
  XOR U7034 ( .A(n6705), .B(n6704), .Z(zout[44]) );
  XNOR U7035 ( .A(n[45]), .B(n6706), .Z(n6707) );
  NANDN U7036 ( .A(n525), .B(n6707), .Z(n6708) );
  XOR U7037 ( .A(n6709), .B(n6708), .Z(zout[45]) );
  XNOR U7038 ( .A(n6711), .B(n6710), .Z(n6712) );
  NANDN U7039 ( .A(n525), .B(n6712), .Z(n6713) );
  XOR U7040 ( .A(n6714), .B(n6713), .Z(zout[46]) );
  XNOR U7041 ( .A(n6716), .B(n6715), .Z(n6717) );
  NANDN U7042 ( .A(n525), .B(n6717), .Z(n6718) );
  XOR U7043 ( .A(n6719), .B(n6718), .Z(zout[47]) );
  XNOR U7044 ( .A(n6721), .B(n6720), .Z(zout[48]) );
  XOR U7045 ( .A(n6723), .B(n6722), .Z(n6724) );
  XNOR U7046 ( .A(n6725), .B(n6724), .Z(zout[49]) );
  XNOR U7047 ( .A(n[4]), .B(n6726), .Z(n6727) );
  NANDN U7048 ( .A(n525), .B(n6727), .Z(n6728) );
  XOR U7049 ( .A(n6729), .B(n6728), .Z(zout[4]) );
  XOR U7050 ( .A(n6731), .B(n6730), .Z(n6732) );
  XNOR U7051 ( .A(n6733), .B(n6732), .Z(zout[50]) );
  XNOR U7052 ( .A(n6735), .B(n6734), .Z(zout[51]) );
  XNOR U7053 ( .A(n6737), .B(n6736), .Z(zout[52]) );
  XOR U7054 ( .A(n6739), .B(n6738), .Z(n6740) );
  XNOR U7055 ( .A(n6741), .B(n6740), .Z(zout[53]) );
  XOR U7056 ( .A(n6743), .B(n6742), .Z(zout[54]) );
  XNOR U7057 ( .A(n6745), .B(n6744), .Z(zout[55]) );
  XNOR U7058 ( .A(n6747), .B(n6746), .Z(zout[56]) );
  XNOR U7059 ( .A(n6749), .B(n6748), .Z(zout[57]) );
  XNOR U7060 ( .A(n6751), .B(n6750), .Z(zout[58]) );
  XNOR U7061 ( .A(n6753), .B(n6752), .Z(zout[59]) );
  AND U7062 ( .A(n[5]), .B(n6814), .Z(n6782) );
  XNOR U7063 ( .A(n6781), .B(n6782), .Z(n6779) );
  NOR U7064 ( .A(n525), .B(n6754), .Z(n6780) );
  XOR U7065 ( .A(n6779), .B(n6780), .Z(zout[5]) );
  XNOR U7066 ( .A(n6756), .B(n6755), .Z(zout[60]) );
  XNOR U7067 ( .A(n6758), .B(n6757), .Z(zout[61]) );
  XNOR U7068 ( .A(n6760), .B(n6759), .Z(zout[62]) );
  XOR U7069 ( .A(n6762), .B(n6761), .Z(zout[63]) );
  XNOR U7070 ( .A(n6764), .B(n6763), .Z(zout[64]) );
  XNOR U7071 ( .A(n6766), .B(n6765), .Z(zout[65]) );
  XOR U7072 ( .A(n6768), .B(n6767), .Z(n6769) );
  XNOR U7073 ( .A(n6770), .B(n6769), .Z(zout[66]) );
  XOR U7074 ( .A(n6772), .B(n6771), .Z(zout[67]) );
  XOR U7075 ( .A(n6774), .B(n6773), .Z(n6775) );
  XNOR U7076 ( .A(n6776), .B(n6775), .Z(zout[68]) );
  XOR U7077 ( .A(n6778), .B(n6777), .Z(zout[69]) );
  OR U7078 ( .A(n6780), .B(n6779), .Z(n6784) );
  OR U7079 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U7080 ( .A(n6784), .B(n6783), .Z(n6786) );
  NANDN U7081 ( .A(n525), .B(n[6]), .Z(n6785) );
  XNOR U7082 ( .A(n6786), .B(n6785), .Z(n6787) );
  XNOR U7083 ( .A(n6788), .B(n6787), .Z(zout[6]) );
  XOR U7084 ( .A(n6790), .B(n6789), .Z(zout[70]) );
  XNOR U7085 ( .A(n6792), .B(n6791), .Z(zout[71]) );
  XNOR U7086 ( .A(n6794), .B(n6793), .Z(zout[72]) );
  XNOR U7087 ( .A(n6796), .B(n6795), .Z(zout[73]) );
  XNOR U7088 ( .A(n6798), .B(n6797), .Z(zout[74]) );
  XOR U7089 ( .A(n6800), .B(n6799), .Z(zout[75]) );
  XNOR U7090 ( .A(n6802), .B(n6801), .Z(zout[76]) );
  XOR U7091 ( .A(n6804), .B(n6803), .Z(n6805) );
  XNOR U7092 ( .A(n6806), .B(n6805), .Z(zout[77]) );
  XNOR U7093 ( .A(n6808), .B(n6807), .Z(zout[78]) );
  XOR U7094 ( .A(n6810), .B(n6809), .Z(n6811) );
  XNOR U7095 ( .A(n6812), .B(n6811), .Z(zout[79]) );
  NOR U7096 ( .A(n525), .B(n6813), .Z(n6838) );
  XNOR U7097 ( .A(n6837), .B(n6838), .Z(n6835) );
  AND U7098 ( .A(n6814), .B(n[7]), .Z(n6836) );
  XOR U7099 ( .A(n6835), .B(n6836), .Z(zout[7]) );
  XNOR U7100 ( .A(n6816), .B(n6815), .Z(zout[80]) );
  XNOR U7101 ( .A(n6818), .B(n6817), .Z(zout[81]) );
  XNOR U7102 ( .A(n6820), .B(n6819), .Z(zout[82]) );
  XNOR U7103 ( .A(n6822), .B(n6821), .Z(zout[83]) );
  XNOR U7104 ( .A(n6824), .B(n6823), .Z(zout[84]) );
  XOR U7105 ( .A(n6826), .B(n6825), .Z(zout[85]) );
  XNOR U7106 ( .A(n6828), .B(n6827), .Z(zout[86]) );
  XNOR U7107 ( .A(n6830), .B(n6829), .Z(zout[87]) );
  XOR U7108 ( .A(n6832), .B(n6831), .Z(zout[88]) );
  XNOR U7109 ( .A(n6834), .B(n6833), .Z(zout[89]) );
  OR U7110 ( .A(n6836), .B(n6835), .Z(n6840) );
  OR U7111 ( .A(n6838), .B(n6837), .Z(n6839) );
  AND U7112 ( .A(n6840), .B(n6839), .Z(n6842) );
  NANDN U7113 ( .A(n525), .B(n[8]), .Z(n6841) );
  XNOR U7114 ( .A(n6842), .B(n6841), .Z(n6843) );
  XNOR U7115 ( .A(n6844), .B(n6843), .Z(zout[8]) );
  XNOR U7116 ( .A(n6846), .B(n6845), .Z(zout[90]) );
  XNOR U7117 ( .A(n6848), .B(n6847), .Z(zout[91]) );
  XNOR U7118 ( .A(n6850), .B(n6849), .Z(zout[92]) );
  XNOR U7119 ( .A(n6852), .B(n6851), .Z(zout[93]) );
  XNOR U7120 ( .A(n6854), .B(n6853), .Z(zout[94]) );
  XOR U7121 ( .A(n6856), .B(n6855), .Z(zout[95]) );
  XNOR U7122 ( .A(n6858), .B(n6857), .Z(zout[96]) );
  XOR U7123 ( .A(n6860), .B(n6859), .Z(n6861) );
  XNOR U7124 ( .A(n6862), .B(n6861), .Z(zout[97]) );
  XOR U7125 ( .A(n6864), .B(n6863), .Z(zout[98]) );
  XOR U7126 ( .A(n6866), .B(n6865), .Z(zout[99]) );
  XNOR U7127 ( .A(n6868), .B(n6867), .Z(n6869) );
  NANDN U7128 ( .A(n525), .B(n6869), .Z(n6870) );
  XOR U7129 ( .A(n6871), .B(n6870), .Z(zout[9]) );
endmodule


module modmult_step_N256_0 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N4, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871;
  assign N4 = y[0];

  NAND U2 ( .A(n[100]), .B(n3946), .Z(n1) );
  XOR U3 ( .A(n3946), .B(n[100]), .Z(n2) );
  NANDN U4 ( .A(n5344), .B(n3950), .Z(n3) );
  XOR U5 ( .A(n3950), .B(n[99]), .Z(n4) );
  NAND U6 ( .A(n[98]), .B(n3954), .Z(n5) );
  XOR U7 ( .A(n3954), .B(n[98]), .Z(n6) );
  NAND U8 ( .A(n[97]), .B(n3958), .Z(n7) );
  XOR U9 ( .A(n3958), .B(n[97]), .Z(n8) );
  XNOR U10 ( .A(n3962), .B(n3963), .Z(n9) );
  NAND U11 ( .A(n9), .B(n2322), .Z(n10) );
  NAND U12 ( .A(n10), .B(n3087), .Z(n11) );
  NAND U13 ( .A(n8), .B(n11), .Z(n12) );
  NAND U14 ( .A(n7), .B(n12), .Z(n13) );
  NAND U15 ( .A(n6), .B(n13), .Z(n14) );
  NAND U16 ( .A(n5), .B(n14), .Z(n15) );
  NAND U17 ( .A(n4), .B(n15), .Z(n16) );
  NAND U18 ( .A(n3), .B(n16), .Z(n17) );
  NAND U19 ( .A(n2), .B(n17), .Z(n18) );
  NAND U20 ( .A(n1), .B(n18), .Z(n2323) );
  XOR U21 ( .A(n3377), .B(n3374), .Z(n19) );
  NAND U22 ( .A(n19), .B(n[240]), .Z(n20) );
  NAND U23 ( .A(n3377), .B(n3374), .Z(n21) );
  AND U24 ( .A(n20), .B(n21), .Z(n3370) );
  NAND U25 ( .A(n6449), .B(n3387), .Z(n22) );
  XOR U26 ( .A(n3387), .B(n6449), .Z(n23) );
  NANDN U27 ( .A(n3390), .B(n23), .Z(n24) );
  NAND U28 ( .A(n22), .B(n24), .Z(n5257) );
  XOR U29 ( .A(n3781), .B(n[137]), .Z(n25) );
  NANDN U30 ( .A(n3778), .B(n25), .Z(n26) );
  NAND U31 ( .A(n3781), .B(n[137]), .Z(n27) );
  AND U32 ( .A(n26), .B(n27), .Z(n3774) );
  XOR U33 ( .A(n3503), .B(n3500), .Z(n28) );
  NAND U34 ( .A(n28), .B(n[207]), .Z(n29) );
  NAND U35 ( .A(n3503), .B(n3500), .Z(n30) );
  AND U36 ( .A(n29), .B(n30), .Z(n3495) );
  NAND U37 ( .A(n3399), .B(n3395), .Z(n31) );
  XOR U38 ( .A(n3395), .B(n3399), .Z(n32) );
  NANDN U39 ( .A(n2872), .B(n32), .Z(n33) );
  NAND U40 ( .A(n31), .B(n33), .Z(n3391) );
  XOR U41 ( .A(n5233), .B(n[230]), .Z(n34) );
  NANDN U42 ( .A(n5230), .B(n34), .Z(n35) );
  NAND U43 ( .A(n5233), .B(n[230]), .Z(n36) );
  AND U44 ( .A(n35), .B(n36), .Z(n3408) );
  XOR U45 ( .A(n3427), .B(n3424), .Z(n37) );
  NAND U46 ( .A(n37), .B(n[226]), .Z(n38) );
  NAND U47 ( .A(n3427), .B(n3424), .Z(n39) );
  AND U48 ( .A(n38), .B(n39), .Z(n3420) );
  XOR U49 ( .A(n3447), .B(n[221]), .Z(n40) );
  NANDN U50 ( .A(n3444), .B(n40), .Z(n41) );
  NAND U51 ( .A(n3447), .B(n[221]), .Z(n42) );
  AND U52 ( .A(n41), .B(n42), .Z(n3440) );
  XOR U53 ( .A(n3463), .B(n[216]), .Z(n43) );
  NANDN U54 ( .A(n3460), .B(n43), .Z(n44) );
  NAND U55 ( .A(n3463), .B(n[216]), .Z(n45) );
  AND U56 ( .A(n44), .B(n45), .Z(n5175) );
  NAND U57 ( .A(n6268), .B(n3485), .Z(n46) );
  XOR U58 ( .A(n3485), .B(n6268), .Z(n47) );
  NANDN U59 ( .A(n2874), .B(n47), .Z(n48) );
  NAND U60 ( .A(n46), .B(n48), .Z(n3481) );
  XOR U61 ( .A(n3542), .B(n[198]), .Z(n49) );
  NANDN U62 ( .A(n3539), .B(n49), .Z(n50) );
  NAND U63 ( .A(n3542), .B(n[198]), .Z(n51) );
  AND U64 ( .A(n50), .B(n51), .Z(n3534) );
  XOR U65 ( .A(n3560), .B(n[194]), .Z(n52) );
  NANDN U66 ( .A(n3557), .B(n52), .Z(n53) );
  NAND U67 ( .A(n3560), .B(n[194]), .Z(n54) );
  AND U68 ( .A(n53), .B(n54), .Z(n3551) );
  XOR U69 ( .A(n3615), .B(n[180]), .Z(n55) );
  NANDN U70 ( .A(n3612), .B(n55), .Z(n56) );
  NAND U71 ( .A(n3615), .B(n[180]), .Z(n57) );
  AND U72 ( .A(n56), .B(n57), .Z(n3608) );
  XOR U73 ( .A(n3685), .B(n[163]), .Z(n58) );
  NANDN U74 ( .A(n3682), .B(n58), .Z(n59) );
  NAND U75 ( .A(n3685), .B(n[163]), .Z(n60) );
  AND U76 ( .A(n59), .B(n60), .Z(n3678) );
  XOR U77 ( .A(n3764), .B(n3761), .Z(n61) );
  NAND U78 ( .A(n61), .B(n[141]), .Z(n62) );
  NAND U79 ( .A(n3764), .B(n3761), .Z(n63) );
  AND U80 ( .A(n62), .B(n63), .Z(n3757) );
  XOR U81 ( .A(n3785), .B(n[136]), .Z(n64) );
  NANDN U82 ( .A(n3782), .B(n64), .Z(n65) );
  NAND U83 ( .A(n3785), .B(n[136]), .Z(n66) );
  AND U84 ( .A(n65), .B(n66), .Z(n3778) );
  XOR U85 ( .A(n3920), .B(n[106]), .Z(n67) );
  NANDN U86 ( .A(n3917), .B(n67), .Z(n68) );
  NAND U87 ( .A(n3920), .B(n[106]), .Z(n69) );
  AND U88 ( .A(n68), .B(n69), .Z(n3913) );
  XOR U89 ( .A(n4010), .B(n[84]), .Z(n70) );
  NANDN U90 ( .A(n4007), .B(n70), .Z(n71) );
  NAND U91 ( .A(n4010), .B(n[84]), .Z(n72) );
  AND U92 ( .A(n71), .B(n72), .Z(n4003) );
  XOR U93 ( .A(n4032), .B(n[79]), .Z(n73) );
  NANDN U94 ( .A(n4029), .B(n73), .Z(n74) );
  NAND U95 ( .A(n4032), .B(n[79]), .Z(n75) );
  AND U96 ( .A(n74), .B(n75), .Z(n4024) );
  XOR U97 ( .A(n3365), .B(n[243]), .Z(n76) );
  NANDN U98 ( .A(n3362), .B(n76), .Z(n77) );
  NAND U99 ( .A(n3365), .B(n[243]), .Z(n78) );
  AND U100 ( .A(n77), .B(n78), .Z(n3357) );
  XOR U101 ( .A(n3386), .B(n[238]), .Z(n79) );
  NANDN U102 ( .A(n3383), .B(n79), .Z(n80) );
  NAND U103 ( .A(n3386), .B(n[238]), .Z(n81) );
  AND U104 ( .A(n80), .B(n81), .Z(n3378) );
  XOR U105 ( .A(n3512), .B(n[205]), .Z(n82) );
  NANDN U106 ( .A(n3509), .B(n82), .Z(n83) );
  NAND U107 ( .A(n3512), .B(n[205]), .Z(n84) );
  AND U108 ( .A(n83), .B(n84), .Z(n3504) );
  XOR U109 ( .A(n3726), .B(n[150]), .Z(n85) );
  NANDN U110 ( .A(n3723), .B(n85), .Z(n86) );
  NAND U111 ( .A(n3726), .B(n[150]), .Z(n87) );
  AND U112 ( .A(n86), .B(n87), .Z(n3719) );
  NAND U113 ( .A(n5344), .B(n3947), .Z(n88) );
  XOR U114 ( .A(n3947), .B(n5344), .Z(n89) );
  NANDN U115 ( .A(n3950), .B(n89), .Z(n90) );
  NAND U116 ( .A(n88), .B(n90), .Z(n3943) );
  XOR U117 ( .A(n3331), .B(n[251]), .Z(n91) );
  NANDN U118 ( .A(n3328), .B(n91), .Z(n92) );
  NAND U119 ( .A(n3331), .B(n[251]), .Z(n93) );
  AND U120 ( .A(n92), .B(n93), .Z(n3323) );
  XOR U121 ( .A(n6436), .B(n6435), .Z(n94) );
  NANDN U122 ( .A(n6434), .B(n94), .Z(n95) );
  NAND U123 ( .A(n6436), .B(n6435), .Z(n96) );
  AND U124 ( .A(n95), .B(n96), .Z(n6438) );
  XOR U125 ( .A(n5924), .B(n5925), .Z(n97) );
  NANDN U126 ( .A(n5923), .B(n97), .Z(n98) );
  NAND U127 ( .A(n5924), .B(n5925), .Z(n99) );
  AND U128 ( .A(n98), .B(n99), .Z(n5927) );
  NAND U129 ( .A(n5621), .B(n5620), .Z(n100) );
  XOR U130 ( .A(n5620), .B(n5621), .Z(n101) );
  NANDN U131 ( .A(n5622), .B(n101), .Z(n102) );
  NAND U132 ( .A(n100), .B(n102), .Z(n5624) );
  XOR U133 ( .A(n4209), .B(n[34]), .Z(n103) );
  NANDN U134 ( .A(n4206), .B(n103), .Z(n104) );
  NAND U135 ( .A(n4209), .B(n[34]), .Z(n105) );
  AND U136 ( .A(n104), .B(n105), .Z(n4428) );
  NAND U137 ( .A(n4399), .B(n4398), .Z(n106) );
  XOR U138 ( .A(n4398), .B(n4399), .Z(n107) );
  NANDN U139 ( .A(n2879), .B(n107), .Z(n108) );
  NAND U140 ( .A(n106), .B(n108), .Z(n4403) );
  NAND U141 ( .A(n[1]), .B(n4296), .Z(n109) );
  XOR U142 ( .A(n4296), .B(n[1]), .Z(n110) );
  NANDN U143 ( .A(n4299), .B(n110), .Z(n111) );
  NAND U144 ( .A(n109), .B(n111), .Z(n4300) );
  XOR U145 ( .A(n[3]), .B(n6676), .Z(n112) );
  NAND U146 ( .A(n112), .B(n6673), .Z(n113) );
  NAND U147 ( .A(n[3]), .B(n6676), .Z(n114) );
  AND U148 ( .A(n113), .B(n114), .Z(n6726) );
  XOR U149 ( .A(n4073), .B(n[69]), .Z(n115) );
  NANDN U150 ( .A(n4070), .B(n115), .Z(n116) );
  NAND U151 ( .A(n4073), .B(n[69]), .Z(n117) );
  AND U152 ( .A(n116), .B(n117), .Z(n4066) );
  XOR U153 ( .A(n3415), .B(n[229]), .Z(n118) );
  NANDN U154 ( .A(n3412), .B(n118), .Z(n119) );
  NAND U155 ( .A(n3415), .B(n[229]), .Z(n120) );
  AND U156 ( .A(n119), .B(n120), .Z(n5230) );
  XOR U157 ( .A(n3435), .B(n[224]), .Z(n121) );
  NANDN U158 ( .A(n3432), .B(n121), .Z(n122) );
  NAND U159 ( .A(n3435), .B(n[224]), .Z(n123) );
  AND U160 ( .A(n122), .B(n123), .Z(n3428) );
  XOR U161 ( .A(n3451), .B(n[220]), .Z(n124) );
  NANDN U162 ( .A(n3448), .B(n124), .Z(n125) );
  NAND U163 ( .A(n3451), .B(n[220]), .Z(n126) );
  AND U164 ( .A(n125), .B(n126), .Z(n3444) );
  XOR U165 ( .A(n5178), .B(n[217]), .Z(n127) );
  NANDN U166 ( .A(n5175), .B(n127), .Z(n128) );
  NAND U167 ( .A(n5178), .B(n[217]), .Z(n129) );
  AND U168 ( .A(n128), .B(n129), .Z(n3456) );
  XOR U169 ( .A(n3471), .B(n3468), .Z(n130) );
  NAND U170 ( .A(n130), .B(n[214]), .Z(n131) );
  NAND U171 ( .A(n3471), .B(n3468), .Z(n132) );
  AND U172 ( .A(n131), .B(n132), .Z(n3464) );
  XOR U173 ( .A(n3546), .B(n[197]), .Z(n133) );
  NANDN U174 ( .A(n3543), .B(n133), .Z(n134) );
  NAND U175 ( .A(n3546), .B(n[197]), .Z(n135) );
  AND U176 ( .A(n134), .B(n135), .Z(n3539) );
  XOR U177 ( .A(n3564), .B(n[193]), .Z(n136) );
  NANDN U178 ( .A(n3561), .B(n136), .Z(n137) );
  NAND U179 ( .A(n3564), .B(n[193]), .Z(n138) );
  AND U180 ( .A(n137), .B(n138), .Z(n3557) );
  XOR U181 ( .A(n3577), .B(n2875), .Z(n139) );
  NANDN U182 ( .A(n3581), .B(n139), .Z(n140) );
  NAND U183 ( .A(n3577), .B(n2875), .Z(n141) );
  AND U184 ( .A(n140), .B(n141), .Z(n3573) );
  XOR U185 ( .A(n5054), .B(n5051), .Z(n142) );
  NAND U186 ( .A(n142), .B(n[185]), .Z(n143) );
  NAND U187 ( .A(n5054), .B(n5051), .Z(n144) );
  AND U188 ( .A(n143), .B(n144), .Z(n3591) );
  XOR U189 ( .A(n3607), .B(n[182]), .Z(n145) );
  NANDN U190 ( .A(n3604), .B(n145), .Z(n146) );
  NAND U191 ( .A(n3607), .B(n[182]), .Z(n147) );
  AND U192 ( .A(n146), .B(n147), .Z(n3599) );
  XOR U193 ( .A(n5026), .B(n[179]), .Z(n148) );
  NANDN U194 ( .A(n5023), .B(n148), .Z(n149) );
  NAND U195 ( .A(n5026), .B(n[179]), .Z(n150) );
  AND U196 ( .A(n149), .B(n150), .Z(n3612) );
  XOR U197 ( .A(n3625), .B(n3628), .Z(n151) );
  NANDN U198 ( .A(n6025), .B(n151), .Z(n152) );
  NAND U199 ( .A(n3625), .B(n3628), .Z(n153) );
  AND U200 ( .A(n152), .B(n153), .Z(n3620) );
  XOR U201 ( .A(n3693), .B(n3690), .Z(n154) );
  NAND U202 ( .A(n154), .B(n[161]), .Z(n155) );
  NAND U203 ( .A(n3693), .B(n3690), .Z(n156) );
  AND U204 ( .A(n155), .B(n156), .Z(n3686) );
  XOR U205 ( .A(n3743), .B(n3740), .Z(n157) );
  NAND U206 ( .A(n157), .B(n[146]), .Z(n158) );
  NAND U207 ( .A(n3743), .B(n3740), .Z(n159) );
  AND U208 ( .A(n158), .B(n159), .Z(n3735) );
  XOR U209 ( .A(n3793), .B(n3790), .Z(n160) );
  NAND U210 ( .A(n160), .B(n[134]), .Z(n161) );
  NAND U211 ( .A(n3793), .B(n3790), .Z(n162) );
  AND U212 ( .A(n161), .B(n162), .Z(n3786) );
  XOR U213 ( .A(n3823), .B(n[127]), .Z(n163) );
  NANDN U214 ( .A(n3820), .B(n163), .Z(n164) );
  NAND U215 ( .A(n3823), .B(n[127]), .Z(n165) );
  AND U216 ( .A(n164), .B(n165), .Z(n3816) );
  XOR U217 ( .A(n3916), .B(n[107]), .Z(n166) );
  NANDN U218 ( .A(n3913), .B(n166), .Z(n167) );
  NAND U219 ( .A(n3916), .B(n[107]), .Z(n168) );
  AND U220 ( .A(n167), .B(n168), .Z(n3908) );
  XOR U221 ( .A(n3928), .B(n3925), .Z(n169) );
  NAND U222 ( .A(n169), .B(n[104]), .Z(n170) );
  NAND U223 ( .A(n3928), .B(n3925), .Z(n171) );
  AND U224 ( .A(n170), .B(n171), .Z(n3921) );
  XOR U225 ( .A(n3993), .B(n3990), .Z(n172) );
  NAND U226 ( .A(n172), .B(n[88]), .Z(n173) );
  NAND U227 ( .A(n3993), .B(n3990), .Z(n174) );
  AND U228 ( .A(n173), .B(n174), .Z(n3986) );
  XOR U229 ( .A(n4014), .B(n[83]), .Z(n175) );
  NANDN U230 ( .A(n4011), .B(n175), .Z(n176) );
  NAND U231 ( .A(n4014), .B(n[83]), .Z(n177) );
  AND U232 ( .A(n176), .B(n177), .Z(n4007) );
  XOR U233 ( .A(n4057), .B(n[73]), .Z(n178) );
  NANDN U234 ( .A(n4054), .B(n178), .Z(n179) );
  NAND U235 ( .A(n4057), .B(n[73]), .Z(n180) );
  AND U236 ( .A(n179), .B(n180), .Z(n4050) );
  ANDN U237 ( .B(n[46]), .A(n4174), .Z(n2989) );
  XOR U238 ( .A(n3343), .B(n3340), .Z(n181) );
  NAND U239 ( .A(n181), .B(n[248]), .Z(n182) );
  NAND U240 ( .A(n3343), .B(n3340), .Z(n183) );
  AND U241 ( .A(n182), .B(n183), .Z(n3336) );
  XOR U242 ( .A(n3373), .B(n[241]), .Z(n184) );
  NANDN U243 ( .A(n3370), .B(n184), .Z(n185) );
  NAND U244 ( .A(n3373), .B(n[241]), .Z(n186) );
  AND U245 ( .A(n185), .B(n186), .Z(n3366) );
  NAND U246 ( .A(n6456), .B(n5257), .Z(n187) );
  XOR U247 ( .A(n5257), .B(n6456), .Z(n188) );
  NANDN U248 ( .A(n5260), .B(n188), .Z(n189) );
  NAND U249 ( .A(n187), .B(n189), .Z(n3383) );
  XOR U250 ( .A(n3403), .B(n[233]), .Z(n190) );
  NANDN U251 ( .A(n3400), .B(n190), .Z(n191) );
  NAND U252 ( .A(n3403), .B(n[233]), .Z(n192) );
  AND U253 ( .A(n191), .B(n192), .Z(n3395) );
  XOR U254 ( .A(n3484), .B(n[211]), .Z(n193) );
  NANDN U255 ( .A(n3481), .B(n193), .Z(n194) );
  NAND U256 ( .A(n3484), .B(n[211]), .Z(n195) );
  AND U257 ( .A(n194), .B(n195), .Z(n3477) );
  XOR U258 ( .A(n3516), .B(n3513), .Z(n196) );
  NAND U259 ( .A(n196), .B(n[204]), .Z(n197) );
  NAND U260 ( .A(n3516), .B(n3513), .Z(n198) );
  AND U261 ( .A(n197), .B(n198), .Z(n3509) );
  XOR U262 ( .A(n3659), .B(n3656), .Z(n199) );
  NAND U263 ( .A(n199), .B(n[169]), .Z(n200) );
  NAND U264 ( .A(n3659), .B(n3656), .Z(n201) );
  AND U265 ( .A(n200), .B(n201), .Z(n3651) );
  XOR U266 ( .A(n3730), .B(n[149]), .Z(n202) );
  NANDN U267 ( .A(n3727), .B(n202), .Z(n203) );
  NAND U268 ( .A(n3730), .B(n[149]), .Z(n204) );
  AND U269 ( .A(n203), .B(n204), .Z(n3723) );
  XOR U270 ( .A(n3777), .B(n[138]), .Z(n205) );
  NANDN U271 ( .A(n3774), .B(n205), .Z(n206) );
  NAND U272 ( .A(n3777), .B(n[138]), .Z(n207) );
  AND U273 ( .A(n206), .B(n207), .Z(n3770) );
  XOR U274 ( .A(n3836), .B(n3833), .Z(n208) );
  NAND U275 ( .A(n208), .B(n[124]), .Z(n209) );
  NAND U276 ( .A(n3836), .B(n3833), .Z(n210) );
  AND U277 ( .A(n209), .B(n210), .Z(n3828) );
  XOR U278 ( .A(n3946), .B(n[100]), .Z(n211) );
  NANDN U279 ( .A(n3943), .B(n211), .Z(n212) );
  NAND U280 ( .A(n3946), .B(n[100]), .Z(n213) );
  AND U281 ( .A(n212), .B(n213), .Z(n3938) );
  XOR U282 ( .A(n3958), .B(n3955), .Z(n214) );
  NAND U283 ( .A(n214), .B(n[97]), .Z(n215) );
  NAND U284 ( .A(n3958), .B(n3955), .Z(n216) );
  AND U285 ( .A(n215), .B(n216), .Z(n3951) );
  XOR U286 ( .A(n4045), .B(n[76]), .Z(n217) );
  NANDN U287 ( .A(n4042), .B(n217), .Z(n218) );
  NAND U288 ( .A(n4045), .B(n[76]), .Z(n219) );
  AND U289 ( .A(n218), .B(n219), .Z(n4037) );
  XOR U290 ( .A(n6776), .B(n6773), .Z(n220) );
  NANDN U291 ( .A(n6774), .B(n220), .Z(n221) );
  NAND U292 ( .A(n6776), .B(n6773), .Z(n222) );
  AND U293 ( .A(n221), .B(n222), .Z(n6778) );
  XOR U294 ( .A(n4086), .B(n[66]), .Z(n223) );
  NAND U295 ( .A(n223), .B(n4083), .Z(n224) );
  NAND U296 ( .A(n4086), .B(n[66]), .Z(n225) );
  AND U297 ( .A(n224), .B(n225), .Z(n4079) );
  XOR U298 ( .A(n3322), .B(n3319), .Z(n226) );
  NAND U299 ( .A(n226), .B(n[253]), .Z(n227) );
  NAND U300 ( .A(n3322), .B(n3319), .Z(n228) );
  AND U301 ( .A(n227), .B(n228), .Z(n3315) );
  NAND U302 ( .A(n6250), .B(n6251), .Z(n229) );
  XOR U303 ( .A(n6251), .B(n6250), .Z(n230) );
  NANDN U304 ( .A(n6249), .B(n230), .Z(n231) );
  NAND U305 ( .A(n229), .B(n231), .Z(n6253) );
  XOR U306 ( .A(n5881), .B(n5880), .Z(n232) );
  NANDN U307 ( .A(n5879), .B(n232), .Z(n233) );
  NAND U308 ( .A(n5881), .B(n5880), .Z(n234) );
  AND U309 ( .A(n233), .B(n234), .Z(n5885) );
  NAND U310 ( .A(n5796), .B(n5797), .Z(n235) );
  XOR U311 ( .A(n5797), .B(n5796), .Z(n236) );
  NANDN U312 ( .A(n5798), .B(n236), .Z(n237) );
  NAND U313 ( .A(n235), .B(n237), .Z(n5803) );
  XOR U314 ( .A(n6810), .B(n6812), .Z(n238) );
  NAND U315 ( .A(n238), .B(n6809), .Z(n239) );
  NAND U316 ( .A(n6810), .B(n6812), .Z(n240) );
  AND U317 ( .A(n239), .B(n240), .Z(n6816) );
  NAND U318 ( .A(n6723), .B(n6725), .Z(n241) );
  XOR U319 ( .A(n6725), .B(n6723), .Z(n242) );
  NAND U320 ( .A(n242), .B(n6722), .Z(n243) );
  NAND U321 ( .A(n241), .B(n243), .Z(n6730) );
  NAND U322 ( .A(n4432), .B(n4428), .Z(n244) );
  XOR U323 ( .A(n4428), .B(n4432), .Z(n245) );
  NANDN U324 ( .A(n4431), .B(n245), .Z(n246) );
  NAND U325 ( .A(n244), .B(n246), .Z(n4202) );
  XOR U326 ( .A(n4217), .B(n4214), .Z(n247) );
  NAND U327 ( .A(n247), .B(n[32]), .Z(n248) );
  NAND U328 ( .A(n4217), .B(n4214), .Z(n249) );
  AND U329 ( .A(n248), .B(n249), .Z(n4210) );
  XOR U330 ( .A(n[28]), .B(n6613), .Z(n250) );
  NAND U331 ( .A(n250), .B(n6610), .Z(n251) );
  NAND U332 ( .A(n[28]), .B(n6613), .Z(n252) );
  AND U333 ( .A(n251), .B(n252), .Z(n6614) );
  XOR U334 ( .A(n4230), .B(n[26]), .Z(n253) );
  NANDN U335 ( .A(n4227), .B(n253), .Z(n254) );
  NAND U336 ( .A(n4230), .B(n[26]), .Z(n255) );
  AND U337 ( .A(n254), .B(n255), .Z(n4398) );
  XNOR U338 ( .A(n6544), .B(n4239), .Z(n256) );
  NANDN U339 ( .A(n4387), .B(n6473), .Z(n257) );
  XOR U340 ( .A(n6473), .B(n[23]), .Z(n258) );
  NAND U341 ( .A(n258), .B(n6537), .Z(n259) );
  NAND U342 ( .A(n257), .B(n259), .Z(n260) );
  NAND U343 ( .A(n256), .B(n260), .Z(n261) );
  NANDN U344 ( .A(n4239), .B(n6544), .Z(n262) );
  AND U345 ( .A(n261), .B(n262), .Z(n6595) );
  XNOR U346 ( .A(n5985), .B(n4266), .Z(n263) );
  NANDN U347 ( .A(n4358), .B(n5918), .Z(n264) );
  XOR U348 ( .A(n5918), .B(n[15]), .Z(n265) );
  NAND U349 ( .A(n265), .B(n5978), .Z(n266) );
  NAND U350 ( .A(n264), .B(n266), .Z(n267) );
  NAND U351 ( .A(n263), .B(n267), .Z(n268) );
  NANDN U352 ( .A(n4266), .B(n5985), .Z(n269) );
  AND U353 ( .A(n268), .B(n269), .Z(n6054) );
  NAND U354 ( .A(n5919), .B(n5920), .Z(n270) );
  XOR U355 ( .A(n5920), .B(n5919), .Z(n271) );
  NAND U356 ( .A(n271), .B(n5921), .Z(n272) );
  NAND U357 ( .A(n270), .B(n272), .Z(n5925) );
  NAND U358 ( .A(n5616), .B(n5617), .Z(n273) );
  XOR U359 ( .A(n5617), .B(n5616), .Z(n274) );
  NANDN U360 ( .A(n5618), .B(n274), .Z(n275) );
  NAND U361 ( .A(n273), .B(n275), .Z(n5620) );
  NAND U362 ( .A(n6698), .B(n6701), .Z(n276) );
  XOR U363 ( .A(n6701), .B(n6698), .Z(n277) );
  NANDN U364 ( .A(n4463), .B(n277), .Z(n278) );
  NAND U365 ( .A(n276), .B(n278), .Z(n6702) );
  NAND U366 ( .A(n6615), .B(n6619), .Z(n279) );
  XOR U367 ( .A(n6619), .B(n6615), .Z(n280) );
  NANDN U368 ( .A(n6616), .B(n280), .Z(n281) );
  NAND U369 ( .A(n279), .B(n281), .Z(n6673) );
  XOR U370 ( .A(n3394), .B(n[235]), .Z(n282) );
  NANDN U371 ( .A(n3391), .B(n282), .Z(n283) );
  NAND U372 ( .A(n3394), .B(n[235]), .Z(n284) );
  AND U373 ( .A(n283), .B(n284), .Z(n3387) );
  XOR U374 ( .A(n3423), .B(n[227]), .Z(n285) );
  NANDN U375 ( .A(n3420), .B(n285), .Z(n286) );
  NAND U376 ( .A(n3423), .B(n[227]), .Z(n287) );
  AND U377 ( .A(n286), .B(n287), .Z(n3416) );
  XOR U378 ( .A(n3439), .B(n3436), .Z(n288) );
  NAND U379 ( .A(n288), .B(n[223]), .Z(n289) );
  NAND U380 ( .A(n3439), .B(n3436), .Z(n290) );
  AND U381 ( .A(n289), .B(n290), .Z(n3432) );
  XOR U382 ( .A(n3455), .B(n3452), .Z(n291) );
  NAND U383 ( .A(n291), .B(n[219]), .Z(n292) );
  NAND U384 ( .A(n3455), .B(n3452), .Z(n293) );
  AND U385 ( .A(n292), .B(n293), .Z(n3448) );
  XOR U386 ( .A(n3467), .B(n[215]), .Z(n294) );
  NANDN U387 ( .A(n3464), .B(n294), .Z(n295) );
  NAND U388 ( .A(n3467), .B(n[215]), .Z(n296) );
  AND U389 ( .A(n295), .B(n296), .Z(n3460) );
  XOR U390 ( .A(n3489), .B(n3492), .Z(n297) );
  NANDN U391 ( .A(n6256), .B(n297), .Z(n298) );
  NAND U392 ( .A(n3489), .B(n3492), .Z(n299) );
  AND U393 ( .A(n298), .B(n299), .Z(n3485) );
  XOR U394 ( .A(n3537), .B(n[199]), .Z(n300) );
  NANDN U395 ( .A(n3534), .B(n300), .Z(n301) );
  NAND U396 ( .A(n3537), .B(n[199]), .Z(n302) );
  AND U397 ( .A(n301), .B(n302), .Z(n3530) );
  XOR U398 ( .A(n3547), .B(n3550), .Z(n303) );
  NANDN U399 ( .A(n6166), .B(n303), .Z(n304) );
  NAND U400 ( .A(n3547), .B(n3550), .Z(n305) );
  AND U401 ( .A(n304), .B(n305), .Z(n3543) );
  XOR U402 ( .A(n3568), .B(n3565), .Z(n306) );
  NAND U403 ( .A(n306), .B(n[192]), .Z(n307) );
  NAND U404 ( .A(n3568), .B(n3565), .Z(n308) );
  AND U405 ( .A(n307), .B(n308), .Z(n3561) );
  XOR U406 ( .A(n3611), .B(n[181]), .Z(n309) );
  NANDN U407 ( .A(n3608), .B(n309), .Z(n310) );
  NAND U408 ( .A(n3611), .B(n[181]), .Z(n311) );
  AND U409 ( .A(n310), .B(n311), .Z(n3604) );
  XOR U410 ( .A(n3616), .B(n3619), .Z(n312) );
  NANDN U411 ( .A(n6039), .B(n312), .Z(n313) );
  NAND U412 ( .A(n3616), .B(n3619), .Z(n314) );
  AND U413 ( .A(n313), .B(n314), .Z(n5023) );
  XOR U414 ( .A(n3636), .B(n3633), .Z(n315) );
  NAND U415 ( .A(n315), .B(n[174]), .Z(n316) );
  NAND U416 ( .A(n3636), .B(n3633), .Z(n317) );
  AND U417 ( .A(n316), .B(n317), .Z(n3629) );
  XOR U418 ( .A(n3689), .B(n[162]), .Z(n318) );
  NANDN U419 ( .A(n3686), .B(n318), .Z(n319) );
  NAND U420 ( .A(n3689), .B(n[162]), .Z(n320) );
  AND U421 ( .A(n319), .B(n320), .Z(n3682) );
  XOR U422 ( .A(n4926), .B(n4923), .Z(n321) );
  NAND U423 ( .A(n321), .B(n[155]), .Z(n322) );
  NAND U424 ( .A(n4926), .B(n4923), .Z(n323) );
  AND U425 ( .A(n322), .B(n323), .Z(n3707) );
  XOR U426 ( .A(n3756), .B(n[143]), .Z(n324) );
  NANDN U427 ( .A(n3753), .B(n324), .Z(n325) );
  NAND U428 ( .A(n3756), .B(n[143]), .Z(n326) );
  AND U429 ( .A(n325), .B(n326), .Z(n3748) );
  XOR U430 ( .A(n3789), .B(n[135]), .Z(n327) );
  NANDN U431 ( .A(n3786), .B(n327), .Z(n328) );
  NAND U432 ( .A(n3789), .B(n[135]), .Z(n329) );
  AND U433 ( .A(n328), .B(n329), .Z(n3782) );
  XOR U434 ( .A(n3802), .B(n3799), .Z(n330) );
  NAND U435 ( .A(n330), .B(n[132]), .Z(n331) );
  NAND U436 ( .A(n3802), .B(n3799), .Z(n332) );
  AND U437 ( .A(n331), .B(n332), .Z(n3794) );
  XOR U438 ( .A(n3815), .B(n3812), .Z(n333) );
  NAND U439 ( .A(n333), .B(n[129]), .Z(n334) );
  NAND U440 ( .A(n3815), .B(n3812), .Z(n335) );
  AND U441 ( .A(n334), .B(n335), .Z(n3807) );
  XOR U442 ( .A(n3827), .B(n3824), .Z(n336) );
  NAND U443 ( .A(n336), .B(n[126]), .Z(n337) );
  NAND U444 ( .A(n3827), .B(n3824), .Z(n338) );
  AND U445 ( .A(n337), .B(n338), .Z(n3820) );
  XOR U446 ( .A(n3924), .B(n[105]), .Z(n339) );
  NANDN U447 ( .A(n3921), .B(n339), .Z(n340) );
  NAND U448 ( .A(n3924), .B(n[105]), .Z(n341) );
  AND U449 ( .A(n340), .B(n341), .Z(n3917) );
  XOR U450 ( .A(n3985), .B(n3982), .Z(n342) );
  NAND U451 ( .A(n342), .B(n[90]), .Z(n343) );
  NAND U452 ( .A(n3985), .B(n3982), .Z(n344) );
  AND U453 ( .A(n343), .B(n344), .Z(n3978) );
  XOR U454 ( .A(n4002), .B(n3999), .Z(n345) );
  NAND U455 ( .A(n345), .B(n[86]), .Z(n346) );
  NAND U456 ( .A(n4002), .B(n3999), .Z(n347) );
  AND U457 ( .A(n346), .B(n347), .Z(n3994) );
  XOR U458 ( .A(n4018), .B(n4015), .Z(n348) );
  NAND U459 ( .A(n348), .B(n[82]), .Z(n349) );
  NAND U460 ( .A(n4018), .B(n4015), .Z(n350) );
  AND U461 ( .A(n349), .B(n350), .Z(n4011) );
  XOR U462 ( .A(n4062), .B(n4065), .Z(n351) );
  NANDN U463 ( .A(n5390), .B(n351), .Z(n352) );
  NAND U464 ( .A(n4062), .B(n4065), .Z(n353) );
  AND U465 ( .A(n352), .B(n353), .Z(n4058) );
  NAND U466 ( .A(n[57]), .B(n4126), .Z(n354) );
  XOR U467 ( .A(n4126), .B(n[57]), .Z(n355) );
  NANDN U468 ( .A(n4123), .B(n355), .Z(n356) );
  NAND U469 ( .A(n354), .B(n356), .Z(n4119) );
  XOR U470 ( .A(n3369), .B(n[242]), .Z(n357) );
  NANDN U471 ( .A(n3366), .B(n357), .Z(n358) );
  NAND U472 ( .A(n3369), .B(n[242]), .Z(n359) );
  AND U473 ( .A(n358), .B(n359), .Z(n3362) );
  NANDN U474 ( .A(n6457), .B(n[237]), .Z(n6459) );
  NAND U475 ( .A(n6439), .B(n6438), .Z(n360) );
  XOR U476 ( .A(n6438), .B(n6439), .Z(n361) );
  NANDN U477 ( .A(n6440), .B(n361), .Z(n362) );
  NAND U478 ( .A(n360), .B(n362), .Z(n6445) );
  XOR U479 ( .A(n3480), .B(n[212]), .Z(n363) );
  NANDN U480 ( .A(n3477), .B(n363), .Z(n364) );
  NAND U481 ( .A(n3480), .B(n[212]), .Z(n365) );
  AND U482 ( .A(n364), .B(n365), .Z(n3472) );
  XOR U483 ( .A(n3524), .B(n3521), .Z(n366) );
  NAND U484 ( .A(n366), .B(n[202]), .Z(n367) );
  NAND U485 ( .A(n3524), .B(n3521), .Z(n368) );
  AND U486 ( .A(n367), .B(n368), .Z(n3517) );
  XOR U487 ( .A(n3594), .B(n[186]), .Z(n369) );
  NANDN U488 ( .A(n3591), .B(n369), .Z(n370) );
  NAND U489 ( .A(n3594), .B(n[186]), .Z(n371) );
  AND U490 ( .A(n370), .B(n371), .Z(n3587) );
  XOR U491 ( .A(n3718), .B(n3715), .Z(n372) );
  NAND U492 ( .A(n372), .B(n[152]), .Z(n373) );
  NAND U493 ( .A(n3718), .B(n3715), .Z(n374) );
  AND U494 ( .A(n373), .B(n374), .Z(n4909) );
  XOR U495 ( .A(n3734), .B(n3731), .Z(n375) );
  NAND U496 ( .A(n375), .B(n[148]), .Z(n376) );
  NAND U497 ( .A(n3734), .B(n3731), .Z(n377) );
  AND U498 ( .A(n376), .B(n377), .Z(n3727) );
  XOR U499 ( .A(n3773), .B(n[139]), .Z(n378) );
  NANDN U500 ( .A(n3770), .B(n378), .Z(n379) );
  NAND U501 ( .A(n3773), .B(n[139]), .Z(n380) );
  AND U502 ( .A(n379), .B(n380), .Z(n3765) );
  XOR U503 ( .A(n3937), .B(n3934), .Z(n381) );
  NAND U504 ( .A(n381), .B(n[102]), .Z(n382) );
  NAND U505 ( .A(n3937), .B(n3934), .Z(n383) );
  AND U506 ( .A(n382), .B(n383), .Z(n3929) );
  XOR U507 ( .A(n3954), .B(n[98]), .Z(n384) );
  NANDN U508 ( .A(n3951), .B(n384), .Z(n385) );
  NAND U509 ( .A(n3954), .B(n[98]), .Z(n386) );
  AND U510 ( .A(n385), .B(n386), .Z(n3947) );
  XOR U511 ( .A(n4036), .B(n4033), .Z(n387) );
  NAND U512 ( .A(n387), .B(n[78]), .Z(n388) );
  NAND U513 ( .A(n4036), .B(n4033), .Z(n389) );
  AND U514 ( .A(n388), .B(n389), .Z(n4029) );
  XOR U515 ( .A(n4049), .B(n[75]), .Z(n390) );
  NANDN U516 ( .A(n4046), .B(n390), .Z(n391) );
  NAND U517 ( .A(n4049), .B(n[75]), .Z(n392) );
  AND U518 ( .A(n391), .B(n392), .Z(n4042) );
  XOR U519 ( .A(n4082), .B(n[67]), .Z(n393) );
  NANDN U520 ( .A(n4079), .B(n393), .Z(n394) );
  NAND U521 ( .A(n4082), .B(n[67]), .Z(n395) );
  AND U522 ( .A(n394), .B(n395), .Z(n4074) );
  XOR U523 ( .A(n4099), .B(n4096), .Z(n396) );
  NAND U524 ( .A(n396), .B(n[63]), .Z(n397) );
  NAND U525 ( .A(n4099), .B(n4096), .Z(n398) );
  AND U526 ( .A(n397), .B(n398), .Z(n4092) );
  XOR U527 ( .A(n4153), .B(n4150), .Z(n399) );
  NAND U528 ( .A(n399), .B(n[51]), .Z(n400) );
  NAND U529 ( .A(n4153), .B(n4150), .Z(n401) );
  AND U530 ( .A(n400), .B(n401), .Z(n4146) );
  XOR U531 ( .A(n3335), .B(n3332), .Z(n402) );
  NAND U532 ( .A(n402), .B(n[250]), .Z(n403) );
  NAND U533 ( .A(n3335), .B(n3332), .Z(n404) );
  AND U534 ( .A(n403), .B(n404), .Z(n3328) );
  XNOR U535 ( .A(n6582), .B(n3318), .Z(n405) );
  NAND U536 ( .A(n[253]), .B(n3322), .Z(n406) );
  XOR U537 ( .A(n3322), .B(n[253]), .Z(n407) );
  XNOR U538 ( .A(n3327), .B(n3326), .Z(n408) );
  NAND U539 ( .A(n2856), .B(n2855), .Z(n409) );
  NAND U540 ( .A(n[251]), .B(n3331), .Z(n410) );
  NAND U541 ( .A(n409), .B(n410), .Z(n411) );
  NAND U542 ( .A(n408), .B(n411), .Z(n412) );
  NAND U543 ( .A(n412), .B(n3300), .Z(n413) );
  NAND U544 ( .A(n407), .B(n413), .Z(n414) );
  NAND U545 ( .A(n406), .B(n414), .Z(n415) );
  NAND U546 ( .A(n405), .B(n415), .Z(n416) );
  AND U547 ( .A(n3303), .B(n416), .Z(n417) );
  NANDN U548 ( .A(n417), .B(n3308), .Z(n418) );
  XNOR U549 ( .A(n3308), .B(n417), .Z(n419) );
  NAND U550 ( .A(n419), .B(n[255]), .Z(n420) );
  NAND U551 ( .A(n418), .B(n420), .Z(n421) );
  ANDN U552 ( .B(n421), .A(n3313), .Z(n422) );
  NANDN U553 ( .A(n3312), .B(n422), .Z(n523) );
  XOR U554 ( .A(n6505), .B(n6504), .Z(n423) );
  NANDN U555 ( .A(n6503), .B(n423), .Z(n424) );
  NAND U556 ( .A(n6505), .B(n6504), .Z(n425) );
  AND U557 ( .A(n424), .B(n425), .Z(n6510) );
  XOR U558 ( .A(n6474), .B(n6475), .Z(n426) );
  NAND U559 ( .A(n426), .B(n6476), .Z(n427) );
  NAND U560 ( .A(n6474), .B(n6475), .Z(n428) );
  AND U561 ( .A(n427), .B(n428), .Z(n6479) );
  XOR U562 ( .A(n3407), .B(n3404), .Z(n429) );
  NAND U563 ( .A(n429), .B(n[232]), .Z(n430) );
  NAND U564 ( .A(n3407), .B(n3404), .Z(n431) );
  AND U565 ( .A(n430), .B(n431), .Z(n3400) );
  NAND U566 ( .A(n6302), .B(n6303), .Z(n432) );
  XOR U567 ( .A(n6303), .B(n6302), .Z(n433) );
  NANDN U568 ( .A(n6304), .B(n433), .Z(n434) );
  NAND U569 ( .A(n432), .B(n434), .Z(n6307) );
  XOR U570 ( .A(n6254), .B(n6255), .Z(n435) );
  NANDN U571 ( .A(n6253), .B(n435), .Z(n436) );
  NAND U572 ( .A(n6254), .B(n6255), .Z(n437) );
  AND U573 ( .A(n436), .B(n437), .Z(n6274) );
  XOR U574 ( .A(n6130), .B(n6131), .Z(n438) );
  NAND U575 ( .A(n438), .B(n6132), .Z(n439) );
  NAND U576 ( .A(n6130), .B(n6131), .Z(n440) );
  AND U577 ( .A(n439), .B(n440), .Z(n6139) );
  NAND U578 ( .A(n5995), .B(n5993), .Z(n441) );
  NANDN U579 ( .A(n5995), .B(n5994), .Z(n442) );
  NANDN U580 ( .A(n5996), .B(n442), .Z(n443) );
  NAND U581 ( .A(n441), .B(n443), .Z(n6002) );
  XOR U582 ( .A(n5928), .B(n5929), .Z(n444) );
  NANDN U583 ( .A(n5927), .B(n444), .Z(n445) );
  NAND U584 ( .A(n5928), .B(n5929), .Z(n446) );
  AND U585 ( .A(n445), .B(n446), .Z(n5933) );
  XOR U586 ( .A(n3702), .B(n3699), .Z(n447) );
  NAND U587 ( .A(n447), .B(n[159]), .Z(n448) );
  NAND U588 ( .A(n3702), .B(n3699), .Z(n449) );
  AND U589 ( .A(n448), .B(n449), .Z(n3694) );
  XOR U590 ( .A(n5863), .B(n5862), .Z(n450) );
  NANDN U591 ( .A(n5861), .B(n450), .Z(n451) );
  NAND U592 ( .A(n5863), .B(n5862), .Z(n452) );
  AND U593 ( .A(n451), .B(n452), .Z(n5868) );
  XOR U594 ( .A(n5696), .B(n5695), .Z(n453) );
  NANDN U595 ( .A(n5694), .B(n453), .Z(n454) );
  NAND U596 ( .A(n5696), .B(n5695), .Z(n455) );
  AND U597 ( .A(n454), .B(n455), .Z(n5699) );
  XOR U598 ( .A(n5666), .B(n5667), .Z(n456) );
  NAND U599 ( .A(n456), .B(n5668), .Z(n457) );
  NAND U600 ( .A(n5666), .B(n5667), .Z(n458) );
  AND U601 ( .A(n457), .B(n458), .Z(n5671) );
  NAND U602 ( .A(n5625), .B(n5624), .Z(n459) );
  XOR U603 ( .A(n5624), .B(n5625), .Z(n460) );
  NANDN U604 ( .A(n5626), .B(n460), .Z(n461) );
  NAND U605 ( .A(n459), .B(n461), .Z(n5629) );
  XOR U606 ( .A(n5569), .B(n5568), .Z(n462) );
  NANDN U607 ( .A(n5567), .B(n462), .Z(n463) );
  NAND U608 ( .A(n5569), .B(n5568), .Z(n464) );
  AND U609 ( .A(n463), .B(n464), .Z(n5572) );
  XOR U610 ( .A(n5551), .B(n5552), .Z(n465) );
  NAND U611 ( .A(n465), .B(n5553), .Z(n466) );
  NAND U612 ( .A(n5551), .B(n5552), .Z(n467) );
  AND U613 ( .A(n466), .B(n467), .Z(n5556) );
  XOR U614 ( .A(n6741), .B(n6738), .Z(n468) );
  NANDN U615 ( .A(n6739), .B(n468), .Z(n469) );
  NAND U616 ( .A(n6741), .B(n6738), .Z(n470) );
  AND U617 ( .A(n469), .B(n470), .Z(n6743) );
  XOR U618 ( .A(n6731), .B(n6730), .Z(n471) );
  NAND U619 ( .A(n471), .B(n6733), .Z(n472) );
  NAND U620 ( .A(n6731), .B(n6730), .Z(n473) );
  AND U621 ( .A(n472), .B(n473), .Z(n6735) );
  XOR U622 ( .A(n4474), .B(n[45]), .Z(n474) );
  NANDN U623 ( .A(n4471), .B(n474), .Z(n475) );
  NAND U624 ( .A(n4474), .B(n[45]), .Z(n476) );
  AND U625 ( .A(n475), .B(n476), .Z(n4171) );
  XOR U626 ( .A(n4213), .B(n[33]), .Z(n477) );
  NANDN U627 ( .A(n4210), .B(n477), .Z(n478) );
  NAND U628 ( .A(n4213), .B(n[33]), .Z(n479) );
  AND U629 ( .A(n478), .B(n479), .Z(n4206) );
  XOR U630 ( .A(n4234), .B(n4231), .Z(n480) );
  NAND U631 ( .A(n480), .B(n[25]), .Z(n481) );
  NAND U632 ( .A(n4234), .B(n4231), .Z(n482) );
  AND U633 ( .A(n481), .B(n482), .Z(n4227) );
  XOR U634 ( .A(n5716), .B(n5719), .Z(n483) );
  NAND U635 ( .A(n483), .B(n[12]), .Z(n484) );
  NAND U636 ( .A(n5716), .B(n5719), .Z(n485) );
  AND U637 ( .A(n484), .B(n485), .Z(n5782) );
  XOR U638 ( .A(n6239), .B(n6240), .Z(n486) );
  NAND U639 ( .A(n486), .B(n6241), .Z(n487) );
  NAND U640 ( .A(n6239), .B(n6240), .Z(n488) );
  AND U641 ( .A(n487), .B(n488), .Z(n6244) );
  NAND U642 ( .A(n5612), .B(n5613), .Z(n489) );
  XOR U643 ( .A(n5613), .B(n5612), .Z(n490) );
  NAND U644 ( .A(n490), .B(n5614), .Z(n491) );
  NAND U645 ( .A(n489), .B(n491), .Z(n5617) );
  XOR U646 ( .A(n6862), .B(n6859), .Z(n492) );
  NANDN U647 ( .A(n6860), .B(n492), .Z(n493) );
  NAND U648 ( .A(n6862), .B(n6859), .Z(n494) );
  AND U649 ( .A(n493), .B(n494), .Z(n6864) );
  XOR U650 ( .A(n6804), .B(n6806), .Z(n495) );
  NAND U651 ( .A(n495), .B(n6803), .Z(n496) );
  NAND U652 ( .A(n6804), .B(n6806), .Z(n497) );
  AND U653 ( .A(n496), .B(n497), .Z(n6807) );
  XOR U654 ( .A(n6770), .B(n6767), .Z(n498) );
  NANDN U655 ( .A(n6768), .B(n498), .Z(n499) );
  NAND U656 ( .A(n6770), .B(n6767), .Z(n500) );
  AND U657 ( .A(n499), .B(n500), .Z(n6772) );
  XOR U658 ( .A(n[44]), .B(n6705), .Z(n501) );
  NAND U659 ( .A(n501), .B(n6702), .Z(n502) );
  NAND U660 ( .A(n[44]), .B(n6705), .Z(n503) );
  AND U661 ( .A(n502), .B(n503), .Z(n6706) );
  XOR U662 ( .A(n[32]), .B(n6640), .Z(n504) );
  NANDN U663 ( .A(n4416), .B(n6630), .Z(n505) );
  XOR U664 ( .A(n6630), .B(n[31]), .Z(n506) );
  NAND U665 ( .A(n506), .B(n6633), .Z(n507) );
  NAND U666 ( .A(n505), .B(n507), .Z(n508) );
  NAND U667 ( .A(n504), .B(n508), .Z(n509) );
  NAND U668 ( .A(n[32]), .B(n6640), .Z(n510) );
  AND U669 ( .A(n509), .B(n510), .Z(n6641) );
  NAND U670 ( .A(n6606), .B(n6609), .Z(n511) );
  XOR U671 ( .A(n6609), .B(n6606), .Z(n512) );
  NANDN U672 ( .A(n4399), .B(n512), .Z(n513) );
  NAND U673 ( .A(n511), .B(n513), .Z(n6610) );
  XOR U674 ( .A(n[21]), .B(n6334), .Z(n514) );
  NAND U675 ( .A(n514), .B(n6331), .Z(n515) );
  NAND U676 ( .A(n[21]), .B(n6334), .Z(n516) );
  AND U677 ( .A(n515), .B(n516), .Z(n6403) );
  XOR U678 ( .A(n6867), .B(n6871), .Z(n517) );
  NANDN U679 ( .A(n6868), .B(n517), .Z(n518) );
  NAND U680 ( .A(n6867), .B(n6871), .Z(n519) );
  AND U681 ( .A(n518), .B(n519), .Z(n5595) );
  NAND U682 ( .A(n6195), .B(n[1]), .Z(n520) );
  XOR U683 ( .A(n[1]), .B(n6195), .Z(n521) );
  NANDN U684 ( .A(n6198), .B(n521), .Z(n522) );
  NAND U685 ( .A(n520), .B(n522), .Z(n6615) );
  IV U686 ( .A(n523), .Z(n524) );
  IV U687 ( .A(n6814), .Z(n525) );
  AND U688 ( .A(N4), .B(xregN_1), .Z(n2880) );
  IV U689 ( .A(n[254]), .Z(n6582) );
  NAND U690 ( .A(y[253]), .B(zin[252]), .Z(n1281) );
  XOR U691 ( .A(zin[252]), .B(y[253]), .Z(n1279) );
  NAND U692 ( .A(y[252]), .B(zin[251]), .Z(n1278) );
  XOR U693 ( .A(zin[251]), .B(y[252]), .Z(n1276) );
  NAND U694 ( .A(y[251]), .B(zin[250]), .Z(n1275) );
  XOR U695 ( .A(zin[250]), .B(y[251]), .Z(n1273) );
  NAND U696 ( .A(y[250]), .B(zin[249]), .Z(n1272) );
  XOR U697 ( .A(zin[249]), .B(y[250]), .Z(n1270) );
  NAND U698 ( .A(y[249]), .B(zin[248]), .Z(n1269) );
  XOR U699 ( .A(zin[248]), .B(y[249]), .Z(n1267) );
  NAND U700 ( .A(y[248]), .B(zin[247]), .Z(n1266) );
  XOR U701 ( .A(zin[247]), .B(y[248]), .Z(n1264) );
  NAND U702 ( .A(y[247]), .B(zin[246]), .Z(n1263) );
  XOR U703 ( .A(zin[246]), .B(y[247]), .Z(n1261) );
  NAND U704 ( .A(y[246]), .B(zin[245]), .Z(n1260) );
  XOR U705 ( .A(zin[245]), .B(y[246]), .Z(n1258) );
  NAND U706 ( .A(y[245]), .B(zin[244]), .Z(n1257) );
  XOR U707 ( .A(zin[244]), .B(y[245]), .Z(n1255) );
  NAND U708 ( .A(y[244]), .B(zin[243]), .Z(n1254) );
  XOR U709 ( .A(zin[243]), .B(y[244]), .Z(n1252) );
  NAND U710 ( .A(y[243]), .B(zin[242]), .Z(n1251) );
  XOR U711 ( .A(zin[242]), .B(y[243]), .Z(n1249) );
  NAND U712 ( .A(y[242]), .B(zin[241]), .Z(n1248) );
  XOR U713 ( .A(zin[241]), .B(y[242]), .Z(n1246) );
  NAND U714 ( .A(y[241]), .B(zin[240]), .Z(n1245) );
  XOR U715 ( .A(zin[240]), .B(y[241]), .Z(n1243) );
  NAND U716 ( .A(y[240]), .B(zin[239]), .Z(n1242) );
  XOR U717 ( .A(zin[239]), .B(y[240]), .Z(n1240) );
  NAND U718 ( .A(y[239]), .B(zin[238]), .Z(n1239) );
  XOR U719 ( .A(zin[238]), .B(y[239]), .Z(n1237) );
  NAND U720 ( .A(y[238]), .B(zin[237]), .Z(n1236) );
  XOR U721 ( .A(zin[237]), .B(y[238]), .Z(n1234) );
  NAND U722 ( .A(y[237]), .B(zin[236]), .Z(n1233) );
  XOR U723 ( .A(zin[236]), .B(y[237]), .Z(n1231) );
  NAND U724 ( .A(y[236]), .B(zin[235]), .Z(n1230) );
  XOR U725 ( .A(zin[235]), .B(y[236]), .Z(n1228) );
  NAND U726 ( .A(y[235]), .B(zin[234]), .Z(n1227) );
  XOR U727 ( .A(zin[234]), .B(y[235]), .Z(n1225) );
  NAND U728 ( .A(y[234]), .B(zin[233]), .Z(n1224) );
  XOR U729 ( .A(zin[233]), .B(y[234]), .Z(n1222) );
  NAND U730 ( .A(y[233]), .B(zin[232]), .Z(n1221) );
  XOR U731 ( .A(zin[232]), .B(y[233]), .Z(n1219) );
  NAND U732 ( .A(y[232]), .B(zin[231]), .Z(n1218) );
  XOR U733 ( .A(zin[231]), .B(y[232]), .Z(n1216) );
  NAND U734 ( .A(y[231]), .B(zin[230]), .Z(n1215) );
  XOR U735 ( .A(zin[230]), .B(y[231]), .Z(n1213) );
  NAND U736 ( .A(y[230]), .B(zin[229]), .Z(n1212) );
  XOR U737 ( .A(zin[229]), .B(y[230]), .Z(n1210) );
  NAND U738 ( .A(y[229]), .B(zin[228]), .Z(n1209) );
  XOR U739 ( .A(zin[228]), .B(y[229]), .Z(n1207) );
  NAND U740 ( .A(y[228]), .B(zin[227]), .Z(n1206) );
  XOR U741 ( .A(zin[227]), .B(y[228]), .Z(n1204) );
  NAND U742 ( .A(y[227]), .B(zin[226]), .Z(n1203) );
  XOR U743 ( .A(zin[226]), .B(y[227]), .Z(n1201) );
  NAND U744 ( .A(y[226]), .B(zin[225]), .Z(n1200) );
  XOR U745 ( .A(zin[225]), .B(y[226]), .Z(n1198) );
  NAND U746 ( .A(y[225]), .B(zin[224]), .Z(n1197) );
  XOR U747 ( .A(zin[224]), .B(y[225]), .Z(n1195) );
  NAND U748 ( .A(y[224]), .B(zin[223]), .Z(n1194) );
  XOR U749 ( .A(zin[223]), .B(y[224]), .Z(n1192) );
  NAND U750 ( .A(y[223]), .B(zin[222]), .Z(n1191) );
  XOR U751 ( .A(zin[222]), .B(y[223]), .Z(n1189) );
  NAND U752 ( .A(y[222]), .B(zin[221]), .Z(n1188) );
  XOR U753 ( .A(zin[221]), .B(y[222]), .Z(n1186) );
  NAND U754 ( .A(y[221]), .B(zin[220]), .Z(n1185) );
  XOR U755 ( .A(zin[220]), .B(y[221]), .Z(n1183) );
  NAND U756 ( .A(y[220]), .B(zin[219]), .Z(n1182) );
  XOR U757 ( .A(zin[219]), .B(y[220]), .Z(n1180) );
  NAND U758 ( .A(y[219]), .B(zin[218]), .Z(n1179) );
  XOR U759 ( .A(zin[218]), .B(y[219]), .Z(n1177) );
  NAND U760 ( .A(y[218]), .B(zin[217]), .Z(n1176) );
  XOR U761 ( .A(zin[217]), .B(y[218]), .Z(n1174) );
  NAND U762 ( .A(y[217]), .B(zin[216]), .Z(n1173) );
  XOR U763 ( .A(zin[216]), .B(y[217]), .Z(n1171) );
  NAND U764 ( .A(y[216]), .B(zin[215]), .Z(n1170) );
  XOR U765 ( .A(zin[215]), .B(y[216]), .Z(n1168) );
  NAND U766 ( .A(y[215]), .B(zin[214]), .Z(n1167) );
  XOR U767 ( .A(zin[214]), .B(y[215]), .Z(n1165) );
  NAND U768 ( .A(y[214]), .B(zin[213]), .Z(n1164) );
  XOR U769 ( .A(zin[213]), .B(y[214]), .Z(n1162) );
  NAND U770 ( .A(y[213]), .B(zin[212]), .Z(n1161) );
  XOR U771 ( .A(zin[212]), .B(y[213]), .Z(n1159) );
  NAND U772 ( .A(y[212]), .B(zin[211]), .Z(n1158) );
  XOR U773 ( .A(zin[211]), .B(y[212]), .Z(n1156) );
  NAND U774 ( .A(y[211]), .B(zin[210]), .Z(n1155) );
  XOR U775 ( .A(zin[210]), .B(y[211]), .Z(n1153) );
  NAND U776 ( .A(y[210]), .B(zin[209]), .Z(n1152) );
  XOR U777 ( .A(zin[209]), .B(y[210]), .Z(n1150) );
  NAND U778 ( .A(y[209]), .B(zin[208]), .Z(n1149) );
  XOR U779 ( .A(zin[208]), .B(y[209]), .Z(n1147) );
  NAND U780 ( .A(y[208]), .B(zin[207]), .Z(n1146) );
  XOR U781 ( .A(zin[207]), .B(y[208]), .Z(n1144) );
  NAND U782 ( .A(y[207]), .B(zin[206]), .Z(n1143) );
  XOR U783 ( .A(zin[206]), .B(y[207]), .Z(n1141) );
  NAND U784 ( .A(y[206]), .B(zin[205]), .Z(n1140) );
  XOR U785 ( .A(zin[205]), .B(y[206]), .Z(n1138) );
  NAND U786 ( .A(y[205]), .B(zin[204]), .Z(n1137) );
  XOR U787 ( .A(zin[204]), .B(y[205]), .Z(n1135) );
  NAND U788 ( .A(y[204]), .B(zin[203]), .Z(n1134) );
  XOR U789 ( .A(zin[203]), .B(y[204]), .Z(n1132) );
  NAND U790 ( .A(y[203]), .B(zin[202]), .Z(n1131) );
  XOR U791 ( .A(zin[202]), .B(y[203]), .Z(n1129) );
  NAND U792 ( .A(y[202]), .B(zin[201]), .Z(n1128) );
  XOR U793 ( .A(zin[201]), .B(y[202]), .Z(n1126) );
  NAND U794 ( .A(y[201]), .B(zin[200]), .Z(n1125) );
  XOR U795 ( .A(zin[200]), .B(y[201]), .Z(n1123) );
  NAND U796 ( .A(y[200]), .B(zin[199]), .Z(n1122) );
  XOR U797 ( .A(zin[199]), .B(y[200]), .Z(n1120) );
  NAND U798 ( .A(y[199]), .B(zin[198]), .Z(n1119) );
  XOR U799 ( .A(zin[198]), .B(y[199]), .Z(n1117) );
  NAND U800 ( .A(y[198]), .B(zin[197]), .Z(n1116) );
  XOR U801 ( .A(zin[197]), .B(y[198]), .Z(n1114) );
  NAND U802 ( .A(y[197]), .B(zin[196]), .Z(n1113) );
  XOR U803 ( .A(zin[196]), .B(y[197]), .Z(n1111) );
  NAND U804 ( .A(y[196]), .B(zin[195]), .Z(n1110) );
  XOR U805 ( .A(zin[195]), .B(y[196]), .Z(n1108) );
  NAND U806 ( .A(y[195]), .B(zin[194]), .Z(n1107) );
  XOR U807 ( .A(zin[194]), .B(y[195]), .Z(n1105) );
  NAND U808 ( .A(y[194]), .B(zin[193]), .Z(n1104) );
  XOR U809 ( .A(zin[193]), .B(y[194]), .Z(n1102) );
  NAND U810 ( .A(y[193]), .B(zin[192]), .Z(n1101) );
  XOR U811 ( .A(zin[192]), .B(y[193]), .Z(n1099) );
  NAND U812 ( .A(y[192]), .B(zin[191]), .Z(n1098) );
  XOR U813 ( .A(zin[191]), .B(y[192]), .Z(n1096) );
  NAND U814 ( .A(y[191]), .B(zin[190]), .Z(n1095) );
  XOR U815 ( .A(zin[190]), .B(y[191]), .Z(n1093) );
  NAND U816 ( .A(y[190]), .B(zin[189]), .Z(n1092) );
  XOR U817 ( .A(zin[189]), .B(y[190]), .Z(n1090) );
  NAND U818 ( .A(y[189]), .B(zin[188]), .Z(n1089) );
  XOR U819 ( .A(zin[188]), .B(y[189]), .Z(n1087) );
  NAND U820 ( .A(y[188]), .B(zin[187]), .Z(n1086) );
  XOR U821 ( .A(zin[187]), .B(y[188]), .Z(n1084) );
  NAND U822 ( .A(y[187]), .B(zin[186]), .Z(n1083) );
  XOR U823 ( .A(zin[186]), .B(y[187]), .Z(n1081) );
  NAND U824 ( .A(y[186]), .B(zin[185]), .Z(n1080) );
  XOR U825 ( .A(zin[185]), .B(y[186]), .Z(n1078) );
  NAND U826 ( .A(y[185]), .B(zin[184]), .Z(n1077) );
  XOR U827 ( .A(zin[184]), .B(y[185]), .Z(n1075) );
  NAND U828 ( .A(y[184]), .B(zin[183]), .Z(n1074) );
  XOR U829 ( .A(zin[183]), .B(y[184]), .Z(n1072) );
  NAND U830 ( .A(y[183]), .B(zin[182]), .Z(n1071) );
  XOR U831 ( .A(zin[182]), .B(y[183]), .Z(n1069) );
  NAND U832 ( .A(y[182]), .B(zin[181]), .Z(n1068) );
  XOR U833 ( .A(zin[181]), .B(y[182]), .Z(n1066) );
  NAND U834 ( .A(y[181]), .B(zin[180]), .Z(n1065) );
  XOR U835 ( .A(zin[180]), .B(y[181]), .Z(n1063) );
  NAND U836 ( .A(y[180]), .B(zin[179]), .Z(n1062) );
  XOR U837 ( .A(zin[179]), .B(y[180]), .Z(n1060) );
  NAND U838 ( .A(y[179]), .B(zin[178]), .Z(n1059) );
  XOR U839 ( .A(zin[178]), .B(y[179]), .Z(n1057) );
  NAND U840 ( .A(y[178]), .B(zin[177]), .Z(n1056) );
  XOR U841 ( .A(zin[177]), .B(y[178]), .Z(n1054) );
  NAND U842 ( .A(y[177]), .B(zin[176]), .Z(n1053) );
  XOR U843 ( .A(zin[176]), .B(y[177]), .Z(n1051) );
  NAND U844 ( .A(y[176]), .B(zin[175]), .Z(n1050) );
  XOR U845 ( .A(zin[175]), .B(y[176]), .Z(n1048) );
  NAND U846 ( .A(y[175]), .B(zin[174]), .Z(n1047) );
  XOR U847 ( .A(zin[174]), .B(y[175]), .Z(n1045) );
  NAND U848 ( .A(y[174]), .B(zin[173]), .Z(n1044) );
  XOR U849 ( .A(zin[173]), .B(y[174]), .Z(n1042) );
  NAND U850 ( .A(y[173]), .B(zin[172]), .Z(n1041) );
  XOR U851 ( .A(zin[172]), .B(y[173]), .Z(n1039) );
  NAND U852 ( .A(y[172]), .B(zin[171]), .Z(n1038) );
  XOR U853 ( .A(zin[171]), .B(y[172]), .Z(n1036) );
  NAND U854 ( .A(y[171]), .B(zin[170]), .Z(n1035) );
  XOR U855 ( .A(zin[170]), .B(y[171]), .Z(n1033) );
  NAND U856 ( .A(y[170]), .B(zin[169]), .Z(n1032) );
  XOR U857 ( .A(zin[169]), .B(y[170]), .Z(n1030) );
  NAND U858 ( .A(y[169]), .B(zin[168]), .Z(n1029) );
  XOR U859 ( .A(zin[168]), .B(y[169]), .Z(n1027) );
  NAND U860 ( .A(y[168]), .B(zin[167]), .Z(n1026) );
  XOR U861 ( .A(zin[167]), .B(y[168]), .Z(n1024) );
  NAND U862 ( .A(y[167]), .B(zin[166]), .Z(n1023) );
  XOR U863 ( .A(zin[166]), .B(y[167]), .Z(n1021) );
  NAND U864 ( .A(y[166]), .B(zin[165]), .Z(n1020) );
  XOR U865 ( .A(zin[165]), .B(y[166]), .Z(n1018) );
  NAND U866 ( .A(y[165]), .B(zin[164]), .Z(n1017) );
  XOR U867 ( .A(zin[164]), .B(y[165]), .Z(n1015) );
  NAND U868 ( .A(y[164]), .B(zin[163]), .Z(n1014) );
  XOR U869 ( .A(zin[163]), .B(y[164]), .Z(n1012) );
  NAND U870 ( .A(y[163]), .B(zin[162]), .Z(n1011) );
  XOR U871 ( .A(zin[162]), .B(y[163]), .Z(n1009) );
  NAND U872 ( .A(y[162]), .B(zin[161]), .Z(n1008) );
  XOR U873 ( .A(zin[161]), .B(y[162]), .Z(n1006) );
  NAND U874 ( .A(y[161]), .B(zin[160]), .Z(n1005) );
  XOR U875 ( .A(zin[160]), .B(y[161]), .Z(n1003) );
  NAND U876 ( .A(y[160]), .B(zin[159]), .Z(n1002) );
  XOR U877 ( .A(zin[159]), .B(y[160]), .Z(n1000) );
  NAND U878 ( .A(y[159]), .B(zin[158]), .Z(n999) );
  XOR U879 ( .A(zin[158]), .B(y[159]), .Z(n997) );
  NAND U880 ( .A(y[158]), .B(zin[157]), .Z(n996) );
  XOR U881 ( .A(zin[157]), .B(y[158]), .Z(n994) );
  NAND U882 ( .A(y[157]), .B(zin[156]), .Z(n993) );
  XOR U883 ( .A(zin[156]), .B(y[157]), .Z(n991) );
  NAND U884 ( .A(y[156]), .B(zin[155]), .Z(n990) );
  XOR U885 ( .A(zin[155]), .B(y[156]), .Z(n988) );
  NAND U886 ( .A(y[155]), .B(zin[154]), .Z(n987) );
  XOR U887 ( .A(zin[154]), .B(y[155]), .Z(n985) );
  NAND U888 ( .A(y[154]), .B(zin[153]), .Z(n984) );
  XOR U889 ( .A(zin[153]), .B(y[154]), .Z(n982) );
  NAND U890 ( .A(y[153]), .B(zin[152]), .Z(n981) );
  XOR U891 ( .A(zin[152]), .B(y[153]), .Z(n979) );
  NAND U892 ( .A(y[152]), .B(zin[151]), .Z(n978) );
  XOR U893 ( .A(zin[151]), .B(y[152]), .Z(n976) );
  NAND U894 ( .A(y[151]), .B(zin[150]), .Z(n975) );
  XOR U895 ( .A(zin[150]), .B(y[151]), .Z(n973) );
  NAND U896 ( .A(y[150]), .B(zin[149]), .Z(n972) );
  XOR U897 ( .A(zin[149]), .B(y[150]), .Z(n970) );
  NAND U898 ( .A(y[149]), .B(zin[148]), .Z(n969) );
  XOR U899 ( .A(zin[148]), .B(y[149]), .Z(n967) );
  NAND U900 ( .A(y[148]), .B(zin[147]), .Z(n966) );
  XOR U901 ( .A(zin[147]), .B(y[148]), .Z(n964) );
  NAND U902 ( .A(y[147]), .B(zin[146]), .Z(n963) );
  XOR U903 ( .A(zin[146]), .B(y[147]), .Z(n961) );
  NAND U904 ( .A(y[146]), .B(zin[145]), .Z(n960) );
  XOR U905 ( .A(zin[145]), .B(y[146]), .Z(n958) );
  NAND U906 ( .A(y[145]), .B(zin[144]), .Z(n957) );
  XOR U907 ( .A(zin[144]), .B(y[145]), .Z(n955) );
  NAND U908 ( .A(y[144]), .B(zin[143]), .Z(n954) );
  XOR U909 ( .A(zin[143]), .B(y[144]), .Z(n952) );
  NAND U910 ( .A(y[143]), .B(zin[142]), .Z(n951) );
  XOR U911 ( .A(zin[142]), .B(y[143]), .Z(n949) );
  NAND U912 ( .A(y[142]), .B(zin[141]), .Z(n948) );
  XOR U913 ( .A(zin[141]), .B(y[142]), .Z(n946) );
  NAND U914 ( .A(y[141]), .B(zin[140]), .Z(n945) );
  XOR U915 ( .A(zin[140]), .B(y[141]), .Z(n943) );
  NAND U916 ( .A(y[140]), .B(zin[139]), .Z(n942) );
  XOR U917 ( .A(zin[139]), .B(y[140]), .Z(n940) );
  NAND U918 ( .A(y[139]), .B(zin[138]), .Z(n939) );
  XOR U919 ( .A(zin[138]), .B(y[139]), .Z(n937) );
  NAND U920 ( .A(y[138]), .B(zin[137]), .Z(n936) );
  XOR U921 ( .A(zin[137]), .B(y[138]), .Z(n934) );
  NAND U922 ( .A(y[137]), .B(zin[136]), .Z(n933) );
  XOR U923 ( .A(zin[136]), .B(y[137]), .Z(n931) );
  NAND U924 ( .A(y[136]), .B(zin[135]), .Z(n930) );
  XOR U925 ( .A(zin[135]), .B(y[136]), .Z(n928) );
  NAND U926 ( .A(y[135]), .B(zin[134]), .Z(n927) );
  XOR U927 ( .A(zin[134]), .B(y[135]), .Z(n925) );
  NAND U928 ( .A(y[134]), .B(zin[133]), .Z(n924) );
  XOR U929 ( .A(zin[133]), .B(y[134]), .Z(n922) );
  NAND U930 ( .A(y[133]), .B(zin[132]), .Z(n921) );
  XOR U931 ( .A(zin[132]), .B(y[133]), .Z(n919) );
  NAND U932 ( .A(y[132]), .B(zin[131]), .Z(n918) );
  XOR U933 ( .A(zin[131]), .B(y[132]), .Z(n916) );
  NAND U934 ( .A(y[131]), .B(zin[130]), .Z(n915) );
  XOR U935 ( .A(zin[130]), .B(y[131]), .Z(n913) );
  NAND U936 ( .A(y[130]), .B(zin[129]), .Z(n912) );
  XOR U937 ( .A(zin[129]), .B(y[130]), .Z(n910) );
  NAND U938 ( .A(y[129]), .B(zin[128]), .Z(n909) );
  XOR U939 ( .A(zin[128]), .B(y[129]), .Z(n907) );
  NAND U940 ( .A(y[128]), .B(zin[127]), .Z(n906) );
  XOR U941 ( .A(zin[127]), .B(y[128]), .Z(n904) );
  NAND U942 ( .A(y[127]), .B(zin[126]), .Z(n903) );
  XOR U943 ( .A(zin[126]), .B(y[127]), .Z(n901) );
  NAND U944 ( .A(y[126]), .B(zin[125]), .Z(n900) );
  XOR U945 ( .A(zin[125]), .B(y[126]), .Z(n898) );
  NAND U946 ( .A(y[125]), .B(zin[124]), .Z(n897) );
  XOR U947 ( .A(zin[124]), .B(y[125]), .Z(n895) );
  NAND U948 ( .A(y[124]), .B(zin[123]), .Z(n894) );
  XOR U949 ( .A(zin[123]), .B(y[124]), .Z(n892) );
  NAND U950 ( .A(y[123]), .B(zin[122]), .Z(n891) );
  XOR U951 ( .A(zin[122]), .B(y[123]), .Z(n889) );
  NAND U952 ( .A(y[122]), .B(zin[121]), .Z(n888) );
  XOR U953 ( .A(zin[121]), .B(y[122]), .Z(n886) );
  NAND U954 ( .A(y[121]), .B(zin[120]), .Z(n885) );
  XOR U955 ( .A(zin[120]), .B(y[121]), .Z(n883) );
  NAND U956 ( .A(y[120]), .B(zin[119]), .Z(n882) );
  XOR U957 ( .A(zin[119]), .B(y[120]), .Z(n880) );
  NAND U958 ( .A(y[119]), .B(zin[118]), .Z(n879) );
  XOR U959 ( .A(zin[118]), .B(y[119]), .Z(n877) );
  NAND U960 ( .A(y[118]), .B(zin[117]), .Z(n876) );
  XOR U961 ( .A(zin[117]), .B(y[118]), .Z(n874) );
  NAND U962 ( .A(y[117]), .B(zin[116]), .Z(n873) );
  XOR U963 ( .A(zin[116]), .B(y[117]), .Z(n871) );
  NAND U964 ( .A(y[116]), .B(zin[115]), .Z(n870) );
  XOR U965 ( .A(zin[115]), .B(y[116]), .Z(n868) );
  NAND U966 ( .A(y[115]), .B(zin[114]), .Z(n867) );
  XOR U967 ( .A(zin[114]), .B(y[115]), .Z(n865) );
  NAND U968 ( .A(y[114]), .B(zin[113]), .Z(n864) );
  XOR U969 ( .A(zin[113]), .B(y[114]), .Z(n862) );
  NAND U970 ( .A(y[113]), .B(zin[112]), .Z(n861) );
  XOR U971 ( .A(zin[112]), .B(y[113]), .Z(n859) );
  NAND U972 ( .A(y[112]), .B(zin[111]), .Z(n858) );
  XOR U973 ( .A(zin[111]), .B(y[112]), .Z(n856) );
  NAND U974 ( .A(y[111]), .B(zin[110]), .Z(n855) );
  XOR U975 ( .A(zin[110]), .B(y[111]), .Z(n853) );
  NAND U976 ( .A(y[110]), .B(zin[109]), .Z(n852) );
  XOR U977 ( .A(zin[109]), .B(y[110]), .Z(n850) );
  NAND U978 ( .A(y[109]), .B(zin[108]), .Z(n849) );
  XOR U979 ( .A(zin[108]), .B(y[109]), .Z(n847) );
  NAND U980 ( .A(y[108]), .B(zin[107]), .Z(n846) );
  XOR U981 ( .A(zin[107]), .B(y[108]), .Z(n844) );
  NAND U982 ( .A(y[107]), .B(zin[106]), .Z(n843) );
  XOR U983 ( .A(zin[106]), .B(y[107]), .Z(n841) );
  NAND U984 ( .A(y[106]), .B(zin[105]), .Z(n840) );
  XOR U985 ( .A(zin[105]), .B(y[106]), .Z(n838) );
  NAND U986 ( .A(y[105]), .B(zin[104]), .Z(n837) );
  XOR U987 ( .A(zin[104]), .B(y[105]), .Z(n835) );
  NAND U988 ( .A(y[104]), .B(zin[103]), .Z(n834) );
  XOR U989 ( .A(zin[103]), .B(y[104]), .Z(n832) );
  NAND U990 ( .A(y[103]), .B(zin[102]), .Z(n831) );
  XOR U991 ( .A(zin[102]), .B(y[103]), .Z(n829) );
  NAND U992 ( .A(y[102]), .B(zin[101]), .Z(n828) );
  XOR U993 ( .A(zin[101]), .B(y[102]), .Z(n826) );
  NAND U994 ( .A(y[101]), .B(zin[100]), .Z(n825) );
  XOR U995 ( .A(zin[100]), .B(y[101]), .Z(n823) );
  NAND U996 ( .A(y[100]), .B(zin[99]), .Z(n822) );
  XOR U997 ( .A(zin[99]), .B(y[100]), .Z(n820) );
  NAND U998 ( .A(zin[98]), .B(y[99]), .Z(n819) );
  XOR U999 ( .A(y[99]), .B(zin[98]), .Z(n817) );
  NAND U1000 ( .A(y[98]), .B(zin[97]), .Z(n816) );
  XOR U1001 ( .A(zin[97]), .B(y[98]), .Z(n814) );
  NAND U1002 ( .A(y[97]), .B(zin[96]), .Z(n813) );
  XOR U1003 ( .A(zin[96]), .B(y[97]), .Z(n811) );
  NAND U1004 ( .A(y[96]), .B(zin[95]), .Z(n810) );
  XOR U1005 ( .A(zin[95]), .B(y[96]), .Z(n808) );
  NAND U1006 ( .A(y[95]), .B(zin[94]), .Z(n807) );
  XOR U1007 ( .A(zin[94]), .B(y[95]), .Z(n805) );
  NAND U1008 ( .A(y[94]), .B(zin[93]), .Z(n804) );
  XOR U1009 ( .A(zin[93]), .B(y[94]), .Z(n802) );
  NAND U1010 ( .A(y[93]), .B(zin[92]), .Z(n801) );
  XOR U1011 ( .A(zin[92]), .B(y[93]), .Z(n799) );
  NAND U1012 ( .A(y[92]), .B(zin[91]), .Z(n798) );
  XOR U1013 ( .A(zin[91]), .B(y[92]), .Z(n796) );
  NAND U1014 ( .A(y[91]), .B(zin[90]), .Z(n795) );
  XOR U1015 ( .A(zin[90]), .B(y[91]), .Z(n793) );
  NAND U1016 ( .A(y[90]), .B(zin[89]), .Z(n792) );
  XOR U1017 ( .A(zin[89]), .B(y[90]), .Z(n790) );
  NAND U1018 ( .A(y[89]), .B(zin[88]), .Z(n789) );
  XOR U1019 ( .A(zin[88]), .B(y[89]), .Z(n787) );
  NAND U1020 ( .A(y[88]), .B(zin[87]), .Z(n786) );
  XOR U1021 ( .A(zin[87]), .B(y[88]), .Z(n784) );
  NAND U1022 ( .A(y[87]), .B(zin[86]), .Z(n783) );
  XOR U1023 ( .A(zin[86]), .B(y[87]), .Z(n781) );
  NAND U1024 ( .A(y[86]), .B(zin[85]), .Z(n780) );
  XOR U1025 ( .A(zin[85]), .B(y[86]), .Z(n778) );
  NAND U1026 ( .A(y[85]), .B(zin[84]), .Z(n777) );
  XOR U1027 ( .A(zin[84]), .B(y[85]), .Z(n775) );
  NAND U1028 ( .A(y[84]), .B(zin[83]), .Z(n774) );
  XOR U1029 ( .A(zin[83]), .B(y[84]), .Z(n772) );
  NAND U1030 ( .A(y[83]), .B(zin[82]), .Z(n771) );
  XOR U1031 ( .A(zin[82]), .B(y[83]), .Z(n769) );
  NAND U1032 ( .A(y[82]), .B(zin[81]), .Z(n768) );
  XOR U1033 ( .A(zin[81]), .B(y[82]), .Z(n766) );
  NAND U1034 ( .A(y[81]), .B(zin[80]), .Z(n765) );
  XOR U1035 ( .A(zin[80]), .B(y[81]), .Z(n763) );
  NAND U1036 ( .A(y[80]), .B(zin[79]), .Z(n762) );
  XOR U1037 ( .A(zin[79]), .B(y[80]), .Z(n760) );
  NAND U1038 ( .A(y[79]), .B(zin[78]), .Z(n759) );
  XOR U1039 ( .A(zin[78]), .B(y[79]), .Z(n757) );
  NAND U1040 ( .A(y[78]), .B(zin[77]), .Z(n756) );
  XOR U1041 ( .A(zin[77]), .B(y[78]), .Z(n754) );
  NAND U1042 ( .A(y[77]), .B(zin[76]), .Z(n753) );
  XOR U1043 ( .A(zin[76]), .B(y[77]), .Z(n751) );
  NAND U1044 ( .A(y[76]), .B(zin[75]), .Z(n750) );
  XOR U1045 ( .A(zin[75]), .B(y[76]), .Z(n748) );
  NAND U1046 ( .A(y[75]), .B(zin[74]), .Z(n747) );
  XOR U1047 ( .A(zin[74]), .B(y[75]), .Z(n745) );
  NAND U1048 ( .A(y[74]), .B(zin[73]), .Z(n744) );
  XOR U1049 ( .A(zin[73]), .B(y[74]), .Z(n742) );
  NAND U1050 ( .A(y[73]), .B(zin[72]), .Z(n741) );
  XOR U1051 ( .A(zin[72]), .B(y[73]), .Z(n739) );
  NAND U1052 ( .A(y[72]), .B(zin[71]), .Z(n738) );
  XOR U1053 ( .A(zin[71]), .B(y[72]), .Z(n736) );
  NAND U1054 ( .A(y[71]), .B(zin[70]), .Z(n735) );
  XOR U1055 ( .A(zin[70]), .B(y[71]), .Z(n733) );
  NAND U1056 ( .A(y[70]), .B(zin[69]), .Z(n732) );
  XOR U1057 ( .A(zin[69]), .B(y[70]), .Z(n730) );
  NAND U1058 ( .A(y[69]), .B(zin[68]), .Z(n729) );
  XOR U1059 ( .A(zin[68]), .B(y[69]), .Z(n727) );
  NAND U1060 ( .A(y[68]), .B(zin[67]), .Z(n726) );
  XOR U1061 ( .A(zin[67]), .B(y[68]), .Z(n724) );
  NAND U1062 ( .A(y[67]), .B(zin[66]), .Z(n723) );
  XOR U1063 ( .A(zin[66]), .B(y[67]), .Z(n721) );
  NAND U1064 ( .A(y[66]), .B(zin[65]), .Z(n720) );
  XOR U1065 ( .A(zin[65]), .B(y[66]), .Z(n718) );
  NAND U1066 ( .A(y[65]), .B(zin[64]), .Z(n717) );
  XOR U1067 ( .A(zin[64]), .B(y[65]), .Z(n715) );
  NAND U1068 ( .A(y[64]), .B(zin[63]), .Z(n714) );
  XOR U1069 ( .A(zin[63]), .B(y[64]), .Z(n712) );
  NAND U1070 ( .A(y[63]), .B(zin[62]), .Z(n711) );
  XOR U1071 ( .A(zin[62]), .B(y[63]), .Z(n709) );
  NAND U1072 ( .A(y[62]), .B(zin[61]), .Z(n708) );
  XOR U1073 ( .A(zin[61]), .B(y[62]), .Z(n706) );
  NAND U1074 ( .A(y[61]), .B(zin[60]), .Z(n705) );
  XOR U1075 ( .A(zin[60]), .B(y[61]), .Z(n703) );
  NAND U1076 ( .A(y[60]), .B(zin[59]), .Z(n702) );
  XOR U1077 ( .A(zin[59]), .B(y[60]), .Z(n700) );
  NAND U1078 ( .A(y[59]), .B(zin[58]), .Z(n699) );
  XOR U1079 ( .A(zin[58]), .B(y[59]), .Z(n697) );
  NAND U1080 ( .A(y[58]), .B(zin[57]), .Z(n696) );
  XOR U1081 ( .A(zin[57]), .B(y[58]), .Z(n694) );
  NAND U1082 ( .A(y[57]), .B(zin[56]), .Z(n693) );
  XOR U1083 ( .A(zin[56]), .B(y[57]), .Z(n691) );
  NAND U1084 ( .A(y[56]), .B(zin[55]), .Z(n690) );
  XOR U1085 ( .A(zin[55]), .B(y[56]), .Z(n688) );
  NAND U1086 ( .A(y[55]), .B(zin[54]), .Z(n687) );
  XOR U1087 ( .A(zin[54]), .B(y[55]), .Z(n685) );
  NAND U1088 ( .A(y[54]), .B(zin[53]), .Z(n684) );
  XOR U1089 ( .A(zin[53]), .B(y[54]), .Z(n682) );
  NAND U1090 ( .A(y[53]), .B(zin[52]), .Z(n681) );
  XOR U1091 ( .A(zin[52]), .B(y[53]), .Z(n679) );
  NAND U1092 ( .A(y[52]), .B(zin[51]), .Z(n678) );
  XOR U1093 ( .A(zin[51]), .B(y[52]), .Z(n676) );
  NAND U1094 ( .A(y[51]), .B(zin[50]), .Z(n675) );
  XOR U1095 ( .A(zin[50]), .B(y[51]), .Z(n673) );
  NAND U1096 ( .A(y[50]), .B(zin[49]), .Z(n672) );
  XOR U1097 ( .A(zin[49]), .B(y[50]), .Z(n670) );
  NAND U1098 ( .A(y[49]), .B(zin[48]), .Z(n669) );
  XOR U1099 ( .A(zin[48]), .B(y[49]), .Z(n667) );
  NAND U1100 ( .A(y[48]), .B(zin[47]), .Z(n666) );
  XOR U1101 ( .A(zin[47]), .B(y[48]), .Z(n664) );
  NAND U1102 ( .A(y[47]), .B(zin[46]), .Z(n663) );
  XOR U1103 ( .A(zin[46]), .B(y[47]), .Z(n661) );
  NAND U1104 ( .A(y[46]), .B(zin[45]), .Z(n660) );
  XOR U1105 ( .A(zin[45]), .B(y[46]), .Z(n658) );
  NAND U1106 ( .A(y[45]), .B(zin[44]), .Z(n657) );
  XOR U1107 ( .A(zin[44]), .B(y[45]), .Z(n655) );
  NAND U1108 ( .A(y[44]), .B(zin[43]), .Z(n654) );
  XOR U1109 ( .A(zin[43]), .B(y[44]), .Z(n652) );
  NAND U1110 ( .A(y[43]), .B(zin[42]), .Z(n651) );
  XOR U1111 ( .A(zin[42]), .B(y[43]), .Z(n649) );
  NAND U1112 ( .A(y[42]), .B(zin[41]), .Z(n648) );
  XOR U1113 ( .A(zin[41]), .B(y[42]), .Z(n646) );
  NAND U1114 ( .A(y[41]), .B(zin[40]), .Z(n645) );
  XOR U1115 ( .A(zin[40]), .B(y[41]), .Z(n643) );
  NAND U1116 ( .A(y[40]), .B(zin[39]), .Z(n642) );
  XOR U1117 ( .A(zin[39]), .B(y[40]), .Z(n640) );
  NAND U1118 ( .A(y[39]), .B(zin[38]), .Z(n639) );
  XOR U1119 ( .A(zin[38]), .B(y[39]), .Z(n637) );
  NAND U1120 ( .A(y[38]), .B(zin[37]), .Z(n636) );
  XOR U1121 ( .A(zin[37]), .B(y[38]), .Z(n634) );
  NAND U1122 ( .A(y[37]), .B(zin[36]), .Z(n633) );
  XOR U1123 ( .A(zin[36]), .B(y[37]), .Z(n631) );
  NAND U1124 ( .A(y[36]), .B(zin[35]), .Z(n630) );
  XOR U1125 ( .A(zin[35]), .B(y[36]), .Z(n628) );
  NAND U1126 ( .A(y[35]), .B(zin[34]), .Z(n627) );
  XOR U1127 ( .A(zin[34]), .B(y[35]), .Z(n625) );
  NAND U1128 ( .A(y[34]), .B(zin[33]), .Z(n624) );
  XOR U1129 ( .A(zin[33]), .B(y[34]), .Z(n622) );
  NAND U1130 ( .A(y[33]), .B(zin[32]), .Z(n621) );
  XOR U1131 ( .A(zin[32]), .B(y[33]), .Z(n619) );
  NAND U1132 ( .A(y[32]), .B(zin[31]), .Z(n618) );
  XOR U1133 ( .A(zin[31]), .B(y[32]), .Z(n616) );
  NAND U1134 ( .A(y[31]), .B(zin[30]), .Z(n615) );
  XOR U1135 ( .A(zin[30]), .B(y[31]), .Z(n613) );
  NAND U1136 ( .A(y[30]), .B(zin[29]), .Z(n612) );
  XOR U1137 ( .A(zin[29]), .B(y[30]), .Z(n610) );
  NAND U1138 ( .A(y[29]), .B(zin[28]), .Z(n609) );
  XOR U1139 ( .A(zin[28]), .B(y[29]), .Z(n607) );
  NAND U1140 ( .A(y[28]), .B(zin[27]), .Z(n606) );
  XOR U1141 ( .A(zin[27]), .B(y[28]), .Z(n604) );
  NAND U1142 ( .A(y[27]), .B(zin[26]), .Z(n603) );
  XOR U1143 ( .A(zin[26]), .B(y[27]), .Z(n601) );
  NAND U1144 ( .A(y[26]), .B(zin[25]), .Z(n600) );
  XOR U1145 ( .A(zin[25]), .B(y[26]), .Z(n598) );
  NAND U1146 ( .A(y[25]), .B(zin[24]), .Z(n597) );
  XOR U1147 ( .A(zin[24]), .B(y[25]), .Z(n595) );
  NAND U1148 ( .A(y[24]), .B(zin[23]), .Z(n594) );
  XOR U1149 ( .A(zin[23]), .B(y[24]), .Z(n592) );
  NAND U1150 ( .A(y[23]), .B(zin[22]), .Z(n591) );
  XOR U1151 ( .A(zin[22]), .B(y[23]), .Z(n589) );
  NAND U1152 ( .A(y[22]), .B(zin[21]), .Z(n588) );
  XOR U1153 ( .A(zin[21]), .B(y[22]), .Z(n586) );
  NAND U1154 ( .A(y[21]), .B(zin[20]), .Z(n585) );
  XOR U1155 ( .A(zin[20]), .B(y[21]), .Z(n583) );
  NAND U1156 ( .A(y[20]), .B(zin[19]), .Z(n582) );
  XOR U1157 ( .A(zin[19]), .B(y[20]), .Z(n580) );
  NAND U1158 ( .A(y[19]), .B(zin[18]), .Z(n579) );
  XOR U1159 ( .A(zin[18]), .B(y[19]), .Z(n577) );
  NAND U1160 ( .A(y[18]), .B(zin[17]), .Z(n576) );
  XOR U1161 ( .A(zin[17]), .B(y[18]), .Z(n574) );
  NAND U1162 ( .A(y[17]), .B(zin[16]), .Z(n573) );
  XOR U1163 ( .A(zin[16]), .B(y[17]), .Z(n571) );
  NAND U1164 ( .A(y[16]), .B(zin[15]), .Z(n570) );
  XOR U1165 ( .A(zin[15]), .B(y[16]), .Z(n568) );
  NAND U1166 ( .A(y[15]), .B(zin[14]), .Z(n567) );
  XOR U1167 ( .A(zin[14]), .B(y[15]), .Z(n565) );
  NAND U1168 ( .A(y[14]), .B(zin[13]), .Z(n564) );
  XOR U1169 ( .A(zin[13]), .B(y[14]), .Z(n562) );
  NAND U1170 ( .A(y[13]), .B(zin[12]), .Z(n561) );
  XOR U1171 ( .A(zin[12]), .B(y[13]), .Z(n559) );
  NAND U1172 ( .A(y[12]), .B(zin[11]), .Z(n558) );
  XOR U1173 ( .A(zin[11]), .B(y[12]), .Z(n556) );
  NAND U1174 ( .A(y[11]), .B(zin[10]), .Z(n555) );
  XOR U1175 ( .A(zin[10]), .B(y[11]), .Z(n553) );
  NAND U1176 ( .A(y[10]), .B(zin[9]), .Z(n552) );
  XOR U1177 ( .A(zin[9]), .B(y[10]), .Z(n550) );
  NAND U1178 ( .A(y[9]), .B(zin[8]), .Z(n549) );
  NAND U1179 ( .A(y[8]), .B(zin[7]), .Z(n546) );
  XOR U1180 ( .A(zin[7]), .B(y[8]), .Z(n544) );
  NAND U1181 ( .A(y[7]), .B(zin[6]), .Z(n543) );
  XOR U1182 ( .A(zin[6]), .B(y[7]), .Z(n541) );
  NAND U1183 ( .A(y[6]), .B(zin[5]), .Z(n540) );
  XOR U1184 ( .A(zin[5]), .B(y[6]), .Z(n538) );
  NAND U1185 ( .A(y[5]), .B(zin[4]), .Z(n537) );
  XOR U1186 ( .A(zin[4]), .B(y[5]), .Z(n535) );
  NAND U1187 ( .A(y[4]), .B(zin[3]), .Z(n534) );
  XOR U1188 ( .A(zin[3]), .B(y[4]), .Z(n532) );
  NAND U1189 ( .A(y[3]), .B(zin[2]), .Z(n531) );
  XOR U1190 ( .A(zin[2]), .B(y[3]), .Z(n529) );
  NAND U1191 ( .A(y[2]), .B(zin[1]), .Z(n528) );
  NAND U1192 ( .A(zin[0]), .B(y[1]), .Z(n2003) );
  XOR U1193 ( .A(zin[1]), .B(y[2]), .Z(n526) );
  NANDN U1194 ( .A(n2003), .B(n526), .Z(n527) );
  NAND U1195 ( .A(n528), .B(n527), .Z(n2000) );
  NAND U1196 ( .A(n529), .B(n2000), .Z(n530) );
  NAND U1197 ( .A(n531), .B(n530), .Z(n1997) );
  NAND U1198 ( .A(n532), .B(n1997), .Z(n533) );
  NAND U1199 ( .A(n534), .B(n533), .Z(n2019) );
  NAND U1200 ( .A(n535), .B(n2019), .Z(n536) );
  NAND U1201 ( .A(n537), .B(n536), .Z(n1994) );
  NAND U1202 ( .A(n538), .B(n1994), .Z(n539) );
  NAND U1203 ( .A(n540), .B(n539), .Z(n1991) );
  NAND U1204 ( .A(n541), .B(n1991), .Z(n542) );
  NAND U1205 ( .A(n543), .B(n542), .Z(n2028) );
  NAND U1206 ( .A(n544), .B(n2028), .Z(n545) );
  AND U1207 ( .A(n546), .B(n545), .Z(n2033) );
  XOR U1208 ( .A(zin[8]), .B(y[9]), .Z(n547) );
  NANDN U1209 ( .A(n2033), .B(n547), .Z(n548) );
  NAND U1210 ( .A(n549), .B(n548), .Z(n2036) );
  NAND U1211 ( .A(n550), .B(n2036), .Z(n551) );
  NAND U1212 ( .A(n552), .B(n551), .Z(n1988) );
  NAND U1213 ( .A(n553), .B(n1988), .Z(n554) );
  NAND U1214 ( .A(n555), .B(n554), .Z(n1984) );
  NAND U1215 ( .A(n556), .B(n1984), .Z(n557) );
  NAND U1216 ( .A(n558), .B(n557), .Z(n1981) );
  NAND U1217 ( .A(n559), .B(n1981), .Z(n560) );
  NAND U1218 ( .A(n561), .B(n560), .Z(n2050) );
  NAND U1219 ( .A(n562), .B(n2050), .Z(n563) );
  NAND U1220 ( .A(n564), .B(n563), .Z(n1978) );
  NAND U1221 ( .A(n565), .B(n1978), .Z(n566) );
  NAND U1222 ( .A(n567), .B(n566), .Z(n1975) );
  NAND U1223 ( .A(n568), .B(n1975), .Z(n569) );
  NAND U1224 ( .A(n570), .B(n569), .Z(n1972) );
  NAND U1225 ( .A(n571), .B(n1972), .Z(n572) );
  NAND U1226 ( .A(n573), .B(n572), .Z(n1969) );
  NAND U1227 ( .A(n574), .B(n1969), .Z(n575) );
  NAND U1228 ( .A(n576), .B(n575), .Z(n1966) );
  NAND U1229 ( .A(n577), .B(n1966), .Z(n578) );
  NAND U1230 ( .A(n579), .B(n578), .Z(n1963) );
  NAND U1231 ( .A(n580), .B(n1963), .Z(n581) );
  NAND U1232 ( .A(n582), .B(n581), .Z(n1960) );
  NAND U1233 ( .A(n583), .B(n1960), .Z(n584) );
  NAND U1234 ( .A(n585), .B(n584), .Z(n1957) );
  NAND U1235 ( .A(n586), .B(n1957), .Z(n587) );
  NAND U1236 ( .A(n588), .B(n587), .Z(n1954) );
  NAND U1237 ( .A(n589), .B(n1954), .Z(n590) );
  NAND U1238 ( .A(n591), .B(n590), .Z(n1951) );
  NAND U1239 ( .A(n592), .B(n1951), .Z(n593) );
  NAND U1240 ( .A(n594), .B(n593), .Z(n1948) );
  NAND U1241 ( .A(n595), .B(n1948), .Z(n596) );
  NAND U1242 ( .A(n597), .B(n596), .Z(n1945) );
  NAND U1243 ( .A(n598), .B(n1945), .Z(n599) );
  NAND U1244 ( .A(n600), .B(n599), .Z(n1942) );
  NAND U1245 ( .A(n601), .B(n1942), .Z(n602) );
  NAND U1246 ( .A(n603), .B(n602), .Z(n1939) );
  NAND U1247 ( .A(n604), .B(n1939), .Z(n605) );
  NAND U1248 ( .A(n606), .B(n605), .Z(n1936) );
  NAND U1249 ( .A(n607), .B(n1936), .Z(n608) );
  NAND U1250 ( .A(n609), .B(n608), .Z(n1933) );
  NAND U1251 ( .A(n610), .B(n1933), .Z(n611) );
  NAND U1252 ( .A(n612), .B(n611), .Z(n1930) );
  NAND U1253 ( .A(n613), .B(n1930), .Z(n614) );
  NAND U1254 ( .A(n615), .B(n614), .Z(n1927) );
  NAND U1255 ( .A(n616), .B(n1927), .Z(n617) );
  NAND U1256 ( .A(n618), .B(n617), .Z(n1924) );
  NAND U1257 ( .A(n619), .B(n1924), .Z(n620) );
  NAND U1258 ( .A(n621), .B(n620), .Z(n1921) );
  NAND U1259 ( .A(n622), .B(n1921), .Z(n623) );
  NAND U1260 ( .A(n624), .B(n623), .Z(n2119) );
  NAND U1261 ( .A(n625), .B(n2119), .Z(n626) );
  NAND U1262 ( .A(n627), .B(n626), .Z(n1918) );
  NAND U1263 ( .A(n628), .B(n1918), .Z(n629) );
  NAND U1264 ( .A(n630), .B(n629), .Z(n1915) );
  NAND U1265 ( .A(n631), .B(n1915), .Z(n632) );
  NAND U1266 ( .A(n633), .B(n632), .Z(n1912) );
  NAND U1267 ( .A(n634), .B(n1912), .Z(n635) );
  NAND U1268 ( .A(n636), .B(n635), .Z(n2134) );
  NAND U1269 ( .A(n637), .B(n2134), .Z(n638) );
  NAND U1270 ( .A(n639), .B(n638), .Z(n1909) );
  NAND U1271 ( .A(n640), .B(n1909), .Z(n641) );
  NAND U1272 ( .A(n642), .B(n641), .Z(n1906) );
  NAND U1273 ( .A(n643), .B(n1906), .Z(n644) );
  NAND U1274 ( .A(n645), .B(n644), .Z(n1903) );
  NAND U1275 ( .A(n646), .B(n1903), .Z(n647) );
  NAND U1276 ( .A(n648), .B(n647), .Z(n1900) );
  NAND U1277 ( .A(n649), .B(n1900), .Z(n650) );
  NAND U1278 ( .A(n651), .B(n650), .Z(n1897) );
  NAND U1279 ( .A(n652), .B(n1897), .Z(n653) );
  NAND U1280 ( .A(n654), .B(n653), .Z(n2149) );
  NAND U1281 ( .A(n655), .B(n2149), .Z(n656) );
  NAND U1282 ( .A(n657), .B(n656), .Z(n1894) );
  NAND U1283 ( .A(n658), .B(n1894), .Z(n659) );
  NAND U1284 ( .A(n660), .B(n659), .Z(n1891) );
  NAND U1285 ( .A(n661), .B(n1891), .Z(n662) );
  NAND U1286 ( .A(n663), .B(n662), .Z(n1888) );
  NAND U1287 ( .A(n664), .B(n1888), .Z(n665) );
  NAND U1288 ( .A(n666), .B(n665), .Z(n1885) );
  NAND U1289 ( .A(n667), .B(n1885), .Z(n668) );
  NAND U1290 ( .A(n669), .B(n668), .Z(n1882) );
  NAND U1291 ( .A(n670), .B(n1882), .Z(n671) );
  NAND U1292 ( .A(n672), .B(n671), .Z(n2167) );
  NAND U1293 ( .A(n673), .B(n2167), .Z(n674) );
  NAND U1294 ( .A(n675), .B(n674), .Z(n1879) );
  NAND U1295 ( .A(n676), .B(n1879), .Z(n677) );
  NAND U1296 ( .A(n678), .B(n677), .Z(n1876) );
  NAND U1297 ( .A(n679), .B(n1876), .Z(n680) );
  NAND U1298 ( .A(n681), .B(n680), .Z(n1873) );
  NAND U1299 ( .A(n682), .B(n1873), .Z(n683) );
  NAND U1300 ( .A(n684), .B(n683), .Z(n1870) );
  NAND U1301 ( .A(n685), .B(n1870), .Z(n686) );
  NAND U1302 ( .A(n687), .B(n686), .Z(n1867) );
  NAND U1303 ( .A(n688), .B(n1867), .Z(n689) );
  NAND U1304 ( .A(n690), .B(n689), .Z(n2186) );
  NAND U1305 ( .A(n691), .B(n2186), .Z(n692) );
  NAND U1306 ( .A(n693), .B(n692), .Z(n1861) );
  NAND U1307 ( .A(n694), .B(n1861), .Z(n695) );
  NAND U1308 ( .A(n696), .B(n695), .Z(n1864) );
  NAND U1309 ( .A(n697), .B(n1864), .Z(n698) );
  NAND U1310 ( .A(n699), .B(n698), .Z(n2197) );
  NAND U1311 ( .A(n700), .B(n2197), .Z(n701) );
  NAND U1312 ( .A(n702), .B(n701), .Z(n1858) );
  NAND U1313 ( .A(n703), .B(n1858), .Z(n704) );
  NAND U1314 ( .A(n705), .B(n704), .Z(n1855) );
  NAND U1315 ( .A(n706), .B(n1855), .Z(n707) );
  NAND U1316 ( .A(n708), .B(n707), .Z(n2206) );
  NAND U1317 ( .A(n709), .B(n2206), .Z(n710) );
  NAND U1318 ( .A(n711), .B(n710), .Z(n1852) );
  NAND U1319 ( .A(n712), .B(n1852), .Z(n713) );
  NAND U1320 ( .A(n714), .B(n713), .Z(n1849) );
  NAND U1321 ( .A(n715), .B(n1849), .Z(n716) );
  NAND U1322 ( .A(n717), .B(n716), .Z(n1846) );
  NAND U1323 ( .A(n718), .B(n1846), .Z(n719) );
  NAND U1324 ( .A(n720), .B(n719), .Z(n1839) );
  NAND U1325 ( .A(n721), .B(n1839), .Z(n722) );
  NAND U1326 ( .A(n723), .B(n722), .Z(n1842) );
  NAND U1327 ( .A(n724), .B(n1842), .Z(n725) );
  NAND U1328 ( .A(n726), .B(n725), .Z(n1836) );
  NAND U1329 ( .A(n727), .B(n1836), .Z(n728) );
  NAND U1330 ( .A(n729), .B(n728), .Z(n1833) );
  NAND U1331 ( .A(n730), .B(n1833), .Z(n731) );
  NAND U1332 ( .A(n732), .B(n731), .Z(n1830) );
  NAND U1333 ( .A(n733), .B(n1830), .Z(n734) );
  NAND U1334 ( .A(n735), .B(n734), .Z(n1827) );
  NAND U1335 ( .A(n736), .B(n1827), .Z(n737) );
  NAND U1336 ( .A(n738), .B(n737), .Z(n1824) );
  NAND U1337 ( .A(n739), .B(n1824), .Z(n740) );
  NAND U1338 ( .A(n741), .B(n740), .Z(n1821) );
  NAND U1339 ( .A(n742), .B(n1821), .Z(n743) );
  NAND U1340 ( .A(n744), .B(n743), .Z(n1818) );
  NAND U1341 ( .A(n745), .B(n1818), .Z(n746) );
  NAND U1342 ( .A(n747), .B(n746), .Z(n1815) );
  NAND U1343 ( .A(n748), .B(n1815), .Z(n749) );
  NAND U1344 ( .A(n750), .B(n749), .Z(n1812) );
  NAND U1345 ( .A(n751), .B(n1812), .Z(n752) );
  NAND U1346 ( .A(n753), .B(n752), .Z(n1809) );
  NAND U1347 ( .A(n754), .B(n1809), .Z(n755) );
  NAND U1348 ( .A(n756), .B(n755), .Z(n1806) );
  NAND U1349 ( .A(n757), .B(n1806), .Z(n758) );
  NAND U1350 ( .A(n759), .B(n758), .Z(n1803) );
  NAND U1351 ( .A(n760), .B(n1803), .Z(n761) );
  NAND U1352 ( .A(n762), .B(n761), .Z(n1800) );
  NAND U1353 ( .A(n763), .B(n1800), .Z(n764) );
  NAND U1354 ( .A(n765), .B(n764), .Z(n1797) );
  NAND U1355 ( .A(n766), .B(n1797), .Z(n767) );
  NAND U1356 ( .A(n768), .B(n767), .Z(n1794) );
  NAND U1357 ( .A(n769), .B(n1794), .Z(n770) );
  NAND U1358 ( .A(n771), .B(n770), .Z(n1791) );
  NAND U1359 ( .A(n772), .B(n1791), .Z(n773) );
  NAND U1360 ( .A(n774), .B(n773), .Z(n1788) );
  NAND U1361 ( .A(n775), .B(n1788), .Z(n776) );
  NAND U1362 ( .A(n777), .B(n776), .Z(n1785) );
  NAND U1363 ( .A(n778), .B(n1785), .Z(n779) );
  NAND U1364 ( .A(n780), .B(n779), .Z(n1782) );
  NAND U1365 ( .A(n781), .B(n1782), .Z(n782) );
  NAND U1366 ( .A(n783), .B(n782), .Z(n1779) );
  NAND U1367 ( .A(n784), .B(n1779), .Z(n785) );
  NAND U1368 ( .A(n786), .B(n785), .Z(n1776) );
  NAND U1369 ( .A(n787), .B(n1776), .Z(n788) );
  NAND U1370 ( .A(n789), .B(n788), .Z(n1773) );
  NAND U1371 ( .A(n790), .B(n1773), .Z(n791) );
  NAND U1372 ( .A(n792), .B(n791), .Z(n1770) );
  NAND U1373 ( .A(n793), .B(n1770), .Z(n794) );
  NAND U1374 ( .A(n795), .B(n794), .Z(n1767) );
  NAND U1375 ( .A(n796), .B(n1767), .Z(n797) );
  NAND U1376 ( .A(n798), .B(n797), .Z(n1764) );
  NAND U1377 ( .A(n799), .B(n1764), .Z(n800) );
  NAND U1378 ( .A(n801), .B(n800), .Z(n1761) );
  NAND U1379 ( .A(n802), .B(n1761), .Z(n803) );
  NAND U1380 ( .A(n804), .B(n803), .Z(n1758) );
  NAND U1381 ( .A(n805), .B(n1758), .Z(n806) );
  NAND U1382 ( .A(n807), .B(n806), .Z(n1755) );
  NAND U1383 ( .A(n808), .B(n1755), .Z(n809) );
  NAND U1384 ( .A(n810), .B(n809), .Z(n1752) );
  NAND U1385 ( .A(n811), .B(n1752), .Z(n812) );
  NAND U1386 ( .A(n813), .B(n812), .Z(n1749) );
  NAND U1387 ( .A(n814), .B(n1749), .Z(n815) );
  NAND U1388 ( .A(n816), .B(n815), .Z(n1746) );
  NAND U1389 ( .A(n817), .B(n1746), .Z(n818) );
  NAND U1390 ( .A(n819), .B(n818), .Z(n1743) );
  NAND U1391 ( .A(n820), .B(n1743), .Z(n821) );
  NAND U1392 ( .A(n822), .B(n821), .Z(n1740) );
  NAND U1393 ( .A(n823), .B(n1740), .Z(n824) );
  NAND U1394 ( .A(n825), .B(n824), .Z(n1737) );
  NAND U1395 ( .A(n826), .B(n1737), .Z(n827) );
  NAND U1396 ( .A(n828), .B(n827), .Z(n1734) );
  NAND U1397 ( .A(n829), .B(n1734), .Z(n830) );
  NAND U1398 ( .A(n831), .B(n830), .Z(n1731) );
  NAND U1399 ( .A(n832), .B(n1731), .Z(n833) );
  NAND U1400 ( .A(n834), .B(n833), .Z(n1728) );
  NAND U1401 ( .A(n835), .B(n1728), .Z(n836) );
  NAND U1402 ( .A(n837), .B(n836), .Z(n1725) );
  NAND U1403 ( .A(n838), .B(n1725), .Z(n839) );
  NAND U1404 ( .A(n840), .B(n839), .Z(n1722) );
  NAND U1405 ( .A(n841), .B(n1722), .Z(n842) );
  NAND U1406 ( .A(n843), .B(n842), .Z(n1719) );
  NAND U1407 ( .A(n844), .B(n1719), .Z(n845) );
  NAND U1408 ( .A(n846), .B(n845), .Z(n1716) );
  NAND U1409 ( .A(n847), .B(n1716), .Z(n848) );
  NAND U1410 ( .A(n849), .B(n848), .Z(n1713) );
  NAND U1411 ( .A(n850), .B(n1713), .Z(n851) );
  NAND U1412 ( .A(n852), .B(n851), .Z(n1710) );
  NAND U1413 ( .A(n853), .B(n1710), .Z(n854) );
  NAND U1414 ( .A(n855), .B(n854), .Z(n1707) );
  NAND U1415 ( .A(n856), .B(n1707), .Z(n857) );
  NAND U1416 ( .A(n858), .B(n857), .Z(n1704) );
  NAND U1417 ( .A(n859), .B(n1704), .Z(n860) );
  NAND U1418 ( .A(n861), .B(n860), .Z(n1701) );
  NAND U1419 ( .A(n862), .B(n1701), .Z(n863) );
  NAND U1420 ( .A(n864), .B(n863), .Z(n1698) );
  NAND U1421 ( .A(n865), .B(n1698), .Z(n866) );
  NAND U1422 ( .A(n867), .B(n866), .Z(n1695) );
  NAND U1423 ( .A(n868), .B(n1695), .Z(n869) );
  NAND U1424 ( .A(n870), .B(n869), .Z(n1692) );
  NAND U1425 ( .A(n871), .B(n1692), .Z(n872) );
  NAND U1426 ( .A(n873), .B(n872), .Z(n1689) );
  NAND U1427 ( .A(n874), .B(n1689), .Z(n875) );
  NAND U1428 ( .A(n876), .B(n875), .Z(n1686) );
  NAND U1429 ( .A(n877), .B(n1686), .Z(n878) );
  NAND U1430 ( .A(n879), .B(n878), .Z(n1683) );
  NAND U1431 ( .A(n880), .B(n1683), .Z(n881) );
  NAND U1432 ( .A(n882), .B(n881), .Z(n1680) );
  NAND U1433 ( .A(n883), .B(n1680), .Z(n884) );
  NAND U1434 ( .A(n885), .B(n884), .Z(n1677) );
  NAND U1435 ( .A(n886), .B(n1677), .Z(n887) );
  NAND U1436 ( .A(n888), .B(n887), .Z(n1674) );
  NAND U1437 ( .A(n889), .B(n1674), .Z(n890) );
  NAND U1438 ( .A(n891), .B(n890), .Z(n1671) );
  NAND U1439 ( .A(n892), .B(n1671), .Z(n893) );
  NAND U1440 ( .A(n894), .B(n893), .Z(n1668) );
  NAND U1441 ( .A(n895), .B(n1668), .Z(n896) );
  NAND U1442 ( .A(n897), .B(n896), .Z(n1665) );
  NAND U1443 ( .A(n898), .B(n1665), .Z(n899) );
  NAND U1444 ( .A(n900), .B(n899), .Z(n1662) );
  NAND U1445 ( .A(n901), .B(n1662), .Z(n902) );
  NAND U1446 ( .A(n903), .B(n902), .Z(n1659) );
  NAND U1447 ( .A(n904), .B(n1659), .Z(n905) );
  NAND U1448 ( .A(n906), .B(n905), .Z(n1656) );
  NAND U1449 ( .A(n907), .B(n1656), .Z(n908) );
  NAND U1450 ( .A(n909), .B(n908), .Z(n1653) );
  NAND U1451 ( .A(n910), .B(n1653), .Z(n911) );
  NAND U1452 ( .A(n912), .B(n911), .Z(n1650) );
  NAND U1453 ( .A(n913), .B(n1650), .Z(n914) );
  NAND U1454 ( .A(n915), .B(n914), .Z(n1647) );
  NAND U1455 ( .A(n916), .B(n1647), .Z(n917) );
  NAND U1456 ( .A(n918), .B(n917), .Z(n1644) );
  NAND U1457 ( .A(n919), .B(n1644), .Z(n920) );
  NAND U1458 ( .A(n921), .B(n920), .Z(n1641) );
  NAND U1459 ( .A(n922), .B(n1641), .Z(n923) );
  NAND U1460 ( .A(n924), .B(n923), .Z(n1638) );
  NAND U1461 ( .A(n925), .B(n1638), .Z(n926) );
  NAND U1462 ( .A(n927), .B(n926), .Z(n1635) );
  NAND U1463 ( .A(n928), .B(n1635), .Z(n929) );
  NAND U1464 ( .A(n930), .B(n929), .Z(n1632) );
  NAND U1465 ( .A(n931), .B(n1632), .Z(n932) );
  NAND U1466 ( .A(n933), .B(n932), .Z(n1629) );
  NAND U1467 ( .A(n934), .B(n1629), .Z(n935) );
  NAND U1468 ( .A(n936), .B(n935), .Z(n1626) );
  NAND U1469 ( .A(n937), .B(n1626), .Z(n938) );
  NAND U1470 ( .A(n939), .B(n938), .Z(n1623) );
  NAND U1471 ( .A(n940), .B(n1623), .Z(n941) );
  NAND U1472 ( .A(n942), .B(n941), .Z(n1620) );
  NAND U1473 ( .A(n943), .B(n1620), .Z(n944) );
  NAND U1474 ( .A(n945), .B(n944), .Z(n1617) );
  NAND U1475 ( .A(n946), .B(n1617), .Z(n947) );
  NAND U1476 ( .A(n948), .B(n947), .Z(n1614) );
  NAND U1477 ( .A(n949), .B(n1614), .Z(n950) );
  NAND U1478 ( .A(n951), .B(n950), .Z(n1611) );
  NAND U1479 ( .A(n952), .B(n1611), .Z(n953) );
  NAND U1480 ( .A(n954), .B(n953), .Z(n1608) );
  NAND U1481 ( .A(n955), .B(n1608), .Z(n956) );
  NAND U1482 ( .A(n957), .B(n956), .Z(n1605) );
  NAND U1483 ( .A(n958), .B(n1605), .Z(n959) );
  NAND U1484 ( .A(n960), .B(n959), .Z(n1602) );
  NAND U1485 ( .A(n961), .B(n1602), .Z(n962) );
  NAND U1486 ( .A(n963), .B(n962), .Z(n1599) );
  NAND U1487 ( .A(n964), .B(n1599), .Z(n965) );
  NAND U1488 ( .A(n966), .B(n965), .Z(n1596) );
  NAND U1489 ( .A(n967), .B(n1596), .Z(n968) );
  NAND U1490 ( .A(n969), .B(n968), .Z(n1593) );
  NAND U1491 ( .A(n970), .B(n1593), .Z(n971) );
  NAND U1492 ( .A(n972), .B(n971), .Z(n1590) );
  NAND U1493 ( .A(n973), .B(n1590), .Z(n974) );
  NAND U1494 ( .A(n975), .B(n974), .Z(n1587) );
  NAND U1495 ( .A(n976), .B(n1587), .Z(n977) );
  NAND U1496 ( .A(n978), .B(n977), .Z(n1584) );
  NAND U1497 ( .A(n979), .B(n1584), .Z(n980) );
  NAND U1498 ( .A(n981), .B(n980), .Z(n1581) );
  NAND U1499 ( .A(n982), .B(n1581), .Z(n983) );
  NAND U1500 ( .A(n984), .B(n983), .Z(n1578) );
  NAND U1501 ( .A(n985), .B(n1578), .Z(n986) );
  NAND U1502 ( .A(n987), .B(n986), .Z(n1575) );
  NAND U1503 ( .A(n988), .B(n1575), .Z(n989) );
  NAND U1504 ( .A(n990), .B(n989), .Z(n1572) );
  NAND U1505 ( .A(n991), .B(n1572), .Z(n992) );
  NAND U1506 ( .A(n993), .B(n992), .Z(n1569) );
  NAND U1507 ( .A(n994), .B(n1569), .Z(n995) );
  NAND U1508 ( .A(n996), .B(n995), .Z(n1566) );
  NAND U1509 ( .A(n997), .B(n1566), .Z(n998) );
  NAND U1510 ( .A(n999), .B(n998), .Z(n1563) );
  NAND U1511 ( .A(n1000), .B(n1563), .Z(n1001) );
  NAND U1512 ( .A(n1002), .B(n1001), .Z(n1560) );
  NAND U1513 ( .A(n1003), .B(n1560), .Z(n1004) );
  NAND U1514 ( .A(n1005), .B(n1004), .Z(n1557) );
  NAND U1515 ( .A(n1006), .B(n1557), .Z(n1007) );
  NAND U1516 ( .A(n1008), .B(n1007), .Z(n1554) );
  NAND U1517 ( .A(n1009), .B(n1554), .Z(n1010) );
  NAND U1518 ( .A(n1011), .B(n1010), .Z(n1551) );
  NAND U1519 ( .A(n1012), .B(n1551), .Z(n1013) );
  NAND U1520 ( .A(n1014), .B(n1013), .Z(n1548) );
  NAND U1521 ( .A(n1015), .B(n1548), .Z(n1016) );
  NAND U1522 ( .A(n1017), .B(n1016), .Z(n1545) );
  NAND U1523 ( .A(n1018), .B(n1545), .Z(n1019) );
  NAND U1524 ( .A(n1020), .B(n1019), .Z(n1542) );
  NAND U1525 ( .A(n1021), .B(n1542), .Z(n1022) );
  NAND U1526 ( .A(n1023), .B(n1022), .Z(n1539) );
  NAND U1527 ( .A(n1024), .B(n1539), .Z(n1025) );
  NAND U1528 ( .A(n1026), .B(n1025), .Z(n1536) );
  NAND U1529 ( .A(n1027), .B(n1536), .Z(n1028) );
  NAND U1530 ( .A(n1029), .B(n1028), .Z(n1533) );
  NAND U1531 ( .A(n1030), .B(n1533), .Z(n1031) );
  NAND U1532 ( .A(n1032), .B(n1031), .Z(n1530) );
  NAND U1533 ( .A(n1033), .B(n1530), .Z(n1034) );
  NAND U1534 ( .A(n1035), .B(n1034), .Z(n1527) );
  NAND U1535 ( .A(n1036), .B(n1527), .Z(n1037) );
  NAND U1536 ( .A(n1038), .B(n1037), .Z(n1524) );
  NAND U1537 ( .A(n1039), .B(n1524), .Z(n1040) );
  NAND U1538 ( .A(n1041), .B(n1040), .Z(n1521) );
  NAND U1539 ( .A(n1042), .B(n1521), .Z(n1043) );
  NAND U1540 ( .A(n1044), .B(n1043), .Z(n1518) );
  NAND U1541 ( .A(n1045), .B(n1518), .Z(n1046) );
  NAND U1542 ( .A(n1047), .B(n1046), .Z(n1515) );
  NAND U1543 ( .A(n1048), .B(n1515), .Z(n1049) );
  NAND U1544 ( .A(n1050), .B(n1049), .Z(n1512) );
  NAND U1545 ( .A(n1051), .B(n1512), .Z(n1052) );
  NAND U1546 ( .A(n1053), .B(n1052), .Z(n1509) );
  NAND U1547 ( .A(n1054), .B(n1509), .Z(n1055) );
  NAND U1548 ( .A(n1056), .B(n1055), .Z(n1506) );
  NAND U1549 ( .A(n1057), .B(n1506), .Z(n1058) );
  NAND U1550 ( .A(n1059), .B(n1058), .Z(n1503) );
  NAND U1551 ( .A(n1060), .B(n1503), .Z(n1061) );
  NAND U1552 ( .A(n1062), .B(n1061), .Z(n1500) );
  NAND U1553 ( .A(n1063), .B(n1500), .Z(n1064) );
  NAND U1554 ( .A(n1065), .B(n1064), .Z(n1497) );
  NAND U1555 ( .A(n1066), .B(n1497), .Z(n1067) );
  NAND U1556 ( .A(n1068), .B(n1067), .Z(n1494) );
  NAND U1557 ( .A(n1069), .B(n1494), .Z(n1070) );
  NAND U1558 ( .A(n1071), .B(n1070), .Z(n1491) );
  NAND U1559 ( .A(n1072), .B(n1491), .Z(n1073) );
  NAND U1560 ( .A(n1074), .B(n1073), .Z(n1488) );
  NAND U1561 ( .A(n1075), .B(n1488), .Z(n1076) );
  NAND U1562 ( .A(n1077), .B(n1076), .Z(n1485) );
  NAND U1563 ( .A(n1078), .B(n1485), .Z(n1079) );
  NAND U1564 ( .A(n1080), .B(n1079), .Z(n1482) );
  NAND U1565 ( .A(n1081), .B(n1482), .Z(n1082) );
  NAND U1566 ( .A(n1083), .B(n1082), .Z(n1479) );
  NAND U1567 ( .A(n1084), .B(n1479), .Z(n1085) );
  NAND U1568 ( .A(n1086), .B(n1085), .Z(n1476) );
  NAND U1569 ( .A(n1087), .B(n1476), .Z(n1088) );
  NAND U1570 ( .A(n1089), .B(n1088), .Z(n1473) );
  NAND U1571 ( .A(n1090), .B(n1473), .Z(n1091) );
  NAND U1572 ( .A(n1092), .B(n1091), .Z(n1470) );
  NAND U1573 ( .A(n1093), .B(n1470), .Z(n1094) );
  NAND U1574 ( .A(n1095), .B(n1094), .Z(n1467) );
  NAND U1575 ( .A(n1096), .B(n1467), .Z(n1097) );
  NAND U1576 ( .A(n1098), .B(n1097), .Z(n1464) );
  NAND U1577 ( .A(n1099), .B(n1464), .Z(n1100) );
  NAND U1578 ( .A(n1101), .B(n1100), .Z(n1461) );
  NAND U1579 ( .A(n1102), .B(n1461), .Z(n1103) );
  NAND U1580 ( .A(n1104), .B(n1103), .Z(n1458) );
  NAND U1581 ( .A(n1105), .B(n1458), .Z(n1106) );
  NAND U1582 ( .A(n1107), .B(n1106), .Z(n1455) );
  NAND U1583 ( .A(n1108), .B(n1455), .Z(n1109) );
  NAND U1584 ( .A(n1110), .B(n1109), .Z(n1452) );
  NAND U1585 ( .A(n1111), .B(n1452), .Z(n1112) );
  NAND U1586 ( .A(n1113), .B(n1112), .Z(n1449) );
  NAND U1587 ( .A(n1114), .B(n1449), .Z(n1115) );
  NAND U1588 ( .A(n1116), .B(n1115), .Z(n1446) );
  NAND U1589 ( .A(n1117), .B(n1446), .Z(n1118) );
  NAND U1590 ( .A(n1119), .B(n1118), .Z(n1443) );
  NAND U1591 ( .A(n1120), .B(n1443), .Z(n1121) );
  NAND U1592 ( .A(n1122), .B(n1121), .Z(n1440) );
  NAND U1593 ( .A(n1123), .B(n1440), .Z(n1124) );
  NAND U1594 ( .A(n1125), .B(n1124), .Z(n1437) );
  NAND U1595 ( .A(n1126), .B(n1437), .Z(n1127) );
  NAND U1596 ( .A(n1128), .B(n1127), .Z(n1434) );
  NAND U1597 ( .A(n1129), .B(n1434), .Z(n1130) );
  NAND U1598 ( .A(n1131), .B(n1130), .Z(n1431) );
  NAND U1599 ( .A(n1132), .B(n1431), .Z(n1133) );
  NAND U1600 ( .A(n1134), .B(n1133), .Z(n1428) );
  NAND U1601 ( .A(n1135), .B(n1428), .Z(n1136) );
  NAND U1602 ( .A(n1137), .B(n1136), .Z(n1425) );
  NAND U1603 ( .A(n1138), .B(n1425), .Z(n1139) );
  NAND U1604 ( .A(n1140), .B(n1139), .Z(n1422) );
  NAND U1605 ( .A(n1141), .B(n1422), .Z(n1142) );
  NAND U1606 ( .A(n1143), .B(n1142), .Z(n1419) );
  NAND U1607 ( .A(n1144), .B(n1419), .Z(n1145) );
  NAND U1608 ( .A(n1146), .B(n1145), .Z(n1416) );
  NAND U1609 ( .A(n1147), .B(n1416), .Z(n1148) );
  NAND U1610 ( .A(n1149), .B(n1148), .Z(n1413) );
  NAND U1611 ( .A(n1150), .B(n1413), .Z(n1151) );
  NAND U1612 ( .A(n1152), .B(n1151), .Z(n1410) );
  NAND U1613 ( .A(n1153), .B(n1410), .Z(n1154) );
  NAND U1614 ( .A(n1155), .B(n1154), .Z(n1407) );
  NAND U1615 ( .A(n1156), .B(n1407), .Z(n1157) );
  NAND U1616 ( .A(n1158), .B(n1157), .Z(n1404) );
  NAND U1617 ( .A(n1159), .B(n1404), .Z(n1160) );
  NAND U1618 ( .A(n1161), .B(n1160), .Z(n1401) );
  NAND U1619 ( .A(n1162), .B(n1401), .Z(n1163) );
  NAND U1620 ( .A(n1164), .B(n1163), .Z(n1398) );
  NAND U1621 ( .A(n1165), .B(n1398), .Z(n1166) );
  NAND U1622 ( .A(n1167), .B(n1166), .Z(n1395) );
  NAND U1623 ( .A(n1168), .B(n1395), .Z(n1169) );
  NAND U1624 ( .A(n1170), .B(n1169), .Z(n1392) );
  NAND U1625 ( .A(n1171), .B(n1392), .Z(n1172) );
  NAND U1626 ( .A(n1173), .B(n1172), .Z(n1389) );
  NAND U1627 ( .A(n1174), .B(n1389), .Z(n1175) );
  NAND U1628 ( .A(n1176), .B(n1175), .Z(n1386) );
  NAND U1629 ( .A(n1177), .B(n1386), .Z(n1178) );
  NAND U1630 ( .A(n1179), .B(n1178), .Z(n1383) );
  NAND U1631 ( .A(n1180), .B(n1383), .Z(n1181) );
  NAND U1632 ( .A(n1182), .B(n1181), .Z(n1380) );
  NAND U1633 ( .A(n1183), .B(n1380), .Z(n1184) );
  NAND U1634 ( .A(n1185), .B(n1184), .Z(n1377) );
  NAND U1635 ( .A(n1186), .B(n1377), .Z(n1187) );
  NAND U1636 ( .A(n1188), .B(n1187), .Z(n1374) );
  NAND U1637 ( .A(n1189), .B(n1374), .Z(n1190) );
  NAND U1638 ( .A(n1191), .B(n1190), .Z(n1371) );
  NAND U1639 ( .A(n1192), .B(n1371), .Z(n1193) );
  NAND U1640 ( .A(n1194), .B(n1193), .Z(n1368) );
  NAND U1641 ( .A(n1195), .B(n1368), .Z(n1196) );
  NAND U1642 ( .A(n1197), .B(n1196), .Z(n1365) );
  NAND U1643 ( .A(n1198), .B(n1365), .Z(n1199) );
  NAND U1644 ( .A(n1200), .B(n1199), .Z(n1362) );
  NAND U1645 ( .A(n1201), .B(n1362), .Z(n1202) );
  NAND U1646 ( .A(n1203), .B(n1202), .Z(n1359) );
  NAND U1647 ( .A(n1204), .B(n1359), .Z(n1205) );
  NAND U1648 ( .A(n1206), .B(n1205), .Z(n1356) );
  NAND U1649 ( .A(n1207), .B(n1356), .Z(n1208) );
  NAND U1650 ( .A(n1209), .B(n1208), .Z(n1353) );
  NAND U1651 ( .A(n1210), .B(n1353), .Z(n1211) );
  NAND U1652 ( .A(n1212), .B(n1211), .Z(n1350) );
  NAND U1653 ( .A(n1213), .B(n1350), .Z(n1214) );
  NAND U1654 ( .A(n1215), .B(n1214), .Z(n1347) );
  NAND U1655 ( .A(n1216), .B(n1347), .Z(n1217) );
  NAND U1656 ( .A(n1218), .B(n1217), .Z(n1344) );
  NAND U1657 ( .A(n1219), .B(n1344), .Z(n1220) );
  NAND U1658 ( .A(n1221), .B(n1220), .Z(n1341) );
  NAND U1659 ( .A(n1222), .B(n1341), .Z(n1223) );
  NAND U1660 ( .A(n1224), .B(n1223), .Z(n1338) );
  NAND U1661 ( .A(n1225), .B(n1338), .Z(n1226) );
  NAND U1662 ( .A(n1227), .B(n1226), .Z(n1335) );
  NAND U1663 ( .A(n1228), .B(n1335), .Z(n1229) );
  NAND U1664 ( .A(n1230), .B(n1229), .Z(n1332) );
  NAND U1665 ( .A(n1231), .B(n1332), .Z(n1232) );
  NAND U1666 ( .A(n1233), .B(n1232), .Z(n1329) );
  NAND U1667 ( .A(n1234), .B(n1329), .Z(n1235) );
  NAND U1668 ( .A(n1236), .B(n1235), .Z(n1326) );
  NAND U1669 ( .A(n1237), .B(n1326), .Z(n1238) );
  NAND U1670 ( .A(n1239), .B(n1238), .Z(n1323) );
  NAND U1671 ( .A(n1240), .B(n1323), .Z(n1241) );
  NAND U1672 ( .A(n1242), .B(n1241), .Z(n1320) );
  NAND U1673 ( .A(n1243), .B(n1320), .Z(n1244) );
  NAND U1674 ( .A(n1245), .B(n1244), .Z(n1317) );
  NAND U1675 ( .A(n1246), .B(n1317), .Z(n1247) );
  NAND U1676 ( .A(n1248), .B(n1247), .Z(n1314) );
  NAND U1677 ( .A(n1249), .B(n1314), .Z(n1250) );
  NAND U1678 ( .A(n1251), .B(n1250), .Z(n1311) );
  NAND U1679 ( .A(n1252), .B(n1311), .Z(n1253) );
  NAND U1680 ( .A(n1254), .B(n1253), .Z(n1308) );
  NAND U1681 ( .A(n1255), .B(n1308), .Z(n1256) );
  NAND U1682 ( .A(n1257), .B(n1256), .Z(n1305) );
  NAND U1683 ( .A(n1258), .B(n1305), .Z(n1259) );
  NAND U1684 ( .A(n1260), .B(n1259), .Z(n1302) );
  NAND U1685 ( .A(n1261), .B(n1302), .Z(n1262) );
  NAND U1686 ( .A(n1263), .B(n1262), .Z(n1299) );
  NAND U1687 ( .A(n1264), .B(n1299), .Z(n1265) );
  NAND U1688 ( .A(n1266), .B(n1265), .Z(n1296) );
  NAND U1689 ( .A(n1267), .B(n1296), .Z(n1268) );
  NAND U1690 ( .A(n1269), .B(n1268), .Z(n1293) );
  NAND U1691 ( .A(n1270), .B(n1293), .Z(n1271) );
  NAND U1692 ( .A(n1272), .B(n1271), .Z(n1290) );
  NAND U1693 ( .A(n1273), .B(n1290), .Z(n1274) );
  NAND U1694 ( .A(n1275), .B(n1274), .Z(n1287) );
  NAND U1695 ( .A(n1276), .B(n1287), .Z(n1277) );
  NAND U1696 ( .A(n1278), .B(n1277), .Z(n1284) );
  NAND U1697 ( .A(n1279), .B(n1284), .Z(n1280) );
  NAND U1698 ( .A(n1281), .B(n1280), .Z(n2857) );
  XOR U1699 ( .A(y[254]), .B(n2857), .Z(n1282) );
  IV U1700 ( .A(xregN_1), .Z(n2868) );
  ANDN U1701 ( .B(n1282), .A(n2868), .Z(n1283) );
  XNOR U1702 ( .A(zin[253]), .B(n1283), .Z(n3318) );
  NANDN U1703 ( .A(n6582), .B(n3318), .Z(n3303) );
  XOR U1704 ( .A(y[253]), .B(n1284), .Z(n1285) );
  ANDN U1705 ( .B(n1285), .A(n2868), .Z(n1286) );
  XNOR U1706 ( .A(zin[252]), .B(n1286), .Z(n3322) );
  IV U1707 ( .A(n[252]), .Z(n3327) );
  XOR U1708 ( .A(y[252]), .B(n1287), .Z(n1288) );
  ANDN U1709 ( .B(n1288), .A(n2868), .Z(n1289) );
  XNOR U1710 ( .A(zin[251]), .B(n1289), .Z(n3326) );
  NANDN U1711 ( .A(n3327), .B(n3326), .Z(n3300) );
  XOR U1712 ( .A(y[251]), .B(n1290), .Z(n1291) );
  ANDN U1713 ( .B(n1291), .A(n2868), .Z(n1292) );
  XNOR U1714 ( .A(zin[250]), .B(n1292), .Z(n3331) );
  XOR U1715 ( .A(n3331), .B(n[251]), .Z(n2856) );
  XOR U1716 ( .A(y[250]), .B(n1293), .Z(n1294) );
  ANDN U1717 ( .B(n1294), .A(n2868), .Z(n1295) );
  XNOR U1718 ( .A(zin[249]), .B(n1295), .Z(n3335) );
  NAND U1719 ( .A(n3335), .B(n[250]), .Z(n2854) );
  XOR U1720 ( .A(n[250]), .B(n3335), .Z(n2852) );
  IV U1721 ( .A(n[249]), .Z(n6534) );
  XOR U1722 ( .A(y[249]), .B(n1296), .Z(n1297) );
  ANDN U1723 ( .B(n1297), .A(n2868), .Z(n1298) );
  XNOR U1724 ( .A(zin[248]), .B(n1298), .Z(n3339) );
  NANDN U1725 ( .A(n6534), .B(n3339), .Z(n3297) );
  XNOR U1726 ( .A(n6534), .B(n3339), .Z(n2849) );
  XOR U1727 ( .A(y[248]), .B(n1299), .Z(n1300) );
  ANDN U1728 ( .B(n1300), .A(n2868), .Z(n1301) );
  XNOR U1729 ( .A(zin[247]), .B(n1301), .Z(n3343) );
  NAND U1730 ( .A(n3343), .B(n[248]), .Z(n2847) );
  XOR U1731 ( .A(n[248]), .B(n3343), .Z(n2845) );
  IV U1732 ( .A(n[247]), .Z(n3348) );
  XOR U1733 ( .A(y[247]), .B(n1302), .Z(n1303) );
  ANDN U1734 ( .B(n1303), .A(n2868), .Z(n1304) );
  XNOR U1735 ( .A(zin[246]), .B(n1304), .Z(n3347) );
  NANDN U1736 ( .A(n3348), .B(n3347), .Z(n3294) );
  XNOR U1737 ( .A(n3348), .B(n3347), .Z(n2842) );
  IV U1738 ( .A(n[246]), .Z(n6514) );
  XOR U1739 ( .A(y[246]), .B(n1305), .Z(n1306) );
  ANDN U1740 ( .B(n1306), .A(n2868), .Z(n1307) );
  XNOR U1741 ( .A(zin[245]), .B(n1307), .Z(n3352) );
  NANDN U1742 ( .A(n6514), .B(n3352), .Z(n3291) );
  XNOR U1743 ( .A(n3352), .B(n6514), .Z(n2839) );
  XOR U1744 ( .A(y[245]), .B(n1308), .Z(n1309) );
  ANDN U1745 ( .B(n1309), .A(n2868), .Z(n1310) );
  XNOR U1746 ( .A(zin[244]), .B(n1310), .Z(n3356) );
  NAND U1747 ( .A(n[245]), .B(n3356), .Z(n3288) );
  XOR U1748 ( .A(n[245]), .B(n3356), .Z(n2836) );
  IV U1749 ( .A(n[244]), .Z(n3361) );
  XOR U1750 ( .A(y[244]), .B(n1311), .Z(n1312) );
  ANDN U1751 ( .B(n1312), .A(n2868), .Z(n1313) );
  XNOR U1752 ( .A(zin[243]), .B(n1313), .Z(n3360) );
  NANDN U1753 ( .A(n3361), .B(n3360), .Z(n3285) );
  XNOR U1754 ( .A(n3360), .B(n3361), .Z(n2833) );
  XOR U1755 ( .A(y[243]), .B(n1314), .Z(n1315) );
  ANDN U1756 ( .B(n1315), .A(n2868), .Z(n1316) );
  XNOR U1757 ( .A(zin[242]), .B(n1316), .Z(n3365) );
  NAND U1758 ( .A(n[243]), .B(n3365), .Z(n2831) );
  XOR U1759 ( .A(n3365), .B(n[243]), .Z(n2829) );
  XOR U1760 ( .A(y[242]), .B(n1317), .Z(n1318) );
  ANDN U1761 ( .B(n1318), .A(n2868), .Z(n1319) );
  XNOR U1762 ( .A(zin[241]), .B(n1319), .Z(n3369) );
  NAND U1763 ( .A(n3369), .B(n[242]), .Z(n2827) );
  XOR U1764 ( .A(n[242]), .B(n3369), .Z(n2825) );
  XOR U1765 ( .A(y[241]), .B(n1320), .Z(n1321) );
  ANDN U1766 ( .B(n1321), .A(n2868), .Z(n1322) );
  XNOR U1767 ( .A(zin[240]), .B(n1322), .Z(n3373) );
  NAND U1768 ( .A(n[241]), .B(n3373), .Z(n2823) );
  XOR U1769 ( .A(n3373), .B(n[241]), .Z(n2821) );
  XOR U1770 ( .A(y[240]), .B(n1323), .Z(n1324) );
  ANDN U1771 ( .B(n1324), .A(n2868), .Z(n1325) );
  XNOR U1772 ( .A(zin[239]), .B(n1325), .Z(n3377) );
  NAND U1773 ( .A(n3377), .B(n[240]), .Z(n2819) );
  XOR U1774 ( .A(n[240]), .B(n3377), .Z(n2817) );
  IV U1775 ( .A(n[239]), .Z(n3382) );
  XOR U1776 ( .A(y[239]), .B(n1326), .Z(n1327) );
  ANDN U1777 ( .B(n1327), .A(n2868), .Z(n1328) );
  XNOR U1778 ( .A(zin[238]), .B(n1328), .Z(n3381) );
  NANDN U1779 ( .A(n3382), .B(n3381), .Z(n3282) );
  XNOR U1780 ( .A(n3382), .B(n3381), .Z(n2814) );
  XOR U1781 ( .A(y[238]), .B(n1329), .Z(n1330) );
  ANDN U1782 ( .B(n1330), .A(n2868), .Z(n1331) );
  XNOR U1783 ( .A(zin[237]), .B(n1331), .Z(n3386) );
  NAND U1784 ( .A(n3386), .B(n[238]), .Z(n2812) );
  XOR U1785 ( .A(n[238]), .B(n3386), .Z(n2810) );
  IV U1786 ( .A(n[237]), .Z(n6456) );
  XOR U1787 ( .A(y[237]), .B(n1332), .Z(n1333) );
  ANDN U1788 ( .B(n1333), .A(n2868), .Z(n1334) );
  XNOR U1789 ( .A(zin[236]), .B(n1334), .Z(n5260) );
  NANDN U1790 ( .A(n6456), .B(n5260), .Z(n2808) );
  XNOR U1791 ( .A(n5260), .B(n6456), .Z(n2806) );
  IV U1792 ( .A(n[236]), .Z(n6449) );
  XOR U1793 ( .A(y[236]), .B(n1335), .Z(n1336) );
  ANDN U1794 ( .B(n1336), .A(n2868), .Z(n1337) );
  XNOR U1795 ( .A(zin[235]), .B(n1337), .Z(n3390) );
  NANDN U1796 ( .A(n6449), .B(n3390), .Z(n2804) );
  XNOR U1797 ( .A(n6449), .B(n3390), .Z(n2802) );
  XOR U1798 ( .A(y[235]), .B(n1338), .Z(n1339) );
  ANDN U1799 ( .B(n1339), .A(n2868), .Z(n1340) );
  XNOR U1800 ( .A(zin[234]), .B(n1340), .Z(n3394) );
  NAND U1801 ( .A(n[235]), .B(n3394), .Z(n2800) );
  XOR U1802 ( .A(n3394), .B(n[235]), .Z(n2798) );
  IV U1803 ( .A(n[234]), .Z(n3399) );
  XOR U1804 ( .A(y[234]), .B(n1341), .Z(n1342) );
  ANDN U1805 ( .B(n1342), .A(n2868), .Z(n1343) );
  XOR U1806 ( .A(zin[233]), .B(n1343), .Z(n3398) );
  IV U1807 ( .A(n3398), .Z(n2872) );
  NANDN U1808 ( .A(n3399), .B(n2872), .Z(n2796) );
  XNOR U1809 ( .A(n3398), .B(n[234]), .Z(n2794) );
  XOR U1810 ( .A(y[233]), .B(n1344), .Z(n1345) );
  ANDN U1811 ( .B(n1345), .A(n2868), .Z(n1346) );
  XNOR U1812 ( .A(zin[232]), .B(n1346), .Z(n3403) );
  NAND U1813 ( .A(n[233]), .B(n3403), .Z(n2792) );
  XOR U1814 ( .A(n3403), .B(n[233]), .Z(n2790) );
  XOR U1815 ( .A(y[232]), .B(n1347), .Z(n1348) );
  ANDN U1816 ( .B(n1348), .A(n2868), .Z(n1349) );
  XNOR U1817 ( .A(zin[231]), .B(n1349), .Z(n3407) );
  NAND U1818 ( .A(n3407), .B(n[232]), .Z(n2788) );
  XOR U1819 ( .A(n[232]), .B(n3407), .Z(n2786) );
  IV U1820 ( .A(n[231]), .Z(n6413) );
  XOR U1821 ( .A(y[231]), .B(n1350), .Z(n1351) );
  ANDN U1822 ( .B(n1351), .A(n2868), .Z(n1352) );
  XNOR U1823 ( .A(zin[230]), .B(n1352), .Z(n3411) );
  NANDN U1824 ( .A(n6413), .B(n3411), .Z(n3279) );
  XNOR U1825 ( .A(n6413), .B(n3411), .Z(n2783) );
  XOR U1826 ( .A(y[230]), .B(n1353), .Z(n1354) );
  ANDN U1827 ( .B(n1354), .A(n2868), .Z(n1355) );
  XNOR U1828 ( .A(zin[229]), .B(n1355), .Z(n5233) );
  NAND U1829 ( .A(n5233), .B(n[230]), .Z(n2781) );
  XOR U1830 ( .A(n[230]), .B(n5233), .Z(n2779) );
  XOR U1831 ( .A(y[229]), .B(n1356), .Z(n1357) );
  ANDN U1832 ( .B(n1357), .A(n2868), .Z(n1358) );
  XNOR U1833 ( .A(zin[228]), .B(n1358), .Z(n3415) );
  NAND U1834 ( .A(n[229]), .B(n3415), .Z(n2777) );
  XOR U1835 ( .A(n3415), .B(n[229]), .Z(n2775) );
  XOR U1836 ( .A(y[228]), .B(n1359), .Z(n1360) );
  ANDN U1837 ( .B(n1360), .A(n2868), .Z(n1361) );
  XOR U1838 ( .A(zin[227]), .B(n1361), .Z(n2873) );
  NANDN U1839 ( .A(n2873), .B(n[228]), .Z(n2773) );
  XNOR U1840 ( .A(n[228]), .B(n2873), .Z(n2771) );
  XOR U1841 ( .A(y[227]), .B(n1362), .Z(n1363) );
  ANDN U1842 ( .B(n1363), .A(n2868), .Z(n1364) );
  XNOR U1843 ( .A(zin[226]), .B(n1364), .Z(n3423) );
  NAND U1844 ( .A(n[227]), .B(n3423), .Z(n2769) );
  XOR U1845 ( .A(n3423), .B(n[227]), .Z(n2767) );
  XOR U1846 ( .A(y[226]), .B(n1365), .Z(n1366) );
  ANDN U1847 ( .B(n1366), .A(n2868), .Z(n1367) );
  XNOR U1848 ( .A(zin[225]), .B(n1367), .Z(n3427) );
  NAND U1849 ( .A(n3427), .B(n[226]), .Z(n2765) );
  XOR U1850 ( .A(n[226]), .B(n3427), .Z(n2763) );
  IV U1851 ( .A(n[225]), .Z(n6376) );
  XOR U1852 ( .A(y[225]), .B(n1368), .Z(n1369) );
  ANDN U1853 ( .B(n1369), .A(n2868), .Z(n1370) );
  XNOR U1854 ( .A(zin[224]), .B(n1370), .Z(n3431) );
  NANDN U1855 ( .A(n6376), .B(n3431), .Z(n3273) );
  XNOR U1856 ( .A(n6376), .B(n3431), .Z(n2760) );
  XOR U1857 ( .A(y[224]), .B(n1371), .Z(n1372) );
  ANDN U1858 ( .B(n1372), .A(n2868), .Z(n1373) );
  XNOR U1859 ( .A(zin[223]), .B(n1373), .Z(n3435) );
  NAND U1860 ( .A(n3435), .B(n[224]), .Z(n2758) );
  XOR U1861 ( .A(n[224]), .B(n3435), .Z(n2756) );
  XOR U1862 ( .A(y[223]), .B(n1374), .Z(n1375) );
  ANDN U1863 ( .B(n1375), .A(n2868), .Z(n1376) );
  XNOR U1864 ( .A(zin[222]), .B(n1376), .Z(n3439) );
  NAND U1865 ( .A(n[223]), .B(n3439), .Z(n2754) );
  XOR U1866 ( .A(n3439), .B(n[223]), .Z(n2752) );
  IV U1867 ( .A(n[222]), .Z(n6357) );
  XOR U1868 ( .A(y[222]), .B(n1377), .Z(n1378) );
  ANDN U1869 ( .B(n1378), .A(n2868), .Z(n1379) );
  XNOR U1870 ( .A(zin[221]), .B(n1379), .Z(n3443) );
  NANDN U1871 ( .A(n6357), .B(n3443), .Z(n3270) );
  XNOR U1872 ( .A(n3443), .B(n6357), .Z(n2749) );
  XOR U1873 ( .A(y[221]), .B(n1380), .Z(n1381) );
  ANDN U1874 ( .B(n1381), .A(n2868), .Z(n1382) );
  XNOR U1875 ( .A(zin[220]), .B(n1382), .Z(n3447) );
  NAND U1876 ( .A(n[221]), .B(n3447), .Z(n2747) );
  XOR U1877 ( .A(n3447), .B(n[221]), .Z(n2745) );
  XOR U1878 ( .A(y[220]), .B(n1383), .Z(n1384) );
  ANDN U1879 ( .B(n1384), .A(n2868), .Z(n1385) );
  XNOR U1880 ( .A(zin[219]), .B(n1385), .Z(n3451) );
  NAND U1881 ( .A(n3451), .B(n[220]), .Z(n2743) );
  XOR U1882 ( .A(n[220]), .B(n3451), .Z(n2741) );
  XOR U1883 ( .A(y[219]), .B(n1386), .Z(n1387) );
  ANDN U1884 ( .B(n1387), .A(n2868), .Z(n1388) );
  XNOR U1885 ( .A(zin[218]), .B(n1388), .Z(n3455) );
  NAND U1886 ( .A(n[219]), .B(n3455), .Z(n2739) );
  XOR U1887 ( .A(n3455), .B(n[219]), .Z(n2737) );
  IV U1888 ( .A(n[218]), .Z(n6317) );
  XOR U1889 ( .A(y[218]), .B(n1389), .Z(n1390) );
  ANDN U1890 ( .B(n1390), .A(n2868), .Z(n1391) );
  XNOR U1891 ( .A(zin[217]), .B(n1391), .Z(n3459) );
  NANDN U1892 ( .A(n6317), .B(n3459), .Z(n3267) );
  XNOR U1893 ( .A(n3459), .B(n6317), .Z(n2734) );
  XOR U1894 ( .A(y[217]), .B(n1392), .Z(n1393) );
  ANDN U1895 ( .B(n1393), .A(n2868), .Z(n1394) );
  XNOR U1896 ( .A(zin[216]), .B(n1394), .Z(n5178) );
  NAND U1897 ( .A(n[217]), .B(n5178), .Z(n2732) );
  XOR U1898 ( .A(n5178), .B(n[217]), .Z(n2730) );
  XOR U1899 ( .A(y[216]), .B(n1395), .Z(n1396) );
  ANDN U1900 ( .B(n1396), .A(n2868), .Z(n1397) );
  XNOR U1901 ( .A(zin[215]), .B(n1397), .Z(n3463) );
  NAND U1902 ( .A(n3463), .B(n[216]), .Z(n2728) );
  XOR U1903 ( .A(n[216]), .B(n3463), .Z(n2726) );
  XOR U1904 ( .A(y[215]), .B(n1398), .Z(n1399) );
  ANDN U1905 ( .B(n1399), .A(n2868), .Z(n1400) );
  XNOR U1906 ( .A(zin[214]), .B(n1400), .Z(n3467) );
  NAND U1907 ( .A(n[215]), .B(n3467), .Z(n2724) );
  XOR U1908 ( .A(n3467), .B(n[215]), .Z(n2722) );
  XOR U1909 ( .A(y[214]), .B(n1401), .Z(n1402) );
  ANDN U1910 ( .B(n1402), .A(n2868), .Z(n1403) );
  XNOR U1911 ( .A(zin[213]), .B(n1403), .Z(n3471) );
  NAND U1912 ( .A(n3471), .B(n[214]), .Z(n2720) );
  XOR U1913 ( .A(n[214]), .B(n3471), .Z(n2718) );
  IV U1914 ( .A(n[213]), .Z(n3476) );
  XOR U1915 ( .A(y[213]), .B(n1404), .Z(n1405) );
  ANDN U1916 ( .B(n1405), .A(n2868), .Z(n1406) );
  XNOR U1917 ( .A(zin[212]), .B(n1406), .Z(n3475) );
  NANDN U1918 ( .A(n3476), .B(n3475), .Z(n3264) );
  XNOR U1919 ( .A(n3476), .B(n3475), .Z(n2715) );
  XOR U1920 ( .A(y[212]), .B(n1407), .Z(n1408) );
  ANDN U1921 ( .B(n1408), .A(n2868), .Z(n1409) );
  XNOR U1922 ( .A(zin[211]), .B(n1409), .Z(n3480) );
  NAND U1923 ( .A(n3480), .B(n[212]), .Z(n2713) );
  XOR U1924 ( .A(n[212]), .B(n3480), .Z(n2711) );
  XOR U1925 ( .A(y[211]), .B(n1410), .Z(n1411) );
  ANDN U1926 ( .B(n1411), .A(n2868), .Z(n1412) );
  XNOR U1927 ( .A(zin[210]), .B(n1412), .Z(n3484) );
  NAND U1928 ( .A(n[211]), .B(n3484), .Z(n2709) );
  XOR U1929 ( .A(n3484), .B(n[211]), .Z(n2707) );
  XOR U1930 ( .A(y[210]), .B(n1413), .Z(n1414) );
  ANDN U1931 ( .B(n1414), .A(n2868), .Z(n1415) );
  XOR U1932 ( .A(zin[209]), .B(n1415), .Z(n3488) );
  NANDN U1933 ( .A(n3488), .B(n[210]), .Z(n2705) );
  IV U1934 ( .A(n[210]), .Z(n6268) );
  IV U1935 ( .A(n3488), .Z(n2874) );
  XNOR U1936 ( .A(n6268), .B(n2874), .Z(n2703) );
  IV U1937 ( .A(n[209]), .Z(n6256) );
  XOR U1938 ( .A(y[209]), .B(n1416), .Z(n1417) );
  ANDN U1939 ( .B(n1417), .A(n2868), .Z(n1418) );
  XNOR U1940 ( .A(zin[208]), .B(n1418), .Z(n3492) );
  NANDN U1941 ( .A(n6256), .B(n3492), .Z(n2701) );
  XNOR U1942 ( .A(n3492), .B(n6256), .Z(n2699) );
  IV U1943 ( .A(n[208]), .Z(n3499) );
  XOR U1944 ( .A(y[208]), .B(n1419), .Z(n1420) );
  ANDN U1945 ( .B(n1420), .A(n2868), .Z(n1421) );
  XNOR U1946 ( .A(zin[207]), .B(n1421), .Z(n3498) );
  NANDN U1947 ( .A(n3499), .B(n3498), .Z(n3261) );
  XNOR U1948 ( .A(n3498), .B(n3499), .Z(n2696) );
  XOR U1949 ( .A(y[207]), .B(n1422), .Z(n1423) );
  ANDN U1950 ( .B(n1423), .A(n2868), .Z(n1424) );
  XNOR U1951 ( .A(zin[206]), .B(n1424), .Z(n3503) );
  NAND U1952 ( .A(n[207]), .B(n3503), .Z(n2694) );
  XOR U1953 ( .A(n3503), .B(n[207]), .Z(n2692) );
  IV U1954 ( .A(n[206]), .Z(n3508) );
  XOR U1955 ( .A(y[206]), .B(n1425), .Z(n1426) );
  ANDN U1956 ( .B(n1426), .A(n2868), .Z(n1427) );
  XNOR U1957 ( .A(zin[205]), .B(n1427), .Z(n3507) );
  NANDN U1958 ( .A(n3508), .B(n3507), .Z(n3258) );
  XNOR U1959 ( .A(n3507), .B(n3508), .Z(n2689) );
  XOR U1960 ( .A(y[205]), .B(n1428), .Z(n1429) );
  ANDN U1961 ( .B(n1429), .A(n2868), .Z(n1430) );
  XNOR U1962 ( .A(zin[204]), .B(n1430), .Z(n3512) );
  NAND U1963 ( .A(n[205]), .B(n3512), .Z(n2687) );
  XOR U1964 ( .A(n3512), .B(n[205]), .Z(n2685) );
  XOR U1965 ( .A(y[204]), .B(n1431), .Z(n1432) );
  ANDN U1966 ( .B(n1432), .A(n2868), .Z(n1433) );
  XNOR U1967 ( .A(zin[203]), .B(n1433), .Z(n3516) );
  NAND U1968 ( .A(n3516), .B(n[204]), .Z(n2683) );
  XOR U1969 ( .A(n[204]), .B(n3516), .Z(n2681) );
  IV U1970 ( .A(n[203]), .Z(n6225) );
  XOR U1971 ( .A(y[203]), .B(n1434), .Z(n1435) );
  ANDN U1972 ( .B(n1435), .A(n2868), .Z(n1436) );
  XNOR U1973 ( .A(zin[202]), .B(n1436), .Z(n3520) );
  NANDN U1974 ( .A(n6225), .B(n3520), .Z(n3255) );
  XNOR U1975 ( .A(n6225), .B(n3520), .Z(n2678) );
  XOR U1976 ( .A(y[202]), .B(n1437), .Z(n1438) );
  ANDN U1977 ( .B(n1438), .A(n2868), .Z(n1439) );
  XNOR U1978 ( .A(zin[201]), .B(n1439), .Z(n3524) );
  NAND U1979 ( .A(n3524), .B(n[202]), .Z(n2676) );
  XOR U1980 ( .A(n[202]), .B(n3524), .Z(n2674) );
  IV U1981 ( .A(n[201]), .Z(n3529) );
  XOR U1982 ( .A(y[201]), .B(n1440), .Z(n1441) );
  ANDN U1983 ( .B(n1441), .A(n2868), .Z(n1442) );
  XNOR U1984 ( .A(zin[200]), .B(n1442), .Z(n3528) );
  NANDN U1985 ( .A(n3529), .B(n3528), .Z(n3252) );
  XNOR U1986 ( .A(n3529), .B(n3528), .Z(n2671) );
  IV U1987 ( .A(n[200]), .Z(n6199) );
  XOR U1988 ( .A(y[200]), .B(n1443), .Z(n1444) );
  ANDN U1989 ( .B(n1444), .A(n2868), .Z(n1445) );
  XNOR U1990 ( .A(zin[199]), .B(n1445), .Z(n3533) );
  NANDN U1991 ( .A(n6199), .B(n3533), .Z(n3249) );
  XNOR U1992 ( .A(n3533), .B(n6199), .Z(n2668) );
  XOR U1993 ( .A(y[199]), .B(n1446), .Z(n1447) );
  ANDN U1994 ( .B(n1447), .A(n2868), .Z(n1448) );
  XNOR U1995 ( .A(zin[198]), .B(n1448), .Z(n3537) );
  NAND U1996 ( .A(n[199]), .B(n3537), .Z(n2666) );
  XOR U1997 ( .A(n3537), .B(n[199]), .Z(n2664) );
  XOR U1998 ( .A(y[198]), .B(n1449), .Z(n1450) );
  ANDN U1999 ( .B(n1450), .A(n2868), .Z(n1451) );
  XNOR U2000 ( .A(zin[197]), .B(n1451), .Z(n3542) );
  NAND U2001 ( .A(n[198]), .B(n3542), .Z(n2662) );
  XOR U2002 ( .A(n3542), .B(n[198]), .Z(n2660) );
  XOR U2003 ( .A(y[197]), .B(n1452), .Z(n1453) );
  ANDN U2004 ( .B(n1453), .A(n2868), .Z(n1454) );
  XNOR U2005 ( .A(zin[196]), .B(n1454), .Z(n3546) );
  NAND U2006 ( .A(n[197]), .B(n3546), .Z(n2658) );
  XOR U2007 ( .A(n3546), .B(n[197]), .Z(n2656) );
  IV U2008 ( .A(n[196]), .Z(n6166) );
  XOR U2009 ( .A(y[196]), .B(n1455), .Z(n1456) );
  ANDN U2010 ( .B(n1456), .A(n2868), .Z(n1457) );
  XNOR U2011 ( .A(zin[195]), .B(n1457), .Z(n3550) );
  NANDN U2012 ( .A(n6166), .B(n3550), .Z(n2654) );
  XNOR U2013 ( .A(n3550), .B(n6166), .Z(n2652) );
  IV U2014 ( .A(n[195]), .Z(n3556) );
  XOR U2015 ( .A(y[195]), .B(n1458), .Z(n1459) );
  ANDN U2016 ( .B(n1459), .A(n2868), .Z(n1460) );
  XNOR U2017 ( .A(zin[194]), .B(n1460), .Z(n3554) );
  NANDN U2018 ( .A(n3556), .B(n3554), .Z(n3246) );
  XNOR U2019 ( .A(n3554), .B(n3556), .Z(n2649) );
  XOR U2020 ( .A(y[194]), .B(n1461), .Z(n1462) );
  ANDN U2021 ( .B(n1462), .A(n2868), .Z(n1463) );
  XNOR U2022 ( .A(zin[193]), .B(n1463), .Z(n3560) );
  NAND U2023 ( .A(n[194]), .B(n3560), .Z(n2647) );
  XOR U2024 ( .A(n3560), .B(n[194]), .Z(n2645) );
  XOR U2025 ( .A(y[193]), .B(n1464), .Z(n1465) );
  ANDN U2026 ( .B(n1465), .A(n2868), .Z(n1466) );
  XNOR U2027 ( .A(zin[192]), .B(n1466), .Z(n3564) );
  NAND U2028 ( .A(n[193]), .B(n3564), .Z(n2643) );
  XOR U2029 ( .A(n3564), .B(n[193]), .Z(n2641) );
  XOR U2030 ( .A(y[192]), .B(n1467), .Z(n1468) );
  ANDN U2031 ( .B(n1468), .A(n2868), .Z(n1469) );
  XNOR U2032 ( .A(zin[191]), .B(n1469), .Z(n3568) );
  NAND U2033 ( .A(n3568), .B(n[192]), .Z(n2639) );
  XOR U2034 ( .A(n[192]), .B(n3568), .Z(n2637) );
  XOR U2035 ( .A(y[191]), .B(n1470), .Z(n1471) );
  ANDN U2036 ( .B(n1471), .A(n2868), .Z(n1472) );
  XNOR U2037 ( .A(zin[190]), .B(n1472), .Z(n3572) );
  NAND U2038 ( .A(n[191]), .B(n3572), .Z(n3243) );
  XOR U2039 ( .A(n[191]), .B(n3572), .Z(n2634) );
  IV U2040 ( .A(n[190]), .Z(n6135) );
  XOR U2041 ( .A(y[190]), .B(n1473), .Z(n1474) );
  ANDN U2042 ( .B(n1474), .A(n2868), .Z(n1475) );
  XNOR U2043 ( .A(zin[189]), .B(n1475), .Z(n3576) );
  NANDN U2044 ( .A(n6135), .B(n3576), .Z(n3240) );
  XNOR U2045 ( .A(n3576), .B(n6135), .Z(n2631) );
  IV U2046 ( .A(n[189]), .Z(n3581) );
  XOR U2047 ( .A(y[189]), .B(n1476), .Z(n1477) );
  ANDN U2048 ( .B(n1477), .A(n2868), .Z(n1478) );
  XOR U2049 ( .A(zin[188]), .B(n1478), .Z(n3580) );
  IV U2050 ( .A(n3580), .Z(n2875) );
  NANDN U2051 ( .A(n3581), .B(n2875), .Z(n2629) );
  XNOR U2052 ( .A(n3580), .B(n[189]), .Z(n2627) );
  IV U2053 ( .A(n[188]), .Z(n3586) );
  XOR U2054 ( .A(y[188]), .B(n1479), .Z(n1480) );
  ANDN U2055 ( .B(n1480), .A(n2868), .Z(n1481) );
  XNOR U2056 ( .A(zin[187]), .B(n1481), .Z(n3585) );
  NANDN U2057 ( .A(n3586), .B(n3585), .Z(n3237) );
  XNOR U2058 ( .A(n3586), .B(n3585), .Z(n2624) );
  IV U2059 ( .A(n[187]), .Z(n6106) );
  XOR U2060 ( .A(y[187]), .B(n1482), .Z(n1483) );
  ANDN U2061 ( .B(n1483), .A(n2868), .Z(n1484) );
  XNOR U2062 ( .A(zin[186]), .B(n1484), .Z(n3590) );
  NANDN U2063 ( .A(n6106), .B(n3590), .Z(n3234) );
  XNOR U2064 ( .A(n6106), .B(n3590), .Z(n2621) );
  XOR U2065 ( .A(y[186]), .B(n1485), .Z(n1486) );
  ANDN U2066 ( .B(n1486), .A(n2868), .Z(n1487) );
  XNOR U2067 ( .A(zin[185]), .B(n1487), .Z(n3594) );
  NAND U2068 ( .A(n3594), .B(n[186]), .Z(n2619) );
  XOR U2069 ( .A(n[186]), .B(n3594), .Z(n2617) );
  XOR U2070 ( .A(y[185]), .B(n1488), .Z(n1489) );
  ANDN U2071 ( .B(n1489), .A(n2868), .Z(n1490) );
  XNOR U2072 ( .A(zin[184]), .B(n1490), .Z(n5054) );
  NAND U2073 ( .A(n[185]), .B(n5054), .Z(n2615) );
  XOR U2074 ( .A(n5054), .B(n[185]), .Z(n2613) );
  IV U2075 ( .A(n[184]), .Z(n6086) );
  XOR U2076 ( .A(y[184]), .B(n1491), .Z(n1492) );
  ANDN U2077 ( .B(n1492), .A(n2868), .Z(n1493) );
  XNOR U2078 ( .A(zin[183]), .B(n1493), .Z(n3598) );
  NANDN U2079 ( .A(n6086), .B(n3598), .Z(n3231) );
  XNOR U2080 ( .A(n3598), .B(n6086), .Z(n2610) );
  IV U2081 ( .A(n[183]), .Z(n3603) );
  XOR U2082 ( .A(y[183]), .B(n1494), .Z(n1495) );
  ANDN U2083 ( .B(n1495), .A(n2868), .Z(n1496) );
  XNOR U2084 ( .A(zin[182]), .B(n1496), .Z(n3602) );
  NANDN U2085 ( .A(n3603), .B(n3602), .Z(n3228) );
  XNOR U2086 ( .A(n3603), .B(n3602), .Z(n2607) );
  XOR U2087 ( .A(y[182]), .B(n1497), .Z(n1498) );
  ANDN U2088 ( .B(n1498), .A(n2868), .Z(n1499) );
  XNOR U2089 ( .A(zin[181]), .B(n1499), .Z(n3607) );
  NAND U2090 ( .A(n[182]), .B(n3607), .Z(n2605) );
  XOR U2091 ( .A(n3607), .B(n[182]), .Z(n2603) );
  XOR U2092 ( .A(y[181]), .B(n1500), .Z(n1501) );
  ANDN U2093 ( .B(n1501), .A(n2868), .Z(n1502) );
  XNOR U2094 ( .A(zin[180]), .B(n1502), .Z(n3611) );
  NAND U2095 ( .A(n3611), .B(n[181]), .Z(n2601) );
  XOR U2096 ( .A(n[181]), .B(n3611), .Z(n2599) );
  XOR U2097 ( .A(y[180]), .B(n1503), .Z(n1504) );
  ANDN U2098 ( .B(n1504), .A(n2868), .Z(n1505) );
  XNOR U2099 ( .A(zin[179]), .B(n1505), .Z(n3615) );
  NAND U2100 ( .A(n[180]), .B(n3615), .Z(n2597) );
  XOR U2101 ( .A(n3615), .B(n[180]), .Z(n2595) );
  XOR U2102 ( .A(y[179]), .B(n1506), .Z(n1507) );
  ANDN U2103 ( .B(n1507), .A(n2868), .Z(n1508) );
  XNOR U2104 ( .A(zin[178]), .B(n1508), .Z(n5026) );
  NAND U2105 ( .A(n[179]), .B(n5026), .Z(n2593) );
  XOR U2106 ( .A(n5026), .B(n[179]), .Z(n2591) );
  IV U2107 ( .A(n[178]), .Z(n6039) );
  XOR U2108 ( .A(y[178]), .B(n1509), .Z(n1510) );
  ANDN U2109 ( .B(n1510), .A(n2868), .Z(n1511) );
  XNOR U2110 ( .A(zin[177]), .B(n1511), .Z(n3619) );
  NANDN U2111 ( .A(n6039), .B(n3619), .Z(n2589) );
  XNOR U2112 ( .A(n3619), .B(n6039), .Z(n2587) );
  IV U2113 ( .A(n[177]), .Z(n6042) );
  XOR U2114 ( .A(y[177]), .B(n1512), .Z(n1513) );
  ANDN U2115 ( .B(n1513), .A(n2868), .Z(n1514) );
  XNOR U2116 ( .A(zin[176]), .B(n1514), .Z(n3623) );
  NANDN U2117 ( .A(n6042), .B(n3623), .Z(n3225) );
  XNOR U2118 ( .A(n3623), .B(n6042), .Z(n2584) );
  IV U2119 ( .A(n[176]), .Z(n6025) );
  XOR U2120 ( .A(y[176]), .B(n1515), .Z(n1516) );
  ANDN U2121 ( .B(n1516), .A(n2868), .Z(n1517) );
  XNOR U2122 ( .A(zin[175]), .B(n1517), .Z(n3628) );
  NANDN U2123 ( .A(n6025), .B(n3628), .Z(n2582) );
  XNOR U2124 ( .A(n3628), .B(n6025), .Z(n2580) );
  IV U2125 ( .A(n[175]), .Z(n6024) );
  XOR U2126 ( .A(y[175]), .B(n1518), .Z(n1519) );
  ANDN U2127 ( .B(n1519), .A(n2868), .Z(n1520) );
  XNOR U2128 ( .A(zin[174]), .B(n1520), .Z(n3632) );
  NANDN U2129 ( .A(n6024), .B(n3632), .Z(n3222) );
  XNOR U2130 ( .A(n6024), .B(n3632), .Z(n2577) );
  XOR U2131 ( .A(y[174]), .B(n1521), .Z(n1522) );
  ANDN U2132 ( .B(n1522), .A(n2868), .Z(n1523) );
  XNOR U2133 ( .A(zin[173]), .B(n1523), .Z(n3636) );
  NAND U2134 ( .A(n[174]), .B(n3636), .Z(n2575) );
  XOR U2135 ( .A(n3636), .B(n[174]), .Z(n2573) );
  IV U2136 ( .A(n[173]), .Z(n3641) );
  XOR U2137 ( .A(y[173]), .B(n1524), .Z(n1525) );
  ANDN U2138 ( .B(n1525), .A(n2868), .Z(n1526) );
  XNOR U2139 ( .A(zin[172]), .B(n1526), .Z(n3640) );
  NANDN U2140 ( .A(n3641), .B(n3640), .Z(n3219) );
  XNOR U2141 ( .A(n3640), .B(n3641), .Z(n2570) );
  IV U2142 ( .A(n[172]), .Z(n3646) );
  XOR U2143 ( .A(y[172]), .B(n1527), .Z(n1528) );
  ANDN U2144 ( .B(n1528), .A(n2868), .Z(n1529) );
  XNOR U2145 ( .A(zin[171]), .B(n1529), .Z(n3645) );
  NANDN U2146 ( .A(n3646), .B(n3645), .Z(n3216) );
  XNOR U2147 ( .A(n3646), .B(n3645), .Z(n2567) );
  IV U2148 ( .A(n[171]), .Z(n5998) );
  XOR U2149 ( .A(y[171]), .B(n1530), .Z(n1531) );
  ANDN U2150 ( .B(n1531), .A(n2868), .Z(n1532) );
  XNOR U2151 ( .A(zin[170]), .B(n1532), .Z(n3650) );
  NANDN U2152 ( .A(n5998), .B(n3650), .Z(n3213) );
  XNOR U2153 ( .A(n3650), .B(n5998), .Z(n2564) );
  IV U2154 ( .A(n[170]), .Z(n3655) );
  XOR U2155 ( .A(y[170]), .B(n1533), .Z(n1534) );
  ANDN U2156 ( .B(n1534), .A(n2868), .Z(n1535) );
  XNOR U2157 ( .A(zin[169]), .B(n1535), .Z(n3654) );
  NANDN U2158 ( .A(n3655), .B(n3654), .Z(n3210) );
  XNOR U2159 ( .A(n3655), .B(n3654), .Z(n2561) );
  XOR U2160 ( .A(y[169]), .B(n1536), .Z(n1537) );
  ANDN U2161 ( .B(n1537), .A(n2868), .Z(n1538) );
  XNOR U2162 ( .A(zin[168]), .B(n1538), .Z(n3659) );
  NAND U2163 ( .A(n3659), .B(n[169]), .Z(n2559) );
  XOR U2164 ( .A(n[169]), .B(n3659), .Z(n2557) );
  IV U2165 ( .A(n[168]), .Z(n3664) );
  XOR U2166 ( .A(y[168]), .B(n1539), .Z(n1540) );
  ANDN U2167 ( .B(n1540), .A(n2868), .Z(n1541) );
  XNOR U2168 ( .A(zin[167]), .B(n1541), .Z(n3663) );
  NANDN U2169 ( .A(n3664), .B(n3663), .Z(n3207) );
  XNOR U2170 ( .A(n3664), .B(n3663), .Z(n2554) );
  XOR U2171 ( .A(y[167]), .B(n1542), .Z(n1543) );
  ANDN U2172 ( .B(n1543), .A(n2868), .Z(n1544) );
  XNOR U2173 ( .A(zin[166]), .B(n1544), .Z(n3668) );
  NAND U2174 ( .A(n[167]), .B(n3668), .Z(n3204) );
  XOR U2175 ( .A(n[167]), .B(n3668), .Z(n2551) );
  IV U2176 ( .A(n[166]), .Z(n3673) );
  XOR U2177 ( .A(y[166]), .B(n1545), .Z(n1546) );
  ANDN U2178 ( .B(n1546), .A(n2868), .Z(n1547) );
  XNOR U2179 ( .A(zin[165]), .B(n1547), .Z(n3672) );
  NANDN U2180 ( .A(n3673), .B(n3672), .Z(n3201) );
  XNOR U2181 ( .A(n3672), .B(n3673), .Z(n2548) );
  XOR U2182 ( .A(y[165]), .B(n1548), .Z(n1549) );
  ANDN U2183 ( .B(n1549), .A(n2868), .Z(n1550) );
  XNOR U2184 ( .A(zin[164]), .B(n1550), .Z(n3677) );
  NAND U2185 ( .A(n[165]), .B(n3677), .Z(n3198) );
  XOR U2186 ( .A(n[165]), .B(n3677), .Z(n2545) );
  IV U2187 ( .A(n[164]), .Z(n5943) );
  XOR U2188 ( .A(y[164]), .B(n1551), .Z(n1552) );
  ANDN U2189 ( .B(n1552), .A(n2868), .Z(n1553) );
  XNOR U2190 ( .A(zin[163]), .B(n1553), .Z(n3681) );
  NANDN U2191 ( .A(n5943), .B(n3681), .Z(n3195) );
  XNOR U2192 ( .A(n3681), .B(n5943), .Z(n2542) );
  XOR U2193 ( .A(y[163]), .B(n1554), .Z(n1555) );
  ANDN U2194 ( .B(n1555), .A(n2868), .Z(n1556) );
  XNOR U2195 ( .A(zin[162]), .B(n1556), .Z(n3685) );
  NAND U2196 ( .A(n[163]), .B(n3685), .Z(n2540) );
  XOR U2197 ( .A(n3685), .B(n[163]), .Z(n2538) );
  XOR U2198 ( .A(y[162]), .B(n1557), .Z(n1558) );
  ANDN U2199 ( .B(n1558), .A(n2868), .Z(n1559) );
  XNOR U2200 ( .A(zin[161]), .B(n1559), .Z(n3689) );
  NAND U2201 ( .A(n3689), .B(n[162]), .Z(n2536) );
  XOR U2202 ( .A(n[162]), .B(n3689), .Z(n2534) );
  XOR U2203 ( .A(y[161]), .B(n1560), .Z(n1561) );
  ANDN U2204 ( .B(n1561), .A(n2868), .Z(n1562) );
  XNOR U2205 ( .A(zin[160]), .B(n1562), .Z(n3693) );
  NAND U2206 ( .A(n[161]), .B(n3693), .Z(n2532) );
  XOR U2207 ( .A(n3693), .B(n[161]), .Z(n2530) );
  IV U2208 ( .A(n[160]), .Z(n3698) );
  XOR U2209 ( .A(y[160]), .B(n1563), .Z(n1564) );
  ANDN U2210 ( .B(n1564), .A(n2868), .Z(n1565) );
  XNOR U2211 ( .A(zin[159]), .B(n1565), .Z(n3697) );
  NANDN U2212 ( .A(n3698), .B(n3697), .Z(n3192) );
  XNOR U2213 ( .A(n3697), .B(n3698), .Z(n2527) );
  XOR U2214 ( .A(y[159]), .B(n1566), .Z(n1567) );
  ANDN U2215 ( .B(n1567), .A(n2868), .Z(n1568) );
  XNOR U2216 ( .A(zin[158]), .B(n1568), .Z(n3702) );
  NAND U2217 ( .A(n[159]), .B(n3702), .Z(n2525) );
  XOR U2218 ( .A(n3702), .B(n[159]), .Z(n2523) );
  IV U2219 ( .A(n[158]), .Z(n5903) );
  XOR U2220 ( .A(y[158]), .B(n1569), .Z(n1570) );
  ANDN U2221 ( .B(n1570), .A(n2868), .Z(n1571) );
  XNOR U2222 ( .A(zin[157]), .B(n1571), .Z(n3706) );
  NANDN U2223 ( .A(n5903), .B(n3706), .Z(n3189) );
  XNOR U2224 ( .A(n3706), .B(n5903), .Z(n2520) );
  IV U2225 ( .A(n[157]), .Z(n4939) );
  XOR U2226 ( .A(y[157]), .B(n1572), .Z(n1573) );
  ANDN U2227 ( .B(n1573), .A(n2868), .Z(n1574) );
  XNOR U2228 ( .A(zin[156]), .B(n1574), .Z(n4937) );
  NANDN U2229 ( .A(n4939), .B(n4937), .Z(n3186) );
  XNOR U2230 ( .A(n4939), .B(n4937), .Z(n2517) );
  IV U2231 ( .A(n[156]), .Z(n5889) );
  XOR U2232 ( .A(y[156]), .B(n1575), .Z(n1576) );
  ANDN U2233 ( .B(n1576), .A(n2868), .Z(n1577) );
  XNOR U2234 ( .A(zin[155]), .B(n1577), .Z(n3710) );
  NANDN U2235 ( .A(n5889), .B(n3710), .Z(n3183) );
  XNOR U2236 ( .A(n3710), .B(n5889), .Z(n2514) );
  XOR U2237 ( .A(y[155]), .B(n1578), .Z(n1579) );
  ANDN U2238 ( .B(n1579), .A(n2868), .Z(n1580) );
  XNOR U2239 ( .A(zin[154]), .B(n1580), .Z(n4926) );
  NAND U2240 ( .A(n[155]), .B(n4926), .Z(n2512) );
  XOR U2241 ( .A(n4926), .B(n[155]), .Z(n2510) );
  XOR U2242 ( .A(y[154]), .B(n1581), .Z(n1582) );
  ANDN U2243 ( .B(n1582), .A(n2868), .Z(n1583) );
  XNOR U2244 ( .A(zin[153]), .B(n1583), .Z(n3714) );
  NAND U2245 ( .A(n[154]), .B(n3714), .Z(n3180) );
  XOR U2246 ( .A(n[154]), .B(n3714), .Z(n2507) );
  IV U2247 ( .A(n[153]), .Z(n4910) );
  XOR U2248 ( .A(y[153]), .B(n1584), .Z(n1585) );
  ANDN U2249 ( .B(n1585), .A(n2868), .Z(n1586) );
  XNOR U2250 ( .A(zin[152]), .B(n1586), .Z(n4913) );
  NANDN U2251 ( .A(n4910), .B(n4913), .Z(n3177) );
  XNOR U2252 ( .A(n4910), .B(n4913), .Z(n2504) );
  XOR U2253 ( .A(y[152]), .B(n1587), .Z(n1588) );
  ANDN U2254 ( .B(n1588), .A(n2868), .Z(n1589) );
  XNOR U2255 ( .A(zin[151]), .B(n1589), .Z(n3718) );
  NAND U2256 ( .A(n[152]), .B(n3718), .Z(n2502) );
  XOR U2257 ( .A(n3718), .B(n[152]), .Z(n2500) );
  XOR U2258 ( .A(y[151]), .B(n1590), .Z(n1591) );
  ANDN U2259 ( .B(n1591), .A(n2868), .Z(n1592) );
  XNOR U2260 ( .A(zin[150]), .B(n1592), .Z(n3722) );
  NAND U2261 ( .A(n[151]), .B(n3722), .Z(n3174) );
  XOR U2262 ( .A(n[151]), .B(n3722), .Z(n2497) );
  XOR U2263 ( .A(y[150]), .B(n1593), .Z(n1594) );
  ANDN U2264 ( .B(n1594), .A(n2868), .Z(n1595) );
  XNOR U2265 ( .A(zin[149]), .B(n1595), .Z(n3726) );
  NAND U2266 ( .A(n3726), .B(n[150]), .Z(n2495) );
  XOR U2267 ( .A(n[150]), .B(n3726), .Z(n2493) );
  XOR U2268 ( .A(y[149]), .B(n1596), .Z(n1597) );
  ANDN U2269 ( .B(n1597), .A(n2868), .Z(n1598) );
  XNOR U2270 ( .A(zin[148]), .B(n1598), .Z(n3730) );
  NAND U2271 ( .A(n[149]), .B(n3730), .Z(n2491) );
  XOR U2272 ( .A(n3730), .B(n[149]), .Z(n2489) );
  XOR U2273 ( .A(y[148]), .B(n1599), .Z(n1600) );
  ANDN U2274 ( .B(n1600), .A(n2868), .Z(n1601) );
  XNOR U2275 ( .A(zin[147]), .B(n1601), .Z(n3734) );
  NAND U2276 ( .A(n3734), .B(n[148]), .Z(n2487) );
  XOR U2277 ( .A(n[148]), .B(n3734), .Z(n2485) );
  IV U2278 ( .A(n[147]), .Z(n3739) );
  XOR U2279 ( .A(y[147]), .B(n1602), .Z(n1603) );
  ANDN U2280 ( .B(n1603), .A(n2868), .Z(n1604) );
  XNOR U2281 ( .A(zin[146]), .B(n1604), .Z(n3738) );
  NANDN U2282 ( .A(n3739), .B(n3738), .Z(n3171) );
  XNOR U2283 ( .A(n3739), .B(n3738), .Z(n2482) );
  XOR U2284 ( .A(y[146]), .B(n1605), .Z(n1606) );
  ANDN U2285 ( .B(n1606), .A(n2868), .Z(n1607) );
  XNOR U2286 ( .A(zin[145]), .B(n1607), .Z(n3743) );
  NAND U2287 ( .A(n[146]), .B(n3743), .Z(n2480) );
  XOR U2288 ( .A(n3743), .B(n[146]), .Z(n2478) );
  XOR U2289 ( .A(y[145]), .B(n1608), .Z(n1609) );
  ANDN U2290 ( .B(n1609), .A(n2868), .Z(n1610) );
  XNOR U2291 ( .A(zin[144]), .B(n1610), .Z(n3747) );
  NAND U2292 ( .A(n[145]), .B(n3747), .Z(n3168) );
  XOR U2293 ( .A(n[145]), .B(n3747), .Z(n2475) );
  IV U2294 ( .A(n[144]), .Z(n3752) );
  XOR U2295 ( .A(y[144]), .B(n1611), .Z(n1612) );
  ANDN U2296 ( .B(n1612), .A(n2868), .Z(n1613) );
  XNOR U2297 ( .A(zin[143]), .B(n1613), .Z(n3751) );
  NANDN U2298 ( .A(n3752), .B(n3751), .Z(n3165) );
  XNOR U2299 ( .A(n3752), .B(n3751), .Z(n2472) );
  XOR U2300 ( .A(y[143]), .B(n1614), .Z(n1615) );
  ANDN U2301 ( .B(n1615), .A(n2868), .Z(n1616) );
  XNOR U2302 ( .A(zin[142]), .B(n1616), .Z(n3756) );
  NAND U2303 ( .A(n[143]), .B(n3756), .Z(n2470) );
  XOR U2304 ( .A(n3756), .B(n[143]), .Z(n2468) );
  XOR U2305 ( .A(y[142]), .B(n1617), .Z(n1618) );
  ANDN U2306 ( .B(n1618), .A(n2868), .Z(n1619) );
  XOR U2307 ( .A(zin[141]), .B(n1619), .Z(n2876) );
  NANDN U2308 ( .A(n2876), .B(n[142]), .Z(n2466) );
  XNOR U2309 ( .A(n[142]), .B(n2876), .Z(n2464) );
  XOR U2310 ( .A(y[141]), .B(n1620), .Z(n1621) );
  ANDN U2311 ( .B(n1621), .A(n2868), .Z(n1622) );
  XNOR U2312 ( .A(zin[140]), .B(n1622), .Z(n3764) );
  NAND U2313 ( .A(n[141]), .B(n3764), .Z(n2462) );
  XOR U2314 ( .A(n3764), .B(n[141]), .Z(n2460) );
  IV U2315 ( .A(n[140]), .Z(n3769) );
  XOR U2316 ( .A(y[140]), .B(n1623), .Z(n1624) );
  ANDN U2317 ( .B(n1624), .A(n2868), .Z(n1625) );
  XNOR U2318 ( .A(zin[139]), .B(n1625), .Z(n3768) );
  NANDN U2319 ( .A(n3769), .B(n3768), .Z(n3159) );
  XNOR U2320 ( .A(n3768), .B(n3769), .Z(n2457) );
  XOR U2321 ( .A(y[139]), .B(n1626), .Z(n1627) );
  ANDN U2322 ( .B(n1627), .A(n2868), .Z(n1628) );
  XNOR U2323 ( .A(zin[138]), .B(n1628), .Z(n3773) );
  NAND U2324 ( .A(n[139]), .B(n3773), .Z(n2455) );
  XOR U2325 ( .A(n3773), .B(n[139]), .Z(n2453) );
  XOR U2326 ( .A(y[138]), .B(n1629), .Z(n1630) );
  ANDN U2327 ( .B(n1630), .A(n2868), .Z(n1631) );
  XNOR U2328 ( .A(zin[137]), .B(n1631), .Z(n3777) );
  NAND U2329 ( .A(n3777), .B(n[138]), .Z(n2451) );
  XOR U2330 ( .A(n[138]), .B(n3777), .Z(n2449) );
  XOR U2331 ( .A(y[137]), .B(n1632), .Z(n1633) );
  ANDN U2332 ( .B(n1633), .A(n2868), .Z(n1634) );
  XNOR U2333 ( .A(zin[136]), .B(n1634), .Z(n3781) );
  NAND U2334 ( .A(n[137]), .B(n3781), .Z(n2447) );
  XOR U2335 ( .A(n3781), .B(n[137]), .Z(n2445) );
  XOR U2336 ( .A(y[136]), .B(n1635), .Z(n1636) );
  ANDN U2337 ( .B(n1636), .A(n2868), .Z(n1637) );
  XNOR U2338 ( .A(zin[135]), .B(n1637), .Z(n3785) );
  NAND U2339 ( .A(n3785), .B(n[136]), .Z(n2443) );
  XOR U2340 ( .A(n[136]), .B(n3785), .Z(n2441) );
  XOR U2341 ( .A(y[135]), .B(n1638), .Z(n1639) );
  ANDN U2342 ( .B(n1639), .A(n2868), .Z(n1640) );
  XNOR U2343 ( .A(zin[134]), .B(n1640), .Z(n3789) );
  NAND U2344 ( .A(n[135]), .B(n3789), .Z(n2439) );
  XOR U2345 ( .A(n3789), .B(n[135]), .Z(n2437) );
  XOR U2346 ( .A(y[134]), .B(n1641), .Z(n1642) );
  ANDN U2347 ( .B(n1642), .A(n2868), .Z(n1643) );
  XNOR U2348 ( .A(zin[133]), .B(n1643), .Z(n3793) );
  NAND U2349 ( .A(n[134]), .B(n3793), .Z(n2435) );
  XOR U2350 ( .A(n3793), .B(n[134]), .Z(n2433) );
  IV U2351 ( .A(n[133]), .Z(n3798) );
  XOR U2352 ( .A(y[133]), .B(n1644), .Z(n1645) );
  ANDN U2353 ( .B(n1645), .A(n2868), .Z(n1646) );
  XNOR U2354 ( .A(zin[132]), .B(n1646), .Z(n3797) );
  NANDN U2355 ( .A(n3798), .B(n3797), .Z(n3156) );
  XNOR U2356 ( .A(n3797), .B(n3798), .Z(n2430) );
  XOR U2357 ( .A(y[132]), .B(n1647), .Z(n1648) );
  ANDN U2358 ( .B(n1648), .A(n2868), .Z(n1649) );
  XNOR U2359 ( .A(zin[131]), .B(n1649), .Z(n3802) );
  NAND U2360 ( .A(n[132]), .B(n3802), .Z(n2428) );
  XOR U2361 ( .A(n3802), .B(n[132]), .Z(n2426) );
  XOR U2362 ( .A(y[131]), .B(n1650), .Z(n1651) );
  ANDN U2363 ( .B(n1651), .A(n2868), .Z(n1652) );
  XNOR U2364 ( .A(zin[130]), .B(n1652), .Z(n3806) );
  NAND U2365 ( .A(n[131]), .B(n3806), .Z(n3153) );
  XOR U2366 ( .A(n[131]), .B(n3806), .Z(n2423) );
  IV U2367 ( .A(n[130]), .Z(n3811) );
  XOR U2368 ( .A(y[130]), .B(n1653), .Z(n1654) );
  ANDN U2369 ( .B(n1654), .A(n2868), .Z(n1655) );
  XNOR U2370 ( .A(zin[129]), .B(n1655), .Z(n3810) );
  NANDN U2371 ( .A(n3811), .B(n3810), .Z(n3150) );
  XNOR U2372 ( .A(n3810), .B(n3811), .Z(n2420) );
  XOR U2373 ( .A(y[129]), .B(n1656), .Z(n1657) );
  ANDN U2374 ( .B(n1657), .A(n2868), .Z(n1658) );
  XNOR U2375 ( .A(zin[128]), .B(n1658), .Z(n3815) );
  NAND U2376 ( .A(n[129]), .B(n3815), .Z(n2418) );
  XOR U2377 ( .A(n3815), .B(n[129]), .Z(n2416) );
  XOR U2378 ( .A(y[128]), .B(n1659), .Z(n1660) );
  ANDN U2379 ( .B(n1660), .A(n2868), .Z(n1661) );
  XNOR U2380 ( .A(zin[127]), .B(n1661), .Z(n3819) );
  NAND U2381 ( .A(n[128]), .B(n3819), .Z(n3147) );
  XOR U2382 ( .A(n[128]), .B(n3819), .Z(n2413) );
  XOR U2383 ( .A(y[127]), .B(n1662), .Z(n1663) );
  ANDN U2384 ( .B(n1663), .A(n2868), .Z(n1664) );
  XNOR U2385 ( .A(zin[126]), .B(n1664), .Z(n3823) );
  NAND U2386 ( .A(n3823), .B(n[127]), .Z(n2411) );
  XOR U2387 ( .A(n[127]), .B(n3823), .Z(n2409) );
  XOR U2388 ( .A(y[126]), .B(n1665), .Z(n1666) );
  ANDN U2389 ( .B(n1666), .A(n2868), .Z(n1667) );
  XNOR U2390 ( .A(zin[125]), .B(n1667), .Z(n3827) );
  NAND U2391 ( .A(n[126]), .B(n3827), .Z(n2407) );
  XOR U2392 ( .A(n3827), .B(n[126]), .Z(n2405) );
  IV U2393 ( .A(n[125]), .Z(n3832) );
  XOR U2394 ( .A(y[125]), .B(n1668), .Z(n1669) );
  ANDN U2395 ( .B(n1669), .A(n2868), .Z(n1670) );
  XNOR U2396 ( .A(zin[124]), .B(n1670), .Z(n3831) );
  NANDN U2397 ( .A(n3832), .B(n3831), .Z(n3144) );
  XNOR U2398 ( .A(n3831), .B(n3832), .Z(n2402) );
  XOR U2399 ( .A(y[124]), .B(n1671), .Z(n1672) );
  ANDN U2400 ( .B(n1672), .A(n2868), .Z(n1673) );
  XNOR U2401 ( .A(zin[123]), .B(n1673), .Z(n3836) );
  NAND U2402 ( .A(n[124]), .B(n3836), .Z(n2400) );
  XOR U2403 ( .A(n3836), .B(n[124]), .Z(n2398) );
  IV U2404 ( .A(n[123]), .Z(n3841) );
  XOR U2405 ( .A(y[123]), .B(n1674), .Z(n1675) );
  ANDN U2406 ( .B(n1675), .A(n2868), .Z(n1676) );
  XNOR U2407 ( .A(zin[122]), .B(n1676), .Z(n3840) );
  NANDN U2408 ( .A(n3841), .B(n3840), .Z(n3141) );
  XNOR U2409 ( .A(n3841), .B(n3840), .Z(n2395) );
  IV U2410 ( .A(n[122]), .Z(n3846) );
  XOR U2411 ( .A(y[122]), .B(n1677), .Z(n1678) );
  ANDN U2412 ( .B(n1678), .A(n2868), .Z(n1679) );
  XNOR U2413 ( .A(zin[121]), .B(n1679), .Z(n3845) );
  NANDN U2414 ( .A(n3846), .B(n3845), .Z(n3138) );
  XNOR U2415 ( .A(n3845), .B(n3846), .Z(n2392) );
  IV U2416 ( .A(n[121]), .Z(n3851) );
  XOR U2417 ( .A(y[121]), .B(n1680), .Z(n1681) );
  ANDN U2418 ( .B(n1681), .A(n2868), .Z(n1682) );
  XNOR U2419 ( .A(zin[120]), .B(n1682), .Z(n3850) );
  NANDN U2420 ( .A(n3851), .B(n3850), .Z(n3135) );
  XNOR U2421 ( .A(n3851), .B(n3850), .Z(n2389) );
  IV U2422 ( .A(n[120]), .Z(n3856) );
  XOR U2423 ( .A(y[120]), .B(n1683), .Z(n1684) );
  ANDN U2424 ( .B(n1684), .A(n2868), .Z(n1685) );
  XNOR U2425 ( .A(zin[119]), .B(n1685), .Z(n3855) );
  NANDN U2426 ( .A(n3856), .B(n3855), .Z(n3132) );
  XNOR U2427 ( .A(n3855), .B(n3856), .Z(n2386) );
  XOR U2428 ( .A(y[119]), .B(n1686), .Z(n1687) );
  ANDN U2429 ( .B(n1687), .A(n2868), .Z(n1688) );
  XNOR U2430 ( .A(zin[118]), .B(n1688), .Z(n3860) );
  NAND U2431 ( .A(n[119]), .B(n3860), .Z(n3129) );
  XOR U2432 ( .A(n[119]), .B(n3860), .Z(n2383) );
  IV U2433 ( .A(n[118]), .Z(n5648) );
  XOR U2434 ( .A(y[118]), .B(n1689), .Z(n1690) );
  ANDN U2435 ( .B(n1690), .A(n2868), .Z(n1691) );
  XNOR U2436 ( .A(zin[117]), .B(n1691), .Z(n3864) );
  NANDN U2437 ( .A(n5648), .B(n3864), .Z(n3126) );
  XNOR U2438 ( .A(n3864), .B(n5648), .Z(n2380) );
  IV U2439 ( .A(n[117]), .Z(n3869) );
  XOR U2440 ( .A(y[117]), .B(n1692), .Z(n1693) );
  ANDN U2441 ( .B(n1693), .A(n2868), .Z(n1694) );
  XNOR U2442 ( .A(zin[116]), .B(n1694), .Z(n3868) );
  NANDN U2443 ( .A(n3869), .B(n3868), .Z(n3123) );
  XNOR U2444 ( .A(n3869), .B(n3868), .Z(n2377) );
  IV U2445 ( .A(n[116]), .Z(n5633) );
  XOR U2446 ( .A(y[116]), .B(n1695), .Z(n1696) );
  ANDN U2447 ( .B(n1696), .A(n2868), .Z(n1697) );
  XNOR U2448 ( .A(zin[115]), .B(n1697), .Z(n3873) );
  NANDN U2449 ( .A(n5633), .B(n3873), .Z(n3120) );
  XNOR U2450 ( .A(n3873), .B(n5633), .Z(n2374) );
  IV U2451 ( .A(n[115]), .Z(n3878) );
  XOR U2452 ( .A(y[115]), .B(n1698), .Z(n1699) );
  ANDN U2453 ( .B(n1699), .A(n2868), .Z(n1700) );
  XNOR U2454 ( .A(zin[114]), .B(n1700), .Z(n3877) );
  NANDN U2455 ( .A(n3878), .B(n3877), .Z(n3117) );
  XNOR U2456 ( .A(n3878), .B(n3877), .Z(n2371) );
  IV U2457 ( .A(n[114]), .Z(n3883) );
  XOR U2458 ( .A(y[114]), .B(n1701), .Z(n1702) );
  ANDN U2459 ( .B(n1702), .A(n2868), .Z(n1703) );
  XNOR U2460 ( .A(zin[113]), .B(n1703), .Z(n3882) );
  NANDN U2461 ( .A(n3883), .B(n3882), .Z(n3114) );
  XNOR U2462 ( .A(n3882), .B(n3883), .Z(n2368) );
  IV U2463 ( .A(n[113]), .Z(n3888) );
  XOR U2464 ( .A(y[113]), .B(n1704), .Z(n1705) );
  ANDN U2465 ( .B(n1705), .A(n2868), .Z(n1706) );
  XNOR U2466 ( .A(zin[112]), .B(n1706), .Z(n3887) );
  NANDN U2467 ( .A(n3888), .B(n3887), .Z(n3111) );
  XNOR U2468 ( .A(n3888), .B(n3887), .Z(n2365) );
  IV U2469 ( .A(n[112]), .Z(n3893) );
  XOR U2470 ( .A(y[112]), .B(n1707), .Z(n1708) );
  ANDN U2471 ( .B(n1708), .A(n2868), .Z(n1709) );
  XNOR U2472 ( .A(zin[111]), .B(n1709), .Z(n3892) );
  NANDN U2473 ( .A(n3893), .B(n3892), .Z(n3108) );
  XNOR U2474 ( .A(n3892), .B(n3893), .Z(n2362) );
  IV U2475 ( .A(n[111]), .Z(n3898) );
  XOR U2476 ( .A(y[111]), .B(n1710), .Z(n1711) );
  ANDN U2477 ( .B(n1711), .A(n2868), .Z(n1712) );
  XNOR U2478 ( .A(zin[110]), .B(n1712), .Z(n3897) );
  NANDN U2479 ( .A(n3898), .B(n3897), .Z(n3105) );
  XNOR U2480 ( .A(n3898), .B(n3897), .Z(n2359) );
  IV U2481 ( .A(n[110]), .Z(n3903) );
  XOR U2482 ( .A(y[110]), .B(n1713), .Z(n1714) );
  ANDN U2483 ( .B(n1714), .A(n2868), .Z(n1715) );
  XNOR U2484 ( .A(zin[109]), .B(n1715), .Z(n3902) );
  NANDN U2485 ( .A(n3903), .B(n3902), .Z(n3102) );
  XNOR U2486 ( .A(n3902), .B(n3903), .Z(n2356) );
  XOR U2487 ( .A(y[109]), .B(n1716), .Z(n1717) );
  ANDN U2488 ( .B(n1717), .A(n2868), .Z(n1718) );
  XNOR U2489 ( .A(zin[108]), .B(n1718), .Z(n3907) );
  NAND U2490 ( .A(n[109]), .B(n3907), .Z(n3099) );
  XOR U2491 ( .A(n[109]), .B(n3907), .Z(n2353) );
  IV U2492 ( .A(n[108]), .Z(n3912) );
  XOR U2493 ( .A(y[108]), .B(n1719), .Z(n1720) );
  ANDN U2494 ( .B(n1720), .A(n2868), .Z(n1721) );
  XNOR U2495 ( .A(zin[107]), .B(n1721), .Z(n3911) );
  NANDN U2496 ( .A(n3912), .B(n3911), .Z(n3096) );
  XNOR U2497 ( .A(n3911), .B(n3912), .Z(n2350) );
  XOR U2498 ( .A(y[107]), .B(n1722), .Z(n1723) );
  ANDN U2499 ( .B(n1723), .A(n2868), .Z(n1724) );
  XNOR U2500 ( .A(zin[106]), .B(n1724), .Z(n3916) );
  NAND U2501 ( .A(n[107]), .B(n3916), .Z(n2348) );
  XOR U2502 ( .A(n3916), .B(n[107]), .Z(n2346) );
  XOR U2503 ( .A(y[106]), .B(n1725), .Z(n1726) );
  ANDN U2504 ( .B(n1726), .A(n2868), .Z(n1727) );
  XNOR U2505 ( .A(zin[105]), .B(n1727), .Z(n3920) );
  NAND U2506 ( .A(n[106]), .B(n3920), .Z(n2344) );
  XOR U2507 ( .A(n3920), .B(n[106]), .Z(n2342) );
  XOR U2508 ( .A(y[105]), .B(n1728), .Z(n1729) );
  ANDN U2509 ( .B(n1729), .A(n2868), .Z(n1730) );
  XNOR U2510 ( .A(zin[104]), .B(n1730), .Z(n3924) );
  NAND U2511 ( .A(n[105]), .B(n3924), .Z(n2340) );
  XOR U2512 ( .A(n3924), .B(n[105]), .Z(n2338) );
  XOR U2513 ( .A(y[104]), .B(n1731), .Z(n1732) );
  ANDN U2514 ( .B(n1732), .A(n2868), .Z(n1733) );
  XNOR U2515 ( .A(zin[103]), .B(n1733), .Z(n3928) );
  NAND U2516 ( .A(n[104]), .B(n3928), .Z(n2336) );
  XOR U2517 ( .A(n3928), .B(n[104]), .Z(n2334) );
  IV U2518 ( .A(n[103]), .Z(n3933) );
  XOR U2519 ( .A(y[103]), .B(n1734), .Z(n1735) );
  ANDN U2520 ( .B(n1735), .A(n2868), .Z(n1736) );
  XNOR U2521 ( .A(zin[102]), .B(n1736), .Z(n3932) );
  NANDN U2522 ( .A(n3933), .B(n3932), .Z(n3093) );
  XNOR U2523 ( .A(n3933), .B(n3932), .Z(n2331) );
  XOR U2524 ( .A(y[102]), .B(n1737), .Z(n1738) );
  ANDN U2525 ( .B(n1738), .A(n2868), .Z(n1739) );
  XNOR U2526 ( .A(zin[101]), .B(n1739), .Z(n3937) );
  NAND U2527 ( .A(n[102]), .B(n3937), .Z(n2329) );
  XOR U2528 ( .A(n3937), .B(n[102]), .Z(n2327) );
  IV U2529 ( .A(n[101]), .Z(n3942) );
  XOR U2530 ( .A(y[101]), .B(n1740), .Z(n1741) );
  ANDN U2531 ( .B(n1741), .A(n2868), .Z(n1742) );
  XNOR U2532 ( .A(zin[100]), .B(n1742), .Z(n3941) );
  NANDN U2533 ( .A(n3942), .B(n3941), .Z(n3090) );
  XNOR U2534 ( .A(n3942), .B(n3941), .Z(n2324) );
  XOR U2535 ( .A(y[100]), .B(n1743), .Z(n1744) );
  ANDN U2536 ( .B(n1744), .A(n2868), .Z(n1745) );
  XNOR U2537 ( .A(zin[99]), .B(n1745), .Z(n3946) );
  IV U2538 ( .A(n[99]), .Z(n5344) );
  XOR U2539 ( .A(y[99]), .B(n1746), .Z(n1747) );
  ANDN U2540 ( .B(n1747), .A(n2868), .Z(n1748) );
  XNOR U2541 ( .A(zin[98]), .B(n1748), .Z(n3950) );
  XOR U2542 ( .A(y[98]), .B(n1749), .Z(n1750) );
  ANDN U2543 ( .B(n1750), .A(n2868), .Z(n1751) );
  XNOR U2544 ( .A(zin[97]), .B(n1751), .Z(n3954) );
  XOR U2545 ( .A(y[97]), .B(n1752), .Z(n1753) );
  ANDN U2546 ( .B(n1753), .A(n2868), .Z(n1754) );
  XNOR U2547 ( .A(zin[96]), .B(n1754), .Z(n3958) );
  IV U2548 ( .A(n[96]), .Z(n3963) );
  XOR U2549 ( .A(y[96]), .B(n1755), .Z(n1756) );
  ANDN U2550 ( .B(n1756), .A(n2868), .Z(n1757) );
  XNOR U2551 ( .A(zin[95]), .B(n1757), .Z(n3962) );
  NANDN U2552 ( .A(n3963), .B(n3962), .Z(n3087) );
  IV U2553 ( .A(n[95]), .Z(n5529) );
  XOR U2554 ( .A(y[95]), .B(n1758), .Z(n1759) );
  ANDN U2555 ( .B(n1759), .A(n2868), .Z(n1760) );
  XNOR U2556 ( .A(zin[94]), .B(n1760), .Z(n3967) );
  NANDN U2557 ( .A(n5529), .B(n3967), .Z(n3084) );
  XNOR U2558 ( .A(n5529), .B(n3967), .Z(n2320) );
  IV U2559 ( .A(n[94]), .Z(n3969) );
  XOR U2560 ( .A(y[94]), .B(n1761), .Z(n1762) );
  ANDN U2561 ( .B(n1762), .A(n2868), .Z(n1763) );
  XNOR U2562 ( .A(zin[93]), .B(n1763), .Z(n3972) );
  NANDN U2563 ( .A(n3969), .B(n3972), .Z(n3081) );
  XNOR U2564 ( .A(n3972), .B(n3969), .Z(n2317) );
  IV U2565 ( .A(n[93]), .Z(n3974) );
  XOR U2566 ( .A(y[93]), .B(n1764), .Z(n1765) );
  ANDN U2567 ( .B(n1765), .A(n2868), .Z(n1766) );
  XNOR U2568 ( .A(zin[92]), .B(n1766), .Z(n3977) );
  NANDN U2569 ( .A(n3974), .B(n3977), .Z(n3078) );
  XNOR U2570 ( .A(n3974), .B(n3977), .Z(n2314) );
  IV U2571 ( .A(n[92]), .Z(n5353) );
  XOR U2572 ( .A(y[92]), .B(n1767), .Z(n1768) );
  ANDN U2573 ( .B(n1768), .A(n2868), .Z(n1769) );
  XNOR U2574 ( .A(zin[91]), .B(n1769), .Z(n4663) );
  NANDN U2575 ( .A(n5353), .B(n4663), .Z(n3075) );
  XNOR U2576 ( .A(n4663), .B(n5353), .Z(n2311) );
  XOR U2577 ( .A(y[91]), .B(n1770), .Z(n1771) );
  ANDN U2578 ( .B(n1771), .A(n2868), .Z(n1772) );
  XNOR U2579 ( .A(zin[90]), .B(n1772), .Z(n3981) );
  NAND U2580 ( .A(n[91]), .B(n3981), .Z(n3072) );
  XOR U2581 ( .A(n[91]), .B(n3981), .Z(n2308) );
  XOR U2582 ( .A(y[90]), .B(n1773), .Z(n1774) );
  ANDN U2583 ( .B(n1774), .A(n2868), .Z(n1775) );
  XNOR U2584 ( .A(zin[89]), .B(n1775), .Z(n3985) );
  NAND U2585 ( .A(n[90]), .B(n3985), .Z(n2306) );
  XOR U2586 ( .A(n3985), .B(n[90]), .Z(n2304) );
  XOR U2587 ( .A(y[89]), .B(n1776), .Z(n1777) );
  ANDN U2588 ( .B(n1777), .A(n2868), .Z(n1778) );
  XNOR U2589 ( .A(zin[88]), .B(n1778), .Z(n3989) );
  NAND U2590 ( .A(n[89]), .B(n3989), .Z(n3069) );
  XOR U2591 ( .A(n[89]), .B(n3989), .Z(n2301) );
  XOR U2592 ( .A(y[88]), .B(n1779), .Z(n1780) );
  ANDN U2593 ( .B(n1780), .A(n2868), .Z(n1781) );
  XNOR U2594 ( .A(zin[87]), .B(n1781), .Z(n3993) );
  NAND U2595 ( .A(n3993), .B(n[88]), .Z(n2299) );
  XOR U2596 ( .A(n[88]), .B(n3993), .Z(n2297) );
  IV U2597 ( .A(n[87]), .Z(n3998) );
  XOR U2598 ( .A(y[87]), .B(n1782), .Z(n1783) );
  ANDN U2599 ( .B(n1783), .A(n2868), .Z(n1784) );
  XNOR U2600 ( .A(zin[86]), .B(n1784), .Z(n3997) );
  NANDN U2601 ( .A(n3998), .B(n3997), .Z(n3066) );
  XNOR U2602 ( .A(n3998), .B(n3997), .Z(n2294) );
  XOR U2603 ( .A(y[86]), .B(n1785), .Z(n1786) );
  ANDN U2604 ( .B(n1786), .A(n2868), .Z(n1787) );
  XNOR U2605 ( .A(zin[85]), .B(n1787), .Z(n4002) );
  NAND U2606 ( .A(n4002), .B(n[86]), .Z(n2292) );
  XOR U2607 ( .A(n[86]), .B(n4002), .Z(n2290) );
  IV U2608 ( .A(n[85]), .Z(n5504) );
  XOR U2609 ( .A(y[85]), .B(n1788), .Z(n1789) );
  ANDN U2610 ( .B(n1789), .A(n2868), .Z(n1790) );
  XNOR U2611 ( .A(zin[84]), .B(n1790), .Z(n4006) );
  NANDN U2612 ( .A(n5504), .B(n4006), .Z(n3063) );
  XNOR U2613 ( .A(n5504), .B(n4006), .Z(n2287) );
  XOR U2614 ( .A(y[84]), .B(n1791), .Z(n1792) );
  ANDN U2615 ( .B(n1792), .A(n2868), .Z(n1793) );
  XNOR U2616 ( .A(zin[83]), .B(n1793), .Z(n4010) );
  NAND U2617 ( .A(n4010), .B(n[84]), .Z(n2285) );
  XOR U2618 ( .A(n[84]), .B(n4010), .Z(n2283) );
  XOR U2619 ( .A(y[83]), .B(n1794), .Z(n1795) );
  ANDN U2620 ( .B(n1795), .A(n2868), .Z(n1796) );
  XNOR U2621 ( .A(zin[82]), .B(n1796), .Z(n4014) );
  NAND U2622 ( .A(n[83]), .B(n4014), .Z(n2281) );
  XOR U2623 ( .A(n4014), .B(n[83]), .Z(n2279) );
  XOR U2624 ( .A(y[82]), .B(n1797), .Z(n1798) );
  ANDN U2625 ( .B(n1798), .A(n2868), .Z(n1799) );
  XNOR U2626 ( .A(zin[81]), .B(n1799), .Z(n4018) );
  NAND U2627 ( .A(n[82]), .B(n4018), .Z(n2277) );
  XOR U2628 ( .A(n4018), .B(n[82]), .Z(n2275) );
  IV U2629 ( .A(n[81]), .Z(n4023) );
  XOR U2630 ( .A(y[81]), .B(n1800), .Z(n1801) );
  ANDN U2631 ( .B(n1801), .A(n2868), .Z(n1802) );
  XNOR U2632 ( .A(zin[80]), .B(n1802), .Z(n4022) );
  NANDN U2633 ( .A(n4023), .B(n4022), .Z(n3060) );
  XNOR U2634 ( .A(n4023), .B(n4022), .Z(n2272) );
  IV U2635 ( .A(n[80]), .Z(n4028) );
  XOR U2636 ( .A(y[80]), .B(n1803), .Z(n1804) );
  ANDN U2637 ( .B(n1804), .A(n2868), .Z(n1805) );
  XNOR U2638 ( .A(zin[79]), .B(n1805), .Z(n4027) );
  NANDN U2639 ( .A(n4028), .B(n4027), .Z(n3057) );
  XNOR U2640 ( .A(n4028), .B(n4027), .Z(n2269) );
  XOR U2641 ( .A(y[79]), .B(n1806), .Z(n1807) );
  ANDN U2642 ( .B(n1807), .A(n2868), .Z(n1808) );
  XNOR U2643 ( .A(zin[78]), .B(n1808), .Z(n4032) );
  NAND U2644 ( .A(n[79]), .B(n4032), .Z(n2267) );
  XOR U2645 ( .A(n4032), .B(n[79]), .Z(n2265) );
  XOR U2646 ( .A(y[78]), .B(n1809), .Z(n1810) );
  ANDN U2647 ( .B(n1810), .A(n2868), .Z(n1811) );
  XNOR U2648 ( .A(zin[77]), .B(n1811), .Z(n4036) );
  NAND U2649 ( .A(n4036), .B(n[78]), .Z(n2263) );
  XOR U2650 ( .A(n[78]), .B(n4036), .Z(n2261) );
  IV U2651 ( .A(n[77]), .Z(n4041) );
  XOR U2652 ( .A(y[77]), .B(n1812), .Z(n1813) );
  ANDN U2653 ( .B(n1813), .A(n2868), .Z(n1814) );
  XNOR U2654 ( .A(zin[76]), .B(n1814), .Z(n4040) );
  NANDN U2655 ( .A(n4041), .B(n4040), .Z(n3054) );
  XNOR U2656 ( .A(n4041), .B(n4040), .Z(n2258) );
  XOR U2657 ( .A(y[76]), .B(n1815), .Z(n1816) );
  ANDN U2658 ( .B(n1816), .A(n2868), .Z(n1817) );
  XNOR U2659 ( .A(zin[75]), .B(n1817), .Z(n4045) );
  NAND U2660 ( .A(n4045), .B(n[76]), .Z(n2256) );
  XOR U2661 ( .A(n[76]), .B(n4045), .Z(n2254) );
  XOR U2662 ( .A(y[75]), .B(n1818), .Z(n1819) );
  ANDN U2663 ( .B(n1819), .A(n2868), .Z(n1820) );
  XNOR U2664 ( .A(zin[74]), .B(n1820), .Z(n4049) );
  NAND U2665 ( .A(n[75]), .B(n4049), .Z(n2252) );
  XOR U2666 ( .A(n4049), .B(n[75]), .Z(n2250) );
  XOR U2667 ( .A(y[74]), .B(n1821), .Z(n1822) );
  ANDN U2668 ( .B(n1822), .A(n2868), .Z(n1823) );
  XOR U2669 ( .A(zin[73]), .B(n1823), .Z(n2877) );
  NANDN U2670 ( .A(n2877), .B(n[74]), .Z(n2248) );
  XNOR U2671 ( .A(n[74]), .B(n2877), .Z(n2246) );
  XOR U2672 ( .A(y[73]), .B(n1824), .Z(n1825) );
  ANDN U2673 ( .B(n1825), .A(n2868), .Z(n1826) );
  XNOR U2674 ( .A(zin[72]), .B(n1826), .Z(n4057) );
  NAND U2675 ( .A(n[73]), .B(n4057), .Z(n2244) );
  XOR U2676 ( .A(n4057), .B(n[73]), .Z(n2242) );
  XOR U2677 ( .A(y[72]), .B(n1827), .Z(n1828) );
  ANDN U2678 ( .B(n1828), .A(n2868), .Z(n1829) );
  XOR U2679 ( .A(zin[71]), .B(n1829), .Z(n2878) );
  NANDN U2680 ( .A(n2878), .B(n[72]), .Z(n2240) );
  XNOR U2681 ( .A(n[72]), .B(n2878), .Z(n2238) );
  IV U2682 ( .A(n[71]), .Z(n5390) );
  XOR U2683 ( .A(y[71]), .B(n1830), .Z(n1831) );
  ANDN U2684 ( .B(n1831), .A(n2868), .Z(n1832) );
  XNOR U2685 ( .A(zin[70]), .B(n1832), .Z(n4065) );
  NANDN U2686 ( .A(n5390), .B(n4065), .Z(n2236) );
  XNOR U2687 ( .A(n4065), .B(n5390), .Z(n2234) );
  IV U2688 ( .A(n[70]), .Z(n5469) );
  XOR U2689 ( .A(y[70]), .B(n1833), .Z(n1834) );
  ANDN U2690 ( .B(n1834), .A(n2868), .Z(n1835) );
  XNOR U2691 ( .A(zin[69]), .B(n1835), .Z(n4069) );
  NANDN U2692 ( .A(n5469), .B(n4069), .Z(n3045) );
  XNOR U2693 ( .A(n4069), .B(n5469), .Z(n2231) );
  XOR U2694 ( .A(y[69]), .B(n1836), .Z(n1837) );
  ANDN U2695 ( .B(n1837), .A(n2868), .Z(n1838) );
  XNOR U2696 ( .A(zin[68]), .B(n1838), .Z(n4073) );
  NAND U2697 ( .A(n[69]), .B(n4073), .Z(n2229) );
  XOR U2698 ( .A(n4073), .B(n[69]), .Z(n2227) );
  XOR U2699 ( .A(y[67]), .B(n1839), .Z(n1840) );
  ANDN U2700 ( .B(n1840), .A(n2868), .Z(n1841) );
  XNOR U2701 ( .A(zin[66]), .B(n1841), .Z(n4082) );
  NAND U2702 ( .A(n[67]), .B(n4082), .Z(n1845) );
  XOR U2703 ( .A(y[68]), .B(n1842), .Z(n1843) );
  ANDN U2704 ( .B(n1843), .A(n2868), .Z(n1844) );
  XNOR U2705 ( .A(zin[67]), .B(n1844), .Z(n4077) );
  AND U2706 ( .A(n4077), .B(n[68]), .Z(n3040) );
  ANDN U2707 ( .B(n1845), .A(n3040), .Z(n2224) );
  XOR U2708 ( .A(n4082), .B(n[67]), .Z(n2222) );
  XOR U2709 ( .A(y[66]), .B(n1846), .Z(n1847) );
  ANDN U2710 ( .B(n1847), .A(n2868), .Z(n1848) );
  XNOR U2711 ( .A(zin[65]), .B(n1848), .Z(n4086) );
  NAND U2712 ( .A(n4086), .B(n[66]), .Z(n2220) );
  XOR U2713 ( .A(n[66]), .B(n4086), .Z(n2218) );
  XOR U2714 ( .A(y[65]), .B(n1849), .Z(n1850) );
  ANDN U2715 ( .B(n1850), .A(n2868), .Z(n1851) );
  XNOR U2716 ( .A(zin[64]), .B(n1851), .Z(n4090) );
  AND U2717 ( .A(n4090), .B(n[65]), .Z(n3037) );
  IV U2718 ( .A(n[65]), .Z(n4091) );
  ANDN U2719 ( .B(n4091), .A(n4090), .Z(n3038) );
  XOR U2720 ( .A(y[64]), .B(n1852), .Z(n1853) );
  ANDN U2721 ( .B(n1853), .A(n2868), .Z(n1854) );
  XOR U2722 ( .A(zin[63]), .B(n1854), .Z(n4095) );
  IV U2723 ( .A(n[64]), .Z(n5399) );
  AND U2724 ( .A(n4095), .B(n5399), .Z(n3036) );
  NOR U2725 ( .A(n3038), .B(n3036), .Z(n2215) );
  XOR U2726 ( .A(y[62]), .B(n1855), .Z(n1856) );
  ANDN U2727 ( .B(n1856), .A(n2868), .Z(n1857) );
  XOR U2728 ( .A(zin[61]), .B(n1857), .Z(n4103) );
  NANDN U2729 ( .A(n[62]), .B(n4103), .Z(n3031) );
  XOR U2730 ( .A(y[61]), .B(n1858), .Z(n1859) );
  ANDN U2731 ( .B(n1859), .A(n2868), .Z(n1860) );
  XOR U2732 ( .A(zin[60]), .B(n1860), .Z(n4107) );
  IV U2733 ( .A(n[61]), .Z(n4108) );
  AND U2734 ( .A(n4107), .B(n4108), .Z(n3030) );
  ANDN U2735 ( .B(n3031), .A(n3030), .Z(n2204) );
  XOR U2736 ( .A(y[58]), .B(n1861), .Z(n1862) );
  ANDN U2737 ( .B(n1862), .A(n2868), .Z(n1863) );
  XOR U2738 ( .A(zin[57]), .B(n1863), .Z(n4122) );
  IV U2739 ( .A(n[58]), .Z(n5411) );
  AND U2740 ( .A(n4122), .B(n5411), .Z(n3019) );
  XOR U2741 ( .A(y[59]), .B(n1864), .Z(n1865) );
  ANDN U2742 ( .B(n1865), .A(n2868), .Z(n1866) );
  XOR U2743 ( .A(zin[58]), .B(n1866), .Z(n4117) );
  IV U2744 ( .A(n[59]), .Z(n4118) );
  AND U2745 ( .A(n4117), .B(n4118), .Z(n3022) );
  NOR U2746 ( .A(n3019), .B(n3022), .Z(n2193) );
  IV U2747 ( .A(n[56]), .Z(n4131) );
  XOR U2748 ( .A(y[56]), .B(n1867), .Z(n1868) );
  ANDN U2749 ( .B(n1868), .A(n2868), .Z(n1869) );
  XNOR U2750 ( .A(zin[55]), .B(n1869), .Z(n4130) );
  ANDN U2751 ( .B(n4131), .A(n4130), .Z(n3018) );
  XOR U2752 ( .A(y[55]), .B(n1870), .Z(n1871) );
  ANDN U2753 ( .B(n1871), .A(n2868), .Z(n1872) );
  XNOR U2754 ( .A(zin[54]), .B(n1872), .Z(n4135) );
  AND U2755 ( .A(n4135), .B(n[55]), .Z(n3013) );
  XOR U2756 ( .A(y[54]), .B(n1873), .Z(n1874) );
  ANDN U2757 ( .B(n1874), .A(n2868), .Z(n1875) );
  XNOR U2758 ( .A(zin[53]), .B(n1875), .Z(n4139) );
  AND U2759 ( .A(n4139), .B(n[54]), .Z(n3010) );
  IV U2760 ( .A(n[54]), .Z(n4140) );
  ANDN U2761 ( .B(n4140), .A(n4139), .Z(n3012) );
  XOR U2762 ( .A(y[53]), .B(n1876), .Z(n1877) );
  ANDN U2763 ( .B(n1877), .A(n2868), .Z(n1878) );
  XOR U2764 ( .A(zin[52]), .B(n1878), .Z(n4144) );
  ANDN U2765 ( .B(n[53]), .A(n4144), .Z(n3009) );
  IV U2766 ( .A(n[53]), .Z(n4145) );
  AND U2767 ( .A(n4144), .B(n4145), .Z(n3007) );
  XOR U2768 ( .A(y[52]), .B(n1879), .Z(n1880) );
  ANDN U2769 ( .B(n1880), .A(n2868), .Z(n1881) );
  XNOR U2770 ( .A(zin[51]), .B(n1881), .Z(n4149) );
  AND U2771 ( .A(n4149), .B(n[52]), .Z(n3006) );
  OR U2772 ( .A(n4149), .B(n[52]), .Z(n3004) );
  XOR U2773 ( .A(y[50]), .B(n1882), .Z(n1883) );
  ANDN U2774 ( .B(n1883), .A(n2868), .Z(n1884) );
  XOR U2775 ( .A(zin[49]), .B(n1884), .Z(n4157) );
  IV U2776 ( .A(n4157), .Z(n2165) );
  NOR U2777 ( .A(n2165), .B(n[50]), .Z(n3001) );
  XOR U2778 ( .A(y[49]), .B(n1885), .Z(n1886) );
  ANDN U2779 ( .B(n1886), .A(n2868), .Z(n1887) );
  XNOR U2780 ( .A(zin[48]), .B(n1887), .Z(n4161) );
  AND U2781 ( .A(n4161), .B(n[49]), .Z(n3000) );
  XOR U2782 ( .A(y[48]), .B(n1888), .Z(n1889) );
  ANDN U2783 ( .B(n1889), .A(n2868), .Z(n1890) );
  XOR U2784 ( .A(zin[47]), .B(n1890), .Z(n4166) );
  ANDN U2785 ( .B(n[48]), .A(n4166), .Z(n2997) );
  XOR U2786 ( .A(y[47]), .B(n1891), .Z(n1892) );
  ANDN U2787 ( .B(n1892), .A(n2868), .Z(n1893) );
  XNOR U2788 ( .A(zin[46]), .B(n1893), .Z(n4170) );
  AND U2789 ( .A(n4170), .B(n[47]), .Z(n2992) );
  IV U2790 ( .A(n[47]), .Z(n6716) );
  NANDN U2791 ( .A(n4170), .B(n6716), .Z(n2994) );
  XOR U2792 ( .A(y[46]), .B(n1894), .Z(n1895) );
  ANDN U2793 ( .B(n1895), .A(n2868), .Z(n1896) );
  XOR U2794 ( .A(zin[45]), .B(n1896), .Z(n4174) );
  IV U2795 ( .A(n[46]), .Z(n6710) );
  AND U2796 ( .A(n4174), .B(n6710), .Z(n2991) );
  ANDN U2797 ( .B(n2994), .A(n2991), .Z(n2158) );
  XOR U2798 ( .A(y[44]), .B(n1897), .Z(n1898) );
  ANDN U2799 ( .B(n1898), .A(n2868), .Z(n1899) );
  XNOR U2800 ( .A(zin[43]), .B(n1899), .Z(n4470) );
  NOR U2801 ( .A(n[44]), .B(n4470), .Z(n2988) );
  XOR U2802 ( .A(y[43]), .B(n1900), .Z(n1901) );
  ANDN U2803 ( .B(n1901), .A(n2868), .Z(n1902) );
  XNOR U2804 ( .A(zin[42]), .B(n1902), .Z(n4466) );
  AND U2805 ( .A(n4466), .B(n[43]), .Z(n2985) );
  XOR U2806 ( .A(y[42]), .B(n1903), .Z(n1904) );
  ANDN U2807 ( .B(n1904), .A(n2868), .Z(n1905) );
  XOR U2808 ( .A(zin[41]), .B(n1905), .Z(n4178) );
  ANDN U2809 ( .B(n[42]), .A(n4178), .Z(n2982) );
  IV U2810 ( .A(n[42]), .Z(n4179) );
  AND U2811 ( .A(n4178), .B(n4179), .Z(n2980) );
  XOR U2812 ( .A(y[41]), .B(n1906), .Z(n1907) );
  ANDN U2813 ( .B(n1907), .A(n2868), .Z(n1908) );
  XOR U2814 ( .A(zin[40]), .B(n1908), .Z(n4183) );
  ANDN U2815 ( .B(n[41]), .A(n4183), .Z(n2979) );
  NANDN U2816 ( .A(n[41]), .B(n4183), .Z(n2977) );
  XOR U2817 ( .A(y[40]), .B(n1909), .Z(n1910) );
  ANDN U2818 ( .B(n1910), .A(n2868), .Z(n1911) );
  XOR U2819 ( .A(zin[39]), .B(n1911), .Z(n4187) );
  IV U2820 ( .A(n[40]), .Z(n4188) );
  AND U2821 ( .A(n4187), .B(n4188), .Z(n2976) );
  ANDN U2822 ( .B(n2977), .A(n2976), .Z(n2141) );
  IV U2823 ( .A(n[38]), .Z(n4197) );
  XOR U2824 ( .A(y[38]), .B(n1912), .Z(n1913) );
  ANDN U2825 ( .B(n1913), .A(n2868), .Z(n1914) );
  XNOR U2826 ( .A(zin[37]), .B(n1914), .Z(n4196) );
  ANDN U2827 ( .B(n4197), .A(n4196), .Z(n2970) );
  XOR U2828 ( .A(y[37]), .B(n1915), .Z(n1916) );
  ANDN U2829 ( .B(n1916), .A(n2868), .Z(n1917) );
  XNOR U2830 ( .A(zin[36]), .B(n1917), .Z(n4201) );
  AND U2831 ( .A(n4201), .B(n[37]), .Z(n2965) );
  XOR U2832 ( .A(y[36]), .B(n1918), .Z(n1919) );
  ANDN U2833 ( .B(n1919), .A(n2868), .Z(n1920) );
  XNOR U2834 ( .A(zin[35]), .B(n1920), .Z(n4205) );
  AND U2835 ( .A(n4205), .B(n[36]), .Z(n2962) );
  XOR U2836 ( .A(y[34]), .B(n1921), .Z(n1922) );
  ANDN U2837 ( .B(n1922), .A(n2868), .Z(n1923) );
  XNOR U2838 ( .A(zin[33]), .B(n1923), .Z(n4209) );
  NAND U2839 ( .A(n[34]), .B(n4209), .Z(n2118) );
  XOR U2840 ( .A(n4209), .B(n[34]), .Z(n2116) );
  XOR U2841 ( .A(y[33]), .B(n1924), .Z(n1925) );
  ANDN U2842 ( .B(n1925), .A(n2868), .Z(n1926) );
  XNOR U2843 ( .A(zin[32]), .B(n1926), .Z(n4213) );
  NAND U2844 ( .A(n[33]), .B(n4213), .Z(n2114) );
  XOR U2845 ( .A(n4213), .B(n[33]), .Z(n2112) );
  XOR U2846 ( .A(y[32]), .B(n1927), .Z(n1928) );
  ANDN U2847 ( .B(n1928), .A(n2868), .Z(n1929) );
  XNOR U2848 ( .A(zin[31]), .B(n1929), .Z(n4217) );
  NAND U2849 ( .A(n4217), .B(n[32]), .Z(n2110) );
  XOR U2850 ( .A(n[32]), .B(n4217), .Z(n2108) );
  IV U2851 ( .A(n[31]), .Z(n4416) );
  XOR U2852 ( .A(y[31]), .B(n1930), .Z(n1931) );
  ANDN U2853 ( .B(n1931), .A(n2868), .Z(n1932) );
  XNOR U2854 ( .A(zin[30]), .B(n1932), .Z(n4419) );
  NANDN U2855 ( .A(n4416), .B(n4419), .Z(n2961) );
  XNOR U2856 ( .A(n4416), .B(n4419), .Z(n2105) );
  IV U2857 ( .A(n[30]), .Z(n4222) );
  XOR U2858 ( .A(y[30]), .B(n1933), .Z(n1934) );
  ANDN U2859 ( .B(n1934), .A(n2868), .Z(n1935) );
  XNOR U2860 ( .A(zin[29]), .B(n1935), .Z(n4221) );
  NANDN U2861 ( .A(n4222), .B(n4221), .Z(n2958) );
  XNOR U2862 ( .A(n4221), .B(n4222), .Z(n2102) );
  IV U2863 ( .A(n[29]), .Z(n4407) );
  XOR U2864 ( .A(y[29]), .B(n1936), .Z(n1937) );
  ANDN U2865 ( .B(n1937), .A(n2868), .Z(n1938) );
  XNOR U2866 ( .A(zin[28]), .B(n1938), .Z(n4226) );
  NANDN U2867 ( .A(n4407), .B(n4226), .Z(n2955) );
  XNOR U2868 ( .A(n4407), .B(n4226), .Z(n2099) );
  XOR U2869 ( .A(y[28]), .B(n1939), .Z(n1940) );
  ANDN U2870 ( .B(n1940), .A(n2868), .Z(n1941) );
  XNOR U2871 ( .A(zin[27]), .B(n1941), .Z(n4406) );
  NAND U2872 ( .A(n[28]), .B(n4406), .Z(n2952) );
  XOR U2873 ( .A(n[28]), .B(n4406), .Z(n2096) );
  IV U2874 ( .A(n[27]), .Z(n4399) );
  XOR U2875 ( .A(y[27]), .B(n1942), .Z(n1943) );
  ANDN U2876 ( .B(n1943), .A(n2868), .Z(n1944) );
  XOR U2877 ( .A(zin[26]), .B(n1944), .Z(n4402) );
  IV U2878 ( .A(n4402), .Z(n2879) );
  NANDN U2879 ( .A(n4399), .B(n2879), .Z(n2094) );
  XNOR U2880 ( .A(n4402), .B(n[27]), .Z(n2092) );
  XOR U2881 ( .A(y[26]), .B(n1945), .Z(n1946) );
  ANDN U2882 ( .B(n1946), .A(n2868), .Z(n1947) );
  XNOR U2883 ( .A(zin[25]), .B(n1947), .Z(n4230) );
  NAND U2884 ( .A(n4230), .B(n[26]), .Z(n2090) );
  XOR U2885 ( .A(n[26]), .B(n4230), .Z(n2088) );
  XOR U2886 ( .A(y[25]), .B(n1948), .Z(n1949) );
  ANDN U2887 ( .B(n1949), .A(n2868), .Z(n1950) );
  XNOR U2888 ( .A(zin[24]), .B(n1950), .Z(n4234) );
  NAND U2889 ( .A(n[25]), .B(n4234), .Z(n2086) );
  XOR U2890 ( .A(n4234), .B(n[25]), .Z(n2084) );
  IV U2891 ( .A(n[24]), .Z(n4239) );
  XOR U2892 ( .A(y[24]), .B(n1951), .Z(n1952) );
  ANDN U2893 ( .B(n1952), .A(n2868), .Z(n1953) );
  XNOR U2894 ( .A(zin[23]), .B(n1953), .Z(n4238) );
  NANDN U2895 ( .A(n4239), .B(n4238), .Z(n2949) );
  XNOR U2896 ( .A(n4238), .B(n4239), .Z(n2081) );
  IV U2897 ( .A(n[23]), .Z(n4387) );
  XOR U2898 ( .A(y[23]), .B(n1954), .Z(n1955) );
  ANDN U2899 ( .B(n1955), .A(n2868), .Z(n1956) );
  XNOR U2900 ( .A(zin[22]), .B(n1956), .Z(n4390) );
  NANDN U2901 ( .A(n4387), .B(n4390), .Z(n2946) );
  XNOR U2902 ( .A(n4387), .B(n4390), .Z(n2078) );
  IV U2903 ( .A(n[22]), .Z(n4382) );
  XOR U2904 ( .A(y[22]), .B(n1957), .Z(n1958) );
  ANDN U2905 ( .B(n1958), .A(n2868), .Z(n1959) );
  XNOR U2906 ( .A(zin[21]), .B(n1959), .Z(n4243) );
  NANDN U2907 ( .A(n4382), .B(n4243), .Z(n2943) );
  XNOR U2908 ( .A(n4243), .B(n4382), .Z(n2075) );
  XOR U2909 ( .A(y[21]), .B(n1960), .Z(n1961) );
  ANDN U2910 ( .B(n1961), .A(n2868), .Z(n1962) );
  XNOR U2911 ( .A(zin[20]), .B(n1962), .Z(n4381) );
  NAND U2912 ( .A(n[21]), .B(n4381), .Z(n2940) );
  XOR U2913 ( .A(n[21]), .B(n4381), .Z(n2072) );
  IV U2914 ( .A(n[20]), .Z(n4248) );
  XOR U2915 ( .A(y[20]), .B(n1963), .Z(n1964) );
  ANDN U2916 ( .B(n1964), .A(n2868), .Z(n1965) );
  XNOR U2917 ( .A(zin[19]), .B(n1965), .Z(n4247) );
  NANDN U2918 ( .A(n4248), .B(n4247), .Z(n2937) );
  XNOR U2919 ( .A(n4247), .B(n4248), .Z(n2069) );
  IV U2920 ( .A(n[19]), .Z(n4370) );
  XOR U2921 ( .A(y[19]), .B(n1966), .Z(n1967) );
  ANDN U2922 ( .B(n1967), .A(n2868), .Z(n1968) );
  XNOR U2923 ( .A(zin[18]), .B(n1968), .Z(n4252) );
  NANDN U2924 ( .A(n4370), .B(n4252), .Z(n2934) );
  XNOR U2925 ( .A(n4370), .B(n4252), .Z(n2066) );
  IV U2926 ( .A(n[18]), .Z(n4257) );
  XOR U2927 ( .A(y[18]), .B(n1969), .Z(n1970) );
  ANDN U2928 ( .B(n1970), .A(n2868), .Z(n1971) );
  XNOR U2929 ( .A(zin[17]), .B(n1971), .Z(n4256) );
  NANDN U2930 ( .A(n4257), .B(n4256), .Z(n2931) );
  XNOR U2931 ( .A(n4257), .B(n4256), .Z(n2063) );
  XOR U2932 ( .A(y[17]), .B(n1972), .Z(n1973) );
  ANDN U2933 ( .B(n1973), .A(n2868), .Z(n1974) );
  XOR U2934 ( .A(zin[16]), .B(n1974), .Z(n4261) );
  ANDN U2935 ( .B(n[17]), .A(n4261), .Z(n2928) );
  XOR U2936 ( .A(y[16]), .B(n1975), .Z(n1976) );
  ANDN U2937 ( .B(n1976), .A(n2868), .Z(n1977) );
  XOR U2938 ( .A(zin[15]), .B(n1977), .Z(n4265) );
  IV U2939 ( .A(n[16]), .Z(n4266) );
  AND U2940 ( .A(n4265), .B(n4266), .Z(n2923) );
  IV U2941 ( .A(n[17]), .Z(n4362) );
  AND U2942 ( .A(n4261), .B(n4362), .Z(n2926) );
  NOR U2943 ( .A(n2923), .B(n2926), .Z(n2060) );
  ANDN U2944 ( .B(n[16]), .A(n4265), .Z(n2925) );
  XOR U2945 ( .A(y[15]), .B(n1978), .Z(n1979) );
  ANDN U2946 ( .B(n1979), .A(n2868), .Z(n1980) );
  XNOR U2947 ( .A(zin[14]), .B(n1980), .Z(n4361) );
  NOR U2948 ( .A(n[15]), .B(n4361), .Z(n2920) );
  XOR U2949 ( .A(y[13]), .B(n1981), .Z(n1982) );
  ANDN U2950 ( .B(n1982), .A(n2868), .Z(n1983) );
  XOR U2951 ( .A(zin[12]), .B(n1983), .Z(n4275) );
  ANDN U2952 ( .B(n[13]), .A(n4275), .Z(n2916) );
  XOR U2953 ( .A(y[12]), .B(n1984), .Z(n1985) );
  ANDN U2954 ( .B(n1985), .A(n2868), .Z(n1986) );
  XOR U2955 ( .A(zin[11]), .B(n1986), .Z(n4348) );
  IV U2956 ( .A(n4348), .Z(n1987) );
  AND U2957 ( .A(n[12]), .B(n1987), .Z(n2913) );
  NOR U2958 ( .A(n1987), .B(n[12]), .Z(n2911) );
  XOR U2959 ( .A(y[11]), .B(n1988), .Z(n1989) );
  ANDN U2960 ( .B(n1989), .A(n2868), .Z(n1990) );
  XOR U2961 ( .A(zin[10]), .B(n1990), .Z(n4341) );
  ANDN U2962 ( .B(n[11]), .A(n4341), .Z(n2910) );
  IV U2963 ( .A(n[11]), .Z(n4337) );
  AND U2964 ( .A(n4341), .B(n4337), .Z(n2908) );
  XOR U2965 ( .A(y[7]), .B(n1991), .Z(n1992) );
  ANDN U2966 ( .B(n1992), .A(n2868), .Z(n1993) );
  XNOR U2967 ( .A(zin[6]), .B(n1993), .Z(n4283) );
  AND U2968 ( .A(n4283), .B(n[7]), .Z(n2896) );
  OR U2969 ( .A(n4283), .B(n[7]), .Z(n2897) );
  XOR U2970 ( .A(y[6]), .B(n1994), .Z(n1995) );
  ANDN U2971 ( .B(n1995), .A(n2868), .Z(n1996) );
  XNOR U2972 ( .A(zin[5]), .B(n1996), .Z(n4287) );
  OR U2973 ( .A(n4287), .B(n[6]), .Z(n2893) );
  AND U2974 ( .A(n2897), .B(n2893), .Z(n2026) );
  XOR U2975 ( .A(y[4]), .B(n1997), .Z(n1998) );
  ANDN U2976 ( .B(n1998), .A(n2868), .Z(n1999) );
  XNOR U2977 ( .A(zin[3]), .B(n1999), .Z(n4295) );
  OR U2978 ( .A(n4295), .B(n[4]), .Z(n2887) );
  XOR U2979 ( .A(y[3]), .B(n2000), .Z(n2001) );
  ANDN U2980 ( .B(n2001), .A(n2868), .Z(n2002) );
  XNOR U2981 ( .A(zin[2]), .B(n2002), .Z(n4307) );
  OR U2982 ( .A(n4307), .B(n[3]), .Z(n2884) );
  AND U2983 ( .A(n2887), .B(n2884), .Z(n2017) );
  IV U2984 ( .A(n[2]), .Z(n6616) );
  XNOR U2985 ( .A(y[2]), .B(n2003), .Z(n2004) );
  ANDN U2986 ( .B(n2004), .A(n2868), .Z(n2005) );
  XNOR U2987 ( .A(zin[1]), .B(n2005), .Z(n4303) );
  NANDN U2988 ( .A(n6616), .B(n4303), .Z(n2014) );
  XNOR U2989 ( .A(n6616), .B(n4303), .Z(n2012) );
  NANDN U2990 ( .A(n[0]), .B(n2880), .Z(n2007) );
  NAND U2991 ( .A(n[1]), .B(n2007), .Z(n2010) );
  NANDN U2992 ( .A(n2868), .B(y[1]), .Z(n2006) );
  XNOR U2993 ( .A(zin[0]), .B(n2006), .Z(n4299) );
  XOR U2994 ( .A(n2007), .B(n[1]), .Z(n2008) );
  NANDN U2995 ( .A(n4299), .B(n2008), .Z(n2009) );
  NAND U2996 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U2997 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2998 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U2999 ( .A(n[3]), .B(n4307), .Z(n2886) );
  NANDN U3000 ( .A(n2015), .B(n2886), .Z(n2016) );
  AND U3001 ( .A(n2017), .B(n2016), .Z(n2018) );
  NAND U3002 ( .A(n[4]), .B(n4295), .Z(n2889) );
  NANDN U3003 ( .A(n2018), .B(n2889), .Z(n2022) );
  XOR U3004 ( .A(y[5]), .B(n2019), .Z(n2020) );
  ANDN U3005 ( .B(n2020), .A(n2868), .Z(n2021) );
  XOR U3006 ( .A(zin[4]), .B(n2021), .Z(n4291) );
  NANDN U3007 ( .A(n[5]), .B(n4291), .Z(n2890) );
  NAND U3008 ( .A(n2022), .B(n2890), .Z(n2023) );
  NAND U3009 ( .A(n[6]), .B(n4287), .Z(n2895) );
  NAND U3010 ( .A(n2023), .B(n2895), .Z(n2024) );
  NANDN U3011 ( .A(n4291), .B(n[5]), .Z(n2892) );
  NANDN U3012 ( .A(n2024), .B(n2892), .Z(n2025) );
  AND U3013 ( .A(n2026), .B(n2025), .Z(n2027) );
  OR U3014 ( .A(n2896), .B(n2027), .Z(n2031) );
  XOR U3015 ( .A(y[8]), .B(n2028), .Z(n2029) );
  ANDN U3016 ( .B(n2029), .A(n2868), .Z(n2030) );
  XOR U3017 ( .A(zin[7]), .B(n2030), .Z(n4279) );
  NANDN U3018 ( .A(n[8]), .B(n4279), .Z(n2900) );
  NAND U3019 ( .A(n2031), .B(n2900), .Z(n2032) );
  ANDN U3020 ( .B(n[8]), .A(n4279), .Z(n2899) );
  ANDN U3021 ( .B(n2032), .A(n2899), .Z(n2040) );
  XNOR U3022 ( .A(y[9]), .B(n2033), .Z(n2034) );
  ANDN U3023 ( .B(n2034), .A(n2868), .Z(n2035) );
  XNOR U3024 ( .A(zin[8]), .B(n2035), .Z(n4329) );
  NANDN U3025 ( .A(n2040), .B(n4329), .Z(n2039) );
  XOR U3026 ( .A(y[10]), .B(n2036), .Z(n2037) );
  ANDN U3027 ( .B(n2037), .A(n2868), .Z(n2038) );
  XNOR U3028 ( .A(zin[9]), .B(n2038), .Z(n4333) );
  AND U3029 ( .A(n4333), .B(n[10]), .Z(n2907) );
  ANDN U3030 ( .B(n2039), .A(n2907), .Z(n2043) );
  IV U3031 ( .A(n[9]), .Z(n6868) );
  XNOR U3032 ( .A(n4329), .B(n2040), .Z(n2041) );
  NANDN U3033 ( .A(n6868), .B(n2041), .Z(n2042) );
  NAND U3034 ( .A(n2043), .B(n2042), .Z(n2044) );
  NOR U3035 ( .A(n[10]), .B(n4333), .Z(n2905) );
  ANDN U3036 ( .B(n2044), .A(n2905), .Z(n2045) );
  NANDN U3037 ( .A(n2908), .B(n2045), .Z(n2046) );
  NANDN U3038 ( .A(n2910), .B(n2046), .Z(n2047) );
  NANDN U3039 ( .A(n2911), .B(n2047), .Z(n2048) );
  NANDN U3040 ( .A(n2913), .B(n2048), .Z(n2049) );
  IV U3041 ( .A(n[13]), .Z(n4349) );
  AND U3042 ( .A(n4275), .B(n4349), .Z(n2914) );
  ANDN U3043 ( .B(n2049), .A(n2914), .Z(n2053) );
  XOR U3044 ( .A(y[14]), .B(n2050), .Z(n2051) );
  ANDN U3045 ( .B(n2051), .A(n2868), .Z(n2052) );
  XOR U3046 ( .A(zin[13]), .B(n2052), .Z(n4270) );
  ANDN U3047 ( .B(n[14]), .A(n4270), .Z(n2919) );
  NOR U3048 ( .A(n2053), .B(n2919), .Z(n2054) );
  NANDN U3049 ( .A(n2916), .B(n2054), .Z(n2055) );
  IV U3050 ( .A(n[14]), .Z(n4271) );
  AND U3051 ( .A(n4270), .B(n4271), .Z(n2917) );
  ANDN U3052 ( .B(n2055), .A(n2917), .Z(n2056) );
  NANDN U3053 ( .A(n2920), .B(n2056), .Z(n2057) );
  AND U3054 ( .A(n4361), .B(n[15]), .Z(n2922) );
  ANDN U3055 ( .B(n2057), .A(n2922), .Z(n2058) );
  NANDN U3056 ( .A(n2925), .B(n2058), .Z(n2059) );
  NAND U3057 ( .A(n2060), .B(n2059), .Z(n2061) );
  NANDN U3058 ( .A(n2928), .B(n2061), .Z(n2062) );
  NAND U3059 ( .A(n2063), .B(n2062), .Z(n2064) );
  NAND U3060 ( .A(n2931), .B(n2064), .Z(n2065) );
  NAND U3061 ( .A(n2066), .B(n2065), .Z(n2067) );
  NAND U3062 ( .A(n2934), .B(n2067), .Z(n2068) );
  NAND U3063 ( .A(n2069), .B(n2068), .Z(n2070) );
  NAND U3064 ( .A(n2937), .B(n2070), .Z(n2071) );
  NAND U3065 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U3066 ( .A(n2940), .B(n2073), .Z(n2074) );
  NAND U3067 ( .A(n2075), .B(n2074), .Z(n2076) );
  NAND U3068 ( .A(n2943), .B(n2076), .Z(n2077) );
  NAND U3069 ( .A(n2078), .B(n2077), .Z(n2079) );
  NAND U3070 ( .A(n2946), .B(n2079), .Z(n2080) );
  NAND U3071 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U3072 ( .A(n2949), .B(n2082), .Z(n2083) );
  NAND U3073 ( .A(n2084), .B(n2083), .Z(n2085) );
  NAND U3074 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U3075 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U3076 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U3077 ( .A(n2092), .B(n2091), .Z(n2093) );
  NAND U3078 ( .A(n2094), .B(n2093), .Z(n2095) );
  NAND U3079 ( .A(n2096), .B(n2095), .Z(n2097) );
  NAND U3080 ( .A(n2952), .B(n2097), .Z(n2098) );
  NAND U3081 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U3082 ( .A(n2955), .B(n2100), .Z(n2101) );
  NAND U3083 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U3084 ( .A(n2958), .B(n2103), .Z(n2104) );
  NAND U3085 ( .A(n2105), .B(n2104), .Z(n2106) );
  NAND U3086 ( .A(n2961), .B(n2106), .Z(n2107) );
  NAND U3087 ( .A(n2108), .B(n2107), .Z(n2109) );
  NAND U3088 ( .A(n2110), .B(n2109), .Z(n2111) );
  NAND U3089 ( .A(n2112), .B(n2111), .Z(n2113) );
  NAND U3090 ( .A(n2114), .B(n2113), .Z(n2115) );
  NAND U3091 ( .A(n2116), .B(n2115), .Z(n2117) );
  AND U3092 ( .A(n2118), .B(n2117), .Z(n2122) );
  XOR U3093 ( .A(y[35]), .B(n2119), .Z(n2120) );
  ANDN U3094 ( .B(n2120), .A(n2868), .Z(n2121) );
  XNOR U3095 ( .A(zin[34]), .B(n2121), .Z(n4431) );
  NANDN U3096 ( .A(n2122), .B(n4431), .Z(n2125) );
  IV U3097 ( .A(n[35]), .Z(n4432) );
  XNOR U3098 ( .A(n4431), .B(n2122), .Z(n2123) );
  NANDN U3099 ( .A(n4432), .B(n2123), .Z(n2124) );
  NAND U3100 ( .A(n2125), .B(n2124), .Z(n2126) );
  IV U3101 ( .A(n[36]), .Z(n6656) );
  ANDN U3102 ( .B(n6656), .A(n4205), .Z(n2964) );
  ANDN U3103 ( .B(n2126), .A(n2964), .Z(n2127) );
  OR U3104 ( .A(n2962), .B(n2127), .Z(n2128) );
  IV U3105 ( .A(n[37]), .Z(n4438) );
  ANDN U3106 ( .B(n4438), .A(n4201), .Z(n2967) );
  ANDN U3107 ( .B(n2128), .A(n2967), .Z(n2129) );
  OR U3108 ( .A(n2965), .B(n2129), .Z(n2130) );
  NANDN U3109 ( .A(n2970), .B(n2130), .Z(n2131) );
  AND U3110 ( .A(n4196), .B(n[38]), .Z(n2968) );
  ANDN U3111 ( .B(n2131), .A(n2968), .Z(n2133) );
  IV U3112 ( .A(n[39]), .Z(n4446) );
  OR U3113 ( .A(n2133), .B(n4446), .Z(n2132) );
  ANDN U3114 ( .B(n[40]), .A(n4187), .Z(n2974) );
  ANDN U3115 ( .B(n2132), .A(n2974), .Z(n2139) );
  XOR U3116 ( .A(n4446), .B(n2133), .Z(n2137) );
  XOR U3117 ( .A(y[39]), .B(n2134), .Z(n2135) );
  ANDN U3118 ( .B(n2135), .A(n2868), .Z(n2136) );
  XNOR U3119 ( .A(zin[38]), .B(n2136), .Z(n4192) );
  NAND U3120 ( .A(n2137), .B(n4192), .Z(n2138) );
  NAND U3121 ( .A(n2139), .B(n2138), .Z(n2140) );
  NAND U3122 ( .A(n2141), .B(n2140), .Z(n2142) );
  NANDN U3123 ( .A(n2979), .B(n2142), .Z(n2143) );
  NANDN U3124 ( .A(n2980), .B(n2143), .Z(n2144) );
  NANDN U3125 ( .A(n2982), .B(n2144), .Z(n2145) );
  NOR U3126 ( .A(n[43]), .B(n4466), .Z(n2983) );
  ANDN U3127 ( .B(n2145), .A(n2983), .Z(n2146) );
  OR U3128 ( .A(n2985), .B(n2146), .Z(n2147) );
  NANDN U3129 ( .A(n2988), .B(n2147), .Z(n2148) );
  AND U3130 ( .A(n4470), .B(n[44]), .Z(n2986) );
  ANDN U3131 ( .B(n2148), .A(n2986), .Z(n2153) );
  XOR U3132 ( .A(y[45]), .B(n2149), .Z(n2150) );
  ANDN U3133 ( .B(n2150), .A(n2868), .Z(n2151) );
  XNOR U3134 ( .A(zin[44]), .B(n2151), .Z(n4474) );
  NANDN U3135 ( .A(n2153), .B(n4474), .Z(n2152) );
  ANDN U3136 ( .B(n2152), .A(n2989), .Z(n2156) );
  XNOR U3137 ( .A(n4474), .B(n2153), .Z(n2154) );
  NAND U3138 ( .A(n[45]), .B(n2154), .Z(n2155) );
  NAND U3139 ( .A(n2156), .B(n2155), .Z(n2157) );
  NAND U3140 ( .A(n2158), .B(n2157), .Z(n2159) );
  NANDN U3141 ( .A(n2992), .B(n2159), .Z(n2160) );
  NANDN U3142 ( .A(n[48]), .B(n4166), .Z(n2995) );
  NAND U3143 ( .A(n2160), .B(n2995), .Z(n2161) );
  NANDN U3144 ( .A(n2997), .B(n2161), .Z(n2162) );
  NOR U3145 ( .A(n[49]), .B(n4161), .Z(n2998) );
  ANDN U3146 ( .B(n2162), .A(n2998), .Z(n2163) );
  OR U3147 ( .A(n3000), .B(n2163), .Z(n2164) );
  NANDN U3148 ( .A(n3001), .B(n2164), .Z(n2166) );
  AND U3149 ( .A(n[50]), .B(n2165), .Z(n3003) );
  ANDN U3150 ( .B(n2166), .A(n3003), .Z(n2170) );
  XOR U3151 ( .A(y[51]), .B(n2167), .Z(n2168) );
  ANDN U3152 ( .B(n2168), .A(n2868), .Z(n2169) );
  XNOR U3153 ( .A(zin[50]), .B(n2169), .Z(n4153) );
  NANDN U3154 ( .A(n2170), .B(n4153), .Z(n2173) );
  XNOR U3155 ( .A(n4153), .B(n2170), .Z(n2171) );
  NAND U3156 ( .A(n[51]), .B(n2171), .Z(n2172) );
  NAND U3157 ( .A(n2173), .B(n2172), .Z(n2174) );
  AND U3158 ( .A(n3004), .B(n2174), .Z(n2175) );
  OR U3159 ( .A(n3006), .B(n2175), .Z(n2176) );
  NANDN U3160 ( .A(n3007), .B(n2176), .Z(n2177) );
  NANDN U3161 ( .A(n3009), .B(n2177), .Z(n2178) );
  NANDN U3162 ( .A(n3012), .B(n2178), .Z(n2179) );
  NANDN U3163 ( .A(n3010), .B(n2179), .Z(n2180) );
  NOR U3164 ( .A(n[55]), .B(n4135), .Z(n3015) );
  ANDN U3165 ( .B(n2180), .A(n3015), .Z(n2181) );
  OR U3166 ( .A(n3013), .B(n2181), .Z(n2182) );
  NANDN U3167 ( .A(n3018), .B(n2182), .Z(n2183) );
  AND U3168 ( .A(n4130), .B(n[56]), .Z(n3016) );
  ANDN U3169 ( .B(n2183), .A(n3016), .Z(n2185) );
  NANDN U3170 ( .A(n2185), .B(n[57]), .Z(n2184) );
  ANDN U3171 ( .B(n[58]), .A(n4122), .Z(n3021) );
  ANDN U3172 ( .B(n2184), .A(n3021), .Z(n2191) );
  XNOR U3173 ( .A(n[57]), .B(n2185), .Z(n2189) );
  XOR U3174 ( .A(y[57]), .B(n2186), .Z(n2187) );
  ANDN U3175 ( .B(n2187), .A(n2868), .Z(n2188) );
  XNOR U3176 ( .A(zin[56]), .B(n2188), .Z(n4126) );
  NAND U3177 ( .A(n2189), .B(n4126), .Z(n2190) );
  NAND U3178 ( .A(n2191), .B(n2190), .Z(n2192) );
  NAND U3179 ( .A(n2193), .B(n2192), .Z(n2194) );
  ANDN U3180 ( .B(n[59]), .A(n4117), .Z(n3024) );
  ANDN U3181 ( .B(n2194), .A(n3024), .Z(n2196) );
  IV U3182 ( .A(n[60]), .Z(n4113) );
  OR U3183 ( .A(n2196), .B(n4113), .Z(n2195) );
  ANDN U3184 ( .B(n[61]), .A(n4107), .Z(n3028) );
  ANDN U3185 ( .B(n2195), .A(n3028), .Z(n2202) );
  XOR U3186 ( .A(n4113), .B(n2196), .Z(n2200) );
  XOR U3187 ( .A(y[60]), .B(n2197), .Z(n2198) );
  ANDN U3188 ( .B(n2198), .A(n2868), .Z(n2199) );
  XNOR U3189 ( .A(zin[59]), .B(n2199), .Z(n4112) );
  NAND U3190 ( .A(n2200), .B(n4112), .Z(n2201) );
  NAND U3191 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U3192 ( .A(n2204), .B(n2203), .Z(n2205) );
  ANDN U3193 ( .B(n[62]), .A(n4103), .Z(n3033) );
  ANDN U3194 ( .B(n2205), .A(n3033), .Z(n2210) );
  XOR U3195 ( .A(y[63]), .B(n2206), .Z(n2207) );
  ANDN U3196 ( .B(n2207), .A(n2868), .Z(n2208) );
  XNOR U3197 ( .A(zin[62]), .B(n2208), .Z(n4099) );
  NANDN U3198 ( .A(n2210), .B(n4099), .Z(n2209) );
  ANDN U3199 ( .B(n[64]), .A(n4095), .Z(n3034) );
  ANDN U3200 ( .B(n2209), .A(n3034), .Z(n2213) );
  XNOR U3201 ( .A(n4099), .B(n2210), .Z(n2211) );
  NAND U3202 ( .A(n[63]), .B(n2211), .Z(n2212) );
  NAND U3203 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U3204 ( .A(n2215), .B(n2214), .Z(n2216) );
  NANDN U3205 ( .A(n3037), .B(n2216), .Z(n2217) );
  NAND U3206 ( .A(n2218), .B(n2217), .Z(n2219) );
  NAND U3207 ( .A(n2220), .B(n2219), .Z(n2221) );
  NAND U3208 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U3209 ( .A(n2224), .B(n2223), .Z(n2225) );
  IV U3210 ( .A(n[68]), .Z(n4078) );
  ANDN U3211 ( .B(n4078), .A(n4077), .Z(n3042) );
  ANDN U3212 ( .B(n2225), .A(n3042), .Z(n2226) );
  NAND U3213 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U3214 ( .A(n2229), .B(n2228), .Z(n2230) );
  NAND U3215 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U3216 ( .A(n3045), .B(n2232), .Z(n2233) );
  NAND U3217 ( .A(n2234), .B(n2233), .Z(n2235) );
  NAND U3218 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U3219 ( .A(n2238), .B(n2237), .Z(n2239) );
  NAND U3220 ( .A(n2240), .B(n2239), .Z(n2241) );
  NAND U3221 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U3222 ( .A(n2244), .B(n2243), .Z(n2245) );
  NAND U3223 ( .A(n2246), .B(n2245), .Z(n2247) );
  NAND U3224 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U3225 ( .A(n2250), .B(n2249), .Z(n2251) );
  NAND U3226 ( .A(n2252), .B(n2251), .Z(n2253) );
  NAND U3227 ( .A(n2254), .B(n2253), .Z(n2255) );
  NAND U3228 ( .A(n2256), .B(n2255), .Z(n2257) );
  NAND U3229 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U3230 ( .A(n3054), .B(n2259), .Z(n2260) );
  NAND U3231 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U3232 ( .A(n2263), .B(n2262), .Z(n2264) );
  NAND U3233 ( .A(n2265), .B(n2264), .Z(n2266) );
  NAND U3234 ( .A(n2267), .B(n2266), .Z(n2268) );
  NAND U3235 ( .A(n2269), .B(n2268), .Z(n2270) );
  NAND U3236 ( .A(n3057), .B(n2270), .Z(n2271) );
  NAND U3237 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U3238 ( .A(n3060), .B(n2273), .Z(n2274) );
  NAND U3239 ( .A(n2275), .B(n2274), .Z(n2276) );
  NAND U3240 ( .A(n2277), .B(n2276), .Z(n2278) );
  NAND U3241 ( .A(n2279), .B(n2278), .Z(n2280) );
  NAND U3242 ( .A(n2281), .B(n2280), .Z(n2282) );
  NAND U3243 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U3244 ( .A(n2285), .B(n2284), .Z(n2286) );
  NAND U3245 ( .A(n2287), .B(n2286), .Z(n2288) );
  NAND U3246 ( .A(n3063), .B(n2288), .Z(n2289) );
  NAND U3247 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U3248 ( .A(n2292), .B(n2291), .Z(n2293) );
  NAND U3249 ( .A(n2294), .B(n2293), .Z(n2295) );
  NAND U3250 ( .A(n3066), .B(n2295), .Z(n2296) );
  NAND U3251 ( .A(n2297), .B(n2296), .Z(n2298) );
  NAND U3252 ( .A(n2299), .B(n2298), .Z(n2300) );
  NAND U3253 ( .A(n2301), .B(n2300), .Z(n2302) );
  NAND U3254 ( .A(n3069), .B(n2302), .Z(n2303) );
  NAND U3255 ( .A(n2304), .B(n2303), .Z(n2305) );
  NAND U3256 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U3257 ( .A(n2308), .B(n2307), .Z(n2309) );
  NAND U3258 ( .A(n3072), .B(n2309), .Z(n2310) );
  NAND U3259 ( .A(n2311), .B(n2310), .Z(n2312) );
  NAND U3260 ( .A(n3075), .B(n2312), .Z(n2313) );
  NAND U3261 ( .A(n2314), .B(n2313), .Z(n2315) );
  NAND U3262 ( .A(n3078), .B(n2315), .Z(n2316) );
  NAND U3263 ( .A(n2317), .B(n2316), .Z(n2318) );
  NAND U3264 ( .A(n3081), .B(n2318), .Z(n2319) );
  NAND U3265 ( .A(n2320), .B(n2319), .Z(n2321) );
  NAND U3266 ( .A(n3084), .B(n2321), .Z(n2322) );
  NAND U3267 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U3268 ( .A(n3090), .B(n2325), .Z(n2326) );
  NAND U3269 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U3270 ( .A(n2329), .B(n2328), .Z(n2330) );
  NAND U3271 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U3272 ( .A(n3093), .B(n2332), .Z(n2333) );
  NAND U3273 ( .A(n2334), .B(n2333), .Z(n2335) );
  NAND U3274 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U3275 ( .A(n2338), .B(n2337), .Z(n2339) );
  NAND U3276 ( .A(n2340), .B(n2339), .Z(n2341) );
  NAND U3277 ( .A(n2342), .B(n2341), .Z(n2343) );
  NAND U3278 ( .A(n2344), .B(n2343), .Z(n2345) );
  NAND U3279 ( .A(n2346), .B(n2345), .Z(n2347) );
  NAND U3280 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U3281 ( .A(n2350), .B(n2349), .Z(n2351) );
  NAND U3282 ( .A(n3096), .B(n2351), .Z(n2352) );
  NAND U3283 ( .A(n2353), .B(n2352), .Z(n2354) );
  NAND U3284 ( .A(n3099), .B(n2354), .Z(n2355) );
  NAND U3285 ( .A(n2356), .B(n2355), .Z(n2357) );
  NAND U3286 ( .A(n3102), .B(n2357), .Z(n2358) );
  NAND U3287 ( .A(n2359), .B(n2358), .Z(n2360) );
  NAND U3288 ( .A(n3105), .B(n2360), .Z(n2361) );
  NAND U3289 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U3290 ( .A(n3108), .B(n2363), .Z(n2364) );
  NAND U3291 ( .A(n2365), .B(n2364), .Z(n2366) );
  NAND U3292 ( .A(n3111), .B(n2366), .Z(n2367) );
  NAND U3293 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U3294 ( .A(n3114), .B(n2369), .Z(n2370) );
  NAND U3295 ( .A(n2371), .B(n2370), .Z(n2372) );
  NAND U3296 ( .A(n3117), .B(n2372), .Z(n2373) );
  NAND U3297 ( .A(n2374), .B(n2373), .Z(n2375) );
  NAND U3298 ( .A(n3120), .B(n2375), .Z(n2376) );
  NAND U3299 ( .A(n2377), .B(n2376), .Z(n2378) );
  NAND U3300 ( .A(n3123), .B(n2378), .Z(n2379) );
  NAND U3301 ( .A(n2380), .B(n2379), .Z(n2381) );
  NAND U3302 ( .A(n3126), .B(n2381), .Z(n2382) );
  NAND U3303 ( .A(n2383), .B(n2382), .Z(n2384) );
  NAND U3304 ( .A(n3129), .B(n2384), .Z(n2385) );
  NAND U3305 ( .A(n2386), .B(n2385), .Z(n2387) );
  NAND U3306 ( .A(n3132), .B(n2387), .Z(n2388) );
  NAND U3307 ( .A(n2389), .B(n2388), .Z(n2390) );
  NAND U3308 ( .A(n3135), .B(n2390), .Z(n2391) );
  NAND U3309 ( .A(n2392), .B(n2391), .Z(n2393) );
  NAND U3310 ( .A(n3138), .B(n2393), .Z(n2394) );
  NAND U3311 ( .A(n2395), .B(n2394), .Z(n2396) );
  NAND U3312 ( .A(n3141), .B(n2396), .Z(n2397) );
  NAND U3313 ( .A(n2398), .B(n2397), .Z(n2399) );
  NAND U3314 ( .A(n2400), .B(n2399), .Z(n2401) );
  NAND U3315 ( .A(n2402), .B(n2401), .Z(n2403) );
  NAND U3316 ( .A(n3144), .B(n2403), .Z(n2404) );
  NAND U3317 ( .A(n2405), .B(n2404), .Z(n2406) );
  NAND U3318 ( .A(n2407), .B(n2406), .Z(n2408) );
  NAND U3319 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U3320 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U3321 ( .A(n2413), .B(n2412), .Z(n2414) );
  NAND U3322 ( .A(n3147), .B(n2414), .Z(n2415) );
  NAND U3323 ( .A(n2416), .B(n2415), .Z(n2417) );
  NAND U3324 ( .A(n2418), .B(n2417), .Z(n2419) );
  NAND U3325 ( .A(n2420), .B(n2419), .Z(n2421) );
  NAND U3326 ( .A(n3150), .B(n2421), .Z(n2422) );
  NAND U3327 ( .A(n2423), .B(n2422), .Z(n2424) );
  NAND U3328 ( .A(n3153), .B(n2424), .Z(n2425) );
  NAND U3329 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U3330 ( .A(n2428), .B(n2427), .Z(n2429) );
  NAND U3331 ( .A(n2430), .B(n2429), .Z(n2431) );
  NAND U3332 ( .A(n3156), .B(n2431), .Z(n2432) );
  NAND U3333 ( .A(n2433), .B(n2432), .Z(n2434) );
  NAND U3334 ( .A(n2435), .B(n2434), .Z(n2436) );
  NAND U3335 ( .A(n2437), .B(n2436), .Z(n2438) );
  NAND U3336 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U3337 ( .A(n2441), .B(n2440), .Z(n2442) );
  NAND U3338 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U3339 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U3340 ( .A(n2447), .B(n2446), .Z(n2448) );
  NAND U3341 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U3342 ( .A(n2451), .B(n2450), .Z(n2452) );
  NAND U3343 ( .A(n2453), .B(n2452), .Z(n2454) );
  NAND U3344 ( .A(n2455), .B(n2454), .Z(n2456) );
  NAND U3345 ( .A(n2457), .B(n2456), .Z(n2458) );
  NAND U3346 ( .A(n3159), .B(n2458), .Z(n2459) );
  NAND U3347 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U3348 ( .A(n2462), .B(n2461), .Z(n2463) );
  NAND U3349 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U3350 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U3351 ( .A(n2468), .B(n2467), .Z(n2469) );
  NAND U3352 ( .A(n2470), .B(n2469), .Z(n2471) );
  NAND U3353 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U3354 ( .A(n3165), .B(n2473), .Z(n2474) );
  NAND U3355 ( .A(n2475), .B(n2474), .Z(n2476) );
  NAND U3356 ( .A(n3168), .B(n2476), .Z(n2477) );
  NAND U3357 ( .A(n2478), .B(n2477), .Z(n2479) );
  NAND U3358 ( .A(n2480), .B(n2479), .Z(n2481) );
  NAND U3359 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U3360 ( .A(n3171), .B(n2483), .Z(n2484) );
  NAND U3361 ( .A(n2485), .B(n2484), .Z(n2486) );
  NAND U3362 ( .A(n2487), .B(n2486), .Z(n2488) );
  NAND U3363 ( .A(n2489), .B(n2488), .Z(n2490) );
  NAND U3364 ( .A(n2491), .B(n2490), .Z(n2492) );
  NAND U3365 ( .A(n2493), .B(n2492), .Z(n2494) );
  NAND U3366 ( .A(n2495), .B(n2494), .Z(n2496) );
  NAND U3367 ( .A(n2497), .B(n2496), .Z(n2498) );
  NAND U3368 ( .A(n3174), .B(n2498), .Z(n2499) );
  NAND U3369 ( .A(n2500), .B(n2499), .Z(n2501) );
  NAND U3370 ( .A(n2502), .B(n2501), .Z(n2503) );
  NAND U3371 ( .A(n2504), .B(n2503), .Z(n2505) );
  NAND U3372 ( .A(n3177), .B(n2505), .Z(n2506) );
  NAND U3373 ( .A(n2507), .B(n2506), .Z(n2508) );
  NAND U3374 ( .A(n3180), .B(n2508), .Z(n2509) );
  NAND U3375 ( .A(n2510), .B(n2509), .Z(n2511) );
  NAND U3376 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U3377 ( .A(n2514), .B(n2513), .Z(n2515) );
  NAND U3378 ( .A(n3183), .B(n2515), .Z(n2516) );
  NAND U3379 ( .A(n2517), .B(n2516), .Z(n2518) );
  NAND U3380 ( .A(n3186), .B(n2518), .Z(n2519) );
  NAND U3381 ( .A(n2520), .B(n2519), .Z(n2521) );
  NAND U3382 ( .A(n3189), .B(n2521), .Z(n2522) );
  NAND U3383 ( .A(n2523), .B(n2522), .Z(n2524) );
  NAND U3384 ( .A(n2525), .B(n2524), .Z(n2526) );
  NAND U3385 ( .A(n2527), .B(n2526), .Z(n2528) );
  NAND U3386 ( .A(n3192), .B(n2528), .Z(n2529) );
  NAND U3387 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U3388 ( .A(n2532), .B(n2531), .Z(n2533) );
  NAND U3389 ( .A(n2534), .B(n2533), .Z(n2535) );
  NAND U3390 ( .A(n2536), .B(n2535), .Z(n2537) );
  NAND U3391 ( .A(n2538), .B(n2537), .Z(n2539) );
  NAND U3392 ( .A(n2540), .B(n2539), .Z(n2541) );
  NAND U3393 ( .A(n2542), .B(n2541), .Z(n2543) );
  NAND U3394 ( .A(n3195), .B(n2543), .Z(n2544) );
  NAND U3395 ( .A(n2545), .B(n2544), .Z(n2546) );
  NAND U3396 ( .A(n3198), .B(n2546), .Z(n2547) );
  NAND U3397 ( .A(n2548), .B(n2547), .Z(n2549) );
  NAND U3398 ( .A(n3201), .B(n2549), .Z(n2550) );
  NAND U3399 ( .A(n2551), .B(n2550), .Z(n2552) );
  NAND U3400 ( .A(n3204), .B(n2552), .Z(n2553) );
  NAND U3401 ( .A(n2554), .B(n2553), .Z(n2555) );
  NAND U3402 ( .A(n3207), .B(n2555), .Z(n2556) );
  NAND U3403 ( .A(n2557), .B(n2556), .Z(n2558) );
  NAND U3404 ( .A(n2559), .B(n2558), .Z(n2560) );
  NAND U3405 ( .A(n2561), .B(n2560), .Z(n2562) );
  NAND U3406 ( .A(n3210), .B(n2562), .Z(n2563) );
  NAND U3407 ( .A(n2564), .B(n2563), .Z(n2565) );
  NAND U3408 ( .A(n3213), .B(n2565), .Z(n2566) );
  NAND U3409 ( .A(n2567), .B(n2566), .Z(n2568) );
  NAND U3410 ( .A(n3216), .B(n2568), .Z(n2569) );
  NAND U3411 ( .A(n2570), .B(n2569), .Z(n2571) );
  NAND U3412 ( .A(n3219), .B(n2571), .Z(n2572) );
  NAND U3413 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U3414 ( .A(n2575), .B(n2574), .Z(n2576) );
  NAND U3415 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U3416 ( .A(n3222), .B(n2578), .Z(n2579) );
  NAND U3417 ( .A(n2580), .B(n2579), .Z(n2581) );
  NAND U3418 ( .A(n2582), .B(n2581), .Z(n2583) );
  NAND U3419 ( .A(n2584), .B(n2583), .Z(n2585) );
  NAND U3420 ( .A(n3225), .B(n2585), .Z(n2586) );
  NAND U3421 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U3422 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U3423 ( .A(n2591), .B(n2590), .Z(n2592) );
  NAND U3424 ( .A(n2593), .B(n2592), .Z(n2594) );
  NAND U3425 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U3426 ( .A(n2597), .B(n2596), .Z(n2598) );
  NAND U3427 ( .A(n2599), .B(n2598), .Z(n2600) );
  NAND U3428 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U3429 ( .A(n2603), .B(n2602), .Z(n2604) );
  NAND U3430 ( .A(n2605), .B(n2604), .Z(n2606) );
  NAND U3431 ( .A(n2607), .B(n2606), .Z(n2608) );
  NAND U3432 ( .A(n3228), .B(n2608), .Z(n2609) );
  NAND U3433 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U3434 ( .A(n3231), .B(n2611), .Z(n2612) );
  NAND U3435 ( .A(n2613), .B(n2612), .Z(n2614) );
  NAND U3436 ( .A(n2615), .B(n2614), .Z(n2616) );
  NAND U3437 ( .A(n2617), .B(n2616), .Z(n2618) );
  NAND U3438 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U3439 ( .A(n2621), .B(n2620), .Z(n2622) );
  NAND U3440 ( .A(n3234), .B(n2622), .Z(n2623) );
  NAND U3441 ( .A(n2624), .B(n2623), .Z(n2625) );
  NAND U3442 ( .A(n3237), .B(n2625), .Z(n2626) );
  NAND U3443 ( .A(n2627), .B(n2626), .Z(n2628) );
  NAND U3444 ( .A(n2629), .B(n2628), .Z(n2630) );
  NAND U3445 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U3446 ( .A(n3240), .B(n2632), .Z(n2633) );
  NAND U3447 ( .A(n2634), .B(n2633), .Z(n2635) );
  NAND U3448 ( .A(n3243), .B(n2635), .Z(n2636) );
  NAND U3449 ( .A(n2637), .B(n2636), .Z(n2638) );
  NAND U3450 ( .A(n2639), .B(n2638), .Z(n2640) );
  NAND U3451 ( .A(n2641), .B(n2640), .Z(n2642) );
  NAND U3452 ( .A(n2643), .B(n2642), .Z(n2644) );
  NAND U3453 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U3454 ( .A(n2647), .B(n2646), .Z(n2648) );
  NAND U3455 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U3456 ( .A(n3246), .B(n2650), .Z(n2651) );
  NAND U3457 ( .A(n2652), .B(n2651), .Z(n2653) );
  NAND U3458 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U3459 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U3460 ( .A(n2658), .B(n2657), .Z(n2659) );
  NAND U3461 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U3462 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U3463 ( .A(n2664), .B(n2663), .Z(n2665) );
  NAND U3464 ( .A(n2666), .B(n2665), .Z(n2667) );
  NAND U3465 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U3466 ( .A(n3249), .B(n2669), .Z(n2670) );
  NAND U3467 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND U3468 ( .A(n3252), .B(n2672), .Z(n2673) );
  NAND U3469 ( .A(n2674), .B(n2673), .Z(n2675) );
  NAND U3470 ( .A(n2676), .B(n2675), .Z(n2677) );
  NAND U3471 ( .A(n2678), .B(n2677), .Z(n2679) );
  NAND U3472 ( .A(n3255), .B(n2679), .Z(n2680) );
  NAND U3473 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U3474 ( .A(n2683), .B(n2682), .Z(n2684) );
  NAND U3475 ( .A(n2685), .B(n2684), .Z(n2686) );
  NAND U3476 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U3477 ( .A(n2689), .B(n2688), .Z(n2690) );
  NAND U3478 ( .A(n3258), .B(n2690), .Z(n2691) );
  NAND U3479 ( .A(n2692), .B(n2691), .Z(n2693) );
  NAND U3480 ( .A(n2694), .B(n2693), .Z(n2695) );
  NAND U3481 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U3482 ( .A(n3261), .B(n2697), .Z(n2698) );
  NAND U3483 ( .A(n2699), .B(n2698), .Z(n2700) );
  NAND U3484 ( .A(n2701), .B(n2700), .Z(n2702) );
  NAND U3485 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U3486 ( .A(n2705), .B(n2704), .Z(n2706) );
  NAND U3487 ( .A(n2707), .B(n2706), .Z(n2708) );
  NAND U3488 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U3489 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U3490 ( .A(n2713), .B(n2712), .Z(n2714) );
  NAND U3491 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U3492 ( .A(n3264), .B(n2716), .Z(n2717) );
  NAND U3493 ( .A(n2718), .B(n2717), .Z(n2719) );
  NAND U3494 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U3495 ( .A(n2722), .B(n2721), .Z(n2723) );
  NAND U3496 ( .A(n2724), .B(n2723), .Z(n2725) );
  NAND U3497 ( .A(n2726), .B(n2725), .Z(n2727) );
  NAND U3498 ( .A(n2728), .B(n2727), .Z(n2729) );
  NAND U3499 ( .A(n2730), .B(n2729), .Z(n2731) );
  NAND U3500 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U3501 ( .A(n2734), .B(n2733), .Z(n2735) );
  NAND U3502 ( .A(n3267), .B(n2735), .Z(n2736) );
  NAND U3503 ( .A(n2737), .B(n2736), .Z(n2738) );
  NAND U3504 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND U3505 ( .A(n2741), .B(n2740), .Z(n2742) );
  NAND U3506 ( .A(n2743), .B(n2742), .Z(n2744) );
  NAND U3507 ( .A(n2745), .B(n2744), .Z(n2746) );
  NAND U3508 ( .A(n2747), .B(n2746), .Z(n2748) );
  NAND U3509 ( .A(n2749), .B(n2748), .Z(n2750) );
  NAND U3510 ( .A(n3270), .B(n2750), .Z(n2751) );
  NAND U3511 ( .A(n2752), .B(n2751), .Z(n2753) );
  NAND U3512 ( .A(n2754), .B(n2753), .Z(n2755) );
  NAND U3513 ( .A(n2756), .B(n2755), .Z(n2757) );
  NAND U3514 ( .A(n2758), .B(n2757), .Z(n2759) );
  NAND U3515 ( .A(n2760), .B(n2759), .Z(n2761) );
  NAND U3516 ( .A(n3273), .B(n2761), .Z(n2762) );
  NAND U3517 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U3518 ( .A(n2765), .B(n2764), .Z(n2766) );
  NAND U3519 ( .A(n2767), .B(n2766), .Z(n2768) );
  NAND U3520 ( .A(n2769), .B(n2768), .Z(n2770) );
  NAND U3521 ( .A(n2771), .B(n2770), .Z(n2772) );
  NAND U3522 ( .A(n2773), .B(n2772), .Z(n2774) );
  NAND U3523 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3524 ( .A(n2777), .B(n2776), .Z(n2778) );
  NAND U3525 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U3526 ( .A(n2781), .B(n2780), .Z(n2782) );
  NAND U3527 ( .A(n2783), .B(n2782), .Z(n2784) );
  NAND U3528 ( .A(n3279), .B(n2784), .Z(n2785) );
  NAND U3529 ( .A(n2786), .B(n2785), .Z(n2787) );
  NAND U3530 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U3531 ( .A(n2790), .B(n2789), .Z(n2791) );
  NAND U3532 ( .A(n2792), .B(n2791), .Z(n2793) );
  NAND U3533 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U3534 ( .A(n2796), .B(n2795), .Z(n2797) );
  NAND U3535 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U3536 ( .A(n2800), .B(n2799), .Z(n2801) );
  NAND U3537 ( .A(n2802), .B(n2801), .Z(n2803) );
  NAND U3538 ( .A(n2804), .B(n2803), .Z(n2805) );
  NAND U3539 ( .A(n2806), .B(n2805), .Z(n2807) );
  NAND U3540 ( .A(n2808), .B(n2807), .Z(n2809) );
  NAND U3541 ( .A(n2810), .B(n2809), .Z(n2811) );
  NAND U3542 ( .A(n2812), .B(n2811), .Z(n2813) );
  NAND U3543 ( .A(n2814), .B(n2813), .Z(n2815) );
  NAND U3544 ( .A(n3282), .B(n2815), .Z(n2816) );
  NAND U3545 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U3546 ( .A(n2819), .B(n2818), .Z(n2820) );
  NAND U3547 ( .A(n2821), .B(n2820), .Z(n2822) );
  NAND U3548 ( .A(n2823), .B(n2822), .Z(n2824) );
  NAND U3549 ( .A(n2825), .B(n2824), .Z(n2826) );
  NAND U3550 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U3551 ( .A(n2829), .B(n2828), .Z(n2830) );
  NAND U3552 ( .A(n2831), .B(n2830), .Z(n2832) );
  NAND U3553 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U3554 ( .A(n3285), .B(n2834), .Z(n2835) );
  NAND U3555 ( .A(n2836), .B(n2835), .Z(n2837) );
  NAND U3556 ( .A(n3288), .B(n2837), .Z(n2838) );
  NAND U3557 ( .A(n2839), .B(n2838), .Z(n2840) );
  NAND U3558 ( .A(n3291), .B(n2840), .Z(n2841) );
  NAND U3559 ( .A(n2842), .B(n2841), .Z(n2843) );
  NAND U3560 ( .A(n3294), .B(n2843), .Z(n2844) );
  NAND U3561 ( .A(n2845), .B(n2844), .Z(n2846) );
  NAND U3562 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U3563 ( .A(n2849), .B(n2848), .Z(n2850) );
  NAND U3564 ( .A(n3297), .B(n2850), .Z(n2851) );
  NAND U3565 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3566 ( .A(n2854), .B(n2853), .Z(n2855) );
  NAND U3567 ( .A(y[254]), .B(zin[253]), .Z(n2860) );
  XOR U3568 ( .A(zin[253]), .B(y[254]), .Z(n2858) );
  NAND U3569 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U3570 ( .A(n2860), .B(n2859), .Z(n2864) );
  XOR U3571 ( .A(y[255]), .B(n2864), .Z(n2861) );
  ANDN U3572 ( .B(n2861), .A(n2868), .Z(n2862) );
  XNOR U3573 ( .A(zin[254]), .B(n2862), .Z(n3308) );
  AND U3574 ( .A(y[255]), .B(zin[254]), .Z(n2866) );
  XOR U3575 ( .A(zin[254]), .B(y[255]), .Z(n2863) );
  AND U3576 ( .A(n2864), .B(n2863), .Z(n2865) );
  OR U3577 ( .A(n2866), .B(n2865), .Z(n2867) );
  NANDN U3578 ( .A(n2868), .B(n2867), .Z(n2870) );
  ANDN U3579 ( .B(zin[255]), .A(n2870), .Z(n2869) );
  XOR U3580 ( .A(n2869), .B(zin[256]), .Z(n3313) );
  XNOR U3581 ( .A(n2870), .B(zin[255]), .Z(n3312) );
  NANDN U3582 ( .A(n524), .B(n[0]), .Z(n2871) );
  XNOR U3583 ( .A(n2880), .B(n2871), .Z(n5342) );
  NOR U3584 ( .A(n[254]), .B(n3318), .Z(n3301) );
  NOR U3585 ( .A(n[252]), .B(n3326), .Z(n3298) );
  NOR U3586 ( .A(n[249]), .B(n3339), .Z(n3295) );
  NOR U3587 ( .A(n[247]), .B(n3347), .Z(n3292) );
  NOR U3588 ( .A(n[246]), .B(n3352), .Z(n3289) );
  NOR U3589 ( .A(n[245]), .B(n3356), .Z(n3286) );
  NOR U3590 ( .A(n[244]), .B(n3360), .Z(n3283) );
  NOR U3591 ( .A(n[239]), .B(n3381), .Z(n3280) );
  NOR U3592 ( .A(n[231]), .B(n3411), .Z(n3277) );
  IV U3593 ( .A(n2873), .Z(n3419) );
  OR U3594 ( .A(n[228]), .B(n3419), .Z(n3276) );
  ANDN U3595 ( .B(n[228]), .A(n2873), .Z(n3274) );
  NOR U3596 ( .A(n[225]), .B(n3431), .Z(n3271) );
  NOR U3597 ( .A(n[222]), .B(n3443), .Z(n3268) );
  NOR U3598 ( .A(n[218]), .B(n3459), .Z(n3265) );
  NOR U3599 ( .A(n[213]), .B(n3475), .Z(n3262) );
  NOR U3600 ( .A(n[208]), .B(n3498), .Z(n3259) );
  NOR U3601 ( .A(n[206]), .B(n3507), .Z(n3256) );
  NOR U3602 ( .A(n[203]), .B(n3520), .Z(n3253) );
  NOR U3603 ( .A(n[201]), .B(n3528), .Z(n3250) );
  NOR U3604 ( .A(n[200]), .B(n3533), .Z(n3247) );
  NOR U3605 ( .A(n[195]), .B(n3554), .Z(n3244) );
  NOR U3606 ( .A(n[191]), .B(n3572), .Z(n3241) );
  NOR U3607 ( .A(n[190]), .B(n3576), .Z(n3238) );
  NOR U3608 ( .A(n[188]), .B(n3585), .Z(n3235) );
  NOR U3609 ( .A(n[187]), .B(n3590), .Z(n3232) );
  NOR U3610 ( .A(n[184]), .B(n3598), .Z(n3229) );
  NOR U3611 ( .A(n[183]), .B(n3602), .Z(n3226) );
  NOR U3612 ( .A(n[177]), .B(n3623), .Z(n3223) );
  NOR U3613 ( .A(n[175]), .B(n3632), .Z(n3220) );
  NOR U3614 ( .A(n[173]), .B(n3640), .Z(n3217) );
  NOR U3615 ( .A(n[172]), .B(n3645), .Z(n3214) );
  NOR U3616 ( .A(n[171]), .B(n3650), .Z(n3211) );
  NOR U3617 ( .A(n[170]), .B(n3654), .Z(n3208) );
  NOR U3618 ( .A(n[168]), .B(n3663), .Z(n3205) );
  NOR U3619 ( .A(n[167]), .B(n3668), .Z(n3202) );
  NOR U3620 ( .A(n[166]), .B(n3672), .Z(n3199) );
  NOR U3621 ( .A(n[165]), .B(n3677), .Z(n3196) );
  NOR U3622 ( .A(n[164]), .B(n3681), .Z(n3193) );
  NOR U3623 ( .A(n[160]), .B(n3697), .Z(n3190) );
  NOR U3624 ( .A(n[158]), .B(n3706), .Z(n3187) );
  NOR U3625 ( .A(n[157]), .B(n4937), .Z(n3184) );
  NOR U3626 ( .A(n[156]), .B(n3710), .Z(n3181) );
  NOR U3627 ( .A(n[154]), .B(n3714), .Z(n3178) );
  NOR U3628 ( .A(n[153]), .B(n4913), .Z(n3175) );
  NOR U3629 ( .A(n[151]), .B(n3722), .Z(n3172) );
  NOR U3630 ( .A(n[147]), .B(n3738), .Z(n3169) );
  NOR U3631 ( .A(n[145]), .B(n3747), .Z(n3166) );
  NOR U3632 ( .A(n[144]), .B(n3751), .Z(n3163) );
  IV U3633 ( .A(n2876), .Z(n3760) );
  OR U3634 ( .A(n[142]), .B(n3760), .Z(n3162) );
  ANDN U3635 ( .B(n[142]), .A(n2876), .Z(n3160) );
  NOR U3636 ( .A(n[140]), .B(n3768), .Z(n3157) );
  NOR U3637 ( .A(n[133]), .B(n3797), .Z(n3154) );
  NOR U3638 ( .A(n[131]), .B(n3806), .Z(n3151) );
  NOR U3639 ( .A(n[130]), .B(n3810), .Z(n3148) );
  NOR U3640 ( .A(n[128]), .B(n3819), .Z(n3145) );
  NOR U3641 ( .A(n[125]), .B(n3831), .Z(n3142) );
  NOR U3642 ( .A(n[123]), .B(n3840), .Z(n3139) );
  NOR U3643 ( .A(n[122]), .B(n3845), .Z(n3136) );
  NOR U3644 ( .A(n[121]), .B(n3850), .Z(n3133) );
  NOR U3645 ( .A(n[120]), .B(n3855), .Z(n3130) );
  NOR U3646 ( .A(n[119]), .B(n3860), .Z(n3127) );
  NOR U3647 ( .A(n[118]), .B(n3864), .Z(n3124) );
  NOR U3648 ( .A(n[117]), .B(n3868), .Z(n3121) );
  NOR U3649 ( .A(n[116]), .B(n3873), .Z(n3118) );
  NOR U3650 ( .A(n[115]), .B(n3877), .Z(n3115) );
  NOR U3651 ( .A(n[114]), .B(n3882), .Z(n3112) );
  NOR U3652 ( .A(n[113]), .B(n3887), .Z(n3109) );
  NOR U3653 ( .A(n[112]), .B(n3892), .Z(n3106) );
  NOR U3654 ( .A(n[111]), .B(n3897), .Z(n3103) );
  NOR U3655 ( .A(n[110]), .B(n3902), .Z(n3100) );
  NOR U3656 ( .A(n[109]), .B(n3907), .Z(n3097) );
  NOR U3657 ( .A(n[108]), .B(n3911), .Z(n3094) );
  NOR U3658 ( .A(n[103]), .B(n3932), .Z(n3091) );
  NOR U3659 ( .A(n[101]), .B(n3941), .Z(n3088) );
  NOR U3660 ( .A(n[96]), .B(n3962), .Z(n3085) );
  NOR U3661 ( .A(n[95]), .B(n3967), .Z(n3082) );
  NOR U3662 ( .A(n[94]), .B(n3972), .Z(n3079) );
  NOR U3663 ( .A(n[93]), .B(n3977), .Z(n3076) );
  NOR U3664 ( .A(n[92]), .B(n4663), .Z(n3073) );
  NOR U3665 ( .A(n[91]), .B(n3981), .Z(n3070) );
  NOR U3666 ( .A(n[89]), .B(n3989), .Z(n3067) );
  NOR U3667 ( .A(n[87]), .B(n3997), .Z(n3064) );
  NOR U3668 ( .A(n[85]), .B(n4006), .Z(n3061) );
  NOR U3669 ( .A(n[81]), .B(n4022), .Z(n3058) );
  NOR U3670 ( .A(n[80]), .B(n4027), .Z(n3055) );
  NOR U3671 ( .A(n[77]), .B(n4040), .Z(n3052) );
  IV U3672 ( .A(n2877), .Z(n4053) );
  OR U3673 ( .A(n[74]), .B(n4053), .Z(n3051) );
  ANDN U3674 ( .B(n[74]), .A(n2877), .Z(n3049) );
  IV U3675 ( .A(n2878), .Z(n4061) );
  OR U3676 ( .A(n[72]), .B(n4061), .Z(n3048) );
  ANDN U3677 ( .B(n[72]), .A(n2878), .Z(n3046) );
  NOR U3678 ( .A(n[70]), .B(n4069), .Z(n3043) );
  NANDN U3679 ( .A(n4113), .B(n4112), .Z(n3027) );
  NOR U3680 ( .A(n[60]), .B(n4112), .Z(n3025) );
  NANDN U3681 ( .A(n4446), .B(n4192), .Z(n2973) );
  NOR U3682 ( .A(n[39]), .B(n4192), .Z(n2971) );
  NOR U3683 ( .A(n[31]), .B(n4419), .Z(n2959) );
  NOR U3684 ( .A(n[30]), .B(n4221), .Z(n2956) );
  NOR U3685 ( .A(n[29]), .B(n4226), .Z(n2953) );
  NOR U3686 ( .A(n[28]), .B(n4406), .Z(n2950) );
  NOR U3687 ( .A(n[24]), .B(n4238), .Z(n2947) );
  NOR U3688 ( .A(n[23]), .B(n4390), .Z(n2944) );
  NOR U3689 ( .A(n[22]), .B(n4243), .Z(n2941) );
  NOR U3690 ( .A(n[21]), .B(n4381), .Z(n2938) );
  NOR U3691 ( .A(n[20]), .B(n4247), .Z(n2935) );
  NOR U3692 ( .A(n[19]), .B(n4252), .Z(n2932) );
  NOR U3693 ( .A(n[18]), .B(n4256), .Z(n2929) );
  NANDN U3694 ( .A(n6868), .B(n4329), .Z(n2904) );
  ANDN U3695 ( .B(n[0]), .A(n2880), .Z(n4296) );
  NANDN U3696 ( .A(n6616), .B(n4300), .Z(n2883) );
  NOR U3697 ( .A(n[2]), .B(n4300), .Z(n2881) );
  NANDN U3698 ( .A(n2881), .B(n4303), .Z(n2882) );
  NAND U3699 ( .A(n2883), .B(n2882), .Z(n4304) );
  NAND U3700 ( .A(n4304), .B(n2884), .Z(n2885) );
  NAND U3701 ( .A(n2886), .B(n2885), .Z(n4292) );
  NAND U3702 ( .A(n4292), .B(n2887), .Z(n2888) );
  NAND U3703 ( .A(n2889), .B(n2888), .Z(n4288) );
  NAND U3704 ( .A(n4288), .B(n2890), .Z(n2891) );
  NAND U3705 ( .A(n2892), .B(n2891), .Z(n4284) );
  NAND U3706 ( .A(n4284), .B(n2893), .Z(n2894) );
  NAND U3707 ( .A(n2895), .B(n2894), .Z(n4280) );
  OR U3708 ( .A(n2896), .B(n4280), .Z(n2898) );
  AND U3709 ( .A(n2898), .B(n2897), .Z(n4276) );
  OR U3710 ( .A(n4276), .B(n2899), .Z(n2901) );
  NAND U3711 ( .A(n2901), .B(n2900), .Z(n4326) );
  NOR U3712 ( .A(n[9]), .B(n4329), .Z(n2902) );
  OR U3713 ( .A(n4326), .B(n2902), .Z(n2903) );
  NAND U3714 ( .A(n2904), .B(n2903), .Z(n4330) );
  NANDN U3715 ( .A(n2905), .B(n4330), .Z(n2906) );
  NANDN U3716 ( .A(n2907), .B(n2906), .Z(n4338) );
  NANDN U3717 ( .A(n2908), .B(n4338), .Z(n2909) );
  NANDN U3718 ( .A(n2910), .B(n2909), .Z(n4345) );
  NANDN U3719 ( .A(n2911), .B(n4345), .Z(n2912) );
  NANDN U3720 ( .A(n2913), .B(n2912), .Z(n4272) );
  NANDN U3721 ( .A(n2914), .B(n4272), .Z(n2915) );
  NANDN U3722 ( .A(n2916), .B(n2915), .Z(n4267) );
  NANDN U3723 ( .A(n2917), .B(n4267), .Z(n2918) );
  NANDN U3724 ( .A(n2919), .B(n2918), .Z(n4357) );
  NANDN U3725 ( .A(n2920), .B(n4357), .Z(n2921) );
  NANDN U3726 ( .A(n2922), .B(n2921), .Z(n4262) );
  NANDN U3727 ( .A(n2923), .B(n4262), .Z(n2924) );
  NANDN U3728 ( .A(n2925), .B(n2924), .Z(n4258) );
  NANDN U3729 ( .A(n2926), .B(n4258), .Z(n2927) );
  NANDN U3730 ( .A(n2928), .B(n2927), .Z(n4253) );
  NANDN U3731 ( .A(n2929), .B(n4253), .Z(n2930) );
  NAND U3732 ( .A(n2931), .B(n2930), .Z(n4249) );
  NANDN U3733 ( .A(n2932), .B(n4249), .Z(n2933) );
  NAND U3734 ( .A(n2934), .B(n2933), .Z(n4244) );
  NANDN U3735 ( .A(n2935), .B(n4244), .Z(n2936) );
  NAND U3736 ( .A(n2937), .B(n2936), .Z(n4378) );
  NANDN U3737 ( .A(n2938), .B(n4378), .Z(n2939) );
  NAND U3738 ( .A(n2940), .B(n2939), .Z(n4240) );
  NANDN U3739 ( .A(n2941), .B(n4240), .Z(n2942) );
  NAND U3740 ( .A(n2943), .B(n2942), .Z(n4386) );
  NANDN U3741 ( .A(n2944), .B(n4386), .Z(n2945) );
  NAND U3742 ( .A(n2946), .B(n2945), .Z(n4235) );
  NANDN U3743 ( .A(n2947), .B(n4235), .Z(n2948) );
  NAND U3744 ( .A(n2949), .B(n2948), .Z(n4231) );
  OR U3745 ( .A(n2950), .B(n4403), .Z(n2951) );
  NAND U3746 ( .A(n2952), .B(n2951), .Z(n4223) );
  NANDN U3747 ( .A(n2953), .B(n4223), .Z(n2954) );
  NAND U3748 ( .A(n2955), .B(n2954), .Z(n4218) );
  NANDN U3749 ( .A(n2956), .B(n4218), .Z(n2957) );
  NAND U3750 ( .A(n2958), .B(n2957), .Z(n4415) );
  NANDN U3751 ( .A(n2959), .B(n4415), .Z(n2960) );
  NAND U3752 ( .A(n2961), .B(n2960), .Z(n4214) );
  NANDN U3753 ( .A(n2962), .B(n4202), .Z(n2963) );
  NANDN U3754 ( .A(n2964), .B(n2963), .Z(n4198) );
  NANDN U3755 ( .A(n2965), .B(n4198), .Z(n2966) );
  NANDN U3756 ( .A(n2967), .B(n2966), .Z(n4193) );
  NANDN U3757 ( .A(n2968), .B(n4193), .Z(n2969) );
  NANDN U3758 ( .A(n2970), .B(n2969), .Z(n4189) );
  OR U3759 ( .A(n2971), .B(n4189), .Z(n2972) );
  NAND U3760 ( .A(n2973), .B(n2972), .Z(n4184) );
  OR U3761 ( .A(n2974), .B(n4184), .Z(n2975) );
  NANDN U3762 ( .A(n2976), .B(n2975), .Z(n4180) );
  NANDN U3763 ( .A(n4180), .B(n2977), .Z(n2978) );
  NANDN U3764 ( .A(n2979), .B(n2978), .Z(n4175) );
  NANDN U3765 ( .A(n2980), .B(n4175), .Z(n2981) );
  NANDN U3766 ( .A(n2982), .B(n2981), .Z(n4462) );
  NANDN U3767 ( .A(n2983), .B(n4462), .Z(n2984) );
  NANDN U3768 ( .A(n2985), .B(n2984), .Z(n4467) );
  OR U3769 ( .A(n2986), .B(n4467), .Z(n2987) );
  NANDN U3770 ( .A(n2988), .B(n2987), .Z(n4471) );
  NANDN U3771 ( .A(n2989), .B(n4171), .Z(n2990) );
  NANDN U3772 ( .A(n2991), .B(n2990), .Z(n4167) );
  NANDN U3773 ( .A(n2992), .B(n4167), .Z(n2993) );
  NAND U3774 ( .A(n2994), .B(n2993), .Z(n4163) );
  NANDN U3775 ( .A(n4163), .B(n2995), .Z(n2996) );
  NANDN U3776 ( .A(n2997), .B(n2996), .Z(n4158) );
  NANDN U3777 ( .A(n2998), .B(n4158), .Z(n2999) );
  NANDN U3778 ( .A(n3000), .B(n2999), .Z(n4154) );
  NANDN U3779 ( .A(n3001), .B(n4154), .Z(n3002) );
  NANDN U3780 ( .A(n3003), .B(n3002), .Z(n4150) );
  NANDN U3781 ( .A(n4146), .B(n3004), .Z(n3005) );
  NANDN U3782 ( .A(n3006), .B(n3005), .Z(n4141) );
  NANDN U3783 ( .A(n3007), .B(n4141), .Z(n3008) );
  NANDN U3784 ( .A(n3009), .B(n3008), .Z(n4136) );
  OR U3785 ( .A(n3010), .B(n4136), .Z(n3011) );
  NANDN U3786 ( .A(n3012), .B(n3011), .Z(n4132) );
  NANDN U3787 ( .A(n3013), .B(n4132), .Z(n3014) );
  NANDN U3788 ( .A(n3015), .B(n3014), .Z(n4127) );
  NANDN U3789 ( .A(n3016), .B(n4127), .Z(n3017) );
  NANDN U3790 ( .A(n3018), .B(n3017), .Z(n4123) );
  NANDN U3791 ( .A(n3019), .B(n4119), .Z(n3020) );
  NANDN U3792 ( .A(n3021), .B(n3020), .Z(n4114) );
  NANDN U3793 ( .A(n3022), .B(n4114), .Z(n3023) );
  NANDN U3794 ( .A(n3024), .B(n3023), .Z(n4109) );
  NANDN U3795 ( .A(n3025), .B(n4109), .Z(n3026) );
  NAND U3796 ( .A(n3027), .B(n3026), .Z(n4104) );
  OR U3797 ( .A(n3028), .B(n4104), .Z(n3029) );
  NANDN U3798 ( .A(n3030), .B(n3029), .Z(n4100) );
  NANDN U3799 ( .A(n4100), .B(n3031), .Z(n3032) );
  NANDN U3800 ( .A(n3033), .B(n3032), .Z(n4096) );
  NANDN U3801 ( .A(n3034), .B(n4092), .Z(n3035) );
  NANDN U3802 ( .A(n3036), .B(n3035), .Z(n4087) );
  NANDN U3803 ( .A(n3037), .B(n4087), .Z(n3039) );
  ANDN U3804 ( .B(n3039), .A(n3038), .Z(n4083) );
  NANDN U3805 ( .A(n3040), .B(n4074), .Z(n3041) );
  NANDN U3806 ( .A(n3042), .B(n3041), .Z(n4070) );
  OR U3807 ( .A(n3043), .B(n4066), .Z(n3044) );
  NAND U3808 ( .A(n3045), .B(n3044), .Z(n4062) );
  NANDN U3809 ( .A(n3046), .B(n4058), .Z(n3047) );
  NAND U3810 ( .A(n3048), .B(n3047), .Z(n4054) );
  NANDN U3811 ( .A(n3049), .B(n4050), .Z(n3050) );
  NAND U3812 ( .A(n3051), .B(n3050), .Z(n4046) );
  OR U3813 ( .A(n3052), .B(n4037), .Z(n3053) );
  NAND U3814 ( .A(n3054), .B(n3053), .Z(n4033) );
  OR U3815 ( .A(n3055), .B(n4024), .Z(n3056) );
  NAND U3816 ( .A(n3057), .B(n3056), .Z(n4019) );
  NANDN U3817 ( .A(n3058), .B(n4019), .Z(n3059) );
  NAND U3818 ( .A(n3060), .B(n3059), .Z(n4015) );
  OR U3819 ( .A(n3061), .B(n4003), .Z(n3062) );
  NAND U3820 ( .A(n3063), .B(n3062), .Z(n3999) );
  OR U3821 ( .A(n3064), .B(n3994), .Z(n3065) );
  NAND U3822 ( .A(n3066), .B(n3065), .Z(n3990) );
  OR U3823 ( .A(n3067), .B(n3986), .Z(n3068) );
  NAND U3824 ( .A(n3069), .B(n3068), .Z(n3982) );
  OR U3825 ( .A(n3070), .B(n3978), .Z(n3071) );
  NAND U3826 ( .A(n3072), .B(n3071), .Z(n4660) );
  NANDN U3827 ( .A(n3073), .B(n4660), .Z(n3074) );
  NAND U3828 ( .A(n3075), .B(n3074), .Z(n3973) );
  NANDN U3829 ( .A(n3076), .B(n3973), .Z(n3077) );
  NAND U3830 ( .A(n3078), .B(n3077), .Z(n3968) );
  NANDN U3831 ( .A(n3079), .B(n3968), .Z(n3080) );
  NAND U3832 ( .A(n3081), .B(n3080), .Z(n3964) );
  NANDN U3833 ( .A(n3082), .B(n3964), .Z(n3083) );
  NAND U3834 ( .A(n3084), .B(n3083), .Z(n3959) );
  NANDN U3835 ( .A(n3085), .B(n3959), .Z(n3086) );
  NAND U3836 ( .A(n3087), .B(n3086), .Z(n3955) );
  OR U3837 ( .A(n3088), .B(n3938), .Z(n3089) );
  NAND U3838 ( .A(n3090), .B(n3089), .Z(n3934) );
  OR U3839 ( .A(n3091), .B(n3929), .Z(n3092) );
  NAND U3840 ( .A(n3093), .B(n3092), .Z(n3925) );
  OR U3841 ( .A(n3094), .B(n3908), .Z(n3095) );
  NAND U3842 ( .A(n3096), .B(n3095), .Z(n3904) );
  NANDN U3843 ( .A(n3097), .B(n3904), .Z(n3098) );
  NAND U3844 ( .A(n3099), .B(n3098), .Z(n3899) );
  NANDN U3845 ( .A(n3100), .B(n3899), .Z(n3101) );
  NAND U3846 ( .A(n3102), .B(n3101), .Z(n3894) );
  NANDN U3847 ( .A(n3103), .B(n3894), .Z(n3104) );
  NAND U3848 ( .A(n3105), .B(n3104), .Z(n3889) );
  NANDN U3849 ( .A(n3106), .B(n3889), .Z(n3107) );
  NAND U3850 ( .A(n3108), .B(n3107), .Z(n3884) );
  NANDN U3851 ( .A(n3109), .B(n3884), .Z(n3110) );
  NAND U3852 ( .A(n3111), .B(n3110), .Z(n3879) );
  NANDN U3853 ( .A(n3112), .B(n3879), .Z(n3113) );
  NAND U3854 ( .A(n3114), .B(n3113), .Z(n3874) );
  NANDN U3855 ( .A(n3115), .B(n3874), .Z(n3116) );
  NAND U3856 ( .A(n3117), .B(n3116), .Z(n3870) );
  NANDN U3857 ( .A(n3118), .B(n3870), .Z(n3119) );
  NAND U3858 ( .A(n3120), .B(n3119), .Z(n3865) );
  NANDN U3859 ( .A(n3121), .B(n3865), .Z(n3122) );
  NAND U3860 ( .A(n3123), .B(n3122), .Z(n3861) );
  NANDN U3861 ( .A(n3124), .B(n3861), .Z(n3125) );
  NAND U3862 ( .A(n3126), .B(n3125), .Z(n3857) );
  NANDN U3863 ( .A(n3127), .B(n3857), .Z(n3128) );
  NAND U3864 ( .A(n3129), .B(n3128), .Z(n3852) );
  NANDN U3865 ( .A(n3130), .B(n3852), .Z(n3131) );
  NAND U3866 ( .A(n3132), .B(n3131), .Z(n3847) );
  NANDN U3867 ( .A(n3133), .B(n3847), .Z(n3134) );
  NAND U3868 ( .A(n3135), .B(n3134), .Z(n3842) );
  NANDN U3869 ( .A(n3136), .B(n3842), .Z(n3137) );
  NAND U3870 ( .A(n3138), .B(n3137), .Z(n3837) );
  NANDN U3871 ( .A(n3139), .B(n3837), .Z(n3140) );
  NAND U3872 ( .A(n3141), .B(n3140), .Z(n3833) );
  OR U3873 ( .A(n3142), .B(n3828), .Z(n3143) );
  NAND U3874 ( .A(n3144), .B(n3143), .Z(n3824) );
  OR U3875 ( .A(n3145), .B(n3816), .Z(n3146) );
  NAND U3876 ( .A(n3147), .B(n3146), .Z(n3812) );
  OR U3877 ( .A(n3148), .B(n3807), .Z(n3149) );
  NAND U3878 ( .A(n3150), .B(n3149), .Z(n3803) );
  NANDN U3879 ( .A(n3151), .B(n3803), .Z(n3152) );
  NAND U3880 ( .A(n3153), .B(n3152), .Z(n3799) );
  OR U3881 ( .A(n3154), .B(n3794), .Z(n3155) );
  NAND U3882 ( .A(n3156), .B(n3155), .Z(n3790) );
  OR U3883 ( .A(n3157), .B(n3765), .Z(n3158) );
  NAND U3884 ( .A(n3159), .B(n3158), .Z(n3761) );
  NANDN U3885 ( .A(n3160), .B(n3757), .Z(n3161) );
  NAND U3886 ( .A(n3162), .B(n3161), .Z(n3753) );
  OR U3887 ( .A(n3163), .B(n3748), .Z(n3164) );
  NAND U3888 ( .A(n3165), .B(n3164), .Z(n3744) );
  NANDN U3889 ( .A(n3166), .B(n3744), .Z(n3167) );
  NAND U3890 ( .A(n3168), .B(n3167), .Z(n3740) );
  OR U3891 ( .A(n3169), .B(n3735), .Z(n3170) );
  NAND U3892 ( .A(n3171), .B(n3170), .Z(n3731) );
  OR U3893 ( .A(n3172), .B(n3719), .Z(n3173) );
  NAND U3894 ( .A(n3174), .B(n3173), .Z(n3715) );
  OR U3895 ( .A(n3175), .B(n4909), .Z(n3176) );
  NAND U3896 ( .A(n3177), .B(n3176), .Z(n3711) );
  NANDN U3897 ( .A(n3178), .B(n3711), .Z(n3179) );
  NAND U3898 ( .A(n3180), .B(n3179), .Z(n4923) );
  OR U3899 ( .A(n3181), .B(n3707), .Z(n3182) );
  NAND U3900 ( .A(n3183), .B(n3182), .Z(n4934) );
  NANDN U3901 ( .A(n3184), .B(n4934), .Z(n3185) );
  NAND U3902 ( .A(n3186), .B(n3185), .Z(n3703) );
  NANDN U3903 ( .A(n3187), .B(n3703), .Z(n3188) );
  NAND U3904 ( .A(n3189), .B(n3188), .Z(n3699) );
  OR U3905 ( .A(n3190), .B(n3694), .Z(n3191) );
  NAND U3906 ( .A(n3192), .B(n3191), .Z(n3690) );
  OR U3907 ( .A(n3193), .B(n3678), .Z(n3194) );
  NAND U3908 ( .A(n3195), .B(n3194), .Z(n3674) );
  NANDN U3909 ( .A(n3196), .B(n3674), .Z(n3197) );
  NAND U3910 ( .A(n3198), .B(n3197), .Z(n3669) );
  NANDN U3911 ( .A(n3199), .B(n3669), .Z(n3200) );
  NAND U3912 ( .A(n3201), .B(n3200), .Z(n3665) );
  NANDN U3913 ( .A(n3202), .B(n3665), .Z(n3203) );
  NAND U3914 ( .A(n3204), .B(n3203), .Z(n3660) );
  NANDN U3915 ( .A(n3205), .B(n3660), .Z(n3206) );
  NAND U3916 ( .A(n3207), .B(n3206), .Z(n3656) );
  OR U3917 ( .A(n3208), .B(n3651), .Z(n3209) );
  NAND U3918 ( .A(n3210), .B(n3209), .Z(n3647) );
  NANDN U3919 ( .A(n3211), .B(n3647), .Z(n3212) );
  NAND U3920 ( .A(n3213), .B(n3212), .Z(n3642) );
  NANDN U3921 ( .A(n3214), .B(n3642), .Z(n3215) );
  NAND U3922 ( .A(n3216), .B(n3215), .Z(n3637) );
  NANDN U3923 ( .A(n3217), .B(n3637), .Z(n3218) );
  NAND U3924 ( .A(n3219), .B(n3218), .Z(n3633) );
  OR U3925 ( .A(n3220), .B(n3629), .Z(n3221) );
  NAND U3926 ( .A(n3222), .B(n3221), .Z(n3625) );
  OR U3927 ( .A(n3223), .B(n3620), .Z(n3224) );
  NAND U3928 ( .A(n3225), .B(n3224), .Z(n3616) );
  OR U3929 ( .A(n3226), .B(n3599), .Z(n3227) );
  NAND U3930 ( .A(n3228), .B(n3227), .Z(n3595) );
  NANDN U3931 ( .A(n3229), .B(n3595), .Z(n3230) );
  NAND U3932 ( .A(n3231), .B(n3230), .Z(n5051) );
  OR U3933 ( .A(n3232), .B(n3587), .Z(n3233) );
  NAND U3934 ( .A(n3234), .B(n3233), .Z(n3582) );
  NANDN U3935 ( .A(n3235), .B(n3582), .Z(n3236) );
  NAND U3936 ( .A(n3237), .B(n3236), .Z(n3577) );
  OR U3937 ( .A(n3238), .B(n3573), .Z(n3239) );
  NAND U3938 ( .A(n3240), .B(n3239), .Z(n3569) );
  NANDN U3939 ( .A(n3241), .B(n3569), .Z(n3242) );
  NAND U3940 ( .A(n3243), .B(n3242), .Z(n3565) );
  OR U3941 ( .A(n3244), .B(n3551), .Z(n3245) );
  NAND U3942 ( .A(n3246), .B(n3245), .Z(n3547) );
  OR U3943 ( .A(n3247), .B(n3530), .Z(n3248) );
  NAND U3944 ( .A(n3249), .B(n3248), .Z(n3525) );
  NANDN U3945 ( .A(n3250), .B(n3525), .Z(n3251) );
  NAND U3946 ( .A(n3252), .B(n3251), .Z(n3521) );
  OR U3947 ( .A(n3253), .B(n3517), .Z(n3254) );
  NAND U3948 ( .A(n3255), .B(n3254), .Z(n3513) );
  OR U3949 ( .A(n3256), .B(n3504), .Z(n3257) );
  NAND U3950 ( .A(n3258), .B(n3257), .Z(n3500) );
  OR U3951 ( .A(n3259), .B(n3495), .Z(n3260) );
  NAND U3952 ( .A(n3261), .B(n3260), .Z(n3489) );
  OR U3953 ( .A(n3262), .B(n3472), .Z(n3263) );
  NAND U3954 ( .A(n3264), .B(n3263), .Z(n3468) );
  OR U3955 ( .A(n3265), .B(n3456), .Z(n3266) );
  NAND U3956 ( .A(n3267), .B(n3266), .Z(n3452) );
  OR U3957 ( .A(n3268), .B(n3440), .Z(n3269) );
  NAND U3958 ( .A(n3270), .B(n3269), .Z(n3436) );
  OR U3959 ( .A(n3271), .B(n3428), .Z(n3272) );
  NAND U3960 ( .A(n3273), .B(n3272), .Z(n3424) );
  NANDN U3961 ( .A(n3274), .B(n3416), .Z(n3275) );
  NAND U3962 ( .A(n3276), .B(n3275), .Z(n3412) );
  OR U3963 ( .A(n3277), .B(n3408), .Z(n3278) );
  NAND U3964 ( .A(n3279), .B(n3278), .Z(n3404) );
  OR U3965 ( .A(n3280), .B(n3378), .Z(n3281) );
  NAND U3966 ( .A(n3282), .B(n3281), .Z(n3374) );
  OR U3967 ( .A(n3283), .B(n3357), .Z(n3284) );
  NAND U3968 ( .A(n3285), .B(n3284), .Z(n3353) );
  NANDN U3969 ( .A(n3286), .B(n3353), .Z(n3287) );
  NAND U3970 ( .A(n3288), .B(n3287), .Z(n3349) );
  NANDN U3971 ( .A(n3289), .B(n3349), .Z(n3290) );
  NAND U3972 ( .A(n3291), .B(n3290), .Z(n3344) );
  NANDN U3973 ( .A(n3292), .B(n3344), .Z(n3293) );
  NAND U3974 ( .A(n3294), .B(n3293), .Z(n3340) );
  OR U3975 ( .A(n3295), .B(n3336), .Z(n3296) );
  NAND U3976 ( .A(n3297), .B(n3296), .Z(n3332) );
  OR U3977 ( .A(n3298), .B(n3323), .Z(n3299) );
  NAND U3978 ( .A(n3300), .B(n3299), .Z(n3319) );
  OR U3979 ( .A(n3301), .B(n3315), .Z(n3302) );
  NAND U3980 ( .A(n3303), .B(n3302), .Z(n3305) );
  XOR U3981 ( .A(n[255]), .B(n3305), .Z(n3304) );
  AND U3982 ( .A(n3304), .B(n523), .Z(n3307) );
  XOR U3983 ( .A(n3308), .B(n3307), .Z(n6580) );
  OR U3984 ( .A(n6580), .B(n[255]), .Z(n3314) );
  NAND U3985 ( .A(n[255]), .B(n3305), .Z(n3306) );
  OR U3986 ( .A(n3306), .B(n524), .Z(n3310) );
  NAND U3987 ( .A(n3308), .B(n3307), .Z(n3309) );
  NAND U3988 ( .A(n3310), .B(n3309), .Z(n3311) );
  XNOR U3989 ( .A(n3312), .B(n3311), .Z(n6594) );
  NANDN U3990 ( .A(n3313), .B(n6594), .Z(n6577) );
  ANDN U3991 ( .B(n3314), .A(n6577), .Z(n5340) );
  XOR U3992 ( .A(n6582), .B(n3315), .Z(n3316) );
  NANDN U3993 ( .A(n524), .B(n3316), .Z(n3317) );
  XNOR U3994 ( .A(n3318), .B(n3317), .Z(n6583) );
  NANDN U3995 ( .A(n6582), .B(n6583), .Z(n5336) );
  XNOR U3996 ( .A(n6582), .B(n6583), .Z(n5334) );
  XOR U3997 ( .A(n[253]), .B(n3319), .Z(n3320) );
  NANDN U3998 ( .A(n524), .B(n3320), .Z(n3321) );
  XNOR U3999 ( .A(n3322), .B(n3321), .Z(n6571) );
  NAND U4000 ( .A(n[253]), .B(n6571), .Z(n5332) );
  XOR U4001 ( .A(n6571), .B(n[253]), .Z(n5330) );
  XOR U4002 ( .A(n3327), .B(n3323), .Z(n3324) );
  NANDN U4003 ( .A(n524), .B(n3324), .Z(n3325) );
  XNOR U4004 ( .A(n3326), .B(n3325), .Z(n6564) );
  NANDN U4005 ( .A(n3327), .B(n6564), .Z(n5328) );
  XNOR U4006 ( .A(n3327), .B(n6564), .Z(n5326) );
  XNOR U4007 ( .A(n[251]), .B(n3328), .Z(n3329) );
  NANDN U4008 ( .A(n524), .B(n3329), .Z(n3330) );
  XNOR U4009 ( .A(n3331), .B(n3330), .Z(n6558) );
  NAND U4010 ( .A(n[251]), .B(n6558), .Z(n5324) );
  XOR U4011 ( .A(n6558), .B(n[251]), .Z(n5322) );
  XOR U4012 ( .A(n[250]), .B(n3332), .Z(n3333) );
  NANDN U4013 ( .A(n524), .B(n3333), .Z(n3334) );
  XNOR U4014 ( .A(n3335), .B(n3334), .Z(n6552) );
  NAND U4015 ( .A(n[250]), .B(n6552), .Z(n5320) );
  XOR U4016 ( .A(n[250]), .B(n6552), .Z(n5318) );
  XOR U4017 ( .A(n6534), .B(n3336), .Z(n3337) );
  NANDN U4018 ( .A(n524), .B(n3337), .Z(n3338) );
  XNOR U4019 ( .A(n3339), .B(n3338), .Z(n6546) );
  NANDN U4020 ( .A(n6534), .B(n6546), .Z(n5316) );
  XNOR U4021 ( .A(n6546), .B(n6534), .Z(n5314) );
  XOR U4022 ( .A(n[248]), .B(n3340), .Z(n3341) );
  NANDN U4023 ( .A(n524), .B(n3341), .Z(n3342) );
  XNOR U4024 ( .A(n3343), .B(n3342), .Z(n6528) );
  NAND U4025 ( .A(n[248]), .B(n6528), .Z(n5312) );
  XOR U4026 ( .A(n[248]), .B(n6528), .Z(n5310) );
  XNOR U4027 ( .A(n3348), .B(n3344), .Z(n3345) );
  NANDN U4028 ( .A(n524), .B(n3345), .Z(n3346) );
  XNOR U4029 ( .A(n3347), .B(n3346), .Z(n6522) );
  NANDN U4030 ( .A(n3348), .B(n6522), .Z(n5308) );
  XNOR U4031 ( .A(n6522), .B(n3348), .Z(n5306) );
  XNOR U4032 ( .A(n6514), .B(n3349), .Z(n3350) );
  NANDN U4033 ( .A(n524), .B(n3350), .Z(n3351) );
  XNOR U4034 ( .A(n3352), .B(n3351), .Z(n6515) );
  NANDN U4035 ( .A(n6514), .B(n6515), .Z(n5304) );
  XNOR U4036 ( .A(n6514), .B(n6515), .Z(n5302) );
  XOR U4037 ( .A(n[245]), .B(n3353), .Z(n3354) );
  NANDN U4038 ( .A(n524), .B(n3354), .Z(n3355) );
  XNOR U4039 ( .A(n3356), .B(n3355), .Z(n6508) );
  NAND U4040 ( .A(n[245]), .B(n6508), .Z(n5300) );
  XOR U4041 ( .A(n6508), .B(n[245]), .Z(n5298) );
  XOR U4042 ( .A(n3361), .B(n3357), .Z(n3358) );
  NANDN U4043 ( .A(n524), .B(n3358), .Z(n3359) );
  XNOR U4044 ( .A(n3360), .B(n3359), .Z(n6503) );
  NANDN U4045 ( .A(n3361), .B(n6503), .Z(n5296) );
  XNOR U4046 ( .A(n3361), .B(n6503), .Z(n5294) );
  XNOR U4047 ( .A(n[243]), .B(n3362), .Z(n3363) );
  NANDN U4048 ( .A(n524), .B(n3363), .Z(n3364) );
  XNOR U4049 ( .A(n3365), .B(n3364), .Z(n6496) );
  NAND U4050 ( .A(n[243]), .B(n6496), .Z(n5292) );
  XOR U4051 ( .A(n6496), .B(n[243]), .Z(n5290) );
  XNOR U4052 ( .A(n[242]), .B(n3366), .Z(n3367) );
  NANDN U4053 ( .A(n524), .B(n3367), .Z(n3368) );
  XNOR U4054 ( .A(n3369), .B(n3368), .Z(n6490) );
  NAND U4055 ( .A(n[242]), .B(n6490), .Z(n5288) );
  XOR U4056 ( .A(n[242]), .B(n6490), .Z(n5286) );
  XNOR U4057 ( .A(n[241]), .B(n3370), .Z(n3371) );
  NANDN U4058 ( .A(n524), .B(n3371), .Z(n3372) );
  XNOR U4059 ( .A(n3373), .B(n3372), .Z(n6483) );
  NAND U4060 ( .A(n[241]), .B(n6483), .Z(n5284) );
  XOR U4061 ( .A(n6483), .B(n[241]), .Z(n5282) );
  XOR U4062 ( .A(n[240]), .B(n3374), .Z(n3375) );
  NANDN U4063 ( .A(n524), .B(n3375), .Z(n3376) );
  XNOR U4064 ( .A(n3377), .B(n3376), .Z(n6477) );
  NAND U4065 ( .A(n[240]), .B(n6477), .Z(n5280) );
  XOR U4066 ( .A(n[240]), .B(n6477), .Z(n5278) );
  XOR U4067 ( .A(n3382), .B(n3378), .Z(n3379) );
  NANDN U4068 ( .A(n524), .B(n3379), .Z(n3380) );
  XNOR U4069 ( .A(n3381), .B(n3380), .Z(n6474) );
  NANDN U4070 ( .A(n3382), .B(n6474), .Z(n5276) );
  XNOR U4071 ( .A(n6474), .B(n3382), .Z(n5274) );
  XNOR U4072 ( .A(n[238]), .B(n3383), .Z(n3384) );
  NANDN U4073 ( .A(n524), .B(n3384), .Z(n3385) );
  XNOR U4074 ( .A(n3386), .B(n3385), .Z(n6466) );
  NAND U4075 ( .A(n[238]), .B(n6466), .Z(n5272) );
  XOR U4076 ( .A(n[238]), .B(n6466), .Z(n5270) );
  XOR U4077 ( .A(n6449), .B(n3387), .Z(n3388) );
  NANDN U4078 ( .A(n524), .B(n3388), .Z(n3389) );
  XOR U4079 ( .A(n3390), .B(n3389), .Z(n5263) );
  IV U4080 ( .A(n5263), .Z(n6450) );
  XNOR U4081 ( .A(n[235]), .B(n3391), .Z(n3392) );
  NANDN U4082 ( .A(n524), .B(n3392), .Z(n3393) );
  XNOR U4083 ( .A(n3394), .B(n3393), .Z(n6443) );
  NAND U4084 ( .A(n[235]), .B(n6443), .Z(n5256) );
  XOR U4085 ( .A(n6443), .B(n[235]), .Z(n5254) );
  XOR U4086 ( .A(n3399), .B(n3395), .Z(n3396) );
  NANDN U4087 ( .A(n524), .B(n3396), .Z(n3397) );
  XOR U4088 ( .A(n3398), .B(n3397), .Z(n6439) );
  NANDN U4089 ( .A(n3399), .B(n6439), .Z(n5252) );
  XNOR U4090 ( .A(n3399), .B(n6439), .Z(n5250) );
  XNOR U4091 ( .A(n[233]), .B(n3400), .Z(n3401) );
  NANDN U4092 ( .A(n524), .B(n3401), .Z(n3402) );
  XNOR U4093 ( .A(n3403), .B(n3402), .Z(n6434) );
  NAND U4094 ( .A(n[233]), .B(n6434), .Z(n5248) );
  XOR U4095 ( .A(n6434), .B(n[233]), .Z(n5246) );
  XOR U4096 ( .A(n[232]), .B(n3404), .Z(n3405) );
  NANDN U4097 ( .A(n524), .B(n3405), .Z(n3406) );
  XNOR U4098 ( .A(n3407), .B(n3406), .Z(n6427) );
  NAND U4099 ( .A(n[232]), .B(n6427), .Z(n5244) );
  XOR U4100 ( .A(n[232]), .B(n6427), .Z(n5242) );
  XOR U4101 ( .A(n6413), .B(n3408), .Z(n3409) );
  NANDN U4102 ( .A(n524), .B(n3409), .Z(n3410) );
  XNOR U4103 ( .A(n3411), .B(n3410), .Z(n6415) );
  OR U4104 ( .A(n6415), .B(n[231]), .Z(n5239) );
  XNOR U4105 ( .A(n[229]), .B(n3412), .Z(n3413) );
  NANDN U4106 ( .A(n524), .B(n3413), .Z(n3414) );
  XNOR U4107 ( .A(n3415), .B(n3414), .Z(n6407) );
  NAND U4108 ( .A(n[229]), .B(n6407), .Z(n5229) );
  XOR U4109 ( .A(n6407), .B(n[229]), .Z(n5227) );
  XNOR U4110 ( .A(n[228]), .B(n3416), .Z(n3417) );
  NANDN U4111 ( .A(n524), .B(n3417), .Z(n3418) );
  XNOR U4112 ( .A(n3419), .B(n3418), .Z(n6397) );
  NAND U4113 ( .A(n[228]), .B(n6397), .Z(n5225) );
  XOR U4114 ( .A(n6397), .B(n[228]), .Z(n5223) );
  XNOR U4115 ( .A(n[227]), .B(n3420), .Z(n3421) );
  NANDN U4116 ( .A(n524), .B(n3421), .Z(n3422) );
  XNOR U4117 ( .A(n3423), .B(n3422), .Z(n6390) );
  NAND U4118 ( .A(n[227]), .B(n6390), .Z(n5221) );
  XOR U4119 ( .A(n[227]), .B(n6390), .Z(n5219) );
  XOR U4120 ( .A(n[226]), .B(n3424), .Z(n3425) );
  NANDN U4121 ( .A(n524), .B(n3425), .Z(n3426) );
  XNOR U4122 ( .A(n3427), .B(n3426), .Z(n6383) );
  NAND U4123 ( .A(n[226]), .B(n6383), .Z(n5217) );
  XOR U4124 ( .A(n6383), .B(n[226]), .Z(n5215) );
  XOR U4125 ( .A(n6376), .B(n3428), .Z(n3429) );
  NANDN U4126 ( .A(n524), .B(n3429), .Z(n3430) );
  XNOR U4127 ( .A(n3431), .B(n3430), .Z(n6377) );
  NANDN U4128 ( .A(n6376), .B(n6377), .Z(n5213) );
  XNOR U4129 ( .A(n6376), .B(n6377), .Z(n5211) );
  XNOR U4130 ( .A(n[224]), .B(n3432), .Z(n3433) );
  NANDN U4131 ( .A(n524), .B(n3433), .Z(n3434) );
  XNOR U4132 ( .A(n3435), .B(n3434), .Z(n6371) );
  NAND U4133 ( .A(n[224]), .B(n6371), .Z(n5209) );
  XOR U4134 ( .A(n6371), .B(n[224]), .Z(n5207) );
  XOR U4135 ( .A(n[223]), .B(n3436), .Z(n3437) );
  NANDN U4136 ( .A(n524), .B(n3437), .Z(n3438) );
  XNOR U4137 ( .A(n3439), .B(n3438), .Z(n6365) );
  NAND U4138 ( .A(n[223]), .B(n6365), .Z(n5205) );
  XOR U4139 ( .A(n[223]), .B(n6365), .Z(n5203) );
  XOR U4140 ( .A(n6357), .B(n3440), .Z(n3441) );
  NANDN U4141 ( .A(n524), .B(n3441), .Z(n3442) );
  XNOR U4142 ( .A(n3443), .B(n3442), .Z(n6358) );
  NANDN U4143 ( .A(n6357), .B(n6358), .Z(n5201) );
  XNOR U4144 ( .A(n6358), .B(n6357), .Z(n5199) );
  XNOR U4145 ( .A(n[221]), .B(n3444), .Z(n3445) );
  NANDN U4146 ( .A(n524), .B(n3445), .Z(n3446) );
  XNOR U4147 ( .A(n3447), .B(n3446), .Z(n6351) );
  NAND U4148 ( .A(n[221]), .B(n6351), .Z(n5197) );
  XOR U4149 ( .A(n6351), .B(n[221]), .Z(n5195) );
  XNOR U4150 ( .A(n[220]), .B(n3448), .Z(n3449) );
  NANDN U4151 ( .A(n524), .B(n3449), .Z(n3450) );
  XNOR U4152 ( .A(n3451), .B(n3450), .Z(n6342) );
  NAND U4153 ( .A(n[220]), .B(n6342), .Z(n5193) );
  XOR U4154 ( .A(n[220]), .B(n6342), .Z(n5191) );
  XOR U4155 ( .A(n[219]), .B(n3452), .Z(n3453) );
  NANDN U4156 ( .A(n524), .B(n3453), .Z(n3454) );
  XNOR U4157 ( .A(n3455), .B(n3454), .Z(n6335) );
  NAND U4158 ( .A(n[219]), .B(n6335), .Z(n5189) );
  XOR U4159 ( .A(n6335), .B(n[219]), .Z(n5187) );
  XOR U4160 ( .A(n6317), .B(n3456), .Z(n3457) );
  NANDN U4161 ( .A(n524), .B(n3457), .Z(n3458) );
  XNOR U4162 ( .A(n3459), .B(n3458), .Z(n6319) );
  NANDN U4163 ( .A(n6317), .B(n6319), .Z(n6326) );
  XNOR U4164 ( .A(n[216]), .B(n3460), .Z(n3461) );
  NANDN U4165 ( .A(n524), .B(n3461), .Z(n3462) );
  XNOR U4166 ( .A(n3463), .B(n3462), .Z(n6311) );
  NAND U4167 ( .A(n[216]), .B(n6311), .Z(n5174) );
  XOR U4168 ( .A(n6311), .B(n[216]), .Z(n5172) );
  XNOR U4169 ( .A(n[215]), .B(n3464), .Z(n3465) );
  NANDN U4170 ( .A(n524), .B(n3465), .Z(n3466) );
  XNOR U4171 ( .A(n3467), .B(n3466), .Z(n6305) );
  NAND U4172 ( .A(n[215]), .B(n6305), .Z(n5170) );
  XOR U4173 ( .A(n[215]), .B(n6305), .Z(n5168) );
  XOR U4174 ( .A(n[214]), .B(n3468), .Z(n3469) );
  NANDN U4175 ( .A(n524), .B(n3469), .Z(n3470) );
  XOR U4176 ( .A(n3471), .B(n3470), .Z(n6302) );
  NANDN U4177 ( .A(n6302), .B(n[214]), .Z(n5166) );
  XNOR U4178 ( .A(n6302), .B(n[214]), .Z(n5164) );
  XOR U4179 ( .A(n3476), .B(n3472), .Z(n3473) );
  NANDN U4180 ( .A(n524), .B(n3473), .Z(n3474) );
  XNOR U4181 ( .A(n3475), .B(n3474), .Z(n6295) );
  NANDN U4182 ( .A(n3476), .B(n6295), .Z(n5162) );
  XNOR U4183 ( .A(n3476), .B(n6295), .Z(n5160) );
  XNOR U4184 ( .A(n[212]), .B(n3477), .Z(n3478) );
  NANDN U4185 ( .A(n524), .B(n3478), .Z(n3479) );
  XNOR U4186 ( .A(n3480), .B(n3479), .Z(n6289) );
  NAND U4187 ( .A(n[212]), .B(n6289), .Z(n5158) );
  XOR U4188 ( .A(n6289), .B(n[212]), .Z(n5156) );
  XNOR U4189 ( .A(n[211]), .B(n3481), .Z(n3482) );
  NANDN U4190 ( .A(n524), .B(n3482), .Z(n3483) );
  XNOR U4191 ( .A(n3484), .B(n3483), .Z(n6283) );
  NAND U4192 ( .A(n[211]), .B(n6283), .Z(n5154) );
  XOR U4193 ( .A(n[211]), .B(n6283), .Z(n5152) );
  XOR U4194 ( .A(n6268), .B(n3485), .Z(n3486) );
  NANDN U4195 ( .A(n524), .B(n3486), .Z(n3487) );
  XOR U4196 ( .A(n3488), .B(n3487), .Z(n6270) );
  ANDN U4197 ( .B(n6270), .A(n6268), .Z(n6278) );
  XNOR U4198 ( .A(n6256), .B(n3489), .Z(n3490) );
  NANDN U4199 ( .A(n524), .B(n3490), .Z(n3491) );
  XOR U4200 ( .A(n3492), .B(n3491), .Z(n6271) );
  NANDN U4201 ( .A(n[209]), .B(n6271), .Z(n3494) );
  NOR U4202 ( .A(n[210]), .B(n6270), .Z(n3493) );
  ANDN U4203 ( .B(n3494), .A(n3493), .Z(n5149) );
  XOR U4204 ( .A(n3499), .B(n3495), .Z(n3496) );
  NANDN U4205 ( .A(n524), .B(n3496), .Z(n3497) );
  XNOR U4206 ( .A(n3498), .B(n3497), .Z(n6254) );
  NANDN U4207 ( .A(n3499), .B(n6254), .Z(n5145) );
  XNOR U4208 ( .A(n3499), .B(n6254), .Z(n5143) );
  XOR U4209 ( .A(n[207]), .B(n3500), .Z(n3501) );
  NANDN U4210 ( .A(n524), .B(n3501), .Z(n3502) );
  XNOR U4211 ( .A(n3503), .B(n3502), .Z(n6249) );
  NAND U4212 ( .A(n[207]), .B(n6249), .Z(n5141) );
  XOR U4213 ( .A(n6249), .B(n[207]), .Z(n5139) );
  XOR U4214 ( .A(n3508), .B(n3504), .Z(n3505) );
  NANDN U4215 ( .A(n524), .B(n3505), .Z(n3506) );
  XNOR U4216 ( .A(n3507), .B(n3506), .Z(n6242) );
  NANDN U4217 ( .A(n3508), .B(n6242), .Z(n5137) );
  XNOR U4218 ( .A(n3508), .B(n6242), .Z(n5135) );
  XNOR U4219 ( .A(n[205]), .B(n3509), .Z(n3510) );
  NANDN U4220 ( .A(n524), .B(n3510), .Z(n3511) );
  XNOR U4221 ( .A(n3512), .B(n3511), .Z(n6239) );
  NAND U4222 ( .A(n[205]), .B(n6239), .Z(n5133) );
  XOR U4223 ( .A(n6239), .B(n[205]), .Z(n5131) );
  XOR U4224 ( .A(n[204]), .B(n3513), .Z(n3514) );
  NANDN U4225 ( .A(n524), .B(n3514), .Z(n3515) );
  XNOR U4226 ( .A(n3516), .B(n3515), .Z(n6232) );
  NAND U4227 ( .A(n[204]), .B(n6232), .Z(n5129) );
  XOR U4228 ( .A(n[204]), .B(n6232), .Z(n5127) );
  XOR U4229 ( .A(n6225), .B(n3517), .Z(n3518) );
  NANDN U4230 ( .A(n524), .B(n3518), .Z(n3519) );
  XNOR U4231 ( .A(n3520), .B(n3519), .Z(n6226) );
  NANDN U4232 ( .A(n6225), .B(n6226), .Z(n5125) );
  XNOR U4233 ( .A(n6226), .B(n6225), .Z(n5123) );
  XOR U4234 ( .A(n[202]), .B(n3521), .Z(n3522) );
  NANDN U4235 ( .A(n524), .B(n3522), .Z(n3523) );
  XNOR U4236 ( .A(n3524), .B(n3523), .Z(n6219) );
  NAND U4237 ( .A(n[202]), .B(n6219), .Z(n5121) );
  XOR U4238 ( .A(n[202]), .B(n6219), .Z(n5119) );
  XNOR U4239 ( .A(n3529), .B(n3525), .Z(n3526) );
  NANDN U4240 ( .A(n524), .B(n3526), .Z(n3527) );
  XNOR U4241 ( .A(n3528), .B(n3527), .Z(n6213) );
  NANDN U4242 ( .A(n3529), .B(n6213), .Z(n5117) );
  XNOR U4243 ( .A(n6213), .B(n3529), .Z(n5115) );
  XOR U4244 ( .A(n6199), .B(n3530), .Z(n3531) );
  NANDN U4245 ( .A(n524), .B(n3531), .Z(n3532) );
  XNOR U4246 ( .A(n3533), .B(n3532), .Z(n6201) );
  NANDN U4247 ( .A(n6199), .B(n6201), .Z(n6208) );
  XNOR U4248 ( .A(n[199]), .B(n3534), .Z(n3535) );
  NANDN U4249 ( .A(n524), .B(n3535), .Z(n3536) );
  XNOR U4250 ( .A(n3537), .B(n3536), .Z(n6202) );
  NAND U4251 ( .A(n[199]), .B(n6202), .Z(n3538) );
  AND U4252 ( .A(n6208), .B(n3538), .Z(n5111) );
  XOR U4253 ( .A(n6202), .B(n[199]), .Z(n5109) );
  XNOR U4254 ( .A(n[198]), .B(n3539), .Z(n3540) );
  NANDN U4255 ( .A(n524), .B(n3540), .Z(n3541) );
  XNOR U4256 ( .A(n3542), .B(n3541), .Z(n6188) );
  NAND U4257 ( .A(n[198]), .B(n6188), .Z(n5107) );
  XOR U4258 ( .A(n[198]), .B(n6188), .Z(n5105) );
  XNOR U4259 ( .A(n[197]), .B(n3543), .Z(n3544) );
  NANDN U4260 ( .A(n524), .B(n3544), .Z(n3545) );
  XNOR U4261 ( .A(n3546), .B(n3545), .Z(n6181) );
  NAND U4262 ( .A(n[197]), .B(n6181), .Z(n5103) );
  XOR U4263 ( .A(n6181), .B(n[197]), .Z(n5101) );
  XNOR U4264 ( .A(n6166), .B(n3547), .Z(n3548) );
  NANDN U4265 ( .A(n524), .B(n3548), .Z(n3549) );
  XNOR U4266 ( .A(n3550), .B(n3549), .Z(n6168) );
  NANDN U4267 ( .A(n6166), .B(n6168), .Z(n6175) );
  XOR U4268 ( .A(n3556), .B(n3551), .Z(n3552) );
  NANDN U4269 ( .A(n524), .B(n3552), .Z(n3553) );
  XNOR U4270 ( .A(n3554), .B(n3553), .Z(n6169) );
  NANDN U4271 ( .A(n3556), .B(n6169), .Z(n3555) );
  AND U4272 ( .A(n6175), .B(n3555), .Z(n5097) );
  XNOR U4273 ( .A(n6169), .B(n3556), .Z(n5095) );
  XNOR U4274 ( .A(n[194]), .B(n3557), .Z(n3558) );
  NANDN U4275 ( .A(n524), .B(n3558), .Z(n3559) );
  XNOR U4276 ( .A(n3560), .B(n3559), .Z(n6160) );
  NAND U4277 ( .A(n[194]), .B(n6160), .Z(n5093) );
  XOR U4278 ( .A(n[194]), .B(n6160), .Z(n5091) );
  XNOR U4279 ( .A(n[193]), .B(n3561), .Z(n3562) );
  NANDN U4280 ( .A(n524), .B(n3562), .Z(n3563) );
  XNOR U4281 ( .A(n3564), .B(n3563), .Z(n6154) );
  NAND U4282 ( .A(n[193]), .B(n6154), .Z(n5089) );
  XOR U4283 ( .A(n6154), .B(n[193]), .Z(n5087) );
  XOR U4284 ( .A(n[192]), .B(n3565), .Z(n3566) );
  NANDN U4285 ( .A(n524), .B(n3566), .Z(n3567) );
  XNOR U4286 ( .A(n3568), .B(n3567), .Z(n6148) );
  NAND U4287 ( .A(n[192]), .B(n6148), .Z(n5085) );
  XOR U4288 ( .A(n[192]), .B(n6148), .Z(n5083) );
  XOR U4289 ( .A(n[191]), .B(n3569), .Z(n3570) );
  NANDN U4290 ( .A(n524), .B(n3570), .Z(n3571) );
  XNOR U4291 ( .A(n3572), .B(n3571), .Z(n6142) );
  NAND U4292 ( .A(n[191]), .B(n6142), .Z(n5081) );
  XOR U4293 ( .A(n6142), .B(n[191]), .Z(n5079) );
  XOR U4294 ( .A(n6135), .B(n3573), .Z(n3574) );
  NANDN U4295 ( .A(n524), .B(n3574), .Z(n3575) );
  XNOR U4296 ( .A(n3576), .B(n3575), .Z(n6136) );
  NANDN U4297 ( .A(n6135), .B(n6136), .Z(n5077) );
  XNOR U4298 ( .A(n6136), .B(n6135), .Z(n5075) );
  XNOR U4299 ( .A(n3581), .B(n3577), .Z(n3578) );
  NANDN U4300 ( .A(n524), .B(n3578), .Z(n3579) );
  XOR U4301 ( .A(n3580), .B(n3579), .Z(n6130) );
  NANDN U4302 ( .A(n3581), .B(n6130), .Z(n5073) );
  XNOR U4303 ( .A(n3581), .B(n6130), .Z(n5071) );
  XNOR U4304 ( .A(n3586), .B(n3582), .Z(n3583) );
  NANDN U4305 ( .A(n524), .B(n3583), .Z(n3584) );
  XNOR U4306 ( .A(n3585), .B(n3584), .Z(n6113) );
  NANDN U4307 ( .A(n3586), .B(n6113), .Z(n5069) );
  XNOR U4308 ( .A(n6113), .B(n3586), .Z(n5067) );
  XOR U4309 ( .A(n6106), .B(n3587), .Z(n3588) );
  NANDN U4310 ( .A(n524), .B(n3588), .Z(n3589) );
  XNOR U4311 ( .A(n3590), .B(n3589), .Z(n6107) );
  NANDN U4312 ( .A(n6106), .B(n6107), .Z(n5065) );
  XNOR U4313 ( .A(n6106), .B(n6107), .Z(n5063) );
  XNOR U4314 ( .A(n[186]), .B(n3591), .Z(n3592) );
  NANDN U4315 ( .A(n524), .B(n3592), .Z(n3593) );
  XNOR U4316 ( .A(n3594), .B(n3593), .Z(n6100) );
  NAND U4317 ( .A(n[186]), .B(n6100), .Z(n5061) );
  XOR U4318 ( .A(n6100), .B(n[186]), .Z(n5059) );
  XNOR U4319 ( .A(n6086), .B(n3595), .Z(n3596) );
  NANDN U4320 ( .A(n524), .B(n3596), .Z(n3597) );
  XNOR U4321 ( .A(n3598), .B(n3597), .Z(n6087) );
  NANDN U4322 ( .A(n6086), .B(n6087), .Z(n5049) );
  XNOR U4323 ( .A(n6086), .B(n6087), .Z(n5047) );
  XOR U4324 ( .A(n3603), .B(n3599), .Z(n3600) );
  NANDN U4325 ( .A(n524), .B(n3600), .Z(n3601) );
  XNOR U4326 ( .A(n3602), .B(n3601), .Z(n6080) );
  NANDN U4327 ( .A(n3603), .B(n6080), .Z(n5045) );
  XNOR U4328 ( .A(n6080), .B(n3603), .Z(n5043) );
  XNOR U4329 ( .A(n[182]), .B(n3604), .Z(n3605) );
  NANDN U4330 ( .A(n524), .B(n3605), .Z(n3606) );
  XNOR U4331 ( .A(n3607), .B(n3606), .Z(n6073) );
  NAND U4332 ( .A(n[182]), .B(n6073), .Z(n5041) );
  XOR U4333 ( .A(n6073), .B(n[182]), .Z(n5039) );
  XNOR U4334 ( .A(n[181]), .B(n3608), .Z(n3609) );
  NANDN U4335 ( .A(n524), .B(n3609), .Z(n3610) );
  XNOR U4336 ( .A(n3611), .B(n3610), .Z(n6067) );
  NAND U4337 ( .A(n[181]), .B(n6067), .Z(n5037) );
  XOR U4338 ( .A(n[181]), .B(n6067), .Z(n5035) );
  XNOR U4339 ( .A(n[180]), .B(n3612), .Z(n3613) );
  NANDN U4340 ( .A(n524), .B(n3613), .Z(n3614) );
  XNOR U4341 ( .A(n3615), .B(n3614), .Z(n6061) );
  NAND U4342 ( .A(n[180]), .B(n6061), .Z(n5033) );
  XOR U4343 ( .A(n6061), .B(n[180]), .Z(n5031) );
  XNOR U4344 ( .A(n6039), .B(n3616), .Z(n3617) );
  NANDN U4345 ( .A(n524), .B(n3617), .Z(n3618) );
  XOR U4346 ( .A(n3619), .B(n3618), .Z(n6041) );
  NANDN U4347 ( .A(n[178]), .B(n6041), .Z(n5021) );
  NANDN U4348 ( .A(n6041), .B(n[178]), .Z(n6049) );
  XOR U4349 ( .A(n6042), .B(n3620), .Z(n3621) );
  NANDN U4350 ( .A(n524), .B(n3621), .Z(n3622) );
  XNOR U4351 ( .A(n3623), .B(n3622), .Z(n6043) );
  NANDN U4352 ( .A(n6042), .B(n6043), .Z(n3624) );
  AND U4353 ( .A(n6049), .B(n3624), .Z(n5019) );
  XNOR U4354 ( .A(n6043), .B(n6042), .Z(n5017) );
  XNOR U4355 ( .A(n6025), .B(n3625), .Z(n3626) );
  NANDN U4356 ( .A(n524), .B(n3626), .Z(n3627) );
  XOR U4357 ( .A(n3628), .B(n3627), .Z(n6033) );
  NANDN U4358 ( .A(n6033), .B(n[176]), .Z(n5015) );
  XNOR U4359 ( .A(n[176]), .B(n6033), .Z(n5013) );
  XOR U4360 ( .A(n6024), .B(n3629), .Z(n3630) );
  NANDN U4361 ( .A(n524), .B(n3630), .Z(n3631) );
  XNOR U4362 ( .A(n3632), .B(n3631), .Z(n6026) );
  NANDN U4363 ( .A(n6024), .B(n6026), .Z(n5011) );
  XNOR U4364 ( .A(n6026), .B(n6024), .Z(n5009) );
  XOR U4365 ( .A(n[174]), .B(n3633), .Z(n3634) );
  NANDN U4366 ( .A(n524), .B(n3634), .Z(n3635) );
  XNOR U4367 ( .A(n3636), .B(n3635), .Z(n6018) );
  NAND U4368 ( .A(n[174]), .B(n6018), .Z(n5007) );
  XOR U4369 ( .A(n[174]), .B(n6018), .Z(n5005) );
  XNOR U4370 ( .A(n3641), .B(n3637), .Z(n3638) );
  NANDN U4371 ( .A(n524), .B(n3638), .Z(n3639) );
  XNOR U4372 ( .A(n3640), .B(n3639), .Z(n6012) );
  NANDN U4373 ( .A(n3641), .B(n6012), .Z(n5003) );
  XNOR U4374 ( .A(n6012), .B(n3641), .Z(n5001) );
  XNOR U4375 ( .A(n3646), .B(n3642), .Z(n3643) );
  NANDN U4376 ( .A(n524), .B(n3643), .Z(n3644) );
  XNOR U4377 ( .A(n3645), .B(n3644), .Z(n6005) );
  NANDN U4378 ( .A(n3646), .B(n6005), .Z(n4999) );
  XNOR U4379 ( .A(n6005), .B(n3646), .Z(n4997) );
  XNOR U4380 ( .A(n5998), .B(n3647), .Z(n3648) );
  NANDN U4381 ( .A(n524), .B(n3648), .Z(n3649) );
  XNOR U4382 ( .A(n3650), .B(n3649), .Z(n5999) );
  NANDN U4383 ( .A(n5998), .B(n5999), .Z(n4995) );
  XNOR U4384 ( .A(n5998), .B(n5999), .Z(n4993) );
  XOR U4385 ( .A(n3655), .B(n3651), .Z(n3652) );
  NANDN U4386 ( .A(n524), .B(n3652), .Z(n3653) );
  XOR U4387 ( .A(n3654), .B(n3653), .Z(n5993) );
  IV U4388 ( .A(n5993), .Z(n5994) );
  NANDN U4389 ( .A(n3655), .B(n5994), .Z(n4991) );
  XNOR U4390 ( .A(n5993), .B(n[170]), .Z(n4989) );
  XOR U4391 ( .A(n[169]), .B(n3656), .Z(n3657) );
  NANDN U4392 ( .A(n524), .B(n3657), .Z(n3658) );
  XNOR U4393 ( .A(n3659), .B(n3658), .Z(n5986) );
  NAND U4394 ( .A(n[169]), .B(n5986), .Z(n4987) );
  XOR U4395 ( .A(n5986), .B(n[169]), .Z(n4985) );
  XNOR U4396 ( .A(n3664), .B(n3660), .Z(n3661) );
  NANDN U4397 ( .A(n524), .B(n3661), .Z(n3662) );
  XNOR U4398 ( .A(n3663), .B(n3662), .Z(n5970) );
  NANDN U4399 ( .A(n3664), .B(n5970), .Z(n4983) );
  XNOR U4400 ( .A(n3664), .B(n5970), .Z(n4981) );
  XOR U4401 ( .A(n[167]), .B(n3665), .Z(n3666) );
  NANDN U4402 ( .A(n524), .B(n3666), .Z(n3667) );
  XNOR U4403 ( .A(n3668), .B(n3667), .Z(n5964) );
  NAND U4404 ( .A(n[167]), .B(n5964), .Z(n4979) );
  XOR U4405 ( .A(n5964), .B(n[167]), .Z(n4977) );
  XNOR U4406 ( .A(n3673), .B(n3669), .Z(n3670) );
  NANDN U4407 ( .A(n524), .B(n3670), .Z(n3671) );
  XNOR U4408 ( .A(n3672), .B(n3671), .Z(n5958) );
  NANDN U4409 ( .A(n3673), .B(n5958), .Z(n4975) );
  XNOR U4410 ( .A(n3673), .B(n5958), .Z(n4973) );
  XOR U4411 ( .A(n[165]), .B(n3674), .Z(n3675) );
  NANDN U4412 ( .A(n524), .B(n3675), .Z(n3676) );
  XNOR U4413 ( .A(n3677), .B(n3676), .Z(n5951) );
  NAND U4414 ( .A(n[165]), .B(n5951), .Z(n4971) );
  XOR U4415 ( .A(n5951), .B(n[165]), .Z(n4969) );
  XOR U4416 ( .A(n5943), .B(n3678), .Z(n3679) );
  NANDN U4417 ( .A(n524), .B(n3679), .Z(n3680) );
  XNOR U4418 ( .A(n3681), .B(n3680), .Z(n5945) );
  NANDN U4419 ( .A(n5943), .B(n5945), .Z(n4967) );
  XNOR U4420 ( .A(n5943), .B(n5945), .Z(n4965) );
  XNOR U4421 ( .A(n[163]), .B(n3682), .Z(n3683) );
  NANDN U4422 ( .A(n524), .B(n3683), .Z(n3684) );
  XNOR U4423 ( .A(n3685), .B(n3684), .Z(n5937) );
  NAND U4424 ( .A(n[163]), .B(n5937), .Z(n4963) );
  XOR U4425 ( .A(n5937), .B(n[163]), .Z(n4961) );
  XNOR U4426 ( .A(n[162]), .B(n3686), .Z(n3687) );
  NANDN U4427 ( .A(n524), .B(n3687), .Z(n3688) );
  XNOR U4428 ( .A(n3689), .B(n3688), .Z(n5931) );
  NAND U4429 ( .A(n[162]), .B(n5931), .Z(n4959) );
  XOR U4430 ( .A(n[162]), .B(n5931), .Z(n4957) );
  XOR U4431 ( .A(n[161]), .B(n3690), .Z(n3691) );
  NANDN U4432 ( .A(n524), .B(n3691), .Z(n3692) );
  XNOR U4433 ( .A(n3693), .B(n3692), .Z(n5928) );
  NAND U4434 ( .A(n[161]), .B(n5928), .Z(n4955) );
  XOR U4435 ( .A(n5928), .B(n[161]), .Z(n4953) );
  XOR U4436 ( .A(n3698), .B(n3694), .Z(n3695) );
  NANDN U4437 ( .A(n524), .B(n3695), .Z(n3696) );
  XNOR U4438 ( .A(n3697), .B(n3696), .Z(n5924) );
  NANDN U4439 ( .A(n3698), .B(n5924), .Z(n4951) );
  XNOR U4440 ( .A(n3698), .B(n5924), .Z(n4949) );
  XOR U4441 ( .A(n[159]), .B(n3699), .Z(n3700) );
  NANDN U4442 ( .A(n524), .B(n3700), .Z(n3701) );
  XNOR U4443 ( .A(n3702), .B(n3701), .Z(n5919) );
  NAND U4444 ( .A(n[159]), .B(n5919), .Z(n4947) );
  XOR U4445 ( .A(n5919), .B(n[159]), .Z(n4945) );
  XNOR U4446 ( .A(n5903), .B(n3703), .Z(n3704) );
  NANDN U4447 ( .A(n524), .B(n3704), .Z(n3705) );
  XNOR U4448 ( .A(n3706), .B(n3705), .Z(n5905) );
  ANDN U4449 ( .B(n5905), .A(n5903), .Z(n5912) );
  XOR U4450 ( .A(n5889), .B(n3707), .Z(n3708) );
  NANDN U4451 ( .A(n524), .B(n3708), .Z(n3709) );
  XOR U4452 ( .A(n3710), .B(n3709), .Z(n5891) );
  NANDN U4453 ( .A(n[156]), .B(n5891), .Z(n4931) );
  NANDN U4454 ( .A(n5891), .B(n[156]), .Z(n5898) );
  XOR U4455 ( .A(n[154]), .B(n3711), .Z(n3712) );
  NANDN U4456 ( .A(n524), .B(n3712), .Z(n3713) );
  XNOR U4457 ( .A(n3714), .B(n3713), .Z(n5883) );
  NAND U4458 ( .A(n[154]), .B(n5883), .Z(n4920) );
  XOR U4459 ( .A(n5883), .B(n[154]), .Z(n4918) );
  XOR U4460 ( .A(n[152]), .B(n3715), .Z(n3716) );
  NANDN U4461 ( .A(n524), .B(n3716), .Z(n3717) );
  XNOR U4462 ( .A(n3718), .B(n3717), .Z(n5872) );
  NAND U4463 ( .A(n[152]), .B(n5872), .Z(n4907) );
  XOR U4464 ( .A(n[152]), .B(n5872), .Z(n4905) );
  XNOR U4465 ( .A(n[151]), .B(n3719), .Z(n3720) );
  NANDN U4466 ( .A(n524), .B(n3720), .Z(n3721) );
  XNOR U4467 ( .A(n3722), .B(n3721), .Z(n5866) );
  NAND U4468 ( .A(n[151]), .B(n5866), .Z(n4903) );
  XOR U4469 ( .A(n5866), .B(n[151]), .Z(n4901) );
  XNOR U4470 ( .A(n[150]), .B(n3723), .Z(n3724) );
  NANDN U4471 ( .A(n524), .B(n3724), .Z(n3725) );
  XNOR U4472 ( .A(n3726), .B(n3725), .Z(n5861) );
  NAND U4473 ( .A(n[150]), .B(n5861), .Z(n4899) );
  XOR U4474 ( .A(n5861), .B(n[150]), .Z(n4897) );
  XNOR U4475 ( .A(n[149]), .B(n3727), .Z(n3728) );
  NANDN U4476 ( .A(n524), .B(n3728), .Z(n3729) );
  XNOR U4477 ( .A(n3730), .B(n3729), .Z(n5854) );
  NAND U4478 ( .A(n[149]), .B(n5854), .Z(n4895) );
  XOR U4479 ( .A(n[149]), .B(n5854), .Z(n4893) );
  XOR U4480 ( .A(n[148]), .B(n3731), .Z(n3732) );
  NANDN U4481 ( .A(n524), .B(n3732), .Z(n3733) );
  XNOR U4482 ( .A(n3734), .B(n3733), .Z(n5838) );
  NAND U4483 ( .A(n[148]), .B(n5838), .Z(n4891) );
  XOR U4484 ( .A(n5838), .B(n[148]), .Z(n4889) );
  XOR U4485 ( .A(n3739), .B(n3735), .Z(n3736) );
  NANDN U4486 ( .A(n524), .B(n3736), .Z(n3737) );
  XNOR U4487 ( .A(n3738), .B(n3737), .Z(n5832) );
  NANDN U4488 ( .A(n3739), .B(n5832), .Z(n4887) );
  XNOR U4489 ( .A(n5832), .B(n3739), .Z(n4885) );
  XOR U4490 ( .A(n[146]), .B(n3740), .Z(n3741) );
  NANDN U4491 ( .A(n524), .B(n3741), .Z(n3742) );
  XNOR U4492 ( .A(n3743), .B(n3742), .Z(n5826) );
  NAND U4493 ( .A(n[146]), .B(n5826), .Z(n4883) );
  XOR U4494 ( .A(n[146]), .B(n5826), .Z(n4881) );
  XOR U4495 ( .A(n[145]), .B(n3744), .Z(n3745) );
  NANDN U4496 ( .A(n524), .B(n3745), .Z(n3746) );
  XNOR U4497 ( .A(n3747), .B(n3746), .Z(n5820) );
  NAND U4498 ( .A(n[145]), .B(n5820), .Z(n4879) );
  XOR U4499 ( .A(n5820), .B(n[145]), .Z(n4877) );
  XOR U4500 ( .A(n3752), .B(n3748), .Z(n3749) );
  NANDN U4501 ( .A(n524), .B(n3749), .Z(n3750) );
  XNOR U4502 ( .A(n3751), .B(n3750), .Z(n5813) );
  NANDN U4503 ( .A(n3752), .B(n5813), .Z(n4875) );
  XNOR U4504 ( .A(n5813), .B(n3752), .Z(n4873) );
  XNOR U4505 ( .A(n[143]), .B(n3753), .Z(n3754) );
  NANDN U4506 ( .A(n524), .B(n3754), .Z(n3755) );
  XNOR U4507 ( .A(n3756), .B(n3755), .Z(n5806) );
  NAND U4508 ( .A(n[143]), .B(n5806), .Z(n4871) );
  XOR U4509 ( .A(n[143]), .B(n5806), .Z(n4869) );
  XNOR U4510 ( .A(n[142]), .B(n3757), .Z(n3758) );
  NANDN U4511 ( .A(n524), .B(n3758), .Z(n3759) );
  XNOR U4512 ( .A(n3760), .B(n3759), .Z(n5800) );
  NAND U4513 ( .A(n[142]), .B(n5800), .Z(n4867) );
  XOR U4514 ( .A(n5800), .B(n[142]), .Z(n4865) );
  XOR U4515 ( .A(n[141]), .B(n3761), .Z(n3762) );
  NANDN U4516 ( .A(n524), .B(n3762), .Z(n3763) );
  XOR U4517 ( .A(n3764), .B(n3763), .Z(n5796) );
  NANDN U4518 ( .A(n5796), .B(n[141]), .Z(n4863) );
  XNOR U4519 ( .A(n[141]), .B(n5796), .Z(n4861) );
  XOR U4520 ( .A(n3769), .B(n3765), .Z(n3766) );
  NANDN U4521 ( .A(n524), .B(n3766), .Z(n3767) );
  XNOR U4522 ( .A(n3768), .B(n3767), .Z(n5789) );
  NANDN U4523 ( .A(n3769), .B(n5789), .Z(n4859) );
  XNOR U4524 ( .A(n5789), .B(n3769), .Z(n4857) );
  XNOR U4525 ( .A(n[139]), .B(n3770), .Z(n3771) );
  NANDN U4526 ( .A(n524), .B(n3771), .Z(n3772) );
  XNOR U4527 ( .A(n3773), .B(n3772), .Z(n5783) );
  NAND U4528 ( .A(n[139]), .B(n5783), .Z(n4855) );
  XOR U4529 ( .A(n5783), .B(n[139]), .Z(n4853) );
  XNOR U4530 ( .A(n[138]), .B(n3774), .Z(n3775) );
  NANDN U4531 ( .A(n524), .B(n3775), .Z(n3776) );
  XNOR U4532 ( .A(n3777), .B(n3776), .Z(n5776) );
  NAND U4533 ( .A(n[138]), .B(n5776), .Z(n4851) );
  XOR U4534 ( .A(n[138]), .B(n5776), .Z(n4849) );
  XNOR U4535 ( .A(n[137]), .B(n3778), .Z(n3779) );
  NANDN U4536 ( .A(n524), .B(n3779), .Z(n3780) );
  XNOR U4537 ( .A(n3781), .B(n3780), .Z(n5770) );
  NAND U4538 ( .A(n[137]), .B(n5770), .Z(n4847) );
  XOR U4539 ( .A(n5770), .B(n[137]), .Z(n4845) );
  XNOR U4540 ( .A(n[136]), .B(n3782), .Z(n3783) );
  NANDN U4541 ( .A(n524), .B(n3783), .Z(n3784) );
  XNOR U4542 ( .A(n3785), .B(n3784), .Z(n5764) );
  NAND U4543 ( .A(n[136]), .B(n5764), .Z(n4843) );
  XOR U4544 ( .A(n[136]), .B(n5764), .Z(n4841) );
  XNOR U4545 ( .A(n[135]), .B(n3786), .Z(n3787) );
  NANDN U4546 ( .A(n524), .B(n3787), .Z(n3788) );
  XNOR U4547 ( .A(n3789), .B(n3788), .Z(n5758) );
  NAND U4548 ( .A(n[135]), .B(n5758), .Z(n4839) );
  XOR U4549 ( .A(n5758), .B(n[135]), .Z(n4837) );
  XOR U4550 ( .A(n[134]), .B(n3790), .Z(n3791) );
  NANDN U4551 ( .A(n524), .B(n3791), .Z(n3792) );
  XNOR U4552 ( .A(n3793), .B(n3792), .Z(n5752) );
  NAND U4553 ( .A(n[134]), .B(n5752), .Z(n4835) );
  XOR U4554 ( .A(n[134]), .B(n5752), .Z(n4833) );
  XOR U4555 ( .A(n3798), .B(n3794), .Z(n3795) );
  NANDN U4556 ( .A(n524), .B(n3795), .Z(n3796) );
  XNOR U4557 ( .A(n3797), .B(n3796), .Z(n5746) );
  NANDN U4558 ( .A(n3798), .B(n5746), .Z(n4831) );
  XNOR U4559 ( .A(n5746), .B(n3798), .Z(n4829) );
  XOR U4560 ( .A(n[132]), .B(n3799), .Z(n3800) );
  NANDN U4561 ( .A(n524), .B(n3800), .Z(n3801) );
  XNOR U4562 ( .A(n3802), .B(n3801), .Z(n5739) );
  NAND U4563 ( .A(n[132]), .B(n5739), .Z(n4827) );
  XOR U4564 ( .A(n[132]), .B(n5739), .Z(n4825) );
  XOR U4565 ( .A(n[131]), .B(n3803), .Z(n3804) );
  NANDN U4566 ( .A(n524), .B(n3804), .Z(n3805) );
  XNOR U4567 ( .A(n3806), .B(n3805), .Z(n5733) );
  NAND U4568 ( .A(n[131]), .B(n5733), .Z(n4823) );
  XOR U4569 ( .A(n5733), .B(n[131]), .Z(n4821) );
  XOR U4570 ( .A(n3811), .B(n3807), .Z(n3808) );
  NANDN U4571 ( .A(n524), .B(n3808), .Z(n3809) );
  XNOR U4572 ( .A(n3810), .B(n3809), .Z(n5727) );
  NANDN U4573 ( .A(n3811), .B(n5727), .Z(n4819) );
  XNOR U4574 ( .A(n3811), .B(n5727), .Z(n4817) );
  XOR U4575 ( .A(n[129]), .B(n3812), .Z(n3813) );
  NANDN U4576 ( .A(n524), .B(n3813), .Z(n3814) );
  XNOR U4577 ( .A(n3815), .B(n3814), .Z(n5720) );
  NAND U4578 ( .A(n[129]), .B(n5720), .Z(n4815) );
  XOR U4579 ( .A(n5720), .B(n[129]), .Z(n4813) );
  XNOR U4580 ( .A(n[128]), .B(n3816), .Z(n3817) );
  NANDN U4581 ( .A(n524), .B(n3817), .Z(n3818) );
  XNOR U4582 ( .A(n3819), .B(n3818), .Z(n5710) );
  NAND U4583 ( .A(n[128]), .B(n5710), .Z(n4811) );
  XOR U4584 ( .A(n5710), .B(n[128]), .Z(n4809) );
  XNOR U4585 ( .A(n[127]), .B(n3820), .Z(n3821) );
  NANDN U4586 ( .A(n524), .B(n3821), .Z(n3822) );
  XNOR U4587 ( .A(n3823), .B(n3822), .Z(n5704) );
  NAND U4588 ( .A(n[127]), .B(n5704), .Z(n4807) );
  XOR U4589 ( .A(n[127]), .B(n5704), .Z(n4805) );
  XOR U4590 ( .A(n[126]), .B(n3824), .Z(n3825) );
  NANDN U4591 ( .A(n524), .B(n3825), .Z(n3826) );
  XNOR U4592 ( .A(n3827), .B(n3826), .Z(n5697) );
  NAND U4593 ( .A(n[126]), .B(n5697), .Z(n4803) );
  XOR U4594 ( .A(n5697), .B(n[126]), .Z(n4801) );
  XOR U4595 ( .A(n3832), .B(n3828), .Z(n3829) );
  NANDN U4596 ( .A(n524), .B(n3829), .Z(n3830) );
  XNOR U4597 ( .A(n3831), .B(n3830), .Z(n5694) );
  NANDN U4598 ( .A(n3832), .B(n5694), .Z(n4799) );
  XNOR U4599 ( .A(n3832), .B(n5694), .Z(n4797) );
  XOR U4600 ( .A(n[124]), .B(n3833), .Z(n3834) );
  NANDN U4601 ( .A(n524), .B(n3834), .Z(n3835) );
  XNOR U4602 ( .A(n3836), .B(n3835), .Z(n5687) );
  NAND U4603 ( .A(n[124]), .B(n5687), .Z(n4795) );
  XOR U4604 ( .A(n5687), .B(n[124]), .Z(n4793) );
  XNOR U4605 ( .A(n3841), .B(n3837), .Z(n3838) );
  NANDN U4606 ( .A(n524), .B(n3838), .Z(n3839) );
  XNOR U4607 ( .A(n3840), .B(n3839), .Z(n5681) );
  NANDN U4608 ( .A(n3841), .B(n5681), .Z(n4791) );
  XNOR U4609 ( .A(n3841), .B(n5681), .Z(n4789) );
  XNOR U4610 ( .A(n3846), .B(n3842), .Z(n3843) );
  NANDN U4611 ( .A(n524), .B(n3843), .Z(n3844) );
  XNOR U4612 ( .A(n3845), .B(n3844), .Z(n5675) );
  NANDN U4613 ( .A(n3846), .B(n5675), .Z(n4787) );
  XNOR U4614 ( .A(n5675), .B(n3846), .Z(n4785) );
  XNOR U4615 ( .A(n3851), .B(n3847), .Z(n3848) );
  NANDN U4616 ( .A(n524), .B(n3848), .Z(n3849) );
  XNOR U4617 ( .A(n3850), .B(n3849), .Z(n5669) );
  NANDN U4618 ( .A(n3851), .B(n5669), .Z(n4783) );
  XNOR U4619 ( .A(n3851), .B(n5669), .Z(n4781) );
  XNOR U4620 ( .A(n3856), .B(n3852), .Z(n3853) );
  NANDN U4621 ( .A(n524), .B(n3853), .Z(n3854) );
  XNOR U4622 ( .A(n3855), .B(n3854), .Z(n5666) );
  NANDN U4623 ( .A(n3856), .B(n5666), .Z(n4779) );
  XNOR U4624 ( .A(n5666), .B(n3856), .Z(n4777) );
  XOR U4625 ( .A(n[119]), .B(n3857), .Z(n3858) );
  NANDN U4626 ( .A(n524), .B(n3858), .Z(n3859) );
  XNOR U4627 ( .A(n3860), .B(n3859), .Z(n5659) );
  NAND U4628 ( .A(n[119]), .B(n5659), .Z(n4775) );
  XOR U4629 ( .A(n5659), .B(n[119]), .Z(n4773) );
  XNOR U4630 ( .A(n5648), .B(n3861), .Z(n3862) );
  NANDN U4631 ( .A(n524), .B(n3862), .Z(n3863) );
  XNOR U4632 ( .A(n3864), .B(n3863), .Z(n5649) );
  NANDN U4633 ( .A(n5648), .B(n5649), .Z(n4771) );
  XNOR U4634 ( .A(n5648), .B(n5649), .Z(n4769) );
  XNOR U4635 ( .A(n3869), .B(n3865), .Z(n3866) );
  NANDN U4636 ( .A(n524), .B(n3866), .Z(n3867) );
  XNOR U4637 ( .A(n3868), .B(n3867), .Z(n5641) );
  NANDN U4638 ( .A(n3869), .B(n5641), .Z(n4767) );
  XNOR U4639 ( .A(n5641), .B(n3869), .Z(n4765) );
  XNOR U4640 ( .A(n5633), .B(n3870), .Z(n3871) );
  NANDN U4641 ( .A(n524), .B(n3871), .Z(n3872) );
  XNOR U4642 ( .A(n3873), .B(n3872), .Z(n5634) );
  NANDN U4643 ( .A(n5633), .B(n5634), .Z(n4763) );
  XNOR U4644 ( .A(n5633), .B(n5634), .Z(n4761) );
  XNOR U4645 ( .A(n3878), .B(n3874), .Z(n3875) );
  NANDN U4646 ( .A(n524), .B(n3875), .Z(n3876) );
  XNOR U4647 ( .A(n3877), .B(n3876), .Z(n5627) );
  NANDN U4648 ( .A(n3878), .B(n5627), .Z(n4759) );
  XNOR U4649 ( .A(n5627), .B(n3878), .Z(n4757) );
  XNOR U4650 ( .A(n3883), .B(n3879), .Z(n3880) );
  NANDN U4651 ( .A(n524), .B(n3880), .Z(n3881) );
  XNOR U4652 ( .A(n3882), .B(n3881), .Z(n5625) );
  NANDN U4653 ( .A(n3883), .B(n5625), .Z(n4755) );
  XNOR U4654 ( .A(n3883), .B(n5625), .Z(n4753) );
  XNOR U4655 ( .A(n3888), .B(n3884), .Z(n3885) );
  NANDN U4656 ( .A(n524), .B(n3885), .Z(n3886) );
  XNOR U4657 ( .A(n3887), .B(n3886), .Z(n5621) );
  NANDN U4658 ( .A(n3888), .B(n5621), .Z(n4751) );
  XNOR U4659 ( .A(n5621), .B(n3888), .Z(n4749) );
  XNOR U4660 ( .A(n3893), .B(n3889), .Z(n3890) );
  NANDN U4661 ( .A(n524), .B(n3890), .Z(n3891) );
  XNOR U4662 ( .A(n3892), .B(n3891), .Z(n5616) );
  NANDN U4663 ( .A(n3893), .B(n5616), .Z(n4747) );
  XNOR U4664 ( .A(n5616), .B(n3893), .Z(n4745) );
  XNOR U4665 ( .A(n3898), .B(n3894), .Z(n3895) );
  NANDN U4666 ( .A(n524), .B(n3895), .Z(n3896) );
  XNOR U4667 ( .A(n3897), .B(n3896), .Z(n5612) );
  NANDN U4668 ( .A(n3898), .B(n5612), .Z(n4743) );
  XNOR U4669 ( .A(n5612), .B(n3898), .Z(n4741) );
  XNOR U4670 ( .A(n3903), .B(n3899), .Z(n3900) );
  NANDN U4671 ( .A(n524), .B(n3900), .Z(n3901) );
  XNOR U4672 ( .A(n3902), .B(n3901), .Z(n5605) );
  NANDN U4673 ( .A(n3903), .B(n5605), .Z(n4739) );
  XNOR U4674 ( .A(n3903), .B(n5605), .Z(n4737) );
  XOR U4675 ( .A(n[109]), .B(n3904), .Z(n3905) );
  NANDN U4676 ( .A(n524), .B(n3905), .Z(n3906) );
  XNOR U4677 ( .A(n3907), .B(n3906), .Z(n5599) );
  NAND U4678 ( .A(n[109]), .B(n5599), .Z(n4735) );
  XOR U4679 ( .A(n5599), .B(n[109]), .Z(n4733) );
  XOR U4680 ( .A(n3912), .B(n3908), .Z(n3909) );
  NANDN U4681 ( .A(n524), .B(n3909), .Z(n3910) );
  XNOR U4682 ( .A(n3911), .B(n3910), .Z(n5589) );
  NANDN U4683 ( .A(n3912), .B(n5589), .Z(n4731) );
  XNOR U4684 ( .A(n3912), .B(n5589), .Z(n4729) );
  XNOR U4685 ( .A(n[107]), .B(n3913), .Z(n3914) );
  NANDN U4686 ( .A(n524), .B(n3914), .Z(n3915) );
  XNOR U4687 ( .A(n3916), .B(n3915), .Z(n5582) );
  NAND U4688 ( .A(n[107]), .B(n5582), .Z(n4727) );
  XOR U4689 ( .A(n5582), .B(n[107]), .Z(n4725) );
  XNOR U4690 ( .A(n[106]), .B(n3917), .Z(n3918) );
  NANDN U4691 ( .A(n524), .B(n3918), .Z(n3919) );
  XNOR U4692 ( .A(n3920), .B(n3919), .Z(n5577) );
  NAND U4693 ( .A(n[106]), .B(n5577), .Z(n4723) );
  XOR U4694 ( .A(n5577), .B(n[106]), .Z(n4721) );
  XNOR U4695 ( .A(n[105]), .B(n3921), .Z(n3922) );
  NANDN U4696 ( .A(n524), .B(n3922), .Z(n3923) );
  XNOR U4697 ( .A(n3924), .B(n3923), .Z(n5570) );
  NAND U4698 ( .A(n[105]), .B(n5570), .Z(n4719) );
  XOR U4699 ( .A(n[105]), .B(n5570), .Z(n4717) );
  XOR U4700 ( .A(n[104]), .B(n3925), .Z(n3926) );
  NANDN U4701 ( .A(n524), .B(n3926), .Z(n3927) );
  XNOR U4702 ( .A(n3928), .B(n3927), .Z(n5567) );
  NAND U4703 ( .A(n[104]), .B(n5567), .Z(n4715) );
  XOR U4704 ( .A(n5567), .B(n[104]), .Z(n4713) );
  XOR U4705 ( .A(n3933), .B(n3929), .Z(n3930) );
  NANDN U4706 ( .A(n524), .B(n3930), .Z(n3931) );
  XNOR U4707 ( .A(n3932), .B(n3931), .Z(n5561) );
  NANDN U4708 ( .A(n3933), .B(n5561), .Z(n4711) );
  XNOR U4709 ( .A(n5561), .B(n3933), .Z(n4709) );
  XOR U4710 ( .A(n[102]), .B(n3934), .Z(n3935) );
  NANDN U4711 ( .A(n524), .B(n3935), .Z(n3936) );
  XNOR U4712 ( .A(n3937), .B(n3936), .Z(n5554) );
  NAND U4713 ( .A(n[102]), .B(n5554), .Z(n4707) );
  XOR U4714 ( .A(n[102]), .B(n5554), .Z(n4705) );
  XOR U4715 ( .A(n3942), .B(n3938), .Z(n3939) );
  NANDN U4716 ( .A(n524), .B(n3939), .Z(n3940) );
  XNOR U4717 ( .A(n3941), .B(n3940), .Z(n5551) );
  NANDN U4718 ( .A(n3942), .B(n5551), .Z(n4703) );
  XNOR U4719 ( .A(n5551), .B(n3942), .Z(n4701) );
  XNOR U4720 ( .A(n[100]), .B(n3943), .Z(n3944) );
  NANDN U4721 ( .A(n524), .B(n3944), .Z(n3945) );
  XNOR U4722 ( .A(n3946), .B(n3945), .Z(n5544) );
  NAND U4723 ( .A(n[100]), .B(n5544), .Z(n4699) );
  XOR U4724 ( .A(n[100]), .B(n5544), .Z(n4697) );
  XOR U4725 ( .A(n5344), .B(n3947), .Z(n3948) );
  NANDN U4726 ( .A(n524), .B(n3948), .Z(n3949) );
  XNOR U4727 ( .A(n3950), .B(n3949), .Z(n6866) );
  NANDN U4728 ( .A(n5344), .B(n6866), .Z(n4695) );
  XNOR U4729 ( .A(n6866), .B(n5344), .Z(n4693) );
  XNOR U4730 ( .A(n[98]), .B(n3951), .Z(n3952) );
  NANDN U4731 ( .A(n524), .B(n3952), .Z(n3953) );
  XNOR U4732 ( .A(n3954), .B(n3953), .Z(n5347) );
  NAND U4733 ( .A(n[98]), .B(n5347), .Z(n4691) );
  XOR U4734 ( .A(n[98]), .B(n5347), .Z(n4689) );
  XOR U4735 ( .A(n[97]), .B(n3955), .Z(n3956) );
  NANDN U4736 ( .A(n524), .B(n3956), .Z(n3957) );
  XNOR U4737 ( .A(n3958), .B(n3957), .Z(n6860) );
  NAND U4738 ( .A(n[97]), .B(n6860), .Z(n4687) );
  XOR U4739 ( .A(n6860), .B(n[97]), .Z(n4685) );
  XNOR U4740 ( .A(n3963), .B(n3959), .Z(n3960) );
  NANDN U4741 ( .A(n524), .B(n3960), .Z(n3961) );
  XNOR U4742 ( .A(n3962), .B(n3961), .Z(n5535) );
  NANDN U4743 ( .A(n3963), .B(n5535), .Z(n4683) );
  XNOR U4744 ( .A(n3963), .B(n5535), .Z(n4681) );
  XNOR U4745 ( .A(n5529), .B(n3964), .Z(n3965) );
  NANDN U4746 ( .A(n524), .B(n3965), .Z(n3966) );
  XNOR U4747 ( .A(n3967), .B(n3966), .Z(n5531) );
  XOR U4748 ( .A(n[95]), .B(n5531), .Z(n4677) );
  XNOR U4749 ( .A(n3969), .B(n3968), .Z(n3970) );
  NANDN U4750 ( .A(n524), .B(n3970), .Z(n3971) );
  XNOR U4751 ( .A(n3972), .B(n3971), .Z(n5350) );
  XNOR U4752 ( .A(n3974), .B(n3973), .Z(n3975) );
  NANDN U4753 ( .A(n524), .B(n3975), .Z(n3976) );
  XNOR U4754 ( .A(n3977), .B(n3976), .Z(n5352) );
  OR U4755 ( .A(n5352), .B(n[93]), .Z(n4671) );
  XOR U4756 ( .A(n5352), .B(n[93]), .Z(n4669) );
  XNOR U4757 ( .A(n[91]), .B(n3978), .Z(n3979) );
  NANDN U4758 ( .A(n524), .B(n3979), .Z(n3980) );
  XNOR U4759 ( .A(n3981), .B(n3980), .Z(n5359) );
  NAND U4760 ( .A(n[91]), .B(n5359), .Z(n4659) );
  XOR U4761 ( .A(n5359), .B(n[91]), .Z(n4657) );
  XOR U4762 ( .A(n[90]), .B(n3982), .Z(n3983) );
  NANDN U4763 ( .A(n524), .B(n3983), .Z(n3984) );
  XNOR U4764 ( .A(n3985), .B(n3984), .Z(n5361) );
  NAND U4765 ( .A(n[90]), .B(n5361), .Z(n4655) );
  XOR U4766 ( .A(n[90]), .B(n5361), .Z(n4653) );
  XNOR U4767 ( .A(n[89]), .B(n3986), .Z(n3987) );
  NANDN U4768 ( .A(n524), .B(n3987), .Z(n3988) );
  XNOR U4769 ( .A(n3989), .B(n3988), .Z(n5364) );
  NAND U4770 ( .A(n[89]), .B(n5364), .Z(n4651) );
  XOR U4771 ( .A(n5364), .B(n[89]), .Z(n4649) );
  XOR U4772 ( .A(n[88]), .B(n3990), .Z(n3991) );
  NANDN U4773 ( .A(n524), .B(n3991), .Z(n3992) );
  XNOR U4774 ( .A(n3993), .B(n3992), .Z(n5514) );
  NAND U4775 ( .A(n[88]), .B(n5514), .Z(n4647) );
  XOR U4776 ( .A(n[88]), .B(n5514), .Z(n4645) );
  XOR U4777 ( .A(n3998), .B(n3994), .Z(n3995) );
  NANDN U4778 ( .A(n524), .B(n3995), .Z(n3996) );
  XNOR U4779 ( .A(n3997), .B(n3996), .Z(n5366) );
  NANDN U4780 ( .A(n3998), .B(n5366), .Z(n4643) );
  XNOR U4781 ( .A(n5366), .B(n3998), .Z(n4641) );
  XOR U4782 ( .A(n[86]), .B(n3999), .Z(n4000) );
  NANDN U4783 ( .A(n524), .B(n4000), .Z(n4001) );
  XNOR U4784 ( .A(n4002), .B(n4001), .Z(n5368) );
  NAND U4785 ( .A(n[86]), .B(n5368), .Z(n4639) );
  XOR U4786 ( .A(n[86]), .B(n5368), .Z(n4637) );
  XOR U4787 ( .A(n5504), .B(n4003), .Z(n4004) );
  NANDN U4788 ( .A(n524), .B(n4004), .Z(n4005) );
  XNOR U4789 ( .A(n4006), .B(n4005), .Z(n5506) );
  NANDN U4790 ( .A(n5504), .B(n5506), .Z(n4635) );
  XNOR U4791 ( .A(n5506), .B(n5504), .Z(n4633) );
  XNOR U4792 ( .A(n[84]), .B(n4007), .Z(n4008) );
  NANDN U4793 ( .A(n524), .B(n4008), .Z(n4009) );
  XNOR U4794 ( .A(n4010), .B(n4009), .Z(n5370) );
  NAND U4795 ( .A(n[84]), .B(n5370), .Z(n4631) );
  XOR U4796 ( .A(n[84]), .B(n5370), .Z(n4629) );
  XNOR U4797 ( .A(n[83]), .B(n4011), .Z(n4012) );
  NANDN U4798 ( .A(n524), .B(n4012), .Z(n4013) );
  XNOR U4799 ( .A(n4014), .B(n4013), .Z(n5372) );
  NAND U4800 ( .A(n[83]), .B(n5372), .Z(n4627) );
  XOR U4801 ( .A(n5372), .B(n[83]), .Z(n4625) );
  XOR U4802 ( .A(n[82]), .B(n4015), .Z(n4016) );
  NANDN U4803 ( .A(n524), .B(n4016), .Z(n4017) );
  XNOR U4804 ( .A(n4018), .B(n4017), .Z(n5375) );
  NAND U4805 ( .A(n[82]), .B(n5375), .Z(n4623) );
  XOR U4806 ( .A(n5375), .B(n[82]), .Z(n4621) );
  XNOR U4807 ( .A(n4023), .B(n4019), .Z(n4020) );
  NANDN U4808 ( .A(n524), .B(n4020), .Z(n4021) );
  XNOR U4809 ( .A(n4022), .B(n4021), .Z(n5377) );
  NANDN U4810 ( .A(n4023), .B(n5377), .Z(n4619) );
  XNOR U4811 ( .A(n4023), .B(n5377), .Z(n4617) );
  XOR U4812 ( .A(n4028), .B(n4024), .Z(n4025) );
  NANDN U4813 ( .A(n524), .B(n4025), .Z(n4026) );
  XNOR U4814 ( .A(n4027), .B(n4026), .Z(n5379) );
  NANDN U4815 ( .A(n4028), .B(n5379), .Z(n4615) );
  XNOR U4816 ( .A(n5379), .B(n4028), .Z(n4613) );
  XNOR U4817 ( .A(n[79]), .B(n4029), .Z(n4030) );
  NANDN U4818 ( .A(n524), .B(n4030), .Z(n4031) );
  XNOR U4819 ( .A(n4032), .B(n4031), .Z(n6810) );
  NAND U4820 ( .A(n[79]), .B(n6810), .Z(n4611) );
  XOR U4821 ( .A(n6810), .B(n[79]), .Z(n4609) );
  XOR U4822 ( .A(n[78]), .B(n4033), .Z(n4034) );
  NANDN U4823 ( .A(n524), .B(n4034), .Z(n4035) );
  XNOR U4824 ( .A(n4036), .B(n4035), .Z(n5381) );
  NAND U4825 ( .A(n[78]), .B(n5381), .Z(n4607) );
  XOR U4826 ( .A(n[78]), .B(n5381), .Z(n4605) );
  XOR U4827 ( .A(n4041), .B(n4037), .Z(n4038) );
  NANDN U4828 ( .A(n524), .B(n4038), .Z(n4039) );
  XNOR U4829 ( .A(n4040), .B(n4039), .Z(n6804) );
  NANDN U4830 ( .A(n4041), .B(n6804), .Z(n4603) );
  XNOR U4831 ( .A(n6804), .B(n4041), .Z(n4601) );
  XNOR U4832 ( .A(n[76]), .B(n4042), .Z(n4043) );
  NANDN U4833 ( .A(n524), .B(n4043), .Z(n4044) );
  XNOR U4834 ( .A(n4045), .B(n4044), .Z(n5383) );
  NAND U4835 ( .A(n[76]), .B(n5383), .Z(n4599) );
  XOR U4836 ( .A(n5383), .B(n[76]), .Z(n4597) );
  XNOR U4837 ( .A(n[75]), .B(n4046), .Z(n4047) );
  NANDN U4838 ( .A(n524), .B(n4047), .Z(n4048) );
  XNOR U4839 ( .A(n4049), .B(n4048), .Z(n5487) );
  NAND U4840 ( .A(n[75]), .B(n5487), .Z(n4595) );
  XOR U4841 ( .A(n[75]), .B(n5487), .Z(n4593) );
  XNOR U4842 ( .A(n[74]), .B(n4050), .Z(n4051) );
  NANDN U4843 ( .A(n524), .B(n4051), .Z(n4052) );
  XNOR U4844 ( .A(n4053), .B(n4052), .Z(n5386) );
  NAND U4845 ( .A(n[74]), .B(n5386), .Z(n4591) );
  XOR U4846 ( .A(n5386), .B(n[74]), .Z(n4589) );
  XNOR U4847 ( .A(n[73]), .B(n4054), .Z(n4055) );
  NANDN U4848 ( .A(n524), .B(n4055), .Z(n4056) );
  XNOR U4849 ( .A(n4057), .B(n4056), .Z(n5388) );
  NAND U4850 ( .A(n[73]), .B(n5388), .Z(n4587) );
  XOR U4851 ( .A(n[73]), .B(n5388), .Z(n4585) );
  XNOR U4852 ( .A(n[72]), .B(n4058), .Z(n4059) );
  NANDN U4853 ( .A(n524), .B(n4059), .Z(n4060) );
  XNOR U4854 ( .A(n4061), .B(n4060), .Z(n5479) );
  NAND U4855 ( .A(n[72]), .B(n5479), .Z(n4583) );
  XOR U4856 ( .A(n5479), .B(n[72]), .Z(n4581) );
  XNOR U4857 ( .A(n5390), .B(n4062), .Z(n4063) );
  NANDN U4858 ( .A(n524), .B(n4063), .Z(n4064) );
  XOR U4859 ( .A(n4065), .B(n4064), .Z(n5475) );
  NANDN U4860 ( .A(n5475), .B(n[71]), .Z(n4579) );
  XOR U4861 ( .A(n5469), .B(n4066), .Z(n4067) );
  NANDN U4862 ( .A(n524), .B(n4067), .Z(n4068) );
  XOR U4863 ( .A(n4069), .B(n4068), .Z(n4573) );
  IV U4864 ( .A(n4573), .Z(n5471) );
  XNOR U4865 ( .A(n[69]), .B(n4070), .Z(n4071) );
  NANDN U4866 ( .A(n524), .B(n4071), .Z(n4072) );
  XNOR U4867 ( .A(n4073), .B(n4072), .Z(n5393) );
  NAND U4868 ( .A(n[69]), .B(n5393), .Z(n4570) );
  XOR U4869 ( .A(n5393), .B(n[69]), .Z(n4568) );
  XOR U4870 ( .A(n4078), .B(n4074), .Z(n4075) );
  NANDN U4871 ( .A(n524), .B(n4075), .Z(n4076) );
  XNOR U4872 ( .A(n4077), .B(n4076), .Z(n6774) );
  NANDN U4873 ( .A(n4078), .B(n6774), .Z(n4566) );
  XNOR U4874 ( .A(n4078), .B(n6774), .Z(n4564) );
  XNOR U4875 ( .A(n[67]), .B(n4079), .Z(n4080) );
  NANDN U4876 ( .A(n524), .B(n4080), .Z(n4081) );
  XNOR U4877 ( .A(n4082), .B(n4081), .Z(n5396) );
  NAND U4878 ( .A(n[67]), .B(n5396), .Z(n4562) );
  XOR U4879 ( .A(n5396), .B(n[67]), .Z(n4560) );
  XOR U4880 ( .A(n[66]), .B(n4083), .Z(n4084) );
  NANDN U4881 ( .A(n524), .B(n4084), .Z(n4085) );
  XNOR U4882 ( .A(n4086), .B(n4085), .Z(n6768) );
  NAND U4883 ( .A(n[66]), .B(n6768), .Z(n4558) );
  XOR U4884 ( .A(n6768), .B(n[66]), .Z(n4556) );
  XOR U4885 ( .A(n4091), .B(n4087), .Z(n4088) );
  NANDN U4886 ( .A(n524), .B(n4088), .Z(n4089) );
  XNOR U4887 ( .A(n4090), .B(n4089), .Z(n5398) );
  NANDN U4888 ( .A(n4091), .B(n5398), .Z(n4554) );
  XNOR U4889 ( .A(n4091), .B(n5398), .Z(n4552) );
  XOR U4890 ( .A(n5399), .B(n4092), .Z(n4093) );
  NANDN U4891 ( .A(n524), .B(n4093), .Z(n4094) );
  XOR U4892 ( .A(n4095), .B(n4094), .Z(n5402) );
  NANDN U4893 ( .A(n5399), .B(n5402), .Z(n4550) );
  XNOR U4894 ( .A(n5402), .B(n5399), .Z(n4548) );
  XOR U4895 ( .A(n[63]), .B(n4096), .Z(n4097) );
  NANDN U4896 ( .A(n524), .B(n4097), .Z(n4098) );
  XNOR U4897 ( .A(n4099), .B(n4098), .Z(n5458) );
  NAND U4898 ( .A(n[63]), .B(n5458), .Z(n4546) );
  XOR U4899 ( .A(n[63]), .B(n5458), .Z(n4544) );
  XNOR U4900 ( .A(n[62]), .B(n4100), .Z(n4101) );
  NANDN U4901 ( .A(n524), .B(n4101), .Z(n4102) );
  XOR U4902 ( .A(n4103), .B(n4102), .Z(n5404) );
  NAND U4903 ( .A(n[62]), .B(n5404), .Z(n4542) );
  XOR U4904 ( .A(n5404), .B(n[62]), .Z(n4540) );
  XNOR U4905 ( .A(n4108), .B(n4104), .Z(n4105) );
  NANDN U4906 ( .A(n524), .B(n4105), .Z(n4106) );
  XOR U4907 ( .A(n4107), .B(n4106), .Z(n5406) );
  NANDN U4908 ( .A(n4108), .B(n5406), .Z(n4538) );
  XNOR U4909 ( .A(n4108), .B(n5406), .Z(n4536) );
  XNOR U4910 ( .A(n4113), .B(n4109), .Z(n4110) );
  NANDN U4911 ( .A(n524), .B(n4110), .Z(n4111) );
  XNOR U4912 ( .A(n4112), .B(n4111), .Z(n5408) );
  NANDN U4913 ( .A(n4113), .B(n5408), .Z(n4534) );
  XNOR U4914 ( .A(n5408), .B(n4113), .Z(n4532) );
  XNOR U4915 ( .A(n4118), .B(n4114), .Z(n4115) );
  NANDN U4916 ( .A(n524), .B(n4115), .Z(n4116) );
  XOR U4917 ( .A(n4117), .B(n4116), .Z(n5410) );
  NANDN U4918 ( .A(n4118), .B(n5410), .Z(n4530) );
  XNOR U4919 ( .A(n4118), .B(n5410), .Z(n4528) );
  XNOR U4920 ( .A(n5411), .B(n4119), .Z(n4120) );
  NANDN U4921 ( .A(n524), .B(n4120), .Z(n4121) );
  XOR U4922 ( .A(n4122), .B(n4121), .Z(n5414) );
  NANDN U4923 ( .A(n5411), .B(n5414), .Z(n4526) );
  XNOR U4924 ( .A(n5414), .B(n5411), .Z(n4524) );
  XNOR U4925 ( .A(n[57]), .B(n4123), .Z(n4124) );
  NANDN U4926 ( .A(n524), .B(n4124), .Z(n4125) );
  XNOR U4927 ( .A(n4126), .B(n4125), .Z(n5417) );
  NAND U4928 ( .A(n[57]), .B(n5417), .Z(n4522) );
  XOR U4929 ( .A(n5417), .B(n[57]), .Z(n4520) );
  XOR U4930 ( .A(n4131), .B(n4127), .Z(n4128) );
  NANDN U4931 ( .A(n524), .B(n4128), .Z(n4129) );
  XNOR U4932 ( .A(n4130), .B(n4129), .Z(n5419) );
  NANDN U4933 ( .A(n4131), .B(n5419), .Z(n4518) );
  XNOR U4934 ( .A(n4131), .B(n5419), .Z(n4516) );
  XNOR U4935 ( .A(n[55]), .B(n4132), .Z(n4133) );
  NANDN U4936 ( .A(n524), .B(n4133), .Z(n4134) );
  XNOR U4937 ( .A(n4135), .B(n4134), .Z(n5421) );
  NAND U4938 ( .A(n[55]), .B(n5421), .Z(n4514) );
  XOR U4939 ( .A(n5421), .B(n[55]), .Z(n4512) );
  XNOR U4940 ( .A(n4140), .B(n4136), .Z(n4137) );
  NANDN U4941 ( .A(n524), .B(n4137), .Z(n4138) );
  XNOR U4942 ( .A(n4139), .B(n4138), .Z(n5423) );
  NANDN U4943 ( .A(n4140), .B(n5423), .Z(n4510) );
  XNOR U4944 ( .A(n4140), .B(n5423), .Z(n4508) );
  XNOR U4945 ( .A(n4145), .B(n4141), .Z(n4142) );
  NANDN U4946 ( .A(n524), .B(n4142), .Z(n4143) );
  XOR U4947 ( .A(n4144), .B(n4143), .Z(n6739) );
  NANDN U4948 ( .A(n4145), .B(n6739), .Z(n4506) );
  XNOR U4949 ( .A(n6739), .B(n4145), .Z(n4504) );
  XNOR U4950 ( .A(n[52]), .B(n4146), .Z(n4147) );
  NANDN U4951 ( .A(n524), .B(n4147), .Z(n4148) );
  XNOR U4952 ( .A(n4149), .B(n4148), .Z(n5426) );
  NAND U4953 ( .A(n5426), .B(n[52]), .Z(n4502) );
  XOR U4954 ( .A(n[52]), .B(n5426), .Z(n4500) );
  XOR U4955 ( .A(n[51]), .B(n4150), .Z(n4151) );
  NANDN U4956 ( .A(n524), .B(n4151), .Z(n4152) );
  XNOR U4957 ( .A(n4153), .B(n4152), .Z(n5428) );
  NAND U4958 ( .A(n[51]), .B(n5428), .Z(n4498) );
  XOR U4959 ( .A(n5428), .B(n[51]), .Z(n4496) );
  XOR U4960 ( .A(n[50]), .B(n4154), .Z(n4155) );
  NANDN U4961 ( .A(n524), .B(n4155), .Z(n4156) );
  XOR U4962 ( .A(n4157), .B(n4156), .Z(n6731) );
  NAND U4963 ( .A(n[50]), .B(n6731), .Z(n4494) );
  XOR U4964 ( .A(n[50]), .B(n6731), .Z(n4492) );
  IV U4965 ( .A(n[49]), .Z(n4162) );
  XNOR U4966 ( .A(n4162), .B(n4158), .Z(n4159) );
  NANDN U4967 ( .A(n524), .B(n4159), .Z(n4160) );
  XNOR U4968 ( .A(n4161), .B(n4160), .Z(n6723) );
  NANDN U4969 ( .A(n4162), .B(n6723), .Z(n4490) );
  XNOR U4970 ( .A(n6723), .B(n4162), .Z(n4488) );
  XNOR U4971 ( .A(n[48]), .B(n4163), .Z(n4164) );
  NANDN U4972 ( .A(n524), .B(n4164), .Z(n4165) );
  XOR U4973 ( .A(n4166), .B(n4165), .Z(n5432) );
  NAND U4974 ( .A(n[48]), .B(n5432), .Z(n4486) );
  XOR U4975 ( .A(n6716), .B(n4167), .Z(n4168) );
  NANDN U4976 ( .A(n524), .B(n4168), .Z(n4169) );
  XNOR U4977 ( .A(n4170), .B(n4169), .Z(n6719) );
  NANDN U4978 ( .A(n6716), .B(n6719), .Z(n4483) );
  XNOR U4979 ( .A(n6716), .B(n6719), .Z(n4481) );
  XOR U4980 ( .A(n6710), .B(n4171), .Z(n4172) );
  NANDN U4981 ( .A(n524), .B(n4172), .Z(n4173) );
  XOR U4982 ( .A(n4174), .B(n4173), .Z(n6714) );
  NANDN U4983 ( .A(n6710), .B(n6714), .Z(n4480) );
  NOR U4984 ( .A(n[46]), .B(n6714), .Z(n4478) );
  XNOR U4985 ( .A(n4179), .B(n4175), .Z(n4176) );
  NANDN U4986 ( .A(n524), .B(n4176), .Z(n4177) );
  XOR U4987 ( .A(n4178), .B(n4177), .Z(n6697) );
  NANDN U4988 ( .A(n4179), .B(n6697), .Z(n4461) );
  XNOR U4989 ( .A(n4179), .B(n6697), .Z(n4459) );
  IV U4990 ( .A(n[41]), .Z(n4454) );
  XOR U4991 ( .A(n4454), .B(n4180), .Z(n4181) );
  NANDN U4992 ( .A(n524), .B(n4181), .Z(n4182) );
  XOR U4993 ( .A(n4183), .B(n4182), .Z(n6690) );
  NANDN U4994 ( .A(n4454), .B(n6690), .Z(n4457) );
  XNOR U4995 ( .A(n4188), .B(n4184), .Z(n4185) );
  NANDN U4996 ( .A(n524), .B(n4185), .Z(n4186) );
  XOR U4997 ( .A(n4187), .B(n4186), .Z(n6686) );
  NANDN U4998 ( .A(n4188), .B(n6686), .Z(n4453) );
  XNOR U4999 ( .A(n4188), .B(n6686), .Z(n4451) );
  XOR U5000 ( .A(n4446), .B(n4189), .Z(n4190) );
  NANDN U5001 ( .A(n524), .B(n4190), .Z(n4191) );
  XNOR U5002 ( .A(n4192), .B(n4191), .Z(n6679) );
  NANDN U5003 ( .A(n4446), .B(n6679), .Z(n4449) );
  XOR U5004 ( .A(n4197), .B(n4193), .Z(n4194) );
  NANDN U5005 ( .A(n524), .B(n4194), .Z(n4195) );
  XNOR U5006 ( .A(n4196), .B(n4195), .Z(n6671) );
  NANDN U5007 ( .A(n4197), .B(n6671), .Z(n4445) );
  XNOR U5008 ( .A(n4197), .B(n6671), .Z(n4443) );
  XOR U5009 ( .A(n4438), .B(n4198), .Z(n4199) );
  NANDN U5010 ( .A(n524), .B(n4199), .Z(n4200) );
  XNOR U5011 ( .A(n4201), .B(n4200), .Z(n6664) );
  NANDN U5012 ( .A(n4438), .B(n6664), .Z(n4441) );
  XOR U5013 ( .A(n6656), .B(n4202), .Z(n4203) );
  NANDN U5014 ( .A(n524), .B(n4203), .Z(n4204) );
  XNOR U5015 ( .A(n4205), .B(n4204), .Z(n6658) );
  NANDN U5016 ( .A(n6656), .B(n6658), .Z(n4437) );
  XNOR U5017 ( .A(n[34]), .B(n4206), .Z(n4207) );
  NANDN U5018 ( .A(n524), .B(n4207), .Z(n4208) );
  XNOR U5019 ( .A(n4209), .B(n4208), .Z(n6648) );
  NAND U5020 ( .A(n[34]), .B(n6648), .Z(n4425) );
  XNOR U5021 ( .A(n[33]), .B(n4210), .Z(n4211) );
  NANDN U5022 ( .A(n524), .B(n4211), .Z(n4212) );
  XNOR U5023 ( .A(n4213), .B(n4212), .Z(n6644) );
  NAND U5024 ( .A(n[33]), .B(n6644), .Z(n4422) );
  XOR U5025 ( .A(n[32]), .B(n4214), .Z(n4215) );
  NANDN U5026 ( .A(n524), .B(n4215), .Z(n4216) );
  XNOR U5027 ( .A(n4217), .B(n4216), .Z(n6640) );
  XNOR U5028 ( .A(n4222), .B(n4218), .Z(n4219) );
  NANDN U5029 ( .A(n524), .B(n4219), .Z(n4220) );
  XNOR U5030 ( .A(n4221), .B(n4220), .Z(n6629) );
  NANDN U5031 ( .A(n4222), .B(n6629), .Z(n4414) );
  XNOR U5032 ( .A(n4222), .B(n6629), .Z(n4412) );
  XNOR U5033 ( .A(n4407), .B(n4223), .Z(n4224) );
  NANDN U5034 ( .A(n524), .B(n4224), .Z(n4225) );
  XNOR U5035 ( .A(n4226), .B(n4225), .Z(n6622) );
  NANDN U5036 ( .A(n4407), .B(n6622), .Z(n4410) );
  XNOR U5037 ( .A(n[26]), .B(n4227), .Z(n4228) );
  NANDN U5038 ( .A(n524), .B(n4228), .Z(n4229) );
  XNOR U5039 ( .A(n4230), .B(n4229), .Z(n6605) );
  NAND U5040 ( .A(n[26]), .B(n6605), .Z(n4397) );
  XOR U5041 ( .A(n[26]), .B(n6605), .Z(n4395) );
  XOR U5042 ( .A(n[25]), .B(n4231), .Z(n4232) );
  NANDN U5043 ( .A(n524), .B(n4232), .Z(n4233) );
  XNOR U5044 ( .A(n4234), .B(n4233), .Z(n6598) );
  NAND U5045 ( .A(n[25]), .B(n6598), .Z(n4393) );
  XNOR U5046 ( .A(n4239), .B(n4235), .Z(n4236) );
  NANDN U5047 ( .A(n524), .B(n4236), .Z(n4237) );
  XNOR U5048 ( .A(n4238), .B(n4237), .Z(n6544) );
  XNOR U5049 ( .A(n4382), .B(n4240), .Z(n4241) );
  NANDN U5050 ( .A(n524), .B(n4241), .Z(n4242) );
  XNOR U5051 ( .A(n4243), .B(n4242), .Z(n6406) );
  NANDN U5052 ( .A(n4382), .B(n6406), .Z(n4385) );
  XNOR U5053 ( .A(n4248), .B(n4244), .Z(n4245) );
  NANDN U5054 ( .A(n524), .B(n4245), .Z(n4246) );
  XNOR U5055 ( .A(n4247), .B(n4246), .Z(n6267) );
  NANDN U5056 ( .A(n4248), .B(n6267), .Z(n4377) );
  XNOR U5057 ( .A(n4248), .B(n6267), .Z(n4375) );
  XNOR U5058 ( .A(n4370), .B(n4249), .Z(n4250) );
  NANDN U5059 ( .A(n524), .B(n4250), .Z(n4251) );
  XNOR U5060 ( .A(n4252), .B(n4251), .Z(n6260) );
  NANDN U5061 ( .A(n4370), .B(n6260), .Z(n4373) );
  XNOR U5062 ( .A(n4257), .B(n4253), .Z(n4254) );
  NANDN U5063 ( .A(n524), .B(n4254), .Z(n4255) );
  XNOR U5064 ( .A(n4256), .B(n4255), .Z(n6129) );
  NANDN U5065 ( .A(n4257), .B(n6129), .Z(n4369) );
  XNOR U5066 ( .A(n4257), .B(n6129), .Z(n4367) );
  XNOR U5067 ( .A(n4362), .B(n4258), .Z(n4259) );
  NANDN U5068 ( .A(n524), .B(n4259), .Z(n4260) );
  XOR U5069 ( .A(n4261), .B(n4260), .Z(n6122) );
  NANDN U5070 ( .A(n4362), .B(n6122), .Z(n4365) );
  XNOR U5071 ( .A(n4266), .B(n4262), .Z(n4263) );
  NANDN U5072 ( .A(n524), .B(n4263), .Z(n4264) );
  XOR U5073 ( .A(n4265), .B(n4264), .Z(n5985) );
  IV U5074 ( .A(n[15]), .Z(n4358) );
  XNOR U5075 ( .A(n4271), .B(n4267), .Z(n4268) );
  NANDN U5076 ( .A(n524), .B(n4268), .Z(n4269) );
  XOR U5077 ( .A(n4270), .B(n4269), .Z(n5853) );
  NANDN U5078 ( .A(n4271), .B(n5853), .Z(n4356) );
  XNOR U5079 ( .A(n4271), .B(n5853), .Z(n4354) );
  XNOR U5080 ( .A(n4349), .B(n4272), .Z(n4273) );
  NANDN U5081 ( .A(n524), .B(n4273), .Z(n4274) );
  XOR U5082 ( .A(n4275), .B(n4274), .Z(n5846) );
  NANDN U5083 ( .A(n4349), .B(n5846), .Z(n4352) );
  XOR U5084 ( .A(n4276), .B(n[8]), .Z(n4277) );
  ANDN U5085 ( .B(n4277), .A(n524), .Z(n4278) );
  XNOR U5086 ( .A(n4279), .B(n4278), .Z(n6844) );
  NAND U5087 ( .A(n6844), .B(n[8]), .Z(n4325) );
  XOR U5088 ( .A(n[8]), .B(n6844), .Z(n4323) );
  IV U5089 ( .A(n[7]), .Z(n4318) );
  XNOR U5090 ( .A(n4318), .B(n4280), .Z(n4281) );
  ANDN U5091 ( .B(n4281), .A(n524), .Z(n4282) );
  XOR U5092 ( .A(n4283), .B(n4282), .Z(n6837) );
  NANDN U5093 ( .A(n4318), .B(n6837), .Z(n4321) );
  XOR U5094 ( .A(n[6]), .B(n4284), .Z(n4285) );
  NANDN U5095 ( .A(n524), .B(n4285), .Z(n4286) );
  XNOR U5096 ( .A(n4287), .B(n4286), .Z(n6788) );
  NAND U5097 ( .A(n[6]), .B(n6788), .Z(n4317) );
  XOR U5098 ( .A(n[6]), .B(n6788), .Z(n4315) );
  XOR U5099 ( .A(n4288), .B(n[5]), .Z(n4289) );
  ANDN U5100 ( .B(n4289), .A(n524), .Z(n4290) );
  XNOR U5101 ( .A(n4291), .B(n4290), .Z(n6781) );
  NAND U5102 ( .A(n[5]), .B(n6781), .Z(n4313) );
  XOR U5103 ( .A(n[4]), .B(n4292), .Z(n4293) );
  NANDN U5104 ( .A(n524), .B(n4293), .Z(n4294) );
  XNOR U5105 ( .A(n4295), .B(n4294), .Z(n6729) );
  NAND U5106 ( .A(n[4]), .B(n6729), .Z(n4310) );
  ANDN U5107 ( .B(n[0]), .A(n5342), .Z(n6195) );
  XOR U5108 ( .A(n[1]), .B(n4296), .Z(n4297) );
  NANDN U5109 ( .A(n524), .B(n4297), .Z(n4298) );
  XNOR U5110 ( .A(n4299), .B(n4298), .Z(n6198) );
  XNOR U5111 ( .A(n4300), .B(n6616), .Z(n4301) );
  ANDN U5112 ( .B(n4301), .A(n524), .Z(n4302) );
  XOR U5113 ( .A(n4303), .B(n4302), .Z(n6619) );
  XOR U5114 ( .A(n[3]), .B(n4304), .Z(n4305) );
  NANDN U5115 ( .A(n524), .B(n4305), .Z(n4306) );
  XNOR U5116 ( .A(n4307), .B(n4306), .Z(n6676) );
  XOR U5117 ( .A(n6729), .B(n[4]), .Z(n4308) );
  NANDN U5118 ( .A(n6726), .B(n4308), .Z(n4309) );
  AND U5119 ( .A(n4310), .B(n4309), .Z(n6754) );
  XOR U5120 ( .A(n6781), .B(n[5]), .Z(n4311) );
  NANDN U5121 ( .A(n6754), .B(n4311), .Z(n4312) );
  NAND U5122 ( .A(n4313), .B(n4312), .Z(n4314) );
  NAND U5123 ( .A(n4315), .B(n4314), .Z(n4316) );
  AND U5124 ( .A(n4317), .B(n4316), .Z(n6813) );
  XNOR U5125 ( .A(n6837), .B(n4318), .Z(n4319) );
  NANDN U5126 ( .A(n6813), .B(n4319), .Z(n4320) );
  NAND U5127 ( .A(n4321), .B(n4320), .Z(n4322) );
  NAND U5128 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U5129 ( .A(n4325), .B(n4324), .Z(n6867) );
  XOR U5130 ( .A(n6868), .B(n4326), .Z(n4327) );
  NANDN U5131 ( .A(n524), .B(n4327), .Z(n4328) );
  XNOR U5132 ( .A(n4329), .B(n4328), .Z(n6871) );
  XOR U5133 ( .A(n[10]), .B(n4330), .Z(n4331) );
  NANDN U5134 ( .A(n524), .B(n4331), .Z(n4332) );
  XNOR U5135 ( .A(n4333), .B(n4332), .Z(n5598) );
  XOR U5136 ( .A(n[10]), .B(n5598), .Z(n4334) );
  NANDN U5137 ( .A(n5595), .B(n4334), .Z(n4336) );
  NAND U5138 ( .A(n5598), .B(n[10]), .Z(n4335) );
  NAND U5139 ( .A(n4336), .B(n4335), .Z(n5655) );
  ANDN U5140 ( .B(n5655), .A(n4337), .Z(n4342) );
  XNOR U5141 ( .A(n4338), .B(n4337), .Z(n4339) );
  ANDN U5142 ( .B(n4339), .A(n524), .Z(n4340) );
  XNOR U5143 ( .A(n4341), .B(n4340), .Z(n5658) );
  OR U5144 ( .A(n4342), .B(n5658), .Z(n4344) );
  NOR U5145 ( .A(n[11]), .B(n5655), .Z(n4343) );
  ANDN U5146 ( .B(n4344), .A(n4343), .Z(n5716) );
  XOR U5147 ( .A(n[12]), .B(n4345), .Z(n4346) );
  NANDN U5148 ( .A(n524), .B(n4346), .Z(n4347) );
  XOR U5149 ( .A(n4348), .B(n4347), .Z(n5719) );
  XNOR U5150 ( .A(n5846), .B(n4349), .Z(n4350) );
  NANDN U5151 ( .A(n5782), .B(n4350), .Z(n4351) );
  NAND U5152 ( .A(n4352), .B(n4351), .Z(n4353) );
  NAND U5153 ( .A(n4354), .B(n4353), .Z(n4355) );
  NAND U5154 ( .A(n4356), .B(n4355), .Z(n5918) );
  XNOR U5155 ( .A(n4358), .B(n4357), .Z(n4359) );
  NANDN U5156 ( .A(n524), .B(n4359), .Z(n4360) );
  XNOR U5157 ( .A(n4361), .B(n4360), .Z(n5978) );
  XNOR U5158 ( .A(n6122), .B(n4362), .Z(n4363) );
  NANDN U5159 ( .A(n6054), .B(n4363), .Z(n4364) );
  NAND U5160 ( .A(n4365), .B(n4364), .Z(n4366) );
  NAND U5161 ( .A(n4367), .B(n4366), .Z(n4368) );
  AND U5162 ( .A(n4369), .B(n4368), .Z(n6194) );
  XNOR U5163 ( .A(n6260), .B(n4370), .Z(n4371) );
  NANDN U5164 ( .A(n6194), .B(n4371), .Z(n4372) );
  NAND U5165 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U5166 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U5167 ( .A(n4377), .B(n4376), .Z(n6331) );
  XOR U5168 ( .A(n[21]), .B(n4378), .Z(n4379) );
  NANDN U5169 ( .A(n524), .B(n4379), .Z(n4380) );
  XNOR U5170 ( .A(n4381), .B(n4380), .Z(n6334) );
  XNOR U5171 ( .A(n6406), .B(n4382), .Z(n4383) );
  NANDN U5172 ( .A(n6403), .B(n4383), .Z(n4384) );
  NAND U5173 ( .A(n4385), .B(n4384), .Z(n6473) );
  XNOR U5174 ( .A(n4387), .B(n4386), .Z(n4388) );
  NANDN U5175 ( .A(n524), .B(n4388), .Z(n4389) );
  XNOR U5176 ( .A(n4390), .B(n4389), .Z(n6537) );
  XOR U5177 ( .A(n6598), .B(n[25]), .Z(n4391) );
  NANDN U5178 ( .A(n6595), .B(n4391), .Z(n4392) );
  NAND U5179 ( .A(n4393), .B(n4392), .Z(n4394) );
  NAND U5180 ( .A(n4395), .B(n4394), .Z(n4396) );
  NAND U5181 ( .A(n4397), .B(n4396), .Z(n6606) );
  XOR U5182 ( .A(n4399), .B(n4398), .Z(n4400) );
  NANDN U5183 ( .A(n524), .B(n4400), .Z(n4401) );
  XOR U5184 ( .A(n4402), .B(n4401), .Z(n6609) );
  XNOR U5185 ( .A(n[28]), .B(n4403), .Z(n4404) );
  NANDN U5186 ( .A(n524), .B(n4404), .Z(n4405) );
  XNOR U5187 ( .A(n4406), .B(n4405), .Z(n6613) );
  XNOR U5188 ( .A(n6622), .B(n4407), .Z(n4408) );
  NANDN U5189 ( .A(n6614), .B(n4408), .Z(n4409) );
  NAND U5190 ( .A(n4410), .B(n4409), .Z(n4411) );
  NAND U5191 ( .A(n4412), .B(n4411), .Z(n4413) );
  NAND U5192 ( .A(n4414), .B(n4413), .Z(n6630) );
  XNOR U5193 ( .A(n4416), .B(n4415), .Z(n4417) );
  NANDN U5194 ( .A(n524), .B(n4417), .Z(n4418) );
  XNOR U5195 ( .A(n4419), .B(n4418), .Z(n6633) );
  XOR U5196 ( .A(n6644), .B(n[33]), .Z(n4420) );
  NANDN U5197 ( .A(n6641), .B(n4420), .Z(n4421) );
  AND U5198 ( .A(n4422), .B(n4421), .Z(n6645) );
  XOR U5199 ( .A(n[34]), .B(n6648), .Z(n4423) );
  NANDN U5200 ( .A(n6645), .B(n4423), .Z(n4424) );
  AND U5201 ( .A(n4425), .B(n4424), .Z(n6649) );
  NANDN U5202 ( .A(n[35]), .B(n6649), .Z(n4427) );
  NOR U5203 ( .A(n[36]), .B(n6658), .Z(n4426) );
  ANDN U5204 ( .B(n4427), .A(n4426), .Z(n4435) );
  XOR U5205 ( .A(n4432), .B(n4428), .Z(n4429) );
  NANDN U5206 ( .A(n524), .B(n4429), .Z(n4430) );
  XNOR U5207 ( .A(n4431), .B(n4430), .Z(n6650) );
  XOR U5208 ( .A(n4432), .B(n6649), .Z(n4433) );
  NANDN U5209 ( .A(n6650), .B(n4433), .Z(n4434) );
  NAND U5210 ( .A(n4435), .B(n4434), .Z(n4436) );
  AND U5211 ( .A(n4437), .B(n4436), .Z(n6661) );
  XNOR U5212 ( .A(n6664), .B(n4438), .Z(n4439) );
  NANDN U5213 ( .A(n6661), .B(n4439), .Z(n4440) );
  NAND U5214 ( .A(n4441), .B(n4440), .Z(n4442) );
  NAND U5215 ( .A(n4443), .B(n4442), .Z(n4444) );
  AND U5216 ( .A(n4445), .B(n4444), .Z(n6672) );
  XNOR U5217 ( .A(n6679), .B(n4446), .Z(n4447) );
  NANDN U5218 ( .A(n6672), .B(n4447), .Z(n4448) );
  NAND U5219 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U5220 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U5221 ( .A(n4453), .B(n4452), .Z(n6687) );
  XNOR U5222 ( .A(n6690), .B(n4454), .Z(n4455) );
  NANDN U5223 ( .A(n6687), .B(n4455), .Z(n4456) );
  NAND U5224 ( .A(n4457), .B(n4456), .Z(n4458) );
  NAND U5225 ( .A(n4459), .B(n4458), .Z(n4460) );
  NAND U5226 ( .A(n4461), .B(n4460), .Z(n6698) );
  IV U5227 ( .A(n[43]), .Z(n4463) );
  XNOR U5228 ( .A(n4463), .B(n4462), .Z(n4464) );
  NANDN U5229 ( .A(n524), .B(n4464), .Z(n4465) );
  XNOR U5230 ( .A(n4466), .B(n4465), .Z(n6701) );
  XOR U5231 ( .A(n[44]), .B(n4467), .Z(n4468) );
  NANDN U5232 ( .A(n524), .B(n4468), .Z(n4469) );
  XNOR U5233 ( .A(n4470), .B(n4469), .Z(n6705) );
  XNOR U5234 ( .A(n[45]), .B(n4471), .Z(n4472) );
  NANDN U5235 ( .A(n524), .B(n4472), .Z(n4473) );
  XNOR U5236 ( .A(n4474), .B(n4473), .Z(n6709) );
  XOR U5237 ( .A(n[45]), .B(n6709), .Z(n4475) );
  NANDN U5238 ( .A(n6706), .B(n4475), .Z(n4477) );
  NAND U5239 ( .A(n[45]), .B(n6709), .Z(n4476) );
  NAND U5240 ( .A(n4477), .B(n4476), .Z(n6711) );
  NANDN U5241 ( .A(n4478), .B(n6711), .Z(n4479) );
  NAND U5242 ( .A(n4480), .B(n4479), .Z(n6715) );
  NAND U5243 ( .A(n4481), .B(n6715), .Z(n4482) );
  AND U5244 ( .A(n4483), .B(n4482), .Z(n5430) );
  XOR U5245 ( .A(n5432), .B(n[48]), .Z(n4484) );
  NANDN U5246 ( .A(n5430), .B(n4484), .Z(n4485) );
  NAND U5247 ( .A(n4486), .B(n4485), .Z(n4487) );
  NAND U5248 ( .A(n4488), .B(n4487), .Z(n4489) );
  NAND U5249 ( .A(n4490), .B(n4489), .Z(n4491) );
  NAND U5250 ( .A(n4492), .B(n4491), .Z(n4493) );
  NAND U5251 ( .A(n4494), .B(n4493), .Z(n4495) );
  NAND U5252 ( .A(n4496), .B(n4495), .Z(n4497) );
  NAND U5253 ( .A(n4498), .B(n4497), .Z(n4499) );
  NAND U5254 ( .A(n4500), .B(n4499), .Z(n4501) );
  NAND U5255 ( .A(n4502), .B(n4501), .Z(n4503) );
  NAND U5256 ( .A(n4504), .B(n4503), .Z(n4505) );
  NAND U5257 ( .A(n4506), .B(n4505), .Z(n4507) );
  NAND U5258 ( .A(n4508), .B(n4507), .Z(n4509) );
  NAND U5259 ( .A(n4510), .B(n4509), .Z(n4511) );
  NAND U5260 ( .A(n4512), .B(n4511), .Z(n4513) );
  NAND U5261 ( .A(n4514), .B(n4513), .Z(n4515) );
  NAND U5262 ( .A(n4516), .B(n4515), .Z(n4517) );
  NAND U5263 ( .A(n4518), .B(n4517), .Z(n4519) );
  NAND U5264 ( .A(n4520), .B(n4519), .Z(n4521) );
  NAND U5265 ( .A(n4522), .B(n4521), .Z(n4523) );
  NAND U5266 ( .A(n4524), .B(n4523), .Z(n4525) );
  NAND U5267 ( .A(n4526), .B(n4525), .Z(n4527) );
  NAND U5268 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U5269 ( .A(n4530), .B(n4529), .Z(n4531) );
  NAND U5270 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U5271 ( .A(n4534), .B(n4533), .Z(n4535) );
  NAND U5272 ( .A(n4536), .B(n4535), .Z(n4537) );
  NAND U5273 ( .A(n4538), .B(n4537), .Z(n4539) );
  NAND U5274 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U5275 ( .A(n4542), .B(n4541), .Z(n4543) );
  NAND U5276 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U5277 ( .A(n4546), .B(n4545), .Z(n4547) );
  NAND U5278 ( .A(n4548), .B(n4547), .Z(n4549) );
  NAND U5279 ( .A(n4550), .B(n4549), .Z(n4551) );
  NAND U5280 ( .A(n4552), .B(n4551), .Z(n4553) );
  NAND U5281 ( .A(n4554), .B(n4553), .Z(n4555) );
  NAND U5282 ( .A(n4556), .B(n4555), .Z(n4557) );
  NAND U5283 ( .A(n4558), .B(n4557), .Z(n4559) );
  NAND U5284 ( .A(n4560), .B(n4559), .Z(n4561) );
  NAND U5285 ( .A(n4562), .B(n4561), .Z(n4563) );
  NAND U5286 ( .A(n4564), .B(n4563), .Z(n4565) );
  NAND U5287 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U5288 ( .A(n4568), .B(n4567), .Z(n4569) );
  AND U5289 ( .A(n4570), .B(n4569), .Z(n4574) );
  NANDN U5290 ( .A(n5471), .B(n4574), .Z(n4572) );
  ANDN U5291 ( .B(n5475), .A(n[71]), .Z(n4571) );
  ANDN U5292 ( .B(n4572), .A(n4571), .Z(n4577) );
  XOR U5293 ( .A(n4574), .B(n4573), .Z(n4575) );
  NANDN U5294 ( .A(n[70]), .B(n4575), .Z(n4576) );
  NAND U5295 ( .A(n4577), .B(n4576), .Z(n4578) );
  NAND U5296 ( .A(n4579), .B(n4578), .Z(n4580) );
  NAND U5297 ( .A(n4581), .B(n4580), .Z(n4582) );
  NAND U5298 ( .A(n4583), .B(n4582), .Z(n4584) );
  NAND U5299 ( .A(n4585), .B(n4584), .Z(n4586) );
  NAND U5300 ( .A(n4587), .B(n4586), .Z(n4588) );
  NAND U5301 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U5302 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U5303 ( .A(n4593), .B(n4592), .Z(n4594) );
  NAND U5304 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U5305 ( .A(n4597), .B(n4596), .Z(n4598) );
  NAND U5306 ( .A(n4599), .B(n4598), .Z(n4600) );
  NAND U5307 ( .A(n4601), .B(n4600), .Z(n4602) );
  NAND U5308 ( .A(n4603), .B(n4602), .Z(n4604) );
  NAND U5309 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U5310 ( .A(n4607), .B(n4606), .Z(n4608) );
  NAND U5311 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U5312 ( .A(n4611), .B(n4610), .Z(n4612) );
  NAND U5313 ( .A(n4613), .B(n4612), .Z(n4614) );
  NAND U5314 ( .A(n4615), .B(n4614), .Z(n4616) );
  NAND U5315 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U5316 ( .A(n4619), .B(n4618), .Z(n4620) );
  NAND U5317 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U5318 ( .A(n4623), .B(n4622), .Z(n4624) );
  NAND U5319 ( .A(n4625), .B(n4624), .Z(n4626) );
  NAND U5320 ( .A(n4627), .B(n4626), .Z(n4628) );
  NAND U5321 ( .A(n4629), .B(n4628), .Z(n4630) );
  NAND U5322 ( .A(n4631), .B(n4630), .Z(n4632) );
  NAND U5323 ( .A(n4633), .B(n4632), .Z(n4634) );
  NAND U5324 ( .A(n4635), .B(n4634), .Z(n4636) );
  NAND U5325 ( .A(n4637), .B(n4636), .Z(n4638) );
  NAND U5326 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U5327 ( .A(n4641), .B(n4640), .Z(n4642) );
  NAND U5328 ( .A(n4643), .B(n4642), .Z(n4644) );
  NAND U5329 ( .A(n4645), .B(n4644), .Z(n4646) );
  NAND U5330 ( .A(n4647), .B(n4646), .Z(n4648) );
  NAND U5331 ( .A(n4649), .B(n4648), .Z(n4650) );
  NAND U5332 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U5333 ( .A(n4653), .B(n4652), .Z(n4654) );
  NAND U5334 ( .A(n4655), .B(n4654), .Z(n4656) );
  NAND U5335 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U5336 ( .A(n4659), .B(n4658), .Z(n4665) );
  XNOR U5337 ( .A(n5353), .B(n4660), .Z(n4661) );
  NANDN U5338 ( .A(n524), .B(n4661), .Z(n4662) );
  XNOR U5339 ( .A(n4663), .B(n4662), .Z(n5356) );
  XNOR U5340 ( .A(n4665), .B(n5356), .Z(n4664) );
  NANDN U5341 ( .A(n5353), .B(n4664), .Z(n4667) );
  NANDN U5342 ( .A(n4665), .B(n5356), .Z(n4666) );
  AND U5343 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U5344 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U5345 ( .A(n4671), .B(n4670), .Z(n4672) );
  OR U5346 ( .A(n5350), .B(n4672), .Z(n4675) );
  XOR U5347 ( .A(n5350), .B(n4672), .Z(n4673) );
  NANDN U5348 ( .A(n[94]), .B(n4673), .Z(n4674) );
  NAND U5349 ( .A(n4675), .B(n4674), .Z(n4676) );
  NAND U5350 ( .A(n4677), .B(n4676), .Z(n4679) );
  NANDN U5351 ( .A(n5531), .B(n5529), .Z(n4678) );
  AND U5352 ( .A(n4679), .B(n4678), .Z(n4680) );
  NAND U5353 ( .A(n4681), .B(n4680), .Z(n4682) );
  NAND U5354 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U5355 ( .A(n4685), .B(n4684), .Z(n4686) );
  NAND U5356 ( .A(n4687), .B(n4686), .Z(n4688) );
  NAND U5357 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U5358 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U5359 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U5360 ( .A(n4695), .B(n4694), .Z(n4696) );
  NAND U5361 ( .A(n4697), .B(n4696), .Z(n4698) );
  NAND U5362 ( .A(n4699), .B(n4698), .Z(n4700) );
  NAND U5363 ( .A(n4701), .B(n4700), .Z(n4702) );
  NAND U5364 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U5365 ( .A(n4705), .B(n4704), .Z(n4706) );
  NAND U5366 ( .A(n4707), .B(n4706), .Z(n4708) );
  NAND U5367 ( .A(n4709), .B(n4708), .Z(n4710) );
  NAND U5368 ( .A(n4711), .B(n4710), .Z(n4712) );
  NAND U5369 ( .A(n4713), .B(n4712), .Z(n4714) );
  NAND U5370 ( .A(n4715), .B(n4714), .Z(n4716) );
  NAND U5371 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U5372 ( .A(n4719), .B(n4718), .Z(n4720) );
  NAND U5373 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U5374 ( .A(n4723), .B(n4722), .Z(n4724) );
  NAND U5375 ( .A(n4725), .B(n4724), .Z(n4726) );
  NAND U5376 ( .A(n4727), .B(n4726), .Z(n4728) );
  NAND U5377 ( .A(n4729), .B(n4728), .Z(n4730) );
  NAND U5378 ( .A(n4731), .B(n4730), .Z(n4732) );
  NAND U5379 ( .A(n4733), .B(n4732), .Z(n4734) );
  NAND U5380 ( .A(n4735), .B(n4734), .Z(n4736) );
  NAND U5381 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U5382 ( .A(n4739), .B(n4738), .Z(n4740) );
  NAND U5383 ( .A(n4741), .B(n4740), .Z(n4742) );
  NAND U5384 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U5385 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U5386 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U5387 ( .A(n4749), .B(n4748), .Z(n4750) );
  NAND U5388 ( .A(n4751), .B(n4750), .Z(n4752) );
  NAND U5389 ( .A(n4753), .B(n4752), .Z(n4754) );
  NAND U5390 ( .A(n4755), .B(n4754), .Z(n4756) );
  NAND U5391 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5392 ( .A(n4759), .B(n4758), .Z(n4760) );
  NAND U5393 ( .A(n4761), .B(n4760), .Z(n4762) );
  NAND U5394 ( .A(n4763), .B(n4762), .Z(n4764) );
  NAND U5395 ( .A(n4765), .B(n4764), .Z(n4766) );
  NAND U5396 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U5397 ( .A(n4769), .B(n4768), .Z(n4770) );
  NAND U5398 ( .A(n4771), .B(n4770), .Z(n4772) );
  NAND U5399 ( .A(n4773), .B(n4772), .Z(n4774) );
  NAND U5400 ( .A(n4775), .B(n4774), .Z(n4776) );
  NAND U5401 ( .A(n4777), .B(n4776), .Z(n4778) );
  NAND U5402 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U5403 ( .A(n4781), .B(n4780), .Z(n4782) );
  NAND U5404 ( .A(n4783), .B(n4782), .Z(n4784) );
  NAND U5405 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U5406 ( .A(n4787), .B(n4786), .Z(n4788) );
  NAND U5407 ( .A(n4789), .B(n4788), .Z(n4790) );
  NAND U5408 ( .A(n4791), .B(n4790), .Z(n4792) );
  NAND U5409 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U5410 ( .A(n4795), .B(n4794), .Z(n4796) );
  NAND U5411 ( .A(n4797), .B(n4796), .Z(n4798) );
  NAND U5412 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U5413 ( .A(n4801), .B(n4800), .Z(n4802) );
  NAND U5414 ( .A(n4803), .B(n4802), .Z(n4804) );
  NAND U5415 ( .A(n4805), .B(n4804), .Z(n4806) );
  NAND U5416 ( .A(n4807), .B(n4806), .Z(n4808) );
  NAND U5417 ( .A(n4809), .B(n4808), .Z(n4810) );
  NAND U5418 ( .A(n4811), .B(n4810), .Z(n4812) );
  NAND U5419 ( .A(n4813), .B(n4812), .Z(n4814) );
  NAND U5420 ( .A(n4815), .B(n4814), .Z(n4816) );
  NAND U5421 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U5422 ( .A(n4819), .B(n4818), .Z(n4820) );
  NAND U5423 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U5424 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U5425 ( .A(n4825), .B(n4824), .Z(n4826) );
  NAND U5426 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5427 ( .A(n4829), .B(n4828), .Z(n4830) );
  NAND U5428 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U5429 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U5430 ( .A(n4835), .B(n4834), .Z(n4836) );
  NAND U5431 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U5432 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U5433 ( .A(n4841), .B(n4840), .Z(n4842) );
  NAND U5434 ( .A(n4843), .B(n4842), .Z(n4844) );
  NAND U5435 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5436 ( .A(n4847), .B(n4846), .Z(n4848) );
  NAND U5437 ( .A(n4849), .B(n4848), .Z(n4850) );
  NAND U5438 ( .A(n4851), .B(n4850), .Z(n4852) );
  NAND U5439 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U5440 ( .A(n4855), .B(n4854), .Z(n4856) );
  NAND U5441 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U5442 ( .A(n4859), .B(n4858), .Z(n4860) );
  NAND U5443 ( .A(n4861), .B(n4860), .Z(n4862) );
  NAND U5444 ( .A(n4863), .B(n4862), .Z(n4864) );
  NAND U5445 ( .A(n4865), .B(n4864), .Z(n4866) );
  NAND U5446 ( .A(n4867), .B(n4866), .Z(n4868) );
  NAND U5447 ( .A(n4869), .B(n4868), .Z(n4870) );
  NAND U5448 ( .A(n4871), .B(n4870), .Z(n4872) );
  NAND U5449 ( .A(n4873), .B(n4872), .Z(n4874) );
  NAND U5450 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U5451 ( .A(n4877), .B(n4876), .Z(n4878) );
  NAND U5452 ( .A(n4879), .B(n4878), .Z(n4880) );
  NAND U5453 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U5454 ( .A(n4883), .B(n4882), .Z(n4884) );
  NAND U5455 ( .A(n4885), .B(n4884), .Z(n4886) );
  NAND U5456 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U5457 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U5458 ( .A(n4891), .B(n4890), .Z(n4892) );
  NAND U5459 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U5460 ( .A(n4895), .B(n4894), .Z(n4896) );
  NAND U5461 ( .A(n4897), .B(n4896), .Z(n4898) );
  NAND U5462 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U5463 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U5464 ( .A(n4903), .B(n4902), .Z(n4904) );
  NAND U5465 ( .A(n4905), .B(n4904), .Z(n4906) );
  AND U5466 ( .A(n4907), .B(n4906), .Z(n4908) );
  OR U5467 ( .A(n4908), .B(n4910), .Z(n4916) );
  XOR U5468 ( .A(n4908), .B(n4910), .Z(n4914) );
  XOR U5469 ( .A(n4910), .B(n4909), .Z(n4911) );
  NANDN U5470 ( .A(n524), .B(n4911), .Z(n4912) );
  XNOR U5471 ( .A(n4913), .B(n4912), .Z(n5879) );
  NAND U5472 ( .A(n4914), .B(n5879), .Z(n4915) );
  NAND U5473 ( .A(n4916), .B(n4915), .Z(n4917) );
  NAND U5474 ( .A(n4918), .B(n4917), .Z(n4919) );
  AND U5475 ( .A(n4920), .B(n4919), .Z(n4922) );
  NANDN U5476 ( .A(n4922), .B(n[155]), .Z(n4921) );
  AND U5477 ( .A(n5898), .B(n4921), .Z(n4929) );
  XNOR U5478 ( .A(n[155]), .B(n4922), .Z(n4927) );
  XOR U5479 ( .A(n[155]), .B(n4923), .Z(n4924) );
  NANDN U5480 ( .A(n524), .B(n4924), .Z(n4925) );
  XNOR U5481 ( .A(n4926), .B(n4925), .Z(n5892) );
  NAND U5482 ( .A(n4927), .B(n5892), .Z(n4928) );
  NAND U5483 ( .A(n4929), .B(n4928), .Z(n4930) );
  NAND U5484 ( .A(n4931), .B(n4930), .Z(n4938) );
  NANDN U5485 ( .A(n[157]), .B(n4938), .Z(n4933) );
  NOR U5486 ( .A(n[158]), .B(n5905), .Z(n4932) );
  ANDN U5487 ( .B(n4933), .A(n4932), .Z(n4942) );
  XNOR U5488 ( .A(n4939), .B(n4934), .Z(n4935) );
  NANDN U5489 ( .A(n524), .B(n4935), .Z(n4936) );
  XNOR U5490 ( .A(n4937), .B(n4936), .Z(n5906) );
  XOR U5491 ( .A(n4939), .B(n4938), .Z(n4940) );
  NANDN U5492 ( .A(n5906), .B(n4940), .Z(n4941) );
  NAND U5493 ( .A(n4942), .B(n4941), .Z(n4943) );
  NANDN U5494 ( .A(n5912), .B(n4943), .Z(n4944) );
  NAND U5495 ( .A(n4945), .B(n4944), .Z(n4946) );
  NAND U5496 ( .A(n4947), .B(n4946), .Z(n4948) );
  NAND U5497 ( .A(n4949), .B(n4948), .Z(n4950) );
  NAND U5498 ( .A(n4951), .B(n4950), .Z(n4952) );
  NAND U5499 ( .A(n4953), .B(n4952), .Z(n4954) );
  NAND U5500 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U5501 ( .A(n4957), .B(n4956), .Z(n4958) );
  NAND U5502 ( .A(n4959), .B(n4958), .Z(n4960) );
  NAND U5503 ( .A(n4961), .B(n4960), .Z(n4962) );
  NAND U5504 ( .A(n4963), .B(n4962), .Z(n4964) );
  NAND U5505 ( .A(n4965), .B(n4964), .Z(n4966) );
  NAND U5506 ( .A(n4967), .B(n4966), .Z(n4968) );
  NAND U5507 ( .A(n4969), .B(n4968), .Z(n4970) );
  NAND U5508 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U5509 ( .A(n4973), .B(n4972), .Z(n4974) );
  NAND U5510 ( .A(n4975), .B(n4974), .Z(n4976) );
  NAND U5511 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5512 ( .A(n4979), .B(n4978), .Z(n4980) );
  NAND U5513 ( .A(n4981), .B(n4980), .Z(n4982) );
  NAND U5514 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5515 ( .A(n4985), .B(n4984), .Z(n4986) );
  NAND U5516 ( .A(n4987), .B(n4986), .Z(n4988) );
  NAND U5517 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U5518 ( .A(n4991), .B(n4990), .Z(n4992) );
  NAND U5519 ( .A(n4993), .B(n4992), .Z(n4994) );
  NAND U5520 ( .A(n4995), .B(n4994), .Z(n4996) );
  NAND U5521 ( .A(n4997), .B(n4996), .Z(n4998) );
  NAND U5522 ( .A(n4999), .B(n4998), .Z(n5000) );
  NAND U5523 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U5524 ( .A(n5003), .B(n5002), .Z(n5004) );
  NAND U5525 ( .A(n5005), .B(n5004), .Z(n5006) );
  NAND U5526 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U5527 ( .A(n5009), .B(n5008), .Z(n5010) );
  NAND U5528 ( .A(n5011), .B(n5010), .Z(n5012) );
  NAND U5529 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U5530 ( .A(n5015), .B(n5014), .Z(n5016) );
  NAND U5531 ( .A(n5017), .B(n5016), .Z(n5018) );
  NAND U5532 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U5533 ( .A(n5021), .B(n5020), .Z(n5022) );
  NANDN U5534 ( .A(n5022), .B(n[179]), .Z(n5029) );
  XNOR U5535 ( .A(n5022), .B(n[179]), .Z(n5027) );
  XNOR U5536 ( .A(n[179]), .B(n5023), .Z(n5024) );
  NANDN U5537 ( .A(n524), .B(n5024), .Z(n5025) );
  XNOR U5538 ( .A(n5026), .B(n5025), .Z(n6055) );
  NAND U5539 ( .A(n5027), .B(n6055), .Z(n5028) );
  NAND U5540 ( .A(n5029), .B(n5028), .Z(n5030) );
  NAND U5541 ( .A(n5031), .B(n5030), .Z(n5032) );
  NAND U5542 ( .A(n5033), .B(n5032), .Z(n5034) );
  NAND U5543 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U5544 ( .A(n5037), .B(n5036), .Z(n5038) );
  NAND U5545 ( .A(n5039), .B(n5038), .Z(n5040) );
  NAND U5546 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U5547 ( .A(n5043), .B(n5042), .Z(n5044) );
  NAND U5548 ( .A(n5045), .B(n5044), .Z(n5046) );
  NAND U5549 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U5550 ( .A(n5049), .B(n5048), .Z(n5050) );
  NANDN U5551 ( .A(n5050), .B(n[185]), .Z(n5057) );
  XNOR U5552 ( .A(n5050), .B(n[185]), .Z(n5055) );
  XOR U5553 ( .A(n[185]), .B(n5051), .Z(n5052) );
  NANDN U5554 ( .A(n524), .B(n5052), .Z(n5053) );
  XNOR U5555 ( .A(n5054), .B(n5053), .Z(n6093) );
  NAND U5556 ( .A(n5055), .B(n6093), .Z(n5056) );
  NAND U5557 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U5558 ( .A(n5059), .B(n5058), .Z(n5060) );
  NAND U5559 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U5560 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U5561 ( .A(n5065), .B(n5064), .Z(n5066) );
  NAND U5562 ( .A(n5067), .B(n5066), .Z(n5068) );
  NAND U5563 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND U5564 ( .A(n5071), .B(n5070), .Z(n5072) );
  NAND U5565 ( .A(n5073), .B(n5072), .Z(n5074) );
  NAND U5566 ( .A(n5075), .B(n5074), .Z(n5076) );
  NAND U5567 ( .A(n5077), .B(n5076), .Z(n5078) );
  NAND U5568 ( .A(n5079), .B(n5078), .Z(n5080) );
  NAND U5569 ( .A(n5081), .B(n5080), .Z(n5082) );
  NAND U5570 ( .A(n5083), .B(n5082), .Z(n5084) );
  NAND U5571 ( .A(n5085), .B(n5084), .Z(n5086) );
  NAND U5572 ( .A(n5087), .B(n5086), .Z(n5088) );
  NAND U5573 ( .A(n5089), .B(n5088), .Z(n5090) );
  NAND U5574 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U5575 ( .A(n5093), .B(n5092), .Z(n5094) );
  NAND U5576 ( .A(n5095), .B(n5094), .Z(n5096) );
  NAND U5577 ( .A(n5097), .B(n5096), .Z(n5099) );
  OR U5578 ( .A(n6168), .B(n[196]), .Z(n5098) );
  AND U5579 ( .A(n5099), .B(n5098), .Z(n5100) );
  NAND U5580 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U5581 ( .A(n5103), .B(n5102), .Z(n5104) );
  NAND U5582 ( .A(n5105), .B(n5104), .Z(n5106) );
  NAND U5583 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U5584 ( .A(n5109), .B(n5108), .Z(n5110) );
  NAND U5585 ( .A(n5111), .B(n5110), .Z(n5113) );
  OR U5586 ( .A(n6201), .B(n[200]), .Z(n5112) );
  AND U5587 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5588 ( .A(n5115), .B(n5114), .Z(n5116) );
  NAND U5589 ( .A(n5117), .B(n5116), .Z(n5118) );
  NAND U5590 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U5591 ( .A(n5121), .B(n5120), .Z(n5122) );
  NAND U5592 ( .A(n5123), .B(n5122), .Z(n5124) );
  NAND U5593 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U5594 ( .A(n5127), .B(n5126), .Z(n5128) );
  NAND U5595 ( .A(n5129), .B(n5128), .Z(n5130) );
  NAND U5596 ( .A(n5131), .B(n5130), .Z(n5132) );
  NAND U5597 ( .A(n5133), .B(n5132), .Z(n5134) );
  NAND U5598 ( .A(n5135), .B(n5134), .Z(n5136) );
  NAND U5599 ( .A(n5137), .B(n5136), .Z(n5138) );
  NAND U5600 ( .A(n5139), .B(n5138), .Z(n5140) );
  NAND U5601 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5602 ( .A(n5143), .B(n5142), .Z(n5144) );
  NAND U5603 ( .A(n5145), .B(n5144), .Z(n5147) );
  XNOR U5604 ( .A(n6271), .B(n[209]), .Z(n5146) );
  NANDN U5605 ( .A(n5147), .B(n5146), .Z(n5148) );
  NAND U5606 ( .A(n5149), .B(n5148), .Z(n5150) );
  NANDN U5607 ( .A(n6278), .B(n5150), .Z(n5151) );
  NAND U5608 ( .A(n5152), .B(n5151), .Z(n5153) );
  NAND U5609 ( .A(n5154), .B(n5153), .Z(n5155) );
  NAND U5610 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U5611 ( .A(n5158), .B(n5157), .Z(n5159) );
  NAND U5612 ( .A(n5160), .B(n5159), .Z(n5161) );
  NAND U5613 ( .A(n5162), .B(n5161), .Z(n5163) );
  NAND U5614 ( .A(n5164), .B(n5163), .Z(n5165) );
  NAND U5615 ( .A(n5166), .B(n5165), .Z(n5167) );
  NAND U5616 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U5617 ( .A(n5170), .B(n5169), .Z(n5171) );
  NAND U5618 ( .A(n5172), .B(n5171), .Z(n5173) );
  AND U5619 ( .A(n5174), .B(n5173), .Z(n5180) );
  XNOR U5620 ( .A(n[217]), .B(n5175), .Z(n5176) );
  NANDN U5621 ( .A(n524), .B(n5176), .Z(n5177) );
  XNOR U5622 ( .A(n5178), .B(n5177), .Z(n6320) );
  NANDN U5623 ( .A(n5180), .B(n6320), .Z(n5179) );
  AND U5624 ( .A(n6326), .B(n5179), .Z(n5183) );
  XNOR U5625 ( .A(n6320), .B(n5180), .Z(n5181) );
  NAND U5626 ( .A(n[217]), .B(n5181), .Z(n5182) );
  NAND U5627 ( .A(n5183), .B(n5182), .Z(n5185) );
  OR U5628 ( .A(n6319), .B(n[218]), .Z(n5184) );
  AND U5629 ( .A(n5185), .B(n5184), .Z(n5186) );
  NAND U5630 ( .A(n5187), .B(n5186), .Z(n5188) );
  NAND U5631 ( .A(n5189), .B(n5188), .Z(n5190) );
  NAND U5632 ( .A(n5191), .B(n5190), .Z(n5192) );
  NAND U5633 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U5634 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U5635 ( .A(n5197), .B(n5196), .Z(n5198) );
  NAND U5636 ( .A(n5199), .B(n5198), .Z(n5200) );
  NAND U5637 ( .A(n5201), .B(n5200), .Z(n5202) );
  NAND U5638 ( .A(n5203), .B(n5202), .Z(n5204) );
  NAND U5639 ( .A(n5205), .B(n5204), .Z(n5206) );
  NAND U5640 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U5641 ( .A(n5209), .B(n5208), .Z(n5210) );
  NAND U5642 ( .A(n5211), .B(n5210), .Z(n5212) );
  NAND U5643 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5644 ( .A(n5215), .B(n5214), .Z(n5216) );
  NAND U5645 ( .A(n5217), .B(n5216), .Z(n5218) );
  NAND U5646 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U5647 ( .A(n5221), .B(n5220), .Z(n5222) );
  NAND U5648 ( .A(n5223), .B(n5222), .Z(n5224) );
  NAND U5649 ( .A(n5225), .B(n5224), .Z(n5226) );
  NAND U5650 ( .A(n5227), .B(n5226), .Z(n5228) );
  AND U5651 ( .A(n5229), .B(n5228), .Z(n5234) );
  XNOR U5652 ( .A(n[230]), .B(n5230), .Z(n5231) );
  NANDN U5653 ( .A(n524), .B(n5231), .Z(n5232) );
  XNOR U5654 ( .A(n5233), .B(n5232), .Z(n6416) );
  NANDN U5655 ( .A(n5234), .B(n6416), .Z(n5237) );
  XNOR U5656 ( .A(n6416), .B(n5234), .Z(n5235) );
  NAND U5657 ( .A(n[230]), .B(n5235), .Z(n5236) );
  NAND U5658 ( .A(n5237), .B(n5236), .Z(n5238) );
  AND U5659 ( .A(n5239), .B(n5238), .Z(n5240) );
  ANDN U5660 ( .B(n6415), .A(n6413), .Z(n6422) );
  OR U5661 ( .A(n5240), .B(n6422), .Z(n5241) );
  NAND U5662 ( .A(n5242), .B(n5241), .Z(n5243) );
  NAND U5663 ( .A(n5244), .B(n5243), .Z(n5245) );
  NAND U5664 ( .A(n5246), .B(n5245), .Z(n5247) );
  NAND U5665 ( .A(n5248), .B(n5247), .Z(n5249) );
  NAND U5666 ( .A(n5250), .B(n5249), .Z(n5251) );
  NAND U5667 ( .A(n5252), .B(n5251), .Z(n5253) );
  NAND U5668 ( .A(n5254), .B(n5253), .Z(n5255) );
  AND U5669 ( .A(n5256), .B(n5255), .Z(n5264) );
  NANDN U5670 ( .A(n6450), .B(n5264), .Z(n5262) );
  XOR U5671 ( .A(n6456), .B(n5257), .Z(n5258) );
  NANDN U5672 ( .A(n524), .B(n5258), .Z(n5259) );
  XOR U5673 ( .A(n5260), .B(n5259), .Z(n6457) );
  ANDN U5674 ( .B(n6457), .A(n[237]), .Z(n5261) );
  ANDN U5675 ( .B(n5262), .A(n5261), .Z(n5267) );
  XOR U5676 ( .A(n5264), .B(n5263), .Z(n5265) );
  NANDN U5677 ( .A(n[236]), .B(n5265), .Z(n5266) );
  NAND U5678 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U5679 ( .A(n5268), .B(n6459), .Z(n5269) );
  NAND U5680 ( .A(n5270), .B(n5269), .Z(n5271) );
  NAND U5681 ( .A(n5272), .B(n5271), .Z(n5273) );
  NAND U5682 ( .A(n5274), .B(n5273), .Z(n5275) );
  NAND U5683 ( .A(n5276), .B(n5275), .Z(n5277) );
  NAND U5684 ( .A(n5278), .B(n5277), .Z(n5279) );
  NAND U5685 ( .A(n5280), .B(n5279), .Z(n5281) );
  NAND U5686 ( .A(n5282), .B(n5281), .Z(n5283) );
  NAND U5687 ( .A(n5284), .B(n5283), .Z(n5285) );
  NAND U5688 ( .A(n5286), .B(n5285), .Z(n5287) );
  NAND U5689 ( .A(n5288), .B(n5287), .Z(n5289) );
  NAND U5690 ( .A(n5290), .B(n5289), .Z(n5291) );
  NAND U5691 ( .A(n5292), .B(n5291), .Z(n5293) );
  NAND U5692 ( .A(n5294), .B(n5293), .Z(n5295) );
  NAND U5693 ( .A(n5296), .B(n5295), .Z(n5297) );
  NAND U5694 ( .A(n5298), .B(n5297), .Z(n5299) );
  NAND U5695 ( .A(n5300), .B(n5299), .Z(n5301) );
  NAND U5696 ( .A(n5302), .B(n5301), .Z(n5303) );
  NAND U5697 ( .A(n5304), .B(n5303), .Z(n5305) );
  NAND U5698 ( .A(n5306), .B(n5305), .Z(n5307) );
  NAND U5699 ( .A(n5308), .B(n5307), .Z(n5309) );
  NAND U5700 ( .A(n5310), .B(n5309), .Z(n5311) );
  NAND U5701 ( .A(n5312), .B(n5311), .Z(n5313) );
  NAND U5702 ( .A(n5314), .B(n5313), .Z(n5315) );
  NAND U5703 ( .A(n5316), .B(n5315), .Z(n5317) );
  NAND U5704 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U5705 ( .A(n5320), .B(n5319), .Z(n5321) );
  NAND U5706 ( .A(n5322), .B(n5321), .Z(n5323) );
  NAND U5707 ( .A(n5324), .B(n5323), .Z(n5325) );
  NAND U5708 ( .A(n5326), .B(n5325), .Z(n5327) );
  NAND U5709 ( .A(n5328), .B(n5327), .Z(n5329) );
  NAND U5710 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5711 ( .A(n5332), .B(n5331), .Z(n5333) );
  NAND U5712 ( .A(n5334), .B(n5333), .Z(n5335) );
  NAND U5713 ( .A(n5336), .B(n5335), .Z(n5338) );
  XOR U5714 ( .A(n[255]), .B(n6580), .Z(n5337) );
  NANDN U5715 ( .A(n5338), .B(n5337), .Z(n5339) );
  NAND U5716 ( .A(n5340), .B(n5339), .Z(n6814) );
  ANDN U5717 ( .B(n[0]), .A(n525), .Z(n5341) );
  XOR U5718 ( .A(n5342), .B(n5341), .Z(zout[0]) );
  NANDN U5719 ( .A(n525), .B(n[100]), .Z(n5343) );
  XOR U5720 ( .A(n5544), .B(n5343), .Z(n5547) );
  NANDN U5721 ( .A(n5344), .B(n6814), .Z(n5541) );
  AND U5722 ( .A(n5347), .B(n[98]), .Z(n5345) );
  NANDN U5723 ( .A(n525), .B(n5345), .Z(n5539) );
  NANDN U5724 ( .A(n525), .B(n[98]), .Z(n5346) );
  XOR U5725 ( .A(n5347), .B(n5346), .Z(n6863) );
  AND U5726 ( .A(n6814), .B(n[96]), .Z(n5534) );
  OR U5727 ( .A(n5534), .B(n5535), .Z(n5537) );
  ANDN U5728 ( .B(n5531), .A(n5529), .Z(n5348) );
  NANDN U5729 ( .A(n525), .B(n5348), .Z(n5533) );
  NANDN U5730 ( .A(n525), .B(n[94]), .Z(n5349) );
  NANDN U5731 ( .A(n5349), .B(n5350), .Z(n5528) );
  XOR U5732 ( .A(n5350), .B(n5349), .Z(n6854) );
  NANDN U5733 ( .A(n525), .B(n[93]), .Z(n5351) );
  NANDN U5734 ( .A(n5351), .B(n5352), .Z(n5526) );
  XOR U5735 ( .A(n5352), .B(n5351), .Z(n6852) );
  ANDN U5736 ( .B(n5356), .A(n5353), .Z(n5354) );
  NANDN U5737 ( .A(n525), .B(n5354), .Z(n5524) );
  NANDN U5738 ( .A(n525), .B(n[92]), .Z(n5355) );
  XOR U5739 ( .A(n5356), .B(n5355), .Z(n6850) );
  AND U5740 ( .A(n5359), .B(n[91]), .Z(n5357) );
  NANDN U5741 ( .A(n525), .B(n5357), .Z(n5522) );
  NANDN U5742 ( .A(n525), .B(n[91]), .Z(n5358) );
  XOR U5743 ( .A(n5359), .B(n5358), .Z(n6848) );
  NANDN U5744 ( .A(n525), .B(n[90]), .Z(n5360) );
  NANDN U5745 ( .A(n5360), .B(n5361), .Z(n5520) );
  XOR U5746 ( .A(n5361), .B(n5360), .Z(n6846) );
  AND U5747 ( .A(n5364), .B(n[89]), .Z(n5362) );
  NANDN U5748 ( .A(n525), .B(n5362), .Z(n5518) );
  NANDN U5749 ( .A(n525), .B(n[89]), .Z(n5363) );
  XOR U5750 ( .A(n5364), .B(n5363), .Z(n6834) );
  NANDN U5751 ( .A(n525), .B(n[87]), .Z(n5365) );
  NANDN U5752 ( .A(n5365), .B(n5366), .Z(n5512) );
  XOR U5753 ( .A(n5366), .B(n5365), .Z(n6830) );
  NANDN U5754 ( .A(n525), .B(n[86]), .Z(n5367) );
  NANDN U5755 ( .A(n5367), .B(n5368), .Z(n5510) );
  XOR U5756 ( .A(n5368), .B(n5367), .Z(n6828) );
  NANDN U5757 ( .A(n525), .B(n[84]), .Z(n5369) );
  NANDN U5758 ( .A(n5369), .B(n5370), .Z(n5503) );
  XOR U5759 ( .A(n5370), .B(n5369), .Z(n6824) );
  NANDN U5760 ( .A(n525), .B(n[83]), .Z(n5371) );
  NANDN U5761 ( .A(n5371), .B(n5372), .Z(n5501) );
  XOR U5762 ( .A(n5372), .B(n5371), .Z(n6822) );
  AND U5763 ( .A(n5375), .B(n[82]), .Z(n5373) );
  NANDN U5764 ( .A(n525), .B(n5373), .Z(n5499) );
  NANDN U5765 ( .A(n525), .B(n[82]), .Z(n5374) );
  XOR U5766 ( .A(n5375), .B(n5374), .Z(n6820) );
  NANDN U5767 ( .A(n525), .B(n[81]), .Z(n5376) );
  NANDN U5768 ( .A(n5376), .B(n5377), .Z(n5497) );
  XOR U5769 ( .A(n5377), .B(n5376), .Z(n6818) );
  NANDN U5770 ( .A(n525), .B(n[80]), .Z(n5378) );
  NANDN U5771 ( .A(n5378), .B(n5379), .Z(n5495) );
  XOR U5772 ( .A(n5379), .B(n5378), .Z(n6815) );
  NANDN U5773 ( .A(n525), .B(n[78]), .Z(n5380) );
  NANDN U5774 ( .A(n5380), .B(n5381), .Z(n5493) );
  XOR U5775 ( .A(n5381), .B(n5380), .Z(n6808) );
  NANDN U5776 ( .A(n525), .B(n[76]), .Z(n5382) );
  NANDN U5777 ( .A(n5382), .B(n5383), .Z(n5491) );
  XOR U5778 ( .A(n5383), .B(n5382), .Z(n6802) );
  AND U5779 ( .A(n5386), .B(n[74]), .Z(n5384) );
  NANDN U5780 ( .A(n525), .B(n5384), .Z(n5485) );
  NANDN U5781 ( .A(n525), .B(n[74]), .Z(n5385) );
  XOR U5782 ( .A(n5386), .B(n5385), .Z(n6798) );
  NANDN U5783 ( .A(n525), .B(n[73]), .Z(n5387) );
  NANDN U5784 ( .A(n5387), .B(n5388), .Z(n5483) );
  XOR U5785 ( .A(n5388), .B(n5387), .Z(n6796) );
  AND U5786 ( .A(n5479), .B(n[72]), .Z(n5389) );
  NANDN U5787 ( .A(n525), .B(n5389), .Z(n5481) );
  NANDN U5788 ( .A(n5390), .B(n6814), .Z(n5474) );
  AND U5789 ( .A(n5475), .B(n5474), .Z(n5477) );
  ANDN U5790 ( .B(n5471), .A(n5469), .Z(n5391) );
  NANDN U5791 ( .A(n525), .B(n5391), .Z(n5473) );
  NANDN U5792 ( .A(n525), .B(n[69]), .Z(n5392) );
  NANDN U5793 ( .A(n5392), .B(n5393), .Z(n5468) );
  XOR U5794 ( .A(n5393), .B(n5392), .Z(n6777) );
  AND U5795 ( .A(n5396), .B(n[67]), .Z(n5394) );
  NANDN U5796 ( .A(n525), .B(n5394), .Z(n5466) );
  NANDN U5797 ( .A(n525), .B(n[67]), .Z(n5395) );
  XOR U5798 ( .A(n5396), .B(n5395), .Z(n6771) );
  NANDN U5799 ( .A(n525), .B(n[65]), .Z(n5397) );
  NANDN U5800 ( .A(n5397), .B(n5398), .Z(n5464) );
  XOR U5801 ( .A(n5398), .B(n5397), .Z(n6766) );
  ANDN U5802 ( .B(n5402), .A(n5399), .Z(n5400) );
  NANDN U5803 ( .A(n525), .B(n5400), .Z(n5462) );
  NANDN U5804 ( .A(n525), .B(n[64]), .Z(n5401) );
  XOR U5805 ( .A(n5402), .B(n5401), .Z(n6764) );
  NANDN U5806 ( .A(n525), .B(n[62]), .Z(n5403) );
  NANDN U5807 ( .A(n5403), .B(n5404), .Z(n5456) );
  XOR U5808 ( .A(n5404), .B(n5403), .Z(n6760) );
  NANDN U5809 ( .A(n525), .B(n[61]), .Z(n5405) );
  NANDN U5810 ( .A(n5405), .B(n5406), .Z(n5454) );
  XOR U5811 ( .A(n5406), .B(n5405), .Z(n6758) );
  NANDN U5812 ( .A(n525), .B(n[60]), .Z(n5407) );
  NANDN U5813 ( .A(n5407), .B(n5408), .Z(n5452) );
  XOR U5814 ( .A(n5408), .B(n5407), .Z(n6756) );
  NANDN U5815 ( .A(n525), .B(n[59]), .Z(n5409) );
  NANDN U5816 ( .A(n5409), .B(n5410), .Z(n5450) );
  XOR U5817 ( .A(n5410), .B(n5409), .Z(n6753) );
  ANDN U5818 ( .B(n5414), .A(n5411), .Z(n5412) );
  NANDN U5819 ( .A(n525), .B(n5412), .Z(n5448) );
  NANDN U5820 ( .A(n525), .B(n[58]), .Z(n5413) );
  XOR U5821 ( .A(n5414), .B(n5413), .Z(n6751) );
  AND U5822 ( .A(n5417), .B(n[57]), .Z(n5415) );
  NANDN U5823 ( .A(n525), .B(n5415), .Z(n5446) );
  NANDN U5824 ( .A(n525), .B(n[57]), .Z(n5416) );
  XOR U5825 ( .A(n5417), .B(n5416), .Z(n6749) );
  NANDN U5826 ( .A(n525), .B(n[56]), .Z(n5418) );
  NANDN U5827 ( .A(n5418), .B(n5419), .Z(n5444) );
  XOR U5828 ( .A(n5419), .B(n5418), .Z(n6747) );
  NANDN U5829 ( .A(n525), .B(n[55]), .Z(n5420) );
  NANDN U5830 ( .A(n5420), .B(n5421), .Z(n5442) );
  XOR U5831 ( .A(n5421), .B(n5420), .Z(n6745) );
  NANDN U5832 ( .A(n525), .B(n[54]), .Z(n5422) );
  NANDN U5833 ( .A(n5422), .B(n5423), .Z(n5440) );
  XOR U5834 ( .A(n5423), .B(n5422), .Z(n6742) );
  AND U5835 ( .A(n5426), .B(n[52]), .Z(n5424) );
  NANDN U5836 ( .A(n525), .B(n5424), .Z(n5438) );
  NANDN U5837 ( .A(n525), .B(n[52]), .Z(n5425) );
  XOR U5838 ( .A(n5426), .B(n5425), .Z(n6737) );
  NANDN U5839 ( .A(n525), .B(n[51]), .Z(n5427) );
  NANDN U5840 ( .A(n5427), .B(n5428), .Z(n5436) );
  XOR U5841 ( .A(n5428), .B(n5427), .Z(n6734) );
  AND U5842 ( .A(n5432), .B(n[48]), .Z(n5429) );
  NANDN U5843 ( .A(n525), .B(n5429), .Z(n5434) );
  OR U5844 ( .A(n5430), .B(n525), .Z(n6721) );
  NANDN U5845 ( .A(n525), .B(n[48]), .Z(n5431) );
  XOR U5846 ( .A(n5432), .B(n5431), .Z(n6720) );
  OR U5847 ( .A(n6721), .B(n6720), .Z(n5433) );
  NAND U5848 ( .A(n5434), .B(n5433), .Z(n6725) );
  AND U5849 ( .A(n6814), .B(n[49]), .Z(n6722) );
  AND U5850 ( .A(n[50]), .B(n6814), .Z(n6733) );
  OR U5851 ( .A(n6734), .B(n6735), .Z(n5435) );
  AND U5852 ( .A(n5436), .B(n5435), .Z(n6736) );
  OR U5853 ( .A(n6737), .B(n6736), .Z(n5437) );
  AND U5854 ( .A(n5438), .B(n5437), .Z(n6738) );
  NANDN U5855 ( .A(n525), .B(n[53]), .Z(n6741) );
  NANDN U5856 ( .A(n6742), .B(n6743), .Z(n5439) );
  AND U5857 ( .A(n5440), .B(n5439), .Z(n6744) );
  OR U5858 ( .A(n6745), .B(n6744), .Z(n5441) );
  AND U5859 ( .A(n5442), .B(n5441), .Z(n6746) );
  OR U5860 ( .A(n6747), .B(n6746), .Z(n5443) );
  AND U5861 ( .A(n5444), .B(n5443), .Z(n6748) );
  OR U5862 ( .A(n6749), .B(n6748), .Z(n5445) );
  AND U5863 ( .A(n5446), .B(n5445), .Z(n6750) );
  OR U5864 ( .A(n6751), .B(n6750), .Z(n5447) );
  AND U5865 ( .A(n5448), .B(n5447), .Z(n6752) );
  OR U5866 ( .A(n6753), .B(n6752), .Z(n5449) );
  AND U5867 ( .A(n5450), .B(n5449), .Z(n6755) );
  OR U5868 ( .A(n6756), .B(n6755), .Z(n5451) );
  AND U5869 ( .A(n5452), .B(n5451), .Z(n6757) );
  OR U5870 ( .A(n6758), .B(n6757), .Z(n5453) );
  AND U5871 ( .A(n5454), .B(n5453), .Z(n6759) );
  OR U5872 ( .A(n6760), .B(n6759), .Z(n5455) );
  NAND U5873 ( .A(n5456), .B(n5455), .Z(n5457) );
  NAND U5874 ( .A(n5457), .B(n5458), .Z(n5460) );
  NANDN U5875 ( .A(n525), .B(n[63]), .Z(n6761) );
  XOR U5876 ( .A(n5458), .B(n5457), .Z(n6762) );
  NANDN U5877 ( .A(n6761), .B(n6762), .Z(n5459) );
  AND U5878 ( .A(n5460), .B(n5459), .Z(n6763) );
  OR U5879 ( .A(n6764), .B(n6763), .Z(n5461) );
  AND U5880 ( .A(n5462), .B(n5461), .Z(n6765) );
  OR U5881 ( .A(n6766), .B(n6765), .Z(n5463) );
  AND U5882 ( .A(n5464), .B(n5463), .Z(n6767) );
  NANDN U5883 ( .A(n525), .B(n[66]), .Z(n6770) );
  NANDN U5884 ( .A(n6771), .B(n6772), .Z(n5465) );
  AND U5885 ( .A(n5466), .B(n5465), .Z(n6773) );
  NANDN U5886 ( .A(n525), .B(n[68]), .Z(n6776) );
  NANDN U5887 ( .A(n6777), .B(n6778), .Z(n5467) );
  AND U5888 ( .A(n5468), .B(n5467), .Z(n6789) );
  NANDN U5889 ( .A(n5469), .B(n6814), .Z(n5470) );
  XNOR U5890 ( .A(n5471), .B(n5470), .Z(n6790) );
  NANDN U5891 ( .A(n6789), .B(n6790), .Z(n5472) );
  NAND U5892 ( .A(n5473), .B(n5472), .Z(n6791) );
  XOR U5893 ( .A(n5475), .B(n5474), .Z(n6792) );
  NANDN U5894 ( .A(n6791), .B(n6792), .Z(n5476) );
  NANDN U5895 ( .A(n5477), .B(n5476), .Z(n6794) );
  NANDN U5896 ( .A(n525), .B(n[72]), .Z(n5478) );
  XOR U5897 ( .A(n5479), .B(n5478), .Z(n6793) );
  OR U5898 ( .A(n6794), .B(n6793), .Z(n5480) );
  AND U5899 ( .A(n5481), .B(n5480), .Z(n6795) );
  OR U5900 ( .A(n6796), .B(n6795), .Z(n5482) );
  AND U5901 ( .A(n5483), .B(n5482), .Z(n6797) );
  OR U5902 ( .A(n6798), .B(n6797), .Z(n5484) );
  NAND U5903 ( .A(n5485), .B(n5484), .Z(n5486) );
  NAND U5904 ( .A(n5486), .B(n5487), .Z(n5489) );
  NANDN U5905 ( .A(n525), .B(n[75]), .Z(n6799) );
  XOR U5906 ( .A(n5487), .B(n5486), .Z(n6800) );
  NANDN U5907 ( .A(n6799), .B(n6800), .Z(n5488) );
  AND U5908 ( .A(n5489), .B(n5488), .Z(n6801) );
  OR U5909 ( .A(n6802), .B(n6801), .Z(n5490) );
  NAND U5910 ( .A(n5491), .B(n5490), .Z(n6806) );
  AND U5911 ( .A(n6814), .B(n[77]), .Z(n6803) );
  OR U5912 ( .A(n6808), .B(n6807), .Z(n5492) );
  NAND U5913 ( .A(n5493), .B(n5492), .Z(n6812) );
  AND U5914 ( .A(n[79]), .B(n6814), .Z(n6809) );
  OR U5915 ( .A(n6815), .B(n6816), .Z(n5494) );
  AND U5916 ( .A(n5495), .B(n5494), .Z(n6817) );
  OR U5917 ( .A(n6818), .B(n6817), .Z(n5496) );
  AND U5918 ( .A(n5497), .B(n5496), .Z(n6819) );
  OR U5919 ( .A(n6820), .B(n6819), .Z(n5498) );
  AND U5920 ( .A(n5499), .B(n5498), .Z(n6821) );
  OR U5921 ( .A(n6822), .B(n6821), .Z(n5500) );
  AND U5922 ( .A(n5501), .B(n5500), .Z(n6823) );
  OR U5923 ( .A(n6824), .B(n6823), .Z(n5502) );
  NAND U5924 ( .A(n5503), .B(n5502), .Z(n5505) );
  NAND U5925 ( .A(n5505), .B(n5506), .Z(n5508) );
  NANDN U5926 ( .A(n5504), .B(n6814), .Z(n6825) );
  XOR U5927 ( .A(n5506), .B(n5505), .Z(n6826) );
  NANDN U5928 ( .A(n6825), .B(n6826), .Z(n5507) );
  AND U5929 ( .A(n5508), .B(n5507), .Z(n6827) );
  OR U5930 ( .A(n6828), .B(n6827), .Z(n5509) );
  AND U5931 ( .A(n5510), .B(n5509), .Z(n6829) );
  OR U5932 ( .A(n6830), .B(n6829), .Z(n5511) );
  NAND U5933 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U5934 ( .A(n5513), .B(n5514), .Z(n5516) );
  NANDN U5935 ( .A(n525), .B(n[88]), .Z(n6831) );
  XOR U5936 ( .A(n5514), .B(n5513), .Z(n6832) );
  NANDN U5937 ( .A(n6831), .B(n6832), .Z(n5515) );
  AND U5938 ( .A(n5516), .B(n5515), .Z(n6833) );
  OR U5939 ( .A(n6834), .B(n6833), .Z(n5517) );
  AND U5940 ( .A(n5518), .B(n5517), .Z(n6845) );
  OR U5941 ( .A(n6846), .B(n6845), .Z(n5519) );
  AND U5942 ( .A(n5520), .B(n5519), .Z(n6847) );
  OR U5943 ( .A(n6848), .B(n6847), .Z(n5521) );
  AND U5944 ( .A(n5522), .B(n5521), .Z(n6849) );
  OR U5945 ( .A(n6850), .B(n6849), .Z(n5523) );
  AND U5946 ( .A(n5524), .B(n5523), .Z(n6851) );
  OR U5947 ( .A(n6852), .B(n6851), .Z(n5525) );
  AND U5948 ( .A(n5526), .B(n5525), .Z(n6853) );
  OR U5949 ( .A(n6854), .B(n6853), .Z(n5527) );
  AND U5950 ( .A(n5528), .B(n5527), .Z(n6855) );
  NANDN U5951 ( .A(n5529), .B(n6814), .Z(n5530) );
  XNOR U5952 ( .A(n5531), .B(n5530), .Z(n6856) );
  NANDN U5953 ( .A(n6855), .B(n6856), .Z(n5532) );
  NAND U5954 ( .A(n5533), .B(n5532), .Z(n6858) );
  XOR U5955 ( .A(n5535), .B(n5534), .Z(n6857) );
  NANDN U5956 ( .A(n6858), .B(n6857), .Z(n5536) );
  NAND U5957 ( .A(n5537), .B(n5536), .Z(n6859) );
  NANDN U5958 ( .A(n525), .B(n[97]), .Z(n6862) );
  NANDN U5959 ( .A(n6863), .B(n6864), .Z(n5538) );
  AND U5960 ( .A(n5539), .B(n5538), .Z(n5540) );
  OR U5961 ( .A(n5541), .B(n5540), .Z(n5543) );
  XNOR U5962 ( .A(n5541), .B(n5540), .Z(n6865) );
  NANDN U5963 ( .A(n6865), .B(n6866), .Z(n5542) );
  AND U5964 ( .A(n5543), .B(n5542), .Z(n5546) );
  XNOR U5965 ( .A(n5547), .B(n5546), .Z(zout[100]) );
  AND U5966 ( .A(n5544), .B(n[100]), .Z(n5545) );
  NANDN U5967 ( .A(n525), .B(n5545), .Z(n5549) );
  OR U5968 ( .A(n5547), .B(n5546), .Z(n5548) );
  NAND U5969 ( .A(n5549), .B(n5548), .Z(n5552) );
  AND U5970 ( .A(n6814), .B(n[101]), .Z(n5553) );
  XOR U5971 ( .A(n5551), .B(n5553), .Z(n5550) );
  XNOR U5972 ( .A(n5552), .B(n5550), .Z(zout[101]) );
  NANDN U5973 ( .A(n525), .B(n[102]), .Z(n5555) );
  XOR U5974 ( .A(n5554), .B(n5555), .Z(n5557) );
  XNOR U5975 ( .A(n5556), .B(n5557), .Z(zout[102]) );
  NANDN U5976 ( .A(n5555), .B(n5554), .Z(n5559) );
  OR U5977 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U5978 ( .A(n5559), .B(n5558), .Z(n5560) );
  XOR U5979 ( .A(n5561), .B(n5560), .Z(n5562) );
  AND U5980 ( .A(n6814), .B(n[103]), .Z(n5563) );
  XNOR U5981 ( .A(n5562), .B(n5563), .Z(zout[103]) );
  NANDN U5982 ( .A(n525), .B(n[104]), .Z(n5569) );
  OR U5983 ( .A(n5561), .B(n5560), .Z(n5565) );
  NANDN U5984 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U5985 ( .A(n5565), .B(n5564), .Z(n5568) );
  XOR U5986 ( .A(n5567), .B(n5568), .Z(n5566) );
  XNOR U5987 ( .A(n5569), .B(n5566), .Z(zout[104]) );
  NANDN U5988 ( .A(n525), .B(n[105]), .Z(n5571) );
  XOR U5989 ( .A(n5570), .B(n5571), .Z(n5573) );
  XOR U5990 ( .A(n5572), .B(n5573), .Z(zout[105]) );
  NANDN U5991 ( .A(n5571), .B(n5570), .Z(n5575) );
  NANDN U5992 ( .A(n5573), .B(n5572), .Z(n5574) );
  NAND U5993 ( .A(n5575), .B(n5574), .Z(n5576) );
  XOR U5994 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U5995 ( .A(n[106]), .B(n6814), .Z(n5579) );
  XNOR U5996 ( .A(n5578), .B(n5579), .Z(zout[106]) );
  OR U5997 ( .A(n5577), .B(n5576), .Z(n5581) );
  NANDN U5998 ( .A(n5579), .B(n5578), .Z(n5580) );
  AND U5999 ( .A(n5581), .B(n5580), .Z(n5583) );
  XOR U6000 ( .A(n5582), .B(n5583), .Z(n5584) );
  NANDN U6001 ( .A(n525), .B(n[107]), .Z(n5585) );
  XOR U6002 ( .A(n5584), .B(n5585), .Z(zout[107]) );
  NANDN U6003 ( .A(n525), .B(n[108]), .Z(n5590) );
  XOR U6004 ( .A(n5589), .B(n5590), .Z(n5592) );
  NAND U6005 ( .A(n5583), .B(n5582), .Z(n5587) );
  NANDN U6006 ( .A(n5585), .B(n5584), .Z(n5586) );
  AND U6007 ( .A(n5587), .B(n5586), .Z(n5591) );
  XNOR U6008 ( .A(n5592), .B(n5591), .Z(zout[108]) );
  NANDN U6009 ( .A(n525), .B(n[109]), .Z(n5588) );
  XOR U6010 ( .A(n5599), .B(n5588), .Z(n5602) );
  NANDN U6011 ( .A(n5590), .B(n5589), .Z(n5594) );
  OR U6012 ( .A(n5592), .B(n5591), .Z(n5593) );
  AND U6013 ( .A(n5594), .B(n5593), .Z(n5601) );
  XNOR U6014 ( .A(n5602), .B(n5601), .Z(zout[109]) );
  XNOR U6015 ( .A(n[10]), .B(n5595), .Z(n5596) );
  NANDN U6016 ( .A(n525), .B(n5596), .Z(n5597) );
  XOR U6017 ( .A(n5598), .B(n5597), .Z(zout[10]) );
  NANDN U6018 ( .A(n525), .B(n[110]), .Z(n5606) );
  XOR U6019 ( .A(n5605), .B(n5606), .Z(n5608) );
  AND U6020 ( .A(n5599), .B(n[109]), .Z(n5600) );
  NANDN U6021 ( .A(n525), .B(n5600), .Z(n5604) );
  OR U6022 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U6023 ( .A(n5604), .B(n5603), .Z(n5607) );
  XNOR U6024 ( .A(n5608), .B(n5607), .Z(zout[110]) );
  NANDN U6025 ( .A(n5606), .B(n5605), .Z(n5610) );
  OR U6026 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U6027 ( .A(n5610), .B(n5609), .Z(n5613) );
  AND U6028 ( .A(n6814), .B(n[111]), .Z(n5614) );
  XOR U6029 ( .A(n5612), .B(n5614), .Z(n5611) );
  XNOR U6030 ( .A(n5613), .B(n5611), .Z(zout[111]) );
  NANDN U6031 ( .A(n525), .B(n[112]), .Z(n5618) );
  XNOR U6032 ( .A(n5616), .B(n5617), .Z(n5615) );
  XNOR U6033 ( .A(n5618), .B(n5615), .Z(zout[112]) );
  NANDN U6034 ( .A(n525), .B(n[113]), .Z(n5622) );
  XNOR U6035 ( .A(n5621), .B(n5620), .Z(n5619) );
  XNOR U6036 ( .A(n5622), .B(n5619), .Z(zout[113]) );
  NANDN U6037 ( .A(n525), .B(n[114]), .Z(n5626) );
  XNOR U6038 ( .A(n5625), .B(n5624), .Z(n5623) );
  XNOR U6039 ( .A(n5626), .B(n5623), .Z(zout[114]) );
  NANDN U6040 ( .A(n525), .B(n[115]), .Z(n5628) );
  XOR U6041 ( .A(n5627), .B(n5628), .Z(n5630) );
  XOR U6042 ( .A(n5629), .B(n5630), .Z(zout[115]) );
  NANDN U6043 ( .A(n5628), .B(n5627), .Z(n5632) );
  NANDN U6044 ( .A(n5630), .B(n5629), .Z(n5631) );
  NAND U6045 ( .A(n5632), .B(n5631), .Z(n5635) );
  XOR U6046 ( .A(n5634), .B(n5635), .Z(n5636) );
  NANDN U6047 ( .A(n5633), .B(n6814), .Z(n5637) );
  XOR U6048 ( .A(n5636), .B(n5637), .Z(zout[116]) );
  NANDN U6049 ( .A(n525), .B(n[117]), .Z(n5642) );
  XOR U6050 ( .A(n5641), .B(n5642), .Z(n5644) );
  NAND U6051 ( .A(n5635), .B(n5634), .Z(n5639) );
  NANDN U6052 ( .A(n5637), .B(n5636), .Z(n5638) );
  AND U6053 ( .A(n5639), .B(n5638), .Z(n5643) );
  XNOR U6054 ( .A(n5644), .B(n5643), .Z(zout[117]) );
  NANDN U6055 ( .A(n5648), .B(n6814), .Z(n5640) );
  XOR U6056 ( .A(n5649), .B(n5640), .Z(n5652) );
  NANDN U6057 ( .A(n5642), .B(n5641), .Z(n5646) );
  OR U6058 ( .A(n5644), .B(n5643), .Z(n5645) );
  AND U6059 ( .A(n5646), .B(n5645), .Z(n5651) );
  XNOR U6060 ( .A(n5652), .B(n5651), .Z(zout[118]) );
  NANDN U6061 ( .A(n525), .B(n[119]), .Z(n5647) );
  XOR U6062 ( .A(n5659), .B(n5647), .Z(n5662) );
  ANDN U6063 ( .B(n5649), .A(n5648), .Z(n5650) );
  NANDN U6064 ( .A(n525), .B(n5650), .Z(n5654) );
  OR U6065 ( .A(n5652), .B(n5651), .Z(n5653) );
  AND U6066 ( .A(n5654), .B(n5653), .Z(n5661) );
  XNOR U6067 ( .A(n5662), .B(n5661), .Z(zout[119]) );
  XOR U6068 ( .A(n[11]), .B(n5655), .Z(n5656) );
  ANDN U6069 ( .B(n5656), .A(n525), .Z(n5657) );
  XNOR U6070 ( .A(n5658), .B(n5657), .Z(zout[11]) );
  AND U6071 ( .A(n5659), .B(n[119]), .Z(n5660) );
  NANDN U6072 ( .A(n525), .B(n5660), .Z(n5664) );
  OR U6073 ( .A(n5662), .B(n5661), .Z(n5663) );
  NAND U6074 ( .A(n5664), .B(n5663), .Z(n5667) );
  AND U6075 ( .A(n6814), .B(n[120]), .Z(n5668) );
  XOR U6076 ( .A(n5666), .B(n5668), .Z(n5665) );
  XNOR U6077 ( .A(n5667), .B(n5665), .Z(zout[120]) );
  NANDN U6078 ( .A(n525), .B(n[121]), .Z(n5670) );
  XOR U6079 ( .A(n5669), .B(n5670), .Z(n5672) );
  XNOR U6080 ( .A(n5671), .B(n5672), .Z(zout[121]) );
  NANDN U6081 ( .A(n525), .B(n[122]), .Z(n5676) );
  XOR U6082 ( .A(n5675), .B(n5676), .Z(n5678) );
  NANDN U6083 ( .A(n5670), .B(n5669), .Z(n5674) );
  OR U6084 ( .A(n5672), .B(n5671), .Z(n5673) );
  AND U6085 ( .A(n5674), .B(n5673), .Z(n5677) );
  XNOR U6086 ( .A(n5678), .B(n5677), .Z(zout[122]) );
  NANDN U6087 ( .A(n525), .B(n[123]), .Z(n5682) );
  XOR U6088 ( .A(n5681), .B(n5682), .Z(n5684) );
  NANDN U6089 ( .A(n5676), .B(n5675), .Z(n5680) );
  OR U6090 ( .A(n5678), .B(n5677), .Z(n5679) );
  AND U6091 ( .A(n5680), .B(n5679), .Z(n5683) );
  XNOR U6092 ( .A(n5684), .B(n5683), .Z(zout[123]) );
  NANDN U6093 ( .A(n525), .B(n[124]), .Z(n5688) );
  XOR U6094 ( .A(n5687), .B(n5688), .Z(n5690) );
  NANDN U6095 ( .A(n5682), .B(n5681), .Z(n5686) );
  OR U6096 ( .A(n5684), .B(n5683), .Z(n5685) );
  AND U6097 ( .A(n5686), .B(n5685), .Z(n5689) );
  XNOR U6098 ( .A(n5690), .B(n5689), .Z(zout[124]) );
  NANDN U6099 ( .A(n525), .B(n[125]), .Z(n5696) );
  NANDN U6100 ( .A(n5688), .B(n5687), .Z(n5692) );
  OR U6101 ( .A(n5690), .B(n5689), .Z(n5691) );
  AND U6102 ( .A(n5692), .B(n5691), .Z(n5695) );
  XOR U6103 ( .A(n5694), .B(n5695), .Z(n5693) );
  XNOR U6104 ( .A(n5696), .B(n5693), .Z(zout[125]) );
  NANDN U6105 ( .A(n525), .B(n[126]), .Z(n5698) );
  XOR U6106 ( .A(n5697), .B(n5698), .Z(n5700) );
  XOR U6107 ( .A(n5699), .B(n5700), .Z(zout[126]) );
  NANDN U6108 ( .A(n525), .B(n[127]), .Z(n5705) );
  XOR U6109 ( .A(n5704), .B(n5705), .Z(n5707) );
  NANDN U6110 ( .A(n5698), .B(n5697), .Z(n5702) );
  NANDN U6111 ( .A(n5700), .B(n5699), .Z(n5701) );
  AND U6112 ( .A(n5702), .B(n5701), .Z(n5706) );
  XNOR U6113 ( .A(n5707), .B(n5706), .Z(zout[127]) );
  NANDN U6114 ( .A(n525), .B(n[128]), .Z(n5703) );
  XOR U6115 ( .A(n5710), .B(n5703), .Z(n5713) );
  NANDN U6116 ( .A(n5705), .B(n5704), .Z(n5709) );
  OR U6117 ( .A(n5707), .B(n5706), .Z(n5708) );
  AND U6118 ( .A(n5709), .B(n5708), .Z(n5712) );
  XNOR U6119 ( .A(n5713), .B(n5712), .Z(zout[128]) );
  NANDN U6120 ( .A(n525), .B(n[129]), .Z(n5721) );
  XOR U6121 ( .A(n5720), .B(n5721), .Z(n5723) );
  AND U6122 ( .A(n5710), .B(n[128]), .Z(n5711) );
  NANDN U6123 ( .A(n525), .B(n5711), .Z(n5715) );
  OR U6124 ( .A(n5713), .B(n5712), .Z(n5714) );
  AND U6125 ( .A(n5715), .B(n5714), .Z(n5722) );
  XNOR U6126 ( .A(n5723), .B(n5722), .Z(zout[129]) );
  XOR U6127 ( .A(n[12]), .B(n5716), .Z(n5717) );
  NANDN U6128 ( .A(n525), .B(n5717), .Z(n5718) );
  XOR U6129 ( .A(n5719), .B(n5718), .Z(zout[12]) );
  NANDN U6130 ( .A(n525), .B(n[130]), .Z(n5728) );
  XOR U6131 ( .A(n5727), .B(n5728), .Z(n5730) );
  NANDN U6132 ( .A(n5721), .B(n5720), .Z(n5725) );
  OR U6133 ( .A(n5723), .B(n5722), .Z(n5724) );
  AND U6134 ( .A(n5725), .B(n5724), .Z(n5729) );
  XNOR U6135 ( .A(n5730), .B(n5729), .Z(zout[130]) );
  NANDN U6136 ( .A(n525), .B(n[131]), .Z(n5726) );
  XOR U6137 ( .A(n5733), .B(n5726), .Z(n5736) );
  NANDN U6138 ( .A(n5728), .B(n5727), .Z(n5732) );
  OR U6139 ( .A(n5730), .B(n5729), .Z(n5731) );
  AND U6140 ( .A(n5732), .B(n5731), .Z(n5735) );
  XNOR U6141 ( .A(n5736), .B(n5735), .Z(zout[131]) );
  NANDN U6142 ( .A(n525), .B(n[132]), .Z(n5740) );
  XOR U6143 ( .A(n5739), .B(n5740), .Z(n5742) );
  AND U6144 ( .A(n5733), .B(n[131]), .Z(n5734) );
  NANDN U6145 ( .A(n525), .B(n5734), .Z(n5738) );
  OR U6146 ( .A(n5736), .B(n5735), .Z(n5737) );
  AND U6147 ( .A(n5738), .B(n5737), .Z(n5741) );
  XNOR U6148 ( .A(n5742), .B(n5741), .Z(zout[132]) );
  NANDN U6149 ( .A(n525), .B(n[133]), .Z(n5747) );
  XOR U6150 ( .A(n5746), .B(n5747), .Z(n5749) );
  NANDN U6151 ( .A(n5740), .B(n5739), .Z(n5744) );
  OR U6152 ( .A(n5742), .B(n5741), .Z(n5743) );
  AND U6153 ( .A(n5744), .B(n5743), .Z(n5748) );
  XNOR U6154 ( .A(n5749), .B(n5748), .Z(zout[133]) );
  NANDN U6155 ( .A(n525), .B(n[134]), .Z(n5745) );
  XOR U6156 ( .A(n5752), .B(n5745), .Z(n5755) );
  NANDN U6157 ( .A(n5747), .B(n5746), .Z(n5751) );
  OR U6158 ( .A(n5749), .B(n5748), .Z(n5750) );
  AND U6159 ( .A(n5751), .B(n5750), .Z(n5754) );
  XNOR U6160 ( .A(n5755), .B(n5754), .Z(zout[134]) );
  NANDN U6161 ( .A(n525), .B(n[135]), .Z(n5759) );
  XOR U6162 ( .A(n5758), .B(n5759), .Z(n5761) );
  AND U6163 ( .A(n5752), .B(n[134]), .Z(n5753) );
  NANDN U6164 ( .A(n525), .B(n5753), .Z(n5757) );
  OR U6165 ( .A(n5755), .B(n5754), .Z(n5756) );
  AND U6166 ( .A(n5757), .B(n5756), .Z(n5760) );
  XNOR U6167 ( .A(n5761), .B(n5760), .Z(zout[135]) );
  NANDN U6168 ( .A(n525), .B(n[136]), .Z(n5765) );
  XOR U6169 ( .A(n5764), .B(n5765), .Z(n5767) );
  NANDN U6170 ( .A(n5759), .B(n5758), .Z(n5763) );
  OR U6171 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U6172 ( .A(n5763), .B(n5762), .Z(n5766) );
  XNOR U6173 ( .A(n5767), .B(n5766), .Z(zout[136]) );
  NANDN U6174 ( .A(n525), .B(n[137]), .Z(n5771) );
  XOR U6175 ( .A(n5770), .B(n5771), .Z(n5773) );
  NANDN U6176 ( .A(n5765), .B(n5764), .Z(n5769) );
  OR U6177 ( .A(n5767), .B(n5766), .Z(n5768) );
  AND U6178 ( .A(n5769), .B(n5768), .Z(n5772) );
  XNOR U6179 ( .A(n5773), .B(n5772), .Z(zout[137]) );
  NANDN U6180 ( .A(n5771), .B(n5770), .Z(n5775) );
  OR U6181 ( .A(n5773), .B(n5772), .Z(n5774) );
  NAND U6182 ( .A(n5775), .B(n5774), .Z(n5777) );
  XOR U6183 ( .A(n5776), .B(n5777), .Z(n5778) );
  NANDN U6184 ( .A(n525), .B(n[138]), .Z(n5779) );
  XOR U6185 ( .A(n5778), .B(n5779), .Z(zout[138]) );
  NAND U6186 ( .A(n5777), .B(n5776), .Z(n5781) );
  NANDN U6187 ( .A(n5779), .B(n5778), .Z(n5780) );
  NAND U6188 ( .A(n5781), .B(n5780), .Z(n5784) );
  XOR U6189 ( .A(n5783), .B(n5784), .Z(n5785) );
  NANDN U6190 ( .A(n525), .B(n[139]), .Z(n5786) );
  XOR U6191 ( .A(n5785), .B(n5786), .Z(zout[139]) );
  AND U6192 ( .A(n6814), .B(n[13]), .Z(n5847) );
  XNOR U6193 ( .A(n5846), .B(n5847), .Z(n5844) );
  NOR U6194 ( .A(n525), .B(n5782), .Z(n5845) );
  XOR U6195 ( .A(n5844), .B(n5845), .Z(zout[13]) );
  NANDN U6196 ( .A(n525), .B(n[140]), .Z(n5790) );
  XOR U6197 ( .A(n5789), .B(n5790), .Z(n5792) );
  NAND U6198 ( .A(n5784), .B(n5783), .Z(n5788) );
  NANDN U6199 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U6200 ( .A(n5788), .B(n5787), .Z(n5791) );
  XNOR U6201 ( .A(n5792), .B(n5791), .Z(zout[140]) );
  AND U6202 ( .A(n[141]), .B(n6814), .Z(n5798) );
  NANDN U6203 ( .A(n5790), .B(n5789), .Z(n5794) );
  OR U6204 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6205 ( .A(n5794), .B(n5793), .Z(n5797) );
  XNOR U6206 ( .A(n5796), .B(n5797), .Z(n5795) );
  XOR U6207 ( .A(n5798), .B(n5795), .Z(zout[141]) );
  NANDN U6208 ( .A(n525), .B(n[142]), .Z(n5799) );
  XOR U6209 ( .A(n5800), .B(n5799), .Z(n5802) );
  XNOR U6210 ( .A(n5803), .B(n5802), .Z(zout[142]) );
  AND U6211 ( .A(n5800), .B(n[142]), .Z(n5801) );
  NANDN U6212 ( .A(n525), .B(n5801), .Z(n5805) );
  OR U6213 ( .A(n5803), .B(n5802), .Z(n5804) );
  NAND U6214 ( .A(n5805), .B(n5804), .Z(n5807) );
  XOR U6215 ( .A(n5806), .B(n5807), .Z(n5808) );
  NANDN U6216 ( .A(n525), .B(n[143]), .Z(n5809) );
  XOR U6217 ( .A(n5808), .B(n5809), .Z(zout[143]) );
  NANDN U6218 ( .A(n525), .B(n[144]), .Z(n5814) );
  XOR U6219 ( .A(n5813), .B(n5814), .Z(n5816) );
  NAND U6220 ( .A(n5807), .B(n5806), .Z(n5811) );
  NANDN U6221 ( .A(n5809), .B(n5808), .Z(n5810) );
  AND U6222 ( .A(n5811), .B(n5810), .Z(n5815) );
  XNOR U6223 ( .A(n5816), .B(n5815), .Z(zout[144]) );
  NANDN U6224 ( .A(n525), .B(n[145]), .Z(n5812) );
  XOR U6225 ( .A(n5820), .B(n5812), .Z(n5823) );
  NANDN U6226 ( .A(n5814), .B(n5813), .Z(n5818) );
  OR U6227 ( .A(n5816), .B(n5815), .Z(n5817) );
  AND U6228 ( .A(n5818), .B(n5817), .Z(n5822) );
  XNOR U6229 ( .A(n5823), .B(n5822), .Z(zout[145]) );
  NANDN U6230 ( .A(n525), .B(n[146]), .Z(n5819) );
  XOR U6231 ( .A(n5826), .B(n5819), .Z(n5829) );
  AND U6232 ( .A(n5820), .B(n[145]), .Z(n5821) );
  NANDN U6233 ( .A(n525), .B(n5821), .Z(n5825) );
  OR U6234 ( .A(n5823), .B(n5822), .Z(n5824) );
  AND U6235 ( .A(n5825), .B(n5824), .Z(n5828) );
  XNOR U6236 ( .A(n5829), .B(n5828), .Z(zout[146]) );
  NANDN U6237 ( .A(n525), .B(n[147]), .Z(n5833) );
  XOR U6238 ( .A(n5832), .B(n5833), .Z(n5835) );
  AND U6239 ( .A(n5826), .B(n[146]), .Z(n5827) );
  NANDN U6240 ( .A(n525), .B(n5827), .Z(n5831) );
  OR U6241 ( .A(n5829), .B(n5828), .Z(n5830) );
  AND U6242 ( .A(n5831), .B(n5830), .Z(n5834) );
  XNOR U6243 ( .A(n5835), .B(n5834), .Z(zout[147]) );
  NANDN U6244 ( .A(n525), .B(n[148]), .Z(n5839) );
  XOR U6245 ( .A(n5838), .B(n5839), .Z(n5841) );
  NANDN U6246 ( .A(n5833), .B(n5832), .Z(n5837) );
  OR U6247 ( .A(n5835), .B(n5834), .Z(n5836) );
  AND U6248 ( .A(n5837), .B(n5836), .Z(n5840) );
  XNOR U6249 ( .A(n5841), .B(n5840), .Z(zout[148]) );
  NANDN U6250 ( .A(n525), .B(n[149]), .Z(n5855) );
  XOR U6251 ( .A(n5854), .B(n5855), .Z(n5857) );
  NANDN U6252 ( .A(n5839), .B(n5838), .Z(n5843) );
  OR U6253 ( .A(n5841), .B(n5840), .Z(n5842) );
  AND U6254 ( .A(n5843), .B(n5842), .Z(n5856) );
  XNOR U6255 ( .A(n5857), .B(n5856), .Z(zout[149]) );
  OR U6256 ( .A(n5845), .B(n5844), .Z(n5849) );
  OR U6257 ( .A(n5847), .B(n5846), .Z(n5848) );
  AND U6258 ( .A(n5849), .B(n5848), .Z(n5851) );
  NANDN U6259 ( .A(n525), .B(n[14]), .Z(n5850) );
  XNOR U6260 ( .A(n5851), .B(n5850), .Z(n5852) );
  XNOR U6261 ( .A(n5853), .B(n5852), .Z(zout[14]) );
  NANDN U6262 ( .A(n525), .B(n[150]), .Z(n5863) );
  NANDN U6263 ( .A(n5855), .B(n5854), .Z(n5859) );
  OR U6264 ( .A(n5857), .B(n5856), .Z(n5858) );
  AND U6265 ( .A(n5859), .B(n5858), .Z(n5862) );
  XOR U6266 ( .A(n5861), .B(n5862), .Z(n5860) );
  XNOR U6267 ( .A(n5863), .B(n5860), .Z(zout[150]) );
  NANDN U6268 ( .A(n525), .B(n[151]), .Z(n5864) );
  XOR U6269 ( .A(n5866), .B(n5864), .Z(n5869) );
  XOR U6270 ( .A(n5868), .B(n5869), .Z(zout[151]) );
  NANDN U6271 ( .A(n525), .B(n[152]), .Z(n5865) );
  XOR U6272 ( .A(n5872), .B(n5865), .Z(n5875) );
  AND U6273 ( .A(n5866), .B(n[151]), .Z(n5867) );
  NANDN U6274 ( .A(n525), .B(n5867), .Z(n5871) );
  NANDN U6275 ( .A(n5869), .B(n5868), .Z(n5870) );
  AND U6276 ( .A(n5871), .B(n5870), .Z(n5874) );
  XNOR U6277 ( .A(n5875), .B(n5874), .Z(zout[152]) );
  NANDN U6278 ( .A(n525), .B(n[153]), .Z(n5881) );
  AND U6279 ( .A(n5872), .B(n[152]), .Z(n5873) );
  NANDN U6280 ( .A(n525), .B(n5873), .Z(n5877) );
  OR U6281 ( .A(n5875), .B(n5874), .Z(n5876) );
  AND U6282 ( .A(n5877), .B(n5876), .Z(n5880) );
  XOR U6283 ( .A(n5879), .B(n5880), .Z(n5878) );
  XNOR U6284 ( .A(n5881), .B(n5878), .Z(zout[153]) );
  NANDN U6285 ( .A(n525), .B(n[154]), .Z(n5882) );
  XOR U6286 ( .A(n5883), .B(n5882), .Z(n5886) );
  XOR U6287 ( .A(n5885), .B(n5886), .Z(zout[154]) );
  NANDN U6288 ( .A(n525), .B(n[155]), .Z(n5893) );
  XOR U6289 ( .A(n5892), .B(n5893), .Z(n5895) );
  AND U6290 ( .A(n5883), .B(n[154]), .Z(n5884) );
  NANDN U6291 ( .A(n525), .B(n5884), .Z(n5888) );
  NANDN U6292 ( .A(n5886), .B(n5885), .Z(n5887) );
  AND U6293 ( .A(n5888), .B(n5887), .Z(n5894) );
  XNOR U6294 ( .A(n5895), .B(n5894), .Z(zout[155]) );
  NANDN U6295 ( .A(n5889), .B(n6814), .Z(n5890) );
  XOR U6296 ( .A(n5891), .B(n5890), .Z(n5899) );
  NANDN U6297 ( .A(n5893), .B(n5892), .Z(n5897) );
  OR U6298 ( .A(n5895), .B(n5894), .Z(n5896) );
  AND U6299 ( .A(n5897), .B(n5896), .Z(n5900) );
  XOR U6300 ( .A(n5899), .B(n5900), .Z(zout[156]) );
  NANDN U6301 ( .A(n525), .B(n[157]), .Z(n5907) );
  XOR U6302 ( .A(n5906), .B(n5907), .Z(n5909) );
  OR U6303 ( .A(n5898), .B(n525), .Z(n5902) );
  NANDN U6304 ( .A(n5900), .B(n5899), .Z(n5901) );
  AND U6305 ( .A(n5902), .B(n5901), .Z(n5908) );
  XNOR U6306 ( .A(n5909), .B(n5908), .Z(zout[157]) );
  NANDN U6307 ( .A(n5903), .B(n6814), .Z(n5904) );
  XNOR U6308 ( .A(n5905), .B(n5904), .Z(n5913) );
  NANDN U6309 ( .A(n5907), .B(n5906), .Z(n5911) );
  OR U6310 ( .A(n5909), .B(n5908), .Z(n5910) );
  AND U6311 ( .A(n5911), .B(n5910), .Z(n5914) );
  XOR U6312 ( .A(n5913), .B(n5914), .Z(zout[158]) );
  NANDN U6313 ( .A(n525), .B(n5912), .Z(n5916) );
  NANDN U6314 ( .A(n5914), .B(n5913), .Z(n5915) );
  NAND U6315 ( .A(n5916), .B(n5915), .Z(n5920) );
  AND U6316 ( .A(n[159]), .B(n6814), .Z(n5921) );
  XOR U6317 ( .A(n5919), .B(n5921), .Z(n5917) );
  XNOR U6318 ( .A(n5920), .B(n5917), .Z(zout[159]) );
  AND U6319 ( .A(n6814), .B(n[15]), .Z(n5979) );
  XNOR U6320 ( .A(n5978), .B(n5979), .Z(n5976) );
  AND U6321 ( .A(n6814), .B(n5918), .Z(n5977) );
  XOR U6322 ( .A(n5976), .B(n5977), .Z(zout[15]) );
  NANDN U6323 ( .A(n525), .B(n[160]), .Z(n5923) );
  XNOR U6324 ( .A(n5924), .B(n5925), .Z(n5922) );
  XNOR U6325 ( .A(n5923), .B(n5922), .Z(zout[160]) );
  AND U6326 ( .A(n[161]), .B(n6814), .Z(n5929) );
  XNOR U6327 ( .A(n5928), .B(n5927), .Z(n5926) );
  XNOR U6328 ( .A(n5929), .B(n5926), .Z(zout[161]) );
  NANDN U6329 ( .A(n525), .B(n[162]), .Z(n5932) );
  XOR U6330 ( .A(n5931), .B(n5932), .Z(n5934) );
  XNOR U6331 ( .A(n5933), .B(n5934), .Z(zout[162]) );
  NANDN U6332 ( .A(n525), .B(n[163]), .Z(n5930) );
  XOR U6333 ( .A(n5937), .B(n5930), .Z(n5940) );
  NANDN U6334 ( .A(n5932), .B(n5931), .Z(n5936) );
  OR U6335 ( .A(n5934), .B(n5933), .Z(n5935) );
  AND U6336 ( .A(n5936), .B(n5935), .Z(n5939) );
  XNOR U6337 ( .A(n5940), .B(n5939), .Z(zout[163]) );
  AND U6338 ( .A(n5937), .B(n[163]), .Z(n5938) );
  NANDN U6339 ( .A(n525), .B(n5938), .Z(n5942) );
  OR U6340 ( .A(n5940), .B(n5939), .Z(n5941) );
  NAND U6341 ( .A(n5942), .B(n5941), .Z(n5946) );
  XOR U6342 ( .A(n5945), .B(n5946), .Z(n5947) );
  NANDN U6343 ( .A(n5943), .B(n6814), .Z(n5948) );
  XOR U6344 ( .A(n5947), .B(n5948), .Z(zout[164]) );
  NANDN U6345 ( .A(n525), .B(n[165]), .Z(n5944) );
  XOR U6346 ( .A(n5951), .B(n5944), .Z(n5954) );
  NAND U6347 ( .A(n5946), .B(n5945), .Z(n5950) );
  NANDN U6348 ( .A(n5948), .B(n5947), .Z(n5949) );
  AND U6349 ( .A(n5950), .B(n5949), .Z(n5953) );
  XNOR U6350 ( .A(n5954), .B(n5953), .Z(zout[165]) );
  NANDN U6351 ( .A(n525), .B(n[166]), .Z(n5959) );
  XOR U6352 ( .A(n5958), .B(n5959), .Z(n5961) );
  AND U6353 ( .A(n5951), .B(n[165]), .Z(n5952) );
  NANDN U6354 ( .A(n525), .B(n5952), .Z(n5956) );
  OR U6355 ( .A(n5954), .B(n5953), .Z(n5955) );
  AND U6356 ( .A(n5956), .B(n5955), .Z(n5960) );
  XNOR U6357 ( .A(n5961), .B(n5960), .Z(zout[166]) );
  NANDN U6358 ( .A(n525), .B(n[167]), .Z(n5957) );
  XOR U6359 ( .A(n5964), .B(n5957), .Z(n5967) );
  NANDN U6360 ( .A(n5959), .B(n5958), .Z(n5963) );
  OR U6361 ( .A(n5961), .B(n5960), .Z(n5962) );
  AND U6362 ( .A(n5963), .B(n5962), .Z(n5966) );
  XNOR U6363 ( .A(n5967), .B(n5966), .Z(zout[167]) );
  NANDN U6364 ( .A(n525), .B(n[168]), .Z(n5971) );
  XOR U6365 ( .A(n5970), .B(n5971), .Z(n5973) );
  AND U6366 ( .A(n5964), .B(n[167]), .Z(n5965) );
  NANDN U6367 ( .A(n525), .B(n5965), .Z(n5969) );
  OR U6368 ( .A(n5967), .B(n5966), .Z(n5968) );
  AND U6369 ( .A(n5969), .B(n5968), .Z(n5972) );
  XNOR U6370 ( .A(n5973), .B(n5972), .Z(zout[168]) );
  NANDN U6371 ( .A(n5971), .B(n5970), .Z(n5975) );
  OR U6372 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U6373 ( .A(n5975), .B(n5974), .Z(n5987) );
  XOR U6374 ( .A(n5986), .B(n5987), .Z(n5988) );
  NANDN U6375 ( .A(n525), .B(n[169]), .Z(n5989) );
  XOR U6376 ( .A(n5988), .B(n5989), .Z(zout[169]) );
  OR U6377 ( .A(n5977), .B(n5976), .Z(n5981) );
  OR U6378 ( .A(n5979), .B(n5978), .Z(n5980) );
  AND U6379 ( .A(n5981), .B(n5980), .Z(n5983) );
  NANDN U6380 ( .A(n525), .B(n[16]), .Z(n5982) );
  XNOR U6381 ( .A(n5983), .B(n5982), .Z(n5984) );
  XNOR U6382 ( .A(n5985), .B(n5984), .Z(zout[16]) );
  AND U6383 ( .A(n6814), .B(n[170]), .Z(n5996) );
  NAND U6384 ( .A(n5987), .B(n5986), .Z(n5991) );
  NANDN U6385 ( .A(n5989), .B(n5988), .Z(n5990) );
  AND U6386 ( .A(n5991), .B(n5990), .Z(n5995) );
  XNOR U6387 ( .A(n5993), .B(n5995), .Z(n5992) );
  XOR U6388 ( .A(n5996), .B(n5992), .Z(zout[170]) );
  NANDN U6389 ( .A(n5998), .B(n6814), .Z(n5997) );
  XOR U6390 ( .A(n5999), .B(n5997), .Z(n6001) );
  XNOR U6391 ( .A(n6002), .B(n6001), .Z(zout[171]) );
  NANDN U6392 ( .A(n525), .B(n[172]), .Z(n6006) );
  XOR U6393 ( .A(n6005), .B(n6006), .Z(n6008) );
  ANDN U6394 ( .B(n5999), .A(n5998), .Z(n6000) );
  NANDN U6395 ( .A(n525), .B(n6000), .Z(n6004) );
  OR U6396 ( .A(n6002), .B(n6001), .Z(n6003) );
  AND U6397 ( .A(n6004), .B(n6003), .Z(n6007) );
  XNOR U6398 ( .A(n6008), .B(n6007), .Z(zout[172]) );
  NANDN U6399 ( .A(n525), .B(n[173]), .Z(n6013) );
  XOR U6400 ( .A(n6012), .B(n6013), .Z(n6015) );
  NANDN U6401 ( .A(n6006), .B(n6005), .Z(n6010) );
  OR U6402 ( .A(n6008), .B(n6007), .Z(n6009) );
  AND U6403 ( .A(n6010), .B(n6009), .Z(n6014) );
  XNOR U6404 ( .A(n6015), .B(n6014), .Z(zout[173]) );
  NANDN U6405 ( .A(n525), .B(n[174]), .Z(n6011) );
  XOR U6406 ( .A(n6018), .B(n6011), .Z(n6021) );
  NANDN U6407 ( .A(n6013), .B(n6012), .Z(n6017) );
  OR U6408 ( .A(n6015), .B(n6014), .Z(n6016) );
  AND U6409 ( .A(n6017), .B(n6016), .Z(n6020) );
  XNOR U6410 ( .A(n6021), .B(n6020), .Z(zout[174]) );
  AND U6411 ( .A(n6018), .B(n[174]), .Z(n6019) );
  NANDN U6412 ( .A(n525), .B(n6019), .Z(n6023) );
  OR U6413 ( .A(n6021), .B(n6020), .Z(n6022) );
  NAND U6414 ( .A(n6023), .B(n6022), .Z(n6027) );
  XOR U6415 ( .A(n6026), .B(n6027), .Z(n6028) );
  NANDN U6416 ( .A(n6024), .B(n6814), .Z(n6029) );
  XOR U6417 ( .A(n6028), .B(n6029), .Z(zout[175]) );
  NANDN U6418 ( .A(n6025), .B(n6814), .Z(n6032) );
  XOR U6419 ( .A(n6033), .B(n6032), .Z(n6034) );
  NAND U6420 ( .A(n6027), .B(n6026), .Z(n6031) );
  NANDN U6421 ( .A(n6029), .B(n6028), .Z(n6030) );
  NAND U6422 ( .A(n6031), .B(n6030), .Z(n6035) );
  XNOR U6423 ( .A(n6034), .B(n6035), .Z(zout[176]) );
  AND U6424 ( .A(n6033), .B(n6032), .Z(n6037) );
  NANDN U6425 ( .A(n6035), .B(n6034), .Z(n6036) );
  NANDN U6426 ( .A(n6037), .B(n6036), .Z(n6046) );
  NANDN U6427 ( .A(n525), .B(n[177]), .Z(n6038) );
  XOR U6428 ( .A(n6043), .B(n6038), .Z(n6045) );
  XNOR U6429 ( .A(n6046), .B(n6045), .Z(zout[177]) );
  NANDN U6430 ( .A(n6039), .B(n6814), .Z(n6040) );
  XOR U6431 ( .A(n6041), .B(n6040), .Z(n6050) );
  ANDN U6432 ( .B(n6043), .A(n6042), .Z(n6044) );
  NANDN U6433 ( .A(n525), .B(n6044), .Z(n6048) );
  OR U6434 ( .A(n6046), .B(n6045), .Z(n6047) );
  AND U6435 ( .A(n6048), .B(n6047), .Z(n6051) );
  XOR U6436 ( .A(n6050), .B(n6051), .Z(zout[178]) );
  NANDN U6437 ( .A(n525), .B(n[179]), .Z(n6056) );
  XOR U6438 ( .A(n6055), .B(n6056), .Z(n6058) );
  OR U6439 ( .A(n6049), .B(n525), .Z(n6053) );
  NANDN U6440 ( .A(n6051), .B(n6050), .Z(n6052) );
  AND U6441 ( .A(n6053), .B(n6052), .Z(n6057) );
  XNOR U6442 ( .A(n6058), .B(n6057), .Z(zout[179]) );
  NOR U6443 ( .A(n525), .B(n6054), .Z(n6123) );
  XNOR U6444 ( .A(n6122), .B(n6123), .Z(n6120) );
  AND U6445 ( .A(n6814), .B(n[17]), .Z(n6121) );
  XOR U6446 ( .A(n6120), .B(n6121), .Z(zout[17]) );
  NANDN U6447 ( .A(n6056), .B(n6055), .Z(n6060) );
  OR U6448 ( .A(n6058), .B(n6057), .Z(n6059) );
  NAND U6449 ( .A(n6060), .B(n6059), .Z(n6062) );
  XOR U6450 ( .A(n6061), .B(n6062), .Z(n6063) );
  NANDN U6451 ( .A(n525), .B(n[180]), .Z(n6064) );
  XOR U6452 ( .A(n6063), .B(n6064), .Z(zout[180]) );
  NANDN U6453 ( .A(n525), .B(n[181]), .Z(n6068) );
  XOR U6454 ( .A(n6067), .B(n6068), .Z(n6070) );
  NAND U6455 ( .A(n6062), .B(n6061), .Z(n6066) );
  NANDN U6456 ( .A(n6064), .B(n6063), .Z(n6065) );
  AND U6457 ( .A(n6066), .B(n6065), .Z(n6069) );
  XNOR U6458 ( .A(n6070), .B(n6069), .Z(zout[181]) );
  NANDN U6459 ( .A(n525), .B(n[182]), .Z(n6074) );
  XOR U6460 ( .A(n6073), .B(n6074), .Z(n6076) );
  NANDN U6461 ( .A(n6068), .B(n6067), .Z(n6072) );
  OR U6462 ( .A(n6070), .B(n6069), .Z(n6071) );
  AND U6463 ( .A(n6072), .B(n6071), .Z(n6075) );
  XNOR U6464 ( .A(n6076), .B(n6075), .Z(zout[182]) );
  NANDN U6465 ( .A(n525), .B(n[183]), .Z(n6081) );
  XOR U6466 ( .A(n6080), .B(n6081), .Z(n6083) );
  NANDN U6467 ( .A(n6074), .B(n6073), .Z(n6078) );
  OR U6468 ( .A(n6076), .B(n6075), .Z(n6077) );
  AND U6469 ( .A(n6078), .B(n6077), .Z(n6082) );
  XNOR U6470 ( .A(n6083), .B(n6082), .Z(zout[183]) );
  NANDN U6471 ( .A(n6086), .B(n6814), .Z(n6079) );
  XOR U6472 ( .A(n6087), .B(n6079), .Z(n6090) );
  NANDN U6473 ( .A(n6081), .B(n6080), .Z(n6085) );
  OR U6474 ( .A(n6083), .B(n6082), .Z(n6084) );
  AND U6475 ( .A(n6085), .B(n6084), .Z(n6089) );
  XNOR U6476 ( .A(n6090), .B(n6089), .Z(zout[184]) );
  ANDN U6477 ( .B(n6087), .A(n6086), .Z(n6088) );
  NANDN U6478 ( .A(n525), .B(n6088), .Z(n6092) );
  OR U6479 ( .A(n6090), .B(n6089), .Z(n6091) );
  NAND U6480 ( .A(n6092), .B(n6091), .Z(n6094) );
  XOR U6481 ( .A(n6093), .B(n6094), .Z(n6095) );
  NANDN U6482 ( .A(n525), .B(n[185]), .Z(n6096) );
  XOR U6483 ( .A(n6095), .B(n6096), .Z(zout[185]) );
  NANDN U6484 ( .A(n525), .B(n[186]), .Z(n6101) );
  XOR U6485 ( .A(n6100), .B(n6101), .Z(n6103) );
  NAND U6486 ( .A(n6094), .B(n6093), .Z(n6098) );
  NANDN U6487 ( .A(n6096), .B(n6095), .Z(n6097) );
  AND U6488 ( .A(n6098), .B(n6097), .Z(n6102) );
  XNOR U6489 ( .A(n6103), .B(n6102), .Z(zout[186]) );
  NANDN U6490 ( .A(n6106), .B(n6814), .Z(n6099) );
  XOR U6491 ( .A(n6107), .B(n6099), .Z(n6110) );
  NANDN U6492 ( .A(n6101), .B(n6100), .Z(n6105) );
  OR U6493 ( .A(n6103), .B(n6102), .Z(n6104) );
  AND U6494 ( .A(n6105), .B(n6104), .Z(n6109) );
  XNOR U6495 ( .A(n6110), .B(n6109), .Z(zout[187]) );
  NANDN U6496 ( .A(n525), .B(n[188]), .Z(n6114) );
  XOR U6497 ( .A(n6113), .B(n6114), .Z(n6116) );
  ANDN U6498 ( .B(n6107), .A(n6106), .Z(n6108) );
  NANDN U6499 ( .A(n525), .B(n6108), .Z(n6112) );
  OR U6500 ( .A(n6110), .B(n6109), .Z(n6111) );
  AND U6501 ( .A(n6112), .B(n6111), .Z(n6115) );
  XNOR U6502 ( .A(n6116), .B(n6115), .Z(zout[188]) );
  NANDN U6503 ( .A(n6114), .B(n6113), .Z(n6118) );
  OR U6504 ( .A(n6116), .B(n6115), .Z(n6117) );
  NAND U6505 ( .A(n6118), .B(n6117), .Z(n6131) );
  AND U6506 ( .A(n6814), .B(n[189]), .Z(n6132) );
  XOR U6507 ( .A(n6130), .B(n6132), .Z(n6119) );
  XNOR U6508 ( .A(n6131), .B(n6119), .Z(zout[189]) );
  OR U6509 ( .A(n6121), .B(n6120), .Z(n6125) );
  OR U6510 ( .A(n6123), .B(n6122), .Z(n6124) );
  AND U6511 ( .A(n6125), .B(n6124), .Z(n6127) );
  NANDN U6512 ( .A(n525), .B(n[18]), .Z(n6126) );
  XNOR U6513 ( .A(n6127), .B(n6126), .Z(n6128) );
  XNOR U6514 ( .A(n6129), .B(n6128), .Z(zout[18]) );
  NANDN U6515 ( .A(n525), .B(n[190]), .Z(n6133) );
  XOR U6516 ( .A(n6136), .B(n6133), .Z(n6138) );
  XNOR U6517 ( .A(n6139), .B(n6138), .Z(zout[190]) );
  NANDN U6518 ( .A(n525), .B(n[191]), .Z(n6134) );
  XOR U6519 ( .A(n6142), .B(n6134), .Z(n6145) );
  ANDN U6520 ( .B(n6136), .A(n6135), .Z(n6137) );
  NANDN U6521 ( .A(n525), .B(n6137), .Z(n6141) );
  OR U6522 ( .A(n6139), .B(n6138), .Z(n6140) );
  AND U6523 ( .A(n6141), .B(n6140), .Z(n6144) );
  XNOR U6524 ( .A(n6145), .B(n6144), .Z(zout[191]) );
  NANDN U6525 ( .A(n525), .B(n[192]), .Z(n6149) );
  XOR U6526 ( .A(n6148), .B(n6149), .Z(n6151) );
  AND U6527 ( .A(n6142), .B(n[191]), .Z(n6143) );
  NANDN U6528 ( .A(n525), .B(n6143), .Z(n6147) );
  OR U6529 ( .A(n6145), .B(n6144), .Z(n6146) );
  AND U6530 ( .A(n6147), .B(n6146), .Z(n6150) );
  XNOR U6531 ( .A(n6151), .B(n6150), .Z(zout[192]) );
  NANDN U6532 ( .A(n525), .B(n[193]), .Z(n6155) );
  XOR U6533 ( .A(n6154), .B(n6155), .Z(n6157) );
  NANDN U6534 ( .A(n6149), .B(n6148), .Z(n6153) );
  OR U6535 ( .A(n6151), .B(n6150), .Z(n6152) );
  AND U6536 ( .A(n6153), .B(n6152), .Z(n6156) );
  XNOR U6537 ( .A(n6157), .B(n6156), .Z(zout[193]) );
  NANDN U6538 ( .A(n525), .B(n[194]), .Z(n6161) );
  XOR U6539 ( .A(n6160), .B(n6161), .Z(n6163) );
  NANDN U6540 ( .A(n6155), .B(n6154), .Z(n6159) );
  OR U6541 ( .A(n6157), .B(n6156), .Z(n6158) );
  AND U6542 ( .A(n6159), .B(n6158), .Z(n6162) );
  XNOR U6543 ( .A(n6163), .B(n6162), .Z(zout[194]) );
  NANDN U6544 ( .A(n525), .B(n[195]), .Z(n6170) );
  XOR U6545 ( .A(n6169), .B(n6170), .Z(n6172) );
  NANDN U6546 ( .A(n6161), .B(n6160), .Z(n6165) );
  OR U6547 ( .A(n6163), .B(n6162), .Z(n6164) );
  AND U6548 ( .A(n6165), .B(n6164), .Z(n6171) );
  XNOR U6549 ( .A(n6172), .B(n6171), .Z(zout[195]) );
  NANDN U6550 ( .A(n6166), .B(n6814), .Z(n6167) );
  XNOR U6551 ( .A(n6168), .B(n6167), .Z(n6176) );
  NANDN U6552 ( .A(n6170), .B(n6169), .Z(n6174) );
  OR U6553 ( .A(n6172), .B(n6171), .Z(n6173) );
  AND U6554 ( .A(n6174), .B(n6173), .Z(n6177) );
  XOR U6555 ( .A(n6176), .B(n6177), .Z(zout[196]) );
  NANDN U6556 ( .A(n525), .B(n[197]), .Z(n6182) );
  XOR U6557 ( .A(n6181), .B(n6182), .Z(n6184) );
  OR U6558 ( .A(n6175), .B(n525), .Z(n6179) );
  NANDN U6559 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U6560 ( .A(n6179), .B(n6178), .Z(n6183) );
  XNOR U6561 ( .A(n6184), .B(n6183), .Z(zout[197]) );
  NANDN U6562 ( .A(n525), .B(n[198]), .Z(n6180) );
  XOR U6563 ( .A(n6188), .B(n6180), .Z(n6191) );
  NANDN U6564 ( .A(n6182), .B(n6181), .Z(n6186) );
  OR U6565 ( .A(n6184), .B(n6183), .Z(n6185) );
  AND U6566 ( .A(n6186), .B(n6185), .Z(n6190) );
  XNOR U6567 ( .A(n6191), .B(n6190), .Z(zout[198]) );
  NANDN U6568 ( .A(n525), .B(n[199]), .Z(n6187) );
  XOR U6569 ( .A(n6202), .B(n6187), .Z(n6205) );
  AND U6570 ( .A(n6188), .B(n[198]), .Z(n6189) );
  NANDN U6571 ( .A(n525), .B(n6189), .Z(n6193) );
  OR U6572 ( .A(n6191), .B(n6190), .Z(n6192) );
  AND U6573 ( .A(n6193), .B(n6192), .Z(n6204) );
  XNOR U6574 ( .A(n6205), .B(n6204), .Z(zout[199]) );
  AND U6575 ( .A(n6814), .B(n[19]), .Z(n6261) );
  XNOR U6576 ( .A(n6260), .B(n6261), .Z(n6258) );
  NOR U6577 ( .A(n525), .B(n6194), .Z(n6259) );
  XOR U6578 ( .A(n6258), .B(n6259), .Z(zout[19]) );
  XOR U6579 ( .A(n[1]), .B(n6195), .Z(n6196) );
  NANDN U6580 ( .A(n525), .B(n6196), .Z(n6197) );
  XNOR U6581 ( .A(n6198), .B(n6197), .Z(zout[1]) );
  NANDN U6582 ( .A(n6199), .B(n6814), .Z(n6200) );
  XNOR U6583 ( .A(n6201), .B(n6200), .Z(n6209) );
  AND U6584 ( .A(n6202), .B(n[199]), .Z(n6203) );
  NANDN U6585 ( .A(n525), .B(n6203), .Z(n6207) );
  OR U6586 ( .A(n6205), .B(n6204), .Z(n6206) );
  AND U6587 ( .A(n6207), .B(n6206), .Z(n6210) );
  XOR U6588 ( .A(n6209), .B(n6210), .Z(zout[200]) );
  NANDN U6589 ( .A(n525), .B(n[201]), .Z(n6214) );
  XOR U6590 ( .A(n6213), .B(n6214), .Z(n6216) );
  OR U6591 ( .A(n6208), .B(n525), .Z(n6212) );
  NANDN U6592 ( .A(n6210), .B(n6209), .Z(n6211) );
  AND U6593 ( .A(n6212), .B(n6211), .Z(n6215) );
  XNOR U6594 ( .A(n6216), .B(n6215), .Z(zout[201]) );
  NANDN U6595 ( .A(n6214), .B(n6213), .Z(n6218) );
  OR U6596 ( .A(n6216), .B(n6215), .Z(n6217) );
  NAND U6597 ( .A(n6218), .B(n6217), .Z(n6220) );
  XOR U6598 ( .A(n6219), .B(n6220), .Z(n6221) );
  NANDN U6599 ( .A(n525), .B(n[202]), .Z(n6222) );
  XOR U6600 ( .A(n6221), .B(n6222), .Z(zout[202]) );
  NAND U6601 ( .A(n6220), .B(n6219), .Z(n6224) );
  NANDN U6602 ( .A(n6222), .B(n6221), .Z(n6223) );
  NAND U6603 ( .A(n6224), .B(n6223), .Z(n6227) );
  XOR U6604 ( .A(n6226), .B(n6227), .Z(n6228) );
  NANDN U6605 ( .A(n6225), .B(n6814), .Z(n6229) );
  XOR U6606 ( .A(n6228), .B(n6229), .Z(zout[203]) );
  NANDN U6607 ( .A(n525), .B(n[204]), .Z(n6233) );
  XOR U6608 ( .A(n6232), .B(n6233), .Z(n6235) );
  NAND U6609 ( .A(n6227), .B(n6226), .Z(n6231) );
  NANDN U6610 ( .A(n6229), .B(n6228), .Z(n6230) );
  AND U6611 ( .A(n6231), .B(n6230), .Z(n6234) );
  XNOR U6612 ( .A(n6235), .B(n6234), .Z(zout[204]) );
  NANDN U6613 ( .A(n6233), .B(n6232), .Z(n6237) );
  OR U6614 ( .A(n6235), .B(n6234), .Z(n6236) );
  NAND U6615 ( .A(n6237), .B(n6236), .Z(n6240) );
  AND U6616 ( .A(n[205]), .B(n6814), .Z(n6241) );
  XOR U6617 ( .A(n6239), .B(n6241), .Z(n6238) );
  XNOR U6618 ( .A(n6240), .B(n6238), .Z(zout[205]) );
  NANDN U6619 ( .A(n525), .B(n[206]), .Z(n6243) );
  XOR U6620 ( .A(n6242), .B(n6243), .Z(n6245) );
  XNOR U6621 ( .A(n6244), .B(n6245), .Z(zout[206]) );
  NANDN U6622 ( .A(n525), .B(n[207]), .Z(n6251) );
  NANDN U6623 ( .A(n6243), .B(n6242), .Z(n6247) );
  OR U6624 ( .A(n6245), .B(n6244), .Z(n6246) );
  AND U6625 ( .A(n6247), .B(n6246), .Z(n6250) );
  XOR U6626 ( .A(n6249), .B(n6250), .Z(n6248) );
  XNOR U6627 ( .A(n6251), .B(n6248), .Z(zout[207]) );
  AND U6628 ( .A(n6814), .B(n[208]), .Z(n6255) );
  XNOR U6629 ( .A(n6254), .B(n6253), .Z(n6252) );
  XNOR U6630 ( .A(n6255), .B(n6252), .Z(zout[208]) );
  NANDN U6631 ( .A(n6256), .B(n6814), .Z(n6257) );
  XOR U6632 ( .A(n6271), .B(n6257), .Z(n6273) );
  XOR U6633 ( .A(n6274), .B(n6273), .Z(zout[209]) );
  OR U6634 ( .A(n6259), .B(n6258), .Z(n6263) );
  OR U6635 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U6636 ( .A(n6263), .B(n6262), .Z(n6265) );
  NANDN U6637 ( .A(n525), .B(n[20]), .Z(n6264) );
  XNOR U6638 ( .A(n6265), .B(n6264), .Z(n6266) );
  XNOR U6639 ( .A(n6267), .B(n6266), .Z(zout[20]) );
  NANDN U6640 ( .A(n6268), .B(n6814), .Z(n6269) );
  XNOR U6641 ( .A(n6270), .B(n6269), .Z(n6279) );
  ANDN U6642 ( .B(n[209]), .A(n6271), .Z(n6272) );
  NANDN U6643 ( .A(n525), .B(n6272), .Z(n6276) );
  NANDN U6644 ( .A(n6274), .B(n6273), .Z(n6275) );
  AND U6645 ( .A(n6276), .B(n6275), .Z(n6280) );
  XOR U6646 ( .A(n6279), .B(n6280), .Z(zout[210]) );
  NANDN U6647 ( .A(n525), .B(n[211]), .Z(n6277) );
  XOR U6648 ( .A(n6283), .B(n6277), .Z(n6286) );
  NANDN U6649 ( .A(n525), .B(n6278), .Z(n6282) );
  NANDN U6650 ( .A(n6280), .B(n6279), .Z(n6281) );
  AND U6651 ( .A(n6282), .B(n6281), .Z(n6285) );
  XNOR U6652 ( .A(n6286), .B(n6285), .Z(zout[211]) );
  NANDN U6653 ( .A(n525), .B(n[212]), .Z(n6290) );
  XOR U6654 ( .A(n6289), .B(n6290), .Z(n6292) );
  AND U6655 ( .A(n6283), .B(n[211]), .Z(n6284) );
  NANDN U6656 ( .A(n525), .B(n6284), .Z(n6288) );
  OR U6657 ( .A(n6286), .B(n6285), .Z(n6287) );
  AND U6658 ( .A(n6288), .B(n6287), .Z(n6291) );
  XNOR U6659 ( .A(n6292), .B(n6291), .Z(zout[212]) );
  NANDN U6660 ( .A(n525), .B(n[213]), .Z(n6296) );
  XOR U6661 ( .A(n6295), .B(n6296), .Z(n6298) );
  NANDN U6662 ( .A(n6290), .B(n6289), .Z(n6294) );
  OR U6663 ( .A(n6292), .B(n6291), .Z(n6293) );
  AND U6664 ( .A(n6294), .B(n6293), .Z(n6297) );
  XNOR U6665 ( .A(n6298), .B(n6297), .Z(zout[213]) );
  AND U6666 ( .A(n[214]), .B(n6814), .Z(n6304) );
  NANDN U6667 ( .A(n6296), .B(n6295), .Z(n6300) );
  OR U6668 ( .A(n6298), .B(n6297), .Z(n6299) );
  AND U6669 ( .A(n6300), .B(n6299), .Z(n6303) );
  XNOR U6670 ( .A(n6302), .B(n6303), .Z(n6301) );
  XOR U6671 ( .A(n6304), .B(n6301), .Z(zout[214]) );
  NANDN U6672 ( .A(n525), .B(n[215]), .Z(n6306) );
  XOR U6673 ( .A(n6305), .B(n6306), .Z(n6308) );
  XNOR U6674 ( .A(n6307), .B(n6308), .Z(zout[215]) );
  NANDN U6675 ( .A(n525), .B(n[216]), .Z(n6312) );
  XOR U6676 ( .A(n6311), .B(n6312), .Z(n6314) );
  NANDN U6677 ( .A(n6306), .B(n6305), .Z(n6310) );
  OR U6678 ( .A(n6308), .B(n6307), .Z(n6309) );
  AND U6679 ( .A(n6310), .B(n6309), .Z(n6313) );
  XNOR U6680 ( .A(n6314), .B(n6313), .Z(zout[216]) );
  NANDN U6681 ( .A(n6312), .B(n6311), .Z(n6316) );
  OR U6682 ( .A(n6314), .B(n6313), .Z(n6315) );
  NAND U6683 ( .A(n6316), .B(n6315), .Z(n6321) );
  XOR U6684 ( .A(n6320), .B(n6321), .Z(n6322) );
  NANDN U6685 ( .A(n525), .B(n[217]), .Z(n6323) );
  XOR U6686 ( .A(n6322), .B(n6323), .Z(zout[217]) );
  NANDN U6687 ( .A(n6317), .B(n6814), .Z(n6318) );
  XNOR U6688 ( .A(n6319), .B(n6318), .Z(n6327) );
  NAND U6689 ( .A(n6321), .B(n6320), .Z(n6325) );
  NANDN U6690 ( .A(n6323), .B(n6322), .Z(n6324) );
  AND U6691 ( .A(n6325), .B(n6324), .Z(n6328) );
  XOR U6692 ( .A(n6327), .B(n6328), .Z(zout[218]) );
  NANDN U6693 ( .A(n525), .B(n[219]), .Z(n6336) );
  XOR U6694 ( .A(n6335), .B(n6336), .Z(n6338) );
  OR U6695 ( .A(n6326), .B(n525), .Z(n6330) );
  NANDN U6696 ( .A(n6328), .B(n6327), .Z(n6329) );
  AND U6697 ( .A(n6330), .B(n6329), .Z(n6337) );
  XNOR U6698 ( .A(n6338), .B(n6337), .Z(zout[219]) );
  XOR U6699 ( .A(n[21]), .B(n6331), .Z(n6332) );
  NANDN U6700 ( .A(n525), .B(n6332), .Z(n6333) );
  XOR U6701 ( .A(n6334), .B(n6333), .Z(zout[21]) );
  NANDN U6702 ( .A(n6336), .B(n6335), .Z(n6340) );
  OR U6703 ( .A(n6338), .B(n6337), .Z(n6339) );
  AND U6704 ( .A(n6340), .B(n6339), .Z(n6347) );
  AND U6705 ( .A(n6342), .B(n[220]), .Z(n6341) );
  NAND U6706 ( .A(n6814), .B(n6341), .Z(n6346) );
  NANDN U6707 ( .A(n525), .B(n[220]), .Z(n6343) );
  ANDN U6708 ( .B(n6343), .A(n6342), .Z(n6349) );
  ANDN U6709 ( .B(n6346), .A(n6349), .Z(n6344) );
  XOR U6710 ( .A(n6347), .B(n6344), .Z(zout[220]) );
  NANDN U6711 ( .A(n525), .B(n[221]), .Z(n6345) );
  XOR U6712 ( .A(n6351), .B(n6345), .Z(n6354) );
  NAND U6713 ( .A(n6347), .B(n6346), .Z(n6348) );
  NANDN U6714 ( .A(n6349), .B(n6348), .Z(n6353) );
  XNOR U6715 ( .A(n6354), .B(n6353), .Z(zout[221]) );
  NANDN U6716 ( .A(n525), .B(n[222]), .Z(n6350) );
  XOR U6717 ( .A(n6358), .B(n6350), .Z(n6361) );
  AND U6718 ( .A(n6351), .B(n[221]), .Z(n6352) );
  NANDN U6719 ( .A(n525), .B(n6352), .Z(n6356) );
  OR U6720 ( .A(n6354), .B(n6353), .Z(n6355) );
  AND U6721 ( .A(n6356), .B(n6355), .Z(n6360) );
  XNOR U6722 ( .A(n6361), .B(n6360), .Z(zout[222]) );
  ANDN U6723 ( .B(n6358), .A(n6357), .Z(n6359) );
  NANDN U6724 ( .A(n525), .B(n6359), .Z(n6363) );
  OR U6725 ( .A(n6361), .B(n6360), .Z(n6362) );
  NAND U6726 ( .A(n6363), .B(n6362), .Z(n6364) );
  XOR U6727 ( .A(n6365), .B(n6364), .Z(n6366) );
  AND U6728 ( .A(n[223]), .B(n6814), .Z(n6367) );
  XNOR U6729 ( .A(n6366), .B(n6367), .Z(zout[223]) );
  OR U6730 ( .A(n6365), .B(n6364), .Z(n6369) );
  NANDN U6731 ( .A(n6367), .B(n6366), .Z(n6368) );
  AND U6732 ( .A(n6369), .B(n6368), .Z(n6370) );
  XOR U6733 ( .A(n6371), .B(n6370), .Z(n6372) );
  AND U6734 ( .A(n[224]), .B(n6814), .Z(n6373) );
  XNOR U6735 ( .A(n6372), .B(n6373), .Z(zout[224]) );
  OR U6736 ( .A(n6371), .B(n6370), .Z(n6375) );
  NANDN U6737 ( .A(n6373), .B(n6372), .Z(n6374) );
  AND U6738 ( .A(n6375), .B(n6374), .Z(n6378) );
  XOR U6739 ( .A(n6377), .B(n6378), .Z(n6379) );
  NANDN U6740 ( .A(n6376), .B(n6814), .Z(n6380) );
  XOR U6741 ( .A(n6379), .B(n6380), .Z(zout[225]) );
  NANDN U6742 ( .A(n525), .B(n[226]), .Z(n6384) );
  XOR U6743 ( .A(n6383), .B(n6384), .Z(n6386) );
  NAND U6744 ( .A(n6378), .B(n6377), .Z(n6382) );
  NANDN U6745 ( .A(n6380), .B(n6379), .Z(n6381) );
  AND U6746 ( .A(n6382), .B(n6381), .Z(n6385) );
  XNOR U6747 ( .A(n6386), .B(n6385), .Z(zout[226]) );
  NANDN U6748 ( .A(n525), .B(n[227]), .Z(n6391) );
  XOR U6749 ( .A(n6390), .B(n6391), .Z(n6393) );
  NANDN U6750 ( .A(n6384), .B(n6383), .Z(n6388) );
  OR U6751 ( .A(n6386), .B(n6385), .Z(n6387) );
  AND U6752 ( .A(n6388), .B(n6387), .Z(n6392) );
  XNOR U6753 ( .A(n6393), .B(n6392), .Z(zout[227]) );
  NANDN U6754 ( .A(n525), .B(n[228]), .Z(n6389) );
  XOR U6755 ( .A(n6397), .B(n6389), .Z(n6400) );
  NANDN U6756 ( .A(n6391), .B(n6390), .Z(n6395) );
  OR U6757 ( .A(n6393), .B(n6392), .Z(n6394) );
  AND U6758 ( .A(n6395), .B(n6394), .Z(n6399) );
  XNOR U6759 ( .A(n6400), .B(n6399), .Z(zout[228]) );
  NANDN U6760 ( .A(n525), .B(n[229]), .Z(n6396) );
  XOR U6761 ( .A(n6407), .B(n6396), .Z(n6410) );
  AND U6762 ( .A(n6397), .B(n[228]), .Z(n6398) );
  NANDN U6763 ( .A(n525), .B(n6398), .Z(n6402) );
  OR U6764 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U6765 ( .A(n6402), .B(n6401), .Z(n6409) );
  XNOR U6766 ( .A(n6410), .B(n6409), .Z(zout[229]) );
  XNOR U6767 ( .A(n[22]), .B(n6403), .Z(n6404) );
  NANDN U6768 ( .A(n525), .B(n6404), .Z(n6405) );
  XOR U6769 ( .A(n6406), .B(n6405), .Z(zout[22]) );
  NANDN U6770 ( .A(n525), .B(n[230]), .Z(n6417) );
  XOR U6771 ( .A(n6416), .B(n6417), .Z(n6419) );
  AND U6772 ( .A(n6407), .B(n[229]), .Z(n6408) );
  NANDN U6773 ( .A(n525), .B(n6408), .Z(n6412) );
  OR U6774 ( .A(n6410), .B(n6409), .Z(n6411) );
  AND U6775 ( .A(n6412), .B(n6411), .Z(n6418) );
  XNOR U6776 ( .A(n6419), .B(n6418), .Z(zout[230]) );
  NANDN U6777 ( .A(n6413), .B(n6814), .Z(n6414) );
  XNOR U6778 ( .A(n6415), .B(n6414), .Z(n6423) );
  NANDN U6779 ( .A(n6417), .B(n6416), .Z(n6421) );
  OR U6780 ( .A(n6419), .B(n6418), .Z(n6420) );
  AND U6781 ( .A(n6421), .B(n6420), .Z(n6424) );
  XOR U6782 ( .A(n6423), .B(n6424), .Z(zout[231]) );
  NANDN U6783 ( .A(n525), .B(n[232]), .Z(n6428) );
  XOR U6784 ( .A(n6427), .B(n6428), .Z(n6430) );
  NANDN U6785 ( .A(n525), .B(n6422), .Z(n6426) );
  NANDN U6786 ( .A(n6424), .B(n6423), .Z(n6425) );
  AND U6787 ( .A(n6426), .B(n6425), .Z(n6429) );
  XNOR U6788 ( .A(n6430), .B(n6429), .Z(zout[232]) );
  NANDN U6789 ( .A(n525), .B(n[233]), .Z(n6436) );
  NANDN U6790 ( .A(n6428), .B(n6427), .Z(n6432) );
  OR U6791 ( .A(n6430), .B(n6429), .Z(n6431) );
  AND U6792 ( .A(n6432), .B(n6431), .Z(n6435) );
  XOR U6793 ( .A(n6434), .B(n6435), .Z(n6433) );
  XNOR U6794 ( .A(n6436), .B(n6433), .Z(zout[233]) );
  NANDN U6795 ( .A(n525), .B(n[234]), .Z(n6440) );
  XNOR U6796 ( .A(n6439), .B(n6438), .Z(n6437) );
  XNOR U6797 ( .A(n6440), .B(n6437), .Z(zout[234]) );
  NANDN U6798 ( .A(n525), .B(n[235]), .Z(n6441) );
  XOR U6799 ( .A(n6443), .B(n6441), .Z(n6446) );
  XOR U6800 ( .A(n6445), .B(n6446), .Z(zout[235]) );
  NANDN U6801 ( .A(n6449), .B(n6814), .Z(n6442) );
  XNOR U6802 ( .A(n6450), .B(n6442), .Z(n6452) );
  AND U6803 ( .A(n6443), .B(n[235]), .Z(n6444) );
  NANDN U6804 ( .A(n525), .B(n6444), .Z(n6448) );
  NANDN U6805 ( .A(n6446), .B(n6445), .Z(n6447) );
  AND U6806 ( .A(n6448), .B(n6447), .Z(n6453) );
  XOR U6807 ( .A(n6452), .B(n6453), .Z(zout[236]) );
  ANDN U6808 ( .B(n6450), .A(n6449), .Z(n6451) );
  NANDN U6809 ( .A(n525), .B(n6451), .Z(n6455) );
  NANDN U6810 ( .A(n6453), .B(n6452), .Z(n6454) );
  NAND U6811 ( .A(n6455), .B(n6454), .Z(n6461) );
  NANDN U6812 ( .A(n6456), .B(n6814), .Z(n6458) );
  AND U6813 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U6814 ( .A(n6459), .B(n6814), .Z(n6463) );
  NANDN U6815 ( .A(n6462), .B(n6463), .Z(n6460) );
  XOR U6816 ( .A(n6461), .B(n6460), .Z(zout[237]) );
  NANDN U6817 ( .A(n6462), .B(n6461), .Z(n6464) );
  AND U6818 ( .A(n6464), .B(n6463), .Z(n6469) );
  NANDN U6819 ( .A(n525), .B(n[238]), .Z(n6465) );
  XOR U6820 ( .A(n6466), .B(n6465), .Z(n6468) );
  XNOR U6821 ( .A(n6469), .B(n6468), .Z(zout[238]) );
  AND U6822 ( .A(n6466), .B(n[238]), .Z(n6467) );
  NANDN U6823 ( .A(n525), .B(n6467), .Z(n6471) );
  OR U6824 ( .A(n6469), .B(n6468), .Z(n6470) );
  NAND U6825 ( .A(n6471), .B(n6470), .Z(n6475) );
  AND U6826 ( .A(n6814), .B(n[239]), .Z(n6476) );
  XOR U6827 ( .A(n6474), .B(n6476), .Z(n6472) );
  XNOR U6828 ( .A(n6475), .B(n6472), .Z(zout[239]) );
  AND U6829 ( .A(n6814), .B(n[23]), .Z(n6538) );
  XNOR U6830 ( .A(n6537), .B(n6538), .Z(n6535) );
  AND U6831 ( .A(n6814), .B(n6473), .Z(n6536) );
  XOR U6832 ( .A(n6535), .B(n6536), .Z(zout[23]) );
  NANDN U6833 ( .A(n525), .B(n[240]), .Z(n6478) );
  XOR U6834 ( .A(n6477), .B(n6478), .Z(n6480) );
  XNOR U6835 ( .A(n6480), .B(n6479), .Z(zout[240]) );
  NANDN U6836 ( .A(n525), .B(n[241]), .Z(n6484) );
  XOR U6837 ( .A(n6483), .B(n6484), .Z(n6486) );
  NANDN U6838 ( .A(n6478), .B(n6477), .Z(n6482) );
  OR U6839 ( .A(n6480), .B(n6479), .Z(n6481) );
  AND U6840 ( .A(n6482), .B(n6481), .Z(n6485) );
  XNOR U6841 ( .A(n6486), .B(n6485), .Z(zout[241]) );
  NANDN U6842 ( .A(n525), .B(n[242]), .Z(n6491) );
  XOR U6843 ( .A(n6490), .B(n6491), .Z(n6493) );
  NANDN U6844 ( .A(n6484), .B(n6483), .Z(n6488) );
  OR U6845 ( .A(n6486), .B(n6485), .Z(n6487) );
  AND U6846 ( .A(n6488), .B(n6487), .Z(n6492) );
  XNOR U6847 ( .A(n6493), .B(n6492), .Z(zout[242]) );
  NANDN U6848 ( .A(n525), .B(n[243]), .Z(n6489) );
  XOR U6849 ( .A(n6496), .B(n6489), .Z(n6499) );
  NANDN U6850 ( .A(n6491), .B(n6490), .Z(n6495) );
  OR U6851 ( .A(n6493), .B(n6492), .Z(n6494) );
  AND U6852 ( .A(n6495), .B(n6494), .Z(n6498) );
  XNOR U6853 ( .A(n6499), .B(n6498), .Z(zout[243]) );
  NANDN U6854 ( .A(n525), .B(n[244]), .Z(n6505) );
  AND U6855 ( .A(n6496), .B(n[243]), .Z(n6497) );
  NANDN U6856 ( .A(n525), .B(n6497), .Z(n6501) );
  OR U6857 ( .A(n6499), .B(n6498), .Z(n6500) );
  AND U6858 ( .A(n6501), .B(n6500), .Z(n6504) );
  XOR U6859 ( .A(n6503), .B(n6504), .Z(n6502) );
  XNOR U6860 ( .A(n6505), .B(n6502), .Z(zout[244]) );
  NANDN U6861 ( .A(n525), .B(n[245]), .Z(n6506) );
  XOR U6862 ( .A(n6508), .B(n6506), .Z(n6511) );
  XOR U6863 ( .A(n6510), .B(n6511), .Z(zout[245]) );
  NANDN U6864 ( .A(n6514), .B(n6814), .Z(n6507) );
  XOR U6865 ( .A(n6515), .B(n6507), .Z(n6518) );
  AND U6866 ( .A(n6508), .B(n[245]), .Z(n6509) );
  NANDN U6867 ( .A(n525), .B(n6509), .Z(n6513) );
  NANDN U6868 ( .A(n6511), .B(n6510), .Z(n6512) );
  AND U6869 ( .A(n6513), .B(n6512), .Z(n6517) );
  XNOR U6870 ( .A(n6518), .B(n6517), .Z(zout[246]) );
  NANDN U6871 ( .A(n525), .B(n[247]), .Z(n6523) );
  XOR U6872 ( .A(n6522), .B(n6523), .Z(n6525) );
  ANDN U6873 ( .B(n6515), .A(n6514), .Z(n6516) );
  NANDN U6874 ( .A(n525), .B(n6516), .Z(n6520) );
  OR U6875 ( .A(n6518), .B(n6517), .Z(n6519) );
  AND U6876 ( .A(n6520), .B(n6519), .Z(n6524) );
  XNOR U6877 ( .A(n6525), .B(n6524), .Z(zout[247]) );
  NANDN U6878 ( .A(n525), .B(n[248]), .Z(n6521) );
  XOR U6879 ( .A(n6528), .B(n6521), .Z(n6531) );
  NANDN U6880 ( .A(n6523), .B(n6522), .Z(n6527) );
  OR U6881 ( .A(n6525), .B(n6524), .Z(n6526) );
  AND U6882 ( .A(n6527), .B(n6526), .Z(n6530) );
  XNOR U6883 ( .A(n6531), .B(n6530), .Z(zout[248]) );
  AND U6884 ( .A(n6528), .B(n[248]), .Z(n6529) );
  NANDN U6885 ( .A(n525), .B(n6529), .Z(n6533) );
  OR U6886 ( .A(n6531), .B(n6530), .Z(n6532) );
  NAND U6887 ( .A(n6533), .B(n6532), .Z(n6547) );
  XOR U6888 ( .A(n6546), .B(n6547), .Z(n6548) );
  NANDN U6889 ( .A(n6534), .B(n6814), .Z(n6549) );
  XOR U6890 ( .A(n6548), .B(n6549), .Z(zout[249]) );
  OR U6891 ( .A(n6536), .B(n6535), .Z(n6540) );
  OR U6892 ( .A(n6538), .B(n6537), .Z(n6539) );
  AND U6893 ( .A(n6540), .B(n6539), .Z(n6542) );
  NANDN U6894 ( .A(n525), .B(n[24]), .Z(n6541) );
  XNOR U6895 ( .A(n6542), .B(n6541), .Z(n6543) );
  XNOR U6896 ( .A(n6544), .B(n6543), .Z(zout[24]) );
  NANDN U6897 ( .A(n525), .B(n[250]), .Z(n6545) );
  XOR U6898 ( .A(n6552), .B(n6545), .Z(n6555) );
  NAND U6899 ( .A(n6547), .B(n6546), .Z(n6551) );
  NANDN U6900 ( .A(n6549), .B(n6548), .Z(n6550) );
  AND U6901 ( .A(n6551), .B(n6550), .Z(n6554) );
  XNOR U6902 ( .A(n6555), .B(n6554), .Z(zout[250]) );
  NANDN U6903 ( .A(n525), .B(n[251]), .Z(n6559) );
  XOR U6904 ( .A(n6558), .B(n6559), .Z(n6561) );
  AND U6905 ( .A(n6552), .B(n[250]), .Z(n6553) );
  NANDN U6906 ( .A(n525), .B(n6553), .Z(n6557) );
  OR U6907 ( .A(n6555), .B(n6554), .Z(n6556) );
  AND U6908 ( .A(n6557), .B(n6556), .Z(n6560) );
  XNOR U6909 ( .A(n6561), .B(n6560), .Z(zout[251]) );
  NANDN U6910 ( .A(n525), .B(n[252]), .Z(n6565) );
  XOR U6911 ( .A(n6564), .B(n6565), .Z(n6567) );
  NANDN U6912 ( .A(n6559), .B(n6558), .Z(n6563) );
  OR U6913 ( .A(n6561), .B(n6560), .Z(n6562) );
  AND U6914 ( .A(n6563), .B(n6562), .Z(n6566) );
  XNOR U6915 ( .A(n6567), .B(n6566), .Z(zout[252]) );
  NANDN U6916 ( .A(n6565), .B(n6564), .Z(n6569) );
  OR U6917 ( .A(n6567), .B(n6566), .Z(n6568) );
  NAND U6918 ( .A(n6569), .B(n6568), .Z(n6572) );
  XOR U6919 ( .A(n6571), .B(n6572), .Z(n6573) );
  NANDN U6920 ( .A(n525), .B(n[253]), .Z(n6574) );
  XOR U6921 ( .A(n6573), .B(n6574), .Z(zout[253]) );
  NANDN U6922 ( .A(n6582), .B(n6814), .Z(n6570) );
  XOR U6923 ( .A(n6583), .B(n6570), .Z(n6586) );
  NAND U6924 ( .A(n6572), .B(n6571), .Z(n6576) );
  NANDN U6925 ( .A(n6574), .B(n6573), .Z(n6575) );
  AND U6926 ( .A(n6576), .B(n6575), .Z(n6585) );
  XNOR U6927 ( .A(n6586), .B(n6585), .Z(zout[254]) );
  AND U6928 ( .A(n6580), .B(n[255]), .Z(n6578) );
  NAND U6929 ( .A(n6578), .B(n6577), .Z(n6592) );
  NANDN U6930 ( .A(n525), .B(n[255]), .Z(n6579) );
  NANDN U6931 ( .A(n6580), .B(n6579), .Z(n6581) );
  NAND U6932 ( .A(n6592), .B(n6581), .Z(n6590) );
  ANDN U6933 ( .B(n6583), .A(n6582), .Z(n6584) );
  NANDN U6934 ( .A(n525), .B(n6584), .Z(n6588) );
  OR U6935 ( .A(n6586), .B(n6585), .Z(n6587) );
  AND U6936 ( .A(n6588), .B(n6587), .Z(n6589) );
  XNOR U6937 ( .A(n6590), .B(n6589), .Z(zout[255]) );
  NOR U6938 ( .A(n6590), .B(n6589), .Z(n6591) );
  ANDN U6939 ( .B(n6592), .A(n6591), .Z(n6593) );
  XOR U6940 ( .A(n6594), .B(n6593), .Z(zout[256]) );
  NOR U6941 ( .A(n525), .B(n6595), .Z(n6599) );
  XNOR U6942 ( .A(n6598), .B(n6599), .Z(n6596) );
  AND U6943 ( .A(n[25]), .B(n6814), .Z(n6597) );
  XOR U6944 ( .A(n6596), .B(n6597), .Z(zout[25]) );
  OR U6945 ( .A(n6597), .B(n6596), .Z(n6601) );
  OR U6946 ( .A(n6599), .B(n6598), .Z(n6600) );
  AND U6947 ( .A(n6601), .B(n6600), .Z(n6603) );
  NANDN U6948 ( .A(n525), .B(n[26]), .Z(n6602) );
  XNOR U6949 ( .A(n6603), .B(n6602), .Z(n6604) );
  XNOR U6950 ( .A(n6605), .B(n6604), .Z(zout[26]) );
  XOR U6951 ( .A(n[27]), .B(n6606), .Z(n6607) );
  NANDN U6952 ( .A(n525), .B(n6607), .Z(n6608) );
  XOR U6953 ( .A(n6609), .B(n6608), .Z(zout[27]) );
  XOR U6954 ( .A(n[28]), .B(n6610), .Z(n6611) );
  NANDN U6955 ( .A(n525), .B(n6611), .Z(n6612) );
  XOR U6956 ( .A(n6613), .B(n6612), .Z(zout[28]) );
  AND U6957 ( .A(n6814), .B(n[29]), .Z(n6623) );
  XNOR U6958 ( .A(n6622), .B(n6623), .Z(n6620) );
  NOR U6959 ( .A(n525), .B(n6614), .Z(n6621) );
  XOR U6960 ( .A(n6620), .B(n6621), .Z(zout[29]) );
  XNOR U6961 ( .A(n6616), .B(n6615), .Z(n6617) );
  NANDN U6962 ( .A(n525), .B(n6617), .Z(n6618) );
  XOR U6963 ( .A(n6619), .B(n6618), .Z(zout[2]) );
  OR U6964 ( .A(n6621), .B(n6620), .Z(n6625) );
  OR U6965 ( .A(n6623), .B(n6622), .Z(n6624) );
  AND U6966 ( .A(n6625), .B(n6624), .Z(n6627) );
  NANDN U6967 ( .A(n525), .B(n[30]), .Z(n6626) );
  XNOR U6968 ( .A(n6627), .B(n6626), .Z(n6628) );
  XNOR U6969 ( .A(n6629), .B(n6628), .Z(zout[30]) );
  AND U6970 ( .A(n6814), .B(n[31]), .Z(n6634) );
  XNOR U6971 ( .A(n6633), .B(n6634), .Z(n6631) );
  AND U6972 ( .A(n6814), .B(n6630), .Z(n6632) );
  XOR U6973 ( .A(n6631), .B(n6632), .Z(zout[31]) );
  OR U6974 ( .A(n6632), .B(n6631), .Z(n6636) );
  OR U6975 ( .A(n6634), .B(n6633), .Z(n6635) );
  AND U6976 ( .A(n6636), .B(n6635), .Z(n6638) );
  NANDN U6977 ( .A(n525), .B(n[32]), .Z(n6637) );
  XNOR U6978 ( .A(n6638), .B(n6637), .Z(n6639) );
  XNOR U6979 ( .A(n6640), .B(n6639), .Z(zout[32]) );
  XNOR U6980 ( .A(n[33]), .B(n6641), .Z(n6642) );
  ANDN U6981 ( .B(n6642), .A(n525), .Z(n6643) );
  XNOR U6982 ( .A(n6644), .B(n6643), .Z(zout[33]) );
  XNOR U6983 ( .A(n[34]), .B(n6645), .Z(n6646) );
  ANDN U6984 ( .B(n6646), .A(n525), .Z(n6647) );
  XNOR U6985 ( .A(n6648), .B(n6647), .Z(zout[34]) );
  ANDN U6986 ( .B(n6814), .A(n6649), .Z(n6651) );
  XOR U6987 ( .A(n6650), .B(n6651), .Z(n6652) );
  AND U6988 ( .A(n6814), .B(n[35]), .Z(n6653) );
  XNOR U6989 ( .A(n6652), .B(n6653), .Z(zout[35]) );
  OR U6990 ( .A(n6651), .B(n6650), .Z(n6655) );
  NANDN U6991 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U6992 ( .A(n6655), .B(n6654), .Z(n6660) );
  NANDN U6993 ( .A(n6656), .B(n6814), .Z(n6657) );
  XNOR U6994 ( .A(n6658), .B(n6657), .Z(n6659) );
  XNOR U6995 ( .A(n6660), .B(n6659), .Z(zout[36]) );
  NOR U6996 ( .A(n525), .B(n6661), .Z(n6665) );
  XNOR U6997 ( .A(n6664), .B(n6665), .Z(n6662) );
  AND U6998 ( .A(n6814), .B(n[37]), .Z(n6663) );
  XOR U6999 ( .A(n6662), .B(n6663), .Z(zout[37]) );
  OR U7000 ( .A(n6663), .B(n6662), .Z(n6667) );
  OR U7001 ( .A(n6665), .B(n6664), .Z(n6666) );
  AND U7002 ( .A(n6667), .B(n6666), .Z(n6669) );
  NANDN U7003 ( .A(n525), .B(n[38]), .Z(n6668) );
  XNOR U7004 ( .A(n6669), .B(n6668), .Z(n6670) );
  XNOR U7005 ( .A(n6671), .B(n6670), .Z(zout[38]) );
  AND U7006 ( .A(n6814), .B(n[39]), .Z(n6680) );
  XNOR U7007 ( .A(n6679), .B(n6680), .Z(n6677) );
  NOR U7008 ( .A(n525), .B(n6672), .Z(n6678) );
  XOR U7009 ( .A(n6677), .B(n6678), .Z(zout[39]) );
  XOR U7010 ( .A(n[3]), .B(n6673), .Z(n6674) );
  NANDN U7011 ( .A(n525), .B(n6674), .Z(n6675) );
  XOR U7012 ( .A(n6676), .B(n6675), .Z(zout[3]) );
  OR U7013 ( .A(n6678), .B(n6677), .Z(n6682) );
  OR U7014 ( .A(n6680), .B(n6679), .Z(n6681) );
  AND U7015 ( .A(n6682), .B(n6681), .Z(n6684) );
  NANDN U7016 ( .A(n525), .B(n[40]), .Z(n6683) );
  XNOR U7017 ( .A(n6684), .B(n6683), .Z(n6685) );
  XNOR U7018 ( .A(n6686), .B(n6685), .Z(zout[40]) );
  AND U7019 ( .A(n6814), .B(n[41]), .Z(n6691) );
  XNOR U7020 ( .A(n6690), .B(n6691), .Z(n6688) );
  NOR U7021 ( .A(n525), .B(n6687), .Z(n6689) );
  XOR U7022 ( .A(n6688), .B(n6689), .Z(zout[41]) );
  OR U7023 ( .A(n6689), .B(n6688), .Z(n6693) );
  OR U7024 ( .A(n6691), .B(n6690), .Z(n6692) );
  AND U7025 ( .A(n6693), .B(n6692), .Z(n6695) );
  NANDN U7026 ( .A(n525), .B(n[42]), .Z(n6694) );
  XNOR U7027 ( .A(n6695), .B(n6694), .Z(n6696) );
  XNOR U7028 ( .A(n6697), .B(n6696), .Z(zout[42]) );
  XOR U7029 ( .A(n[43]), .B(n6698), .Z(n6699) );
  NANDN U7030 ( .A(n525), .B(n6699), .Z(n6700) );
  XOR U7031 ( .A(n6701), .B(n6700), .Z(zout[43]) );
  XOR U7032 ( .A(n[44]), .B(n6702), .Z(n6703) );
  NANDN U7033 ( .A(n525), .B(n6703), .Z(n6704) );
  XOR U7034 ( .A(n6705), .B(n6704), .Z(zout[44]) );
  XNOR U7035 ( .A(n[45]), .B(n6706), .Z(n6707) );
  NANDN U7036 ( .A(n525), .B(n6707), .Z(n6708) );
  XOR U7037 ( .A(n6709), .B(n6708), .Z(zout[45]) );
  XNOR U7038 ( .A(n6711), .B(n6710), .Z(n6712) );
  NANDN U7039 ( .A(n525), .B(n6712), .Z(n6713) );
  XOR U7040 ( .A(n6714), .B(n6713), .Z(zout[46]) );
  XNOR U7041 ( .A(n6716), .B(n6715), .Z(n6717) );
  NANDN U7042 ( .A(n525), .B(n6717), .Z(n6718) );
  XOR U7043 ( .A(n6719), .B(n6718), .Z(zout[47]) );
  XNOR U7044 ( .A(n6721), .B(n6720), .Z(zout[48]) );
  XOR U7045 ( .A(n6723), .B(n6722), .Z(n6724) );
  XNOR U7046 ( .A(n6725), .B(n6724), .Z(zout[49]) );
  XNOR U7047 ( .A(n[4]), .B(n6726), .Z(n6727) );
  NANDN U7048 ( .A(n525), .B(n6727), .Z(n6728) );
  XOR U7049 ( .A(n6729), .B(n6728), .Z(zout[4]) );
  XOR U7050 ( .A(n6731), .B(n6730), .Z(n6732) );
  XNOR U7051 ( .A(n6733), .B(n6732), .Z(zout[50]) );
  XNOR U7052 ( .A(n6735), .B(n6734), .Z(zout[51]) );
  XNOR U7053 ( .A(n6737), .B(n6736), .Z(zout[52]) );
  XOR U7054 ( .A(n6739), .B(n6738), .Z(n6740) );
  XNOR U7055 ( .A(n6741), .B(n6740), .Z(zout[53]) );
  XOR U7056 ( .A(n6743), .B(n6742), .Z(zout[54]) );
  XNOR U7057 ( .A(n6745), .B(n6744), .Z(zout[55]) );
  XNOR U7058 ( .A(n6747), .B(n6746), .Z(zout[56]) );
  XNOR U7059 ( .A(n6749), .B(n6748), .Z(zout[57]) );
  XNOR U7060 ( .A(n6751), .B(n6750), .Z(zout[58]) );
  XNOR U7061 ( .A(n6753), .B(n6752), .Z(zout[59]) );
  AND U7062 ( .A(n[5]), .B(n6814), .Z(n6782) );
  XNOR U7063 ( .A(n6781), .B(n6782), .Z(n6779) );
  NOR U7064 ( .A(n525), .B(n6754), .Z(n6780) );
  XOR U7065 ( .A(n6779), .B(n6780), .Z(zout[5]) );
  XNOR U7066 ( .A(n6756), .B(n6755), .Z(zout[60]) );
  XNOR U7067 ( .A(n6758), .B(n6757), .Z(zout[61]) );
  XNOR U7068 ( .A(n6760), .B(n6759), .Z(zout[62]) );
  XOR U7069 ( .A(n6762), .B(n6761), .Z(zout[63]) );
  XNOR U7070 ( .A(n6764), .B(n6763), .Z(zout[64]) );
  XNOR U7071 ( .A(n6766), .B(n6765), .Z(zout[65]) );
  XOR U7072 ( .A(n6768), .B(n6767), .Z(n6769) );
  XNOR U7073 ( .A(n6770), .B(n6769), .Z(zout[66]) );
  XOR U7074 ( .A(n6772), .B(n6771), .Z(zout[67]) );
  XOR U7075 ( .A(n6774), .B(n6773), .Z(n6775) );
  XNOR U7076 ( .A(n6776), .B(n6775), .Z(zout[68]) );
  XOR U7077 ( .A(n6778), .B(n6777), .Z(zout[69]) );
  OR U7078 ( .A(n6780), .B(n6779), .Z(n6784) );
  OR U7079 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U7080 ( .A(n6784), .B(n6783), .Z(n6786) );
  NANDN U7081 ( .A(n525), .B(n[6]), .Z(n6785) );
  XNOR U7082 ( .A(n6786), .B(n6785), .Z(n6787) );
  XNOR U7083 ( .A(n6788), .B(n6787), .Z(zout[6]) );
  XOR U7084 ( .A(n6790), .B(n6789), .Z(zout[70]) );
  XNOR U7085 ( .A(n6792), .B(n6791), .Z(zout[71]) );
  XNOR U7086 ( .A(n6794), .B(n6793), .Z(zout[72]) );
  XNOR U7087 ( .A(n6796), .B(n6795), .Z(zout[73]) );
  XNOR U7088 ( .A(n6798), .B(n6797), .Z(zout[74]) );
  XOR U7089 ( .A(n6800), .B(n6799), .Z(zout[75]) );
  XNOR U7090 ( .A(n6802), .B(n6801), .Z(zout[76]) );
  XOR U7091 ( .A(n6804), .B(n6803), .Z(n6805) );
  XNOR U7092 ( .A(n6806), .B(n6805), .Z(zout[77]) );
  XNOR U7093 ( .A(n6808), .B(n6807), .Z(zout[78]) );
  XOR U7094 ( .A(n6810), .B(n6809), .Z(n6811) );
  XNOR U7095 ( .A(n6812), .B(n6811), .Z(zout[79]) );
  NOR U7096 ( .A(n525), .B(n6813), .Z(n6838) );
  XNOR U7097 ( .A(n6837), .B(n6838), .Z(n6835) );
  AND U7098 ( .A(n6814), .B(n[7]), .Z(n6836) );
  XOR U7099 ( .A(n6835), .B(n6836), .Z(zout[7]) );
  XNOR U7100 ( .A(n6816), .B(n6815), .Z(zout[80]) );
  XNOR U7101 ( .A(n6818), .B(n6817), .Z(zout[81]) );
  XNOR U7102 ( .A(n6820), .B(n6819), .Z(zout[82]) );
  XNOR U7103 ( .A(n6822), .B(n6821), .Z(zout[83]) );
  XNOR U7104 ( .A(n6824), .B(n6823), .Z(zout[84]) );
  XOR U7105 ( .A(n6826), .B(n6825), .Z(zout[85]) );
  XNOR U7106 ( .A(n6828), .B(n6827), .Z(zout[86]) );
  XNOR U7107 ( .A(n6830), .B(n6829), .Z(zout[87]) );
  XOR U7108 ( .A(n6832), .B(n6831), .Z(zout[88]) );
  XNOR U7109 ( .A(n6834), .B(n6833), .Z(zout[89]) );
  OR U7110 ( .A(n6836), .B(n6835), .Z(n6840) );
  OR U7111 ( .A(n6838), .B(n6837), .Z(n6839) );
  AND U7112 ( .A(n6840), .B(n6839), .Z(n6842) );
  NANDN U7113 ( .A(n525), .B(n[8]), .Z(n6841) );
  XNOR U7114 ( .A(n6842), .B(n6841), .Z(n6843) );
  XNOR U7115 ( .A(n6844), .B(n6843), .Z(zout[8]) );
  XNOR U7116 ( .A(n6846), .B(n6845), .Z(zout[90]) );
  XNOR U7117 ( .A(n6848), .B(n6847), .Z(zout[91]) );
  XNOR U7118 ( .A(n6850), .B(n6849), .Z(zout[92]) );
  XNOR U7119 ( .A(n6852), .B(n6851), .Z(zout[93]) );
  XNOR U7120 ( .A(n6854), .B(n6853), .Z(zout[94]) );
  XOR U7121 ( .A(n6856), .B(n6855), .Z(zout[95]) );
  XNOR U7122 ( .A(n6858), .B(n6857), .Z(zout[96]) );
  XOR U7123 ( .A(n6860), .B(n6859), .Z(n6861) );
  XNOR U7124 ( .A(n6862), .B(n6861), .Z(zout[97]) );
  XOR U7125 ( .A(n6864), .B(n6863), .Z(zout[98]) );
  XOR U7126 ( .A(n6866), .B(n6865), .Z(zout[99]) );
  XNOR U7127 ( .A(n6868), .B(n6867), .Z(n6869) );
  NANDN U7128 ( .A(n525), .B(n6869), .Z(n6870) );
  XOR U7129 ( .A(n6871), .B(n6870), .Z(zout[9]) );
endmodule


module modexp_2N_NN_N256_CC65536 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, \modmult_1/xreg[255] ,
         \modmult_1/xreg[254] , \modmult_1/xreg[253] , \modmult_1/xreg[252] ,
         \modmult_1/xreg[251] , \modmult_1/xreg[250] , \modmult_1/xreg[249] ,
         \modmult_1/xreg[248] , \modmult_1/xreg[247] , \modmult_1/xreg[246] ,
         \modmult_1/xreg[245] , \modmult_1/xreg[244] , \modmult_1/xreg[243] ,
         \modmult_1/xreg[242] , \modmult_1/xreg[241] , \modmult_1/xreg[240] ,
         \modmult_1/xreg[239] , \modmult_1/xreg[238] , \modmult_1/xreg[237] ,
         \modmult_1/xreg[236] , \modmult_1/xreg[235] , \modmult_1/xreg[234] ,
         \modmult_1/xreg[233] , \modmult_1/xreg[232] , \modmult_1/xreg[231] ,
         \modmult_1/xreg[230] , \modmult_1/xreg[229] , \modmult_1/xreg[228] ,
         \modmult_1/xreg[227] , \modmult_1/xreg[226] , \modmult_1/xreg[225] ,
         \modmult_1/xreg[224] , \modmult_1/xreg[223] , \modmult_1/xreg[222] ,
         \modmult_1/xreg[221] , \modmult_1/xreg[220] , \modmult_1/xreg[219] ,
         \modmult_1/xreg[218] , \modmult_1/xreg[217] , \modmult_1/xreg[216] ,
         \modmult_1/xreg[215] , \modmult_1/xreg[214] , \modmult_1/xreg[213] ,
         \modmult_1/xreg[212] , \modmult_1/xreg[211] , \modmult_1/xreg[210] ,
         \modmult_1/xreg[209] , \modmult_1/xreg[208] , \modmult_1/xreg[207] ,
         \modmult_1/xreg[206] , \modmult_1/xreg[205] , \modmult_1/xreg[204] ,
         \modmult_1/xreg[203] , \modmult_1/xreg[202] , \modmult_1/xreg[201] ,
         \modmult_1/xreg[200] , \modmult_1/xreg[199] , \modmult_1/xreg[198] ,
         \modmult_1/xreg[197] , \modmult_1/xreg[196] , \modmult_1/xreg[195] ,
         \modmult_1/xreg[194] , \modmult_1/xreg[193] , \modmult_1/xreg[192] ,
         \modmult_1/xreg[191] , \modmult_1/xreg[190] , \modmult_1/xreg[189] ,
         \modmult_1/xreg[188] , \modmult_1/xreg[187] , \modmult_1/xreg[186] ,
         \modmult_1/xreg[185] , \modmult_1/xreg[184] , \modmult_1/xreg[183] ,
         \modmult_1/xreg[182] , \modmult_1/xreg[181] , \modmult_1/xreg[180] ,
         \modmult_1/xreg[179] , \modmult_1/xreg[178] , \modmult_1/xreg[177] ,
         \modmult_1/xreg[176] , \modmult_1/xreg[175] , \modmult_1/xreg[174] ,
         \modmult_1/xreg[173] , \modmult_1/xreg[172] , \modmult_1/xreg[171] ,
         \modmult_1/xreg[170] , \modmult_1/xreg[169] , \modmult_1/xreg[168] ,
         \modmult_1/xreg[167] , \modmult_1/xreg[166] , \modmult_1/xreg[165] ,
         \modmult_1/xreg[164] , \modmult_1/xreg[163] , \modmult_1/xreg[162] ,
         \modmult_1/xreg[161] , \modmult_1/xreg[160] , \modmult_1/xreg[159] ,
         \modmult_1/xreg[158] , \modmult_1/xreg[157] , \modmult_1/xreg[156] ,
         \modmult_1/xreg[155] , \modmult_1/xreg[154] , \modmult_1/xreg[153] ,
         \modmult_1/xreg[152] , \modmult_1/xreg[151] , \modmult_1/xreg[150] ,
         \modmult_1/xreg[149] , \modmult_1/xreg[148] , \modmult_1/xreg[147] ,
         \modmult_1/xreg[146] , \modmult_1/xreg[145] , \modmult_1/xreg[144] ,
         \modmult_1/xreg[143] , \modmult_1/xreg[142] , \modmult_1/xreg[141] ,
         \modmult_1/xreg[140] , \modmult_1/xreg[139] , \modmult_1/xreg[138] ,
         \modmult_1/xreg[137] , \modmult_1/xreg[136] , \modmult_1/xreg[135] ,
         \modmult_1/xreg[134] , \modmult_1/xreg[133] , \modmult_1/xreg[132] ,
         \modmult_1/xreg[131] , \modmult_1/xreg[130] , \modmult_1/xreg[129] ,
         \modmult_1/xreg[128] , \modmult_1/xreg[127] , \modmult_1/xreg[126] ,
         \modmult_1/xreg[125] , \modmult_1/xreg[124] , \modmult_1/xreg[123] ,
         \modmult_1/xreg[122] , \modmult_1/xreg[121] , \modmult_1/xreg[120] ,
         \modmult_1/xreg[119] , \modmult_1/xreg[118] , \modmult_1/xreg[117] ,
         \modmult_1/xreg[116] , \modmult_1/xreg[115] , \modmult_1/xreg[114] ,
         \modmult_1/xreg[113] , \modmult_1/xreg[112] , \modmult_1/xreg[111] ,
         \modmult_1/xreg[110] , \modmult_1/xreg[109] , \modmult_1/xreg[108] ,
         \modmult_1/xreg[107] , \modmult_1/xreg[106] , \modmult_1/xreg[105] ,
         \modmult_1/xreg[104] , \modmult_1/xreg[103] , \modmult_1/xreg[102] ,
         \modmult_1/xreg[101] , \modmult_1/xreg[100] , \modmult_1/xreg[99] ,
         \modmult_1/xreg[98] , \modmult_1/xreg[97] , \modmult_1/xreg[96] ,
         \modmult_1/xreg[95] , \modmult_1/xreg[94] , \modmult_1/xreg[93] ,
         \modmult_1/xreg[92] , \modmult_1/xreg[91] , \modmult_1/xreg[90] ,
         \modmult_1/xreg[89] , \modmult_1/xreg[88] , \modmult_1/xreg[87] ,
         \modmult_1/xreg[86] , \modmult_1/xreg[85] , \modmult_1/xreg[84] ,
         \modmult_1/xreg[83] , \modmult_1/xreg[82] , \modmult_1/xreg[81] ,
         \modmult_1/xreg[80] , \modmult_1/xreg[79] , \modmult_1/xreg[78] ,
         \modmult_1/xreg[77] , \modmult_1/xreg[76] , \modmult_1/xreg[75] ,
         \modmult_1/xreg[74] , \modmult_1/xreg[73] , \modmult_1/xreg[72] ,
         \modmult_1/xreg[71] , \modmult_1/xreg[70] , \modmult_1/xreg[69] ,
         \modmult_1/xreg[68] , \modmult_1/xreg[67] , \modmult_1/xreg[66] ,
         \modmult_1/xreg[65] , \modmult_1/xreg[64] , \modmult_1/xreg[63] ,
         \modmult_1/xreg[62] , \modmult_1/xreg[61] , \modmult_1/xreg[60] ,
         \modmult_1/xreg[59] , \modmult_1/xreg[58] , \modmult_1/xreg[57] ,
         \modmult_1/xreg[56] , \modmult_1/xreg[55] , \modmult_1/xreg[54] ,
         \modmult_1/xreg[53] , \modmult_1/xreg[52] , \modmult_1/xreg[51] ,
         \modmult_1/xreg[50] , \modmult_1/xreg[49] , \modmult_1/xreg[48] ,
         \modmult_1/xreg[47] , \modmult_1/xreg[46] , \modmult_1/xreg[45] ,
         \modmult_1/xreg[44] , \modmult_1/xreg[43] , \modmult_1/xreg[42] ,
         \modmult_1/xreg[41] , \modmult_1/xreg[40] , \modmult_1/xreg[39] ,
         \modmult_1/xreg[38] , \modmult_1/xreg[37] , \modmult_1/xreg[36] ,
         \modmult_1/xreg[35] , \modmult_1/xreg[34] , \modmult_1/xreg[33] ,
         \modmult_1/xreg[32] , \modmult_1/xreg[31] , \modmult_1/xreg[30] ,
         \modmult_1/xreg[29] , \modmult_1/xreg[28] , \modmult_1/xreg[27] ,
         \modmult_1/xreg[26] , \modmult_1/xreg[25] , \modmult_1/xreg[24] ,
         \modmult_1/xreg[23] , \modmult_1/xreg[22] , \modmult_1/xreg[21] ,
         \modmult_1/xreg[20] , \modmult_1/xreg[19] , \modmult_1/xreg[18] ,
         \modmult_1/xreg[17] , \modmult_1/xreg[16] , \modmult_1/xreg[15] ,
         \modmult_1/xreg[14] , \modmult_1/xreg[13] , \modmult_1/xreg[12] ,
         \modmult_1/xreg[11] , \modmult_1/xreg[10] , \modmult_1/xreg[9] ,
         \modmult_1/xreg[8] , \modmult_1/xreg[7] , \modmult_1/xreg[6] ,
         \modmult_1/xreg[5] , \modmult_1/xreg[4] , \modmult_1/xreg[3] ,
         \modmult_1/xreg[2] , \modmult_1/xin[255] , \modmult_1/xin[254] ,
         \modmult_1/xin[253] , \modmult_1/xin[252] , \modmult_1/xin[251] ,
         \modmult_1/xin[250] , \modmult_1/xin[249] , \modmult_1/xin[248] ,
         \modmult_1/xin[247] , \modmult_1/xin[246] , \modmult_1/xin[245] ,
         \modmult_1/xin[244] , \modmult_1/xin[243] , \modmult_1/xin[242] ,
         \modmult_1/xin[241] , \modmult_1/xin[240] , \modmult_1/xin[239] ,
         \modmult_1/xin[238] , \modmult_1/xin[237] , \modmult_1/xin[236] ,
         \modmult_1/xin[235] , \modmult_1/xin[234] , \modmult_1/xin[233] ,
         \modmult_1/xin[232] , \modmult_1/xin[231] , \modmult_1/xin[230] ,
         \modmult_1/xin[229] , \modmult_1/xin[228] , \modmult_1/xin[227] ,
         \modmult_1/xin[226] , \modmult_1/xin[225] , \modmult_1/xin[224] ,
         \modmult_1/xin[223] , \modmult_1/xin[222] , \modmult_1/xin[221] ,
         \modmult_1/xin[220] , \modmult_1/xin[219] , \modmult_1/xin[218] ,
         \modmult_1/xin[217] , \modmult_1/xin[216] , \modmult_1/xin[215] ,
         \modmult_1/xin[214] , \modmult_1/xin[213] , \modmult_1/xin[212] ,
         \modmult_1/xin[211] , \modmult_1/xin[210] , \modmult_1/xin[209] ,
         \modmult_1/xin[208] , \modmult_1/xin[207] , \modmult_1/xin[206] ,
         \modmult_1/xin[205] , \modmult_1/xin[204] , \modmult_1/xin[203] ,
         \modmult_1/xin[202] , \modmult_1/xin[201] , \modmult_1/xin[200] ,
         \modmult_1/xin[199] , \modmult_1/xin[198] , \modmult_1/xin[197] ,
         \modmult_1/xin[196] , \modmult_1/xin[195] , \modmult_1/xin[194] ,
         \modmult_1/xin[193] , \modmult_1/xin[192] , \modmult_1/xin[191] ,
         \modmult_1/xin[190] , \modmult_1/xin[189] , \modmult_1/xin[188] ,
         \modmult_1/xin[187] , \modmult_1/xin[186] , \modmult_1/xin[185] ,
         \modmult_1/xin[184] , \modmult_1/xin[183] , \modmult_1/xin[182] ,
         \modmult_1/xin[181] , \modmult_1/xin[180] , \modmult_1/xin[179] ,
         \modmult_1/xin[178] , \modmult_1/xin[177] , \modmult_1/xin[176] ,
         \modmult_1/xin[175] , \modmult_1/xin[174] , \modmult_1/xin[173] ,
         \modmult_1/xin[172] , \modmult_1/xin[171] , \modmult_1/xin[170] ,
         \modmult_1/xin[169] , \modmult_1/xin[168] , \modmult_1/xin[167] ,
         \modmult_1/xin[166] , \modmult_1/xin[165] , \modmult_1/xin[164] ,
         \modmult_1/xin[163] , \modmult_1/xin[162] , \modmult_1/xin[161] ,
         \modmult_1/xin[160] , \modmult_1/xin[159] , \modmult_1/xin[158] ,
         \modmult_1/xin[157] , \modmult_1/xin[156] , \modmult_1/xin[155] ,
         \modmult_1/xin[154] , \modmult_1/xin[153] , \modmult_1/xin[152] ,
         \modmult_1/xin[151] , \modmult_1/xin[150] , \modmult_1/xin[149] ,
         \modmult_1/xin[148] , \modmult_1/xin[147] , \modmult_1/xin[146] ,
         \modmult_1/xin[145] , \modmult_1/xin[144] , \modmult_1/xin[143] ,
         \modmult_1/xin[142] , \modmult_1/xin[141] , \modmult_1/xin[140] ,
         \modmult_1/xin[139] , \modmult_1/xin[138] , \modmult_1/xin[137] ,
         \modmult_1/xin[136] , \modmult_1/xin[135] , \modmult_1/xin[134] ,
         \modmult_1/xin[133] , \modmult_1/xin[132] , \modmult_1/xin[131] ,
         \modmult_1/xin[130] , \modmult_1/xin[129] , \modmult_1/xin[128] ,
         \modmult_1/xin[127] , \modmult_1/xin[126] , \modmult_1/xin[125] ,
         \modmult_1/xin[124] , \modmult_1/xin[123] , \modmult_1/xin[122] ,
         \modmult_1/xin[121] , \modmult_1/xin[120] , \modmult_1/xin[119] ,
         \modmult_1/xin[118] , \modmult_1/xin[117] , \modmult_1/xin[116] ,
         \modmult_1/xin[115] , \modmult_1/xin[114] , \modmult_1/xin[113] ,
         \modmult_1/xin[112] , \modmult_1/xin[111] , \modmult_1/xin[110] ,
         \modmult_1/xin[109] , \modmult_1/xin[108] , \modmult_1/xin[107] ,
         \modmult_1/xin[106] , \modmult_1/xin[105] , \modmult_1/xin[104] ,
         \modmult_1/xin[103] , \modmult_1/xin[102] , \modmult_1/xin[101] ,
         \modmult_1/xin[100] , \modmult_1/xin[99] , \modmult_1/xin[98] ,
         \modmult_1/xin[97] , \modmult_1/xin[96] , \modmult_1/xin[95] ,
         \modmult_1/xin[94] , \modmult_1/xin[93] , \modmult_1/xin[92] ,
         \modmult_1/xin[91] , \modmult_1/xin[90] , \modmult_1/xin[89] ,
         \modmult_1/xin[88] , \modmult_1/xin[87] , \modmult_1/xin[86] ,
         \modmult_1/xin[85] , \modmult_1/xin[84] , \modmult_1/xin[83] ,
         \modmult_1/xin[82] , \modmult_1/xin[81] , \modmult_1/xin[80] ,
         \modmult_1/xin[79] , \modmult_1/xin[78] , \modmult_1/xin[77] ,
         \modmult_1/xin[76] , \modmult_1/xin[75] , \modmult_1/xin[74] ,
         \modmult_1/xin[73] , \modmult_1/xin[72] , \modmult_1/xin[71] ,
         \modmult_1/xin[70] , \modmult_1/xin[69] , \modmult_1/xin[68] ,
         \modmult_1/xin[67] , \modmult_1/xin[66] , \modmult_1/xin[65] ,
         \modmult_1/xin[64] , \modmult_1/xin[63] , \modmult_1/xin[62] ,
         \modmult_1/xin[61] , \modmult_1/xin[60] , \modmult_1/xin[59] ,
         \modmult_1/xin[58] , \modmult_1/xin[57] , \modmult_1/xin[56] ,
         \modmult_1/xin[55] , \modmult_1/xin[54] , \modmult_1/xin[53] ,
         \modmult_1/xin[52] , \modmult_1/xin[51] , \modmult_1/xin[50] ,
         \modmult_1/xin[49] , \modmult_1/xin[48] , \modmult_1/xin[47] ,
         \modmult_1/xin[46] , \modmult_1/xin[45] , \modmult_1/xin[44] ,
         \modmult_1/xin[43] , \modmult_1/xin[42] , \modmult_1/xin[41] ,
         \modmult_1/xin[40] , \modmult_1/xin[39] , \modmult_1/xin[38] ,
         \modmult_1/xin[37] , \modmult_1/xin[36] , \modmult_1/xin[35] ,
         \modmult_1/xin[34] , \modmult_1/xin[33] , \modmult_1/xin[32] ,
         \modmult_1/xin[31] , \modmult_1/xin[30] , \modmult_1/xin[29] ,
         \modmult_1/xin[28] , \modmult_1/xin[27] , \modmult_1/xin[26] ,
         \modmult_1/xin[25] , \modmult_1/xin[24] , \modmult_1/xin[23] ,
         \modmult_1/xin[22] , \modmult_1/xin[21] , \modmult_1/xin[20] ,
         \modmult_1/xin[19] , \modmult_1/xin[18] , \modmult_1/xin[17] ,
         \modmult_1/xin[16] , \modmult_1/xin[15] , \modmult_1/xin[14] ,
         \modmult_1/xin[13] , \modmult_1/xin[12] , \modmult_1/xin[11] ,
         \modmult_1/xin[10] , \modmult_1/xin[9] , \modmult_1/xin[8] ,
         \modmult_1/xin[7] , \modmult_1/xin[6] , \modmult_1/xin[5] ,
         \modmult_1/xin[4] , \modmult_1/xin[3] , \modmult_1/xin[2] ,
         \modmult_1/xin[1] , \modmult_1/xin[0] , \modmult_1/zin[1][256] ,
         \modmult_1/zin[1][255] , \modmult_1/zin[1][254] ,
         \modmult_1/zin[1][253] , \modmult_1/zin[1][252] ,
         \modmult_1/zin[1][251] , \modmult_1/zin[1][250] ,
         \modmult_1/zin[1][249] , \modmult_1/zin[1][248] ,
         \modmult_1/zin[1][247] , \modmult_1/zin[1][246] ,
         \modmult_1/zin[1][245] , \modmult_1/zin[1][244] ,
         \modmult_1/zin[1][243] , \modmult_1/zin[1][242] ,
         \modmult_1/zin[1][241] , \modmult_1/zin[1][240] ,
         \modmult_1/zin[1][239] , \modmult_1/zin[1][238] ,
         \modmult_1/zin[1][237] , \modmult_1/zin[1][236] ,
         \modmult_1/zin[1][235] , \modmult_1/zin[1][234] ,
         \modmult_1/zin[1][233] , \modmult_1/zin[1][232] ,
         \modmult_1/zin[1][231] , \modmult_1/zin[1][230] ,
         \modmult_1/zin[1][229] , \modmult_1/zin[1][228] ,
         \modmult_1/zin[1][227] , \modmult_1/zin[1][226] ,
         \modmult_1/zin[1][225] , \modmult_1/zin[1][224] ,
         \modmult_1/zin[1][223] , \modmult_1/zin[1][222] ,
         \modmult_1/zin[1][221] , \modmult_1/zin[1][220] ,
         \modmult_1/zin[1][219] , \modmult_1/zin[1][218] ,
         \modmult_1/zin[1][217] , \modmult_1/zin[1][216] ,
         \modmult_1/zin[1][215] , \modmult_1/zin[1][214] ,
         \modmult_1/zin[1][213] , \modmult_1/zin[1][212] ,
         \modmult_1/zin[1][211] , \modmult_1/zin[1][210] ,
         \modmult_1/zin[1][209] , \modmult_1/zin[1][208] ,
         \modmult_1/zin[1][207] , \modmult_1/zin[1][206] ,
         \modmult_1/zin[1][205] , \modmult_1/zin[1][204] ,
         \modmult_1/zin[1][203] , \modmult_1/zin[1][202] ,
         \modmult_1/zin[1][201] , \modmult_1/zin[1][200] ,
         \modmult_1/zin[1][199] , \modmult_1/zin[1][198] ,
         \modmult_1/zin[1][197] , \modmult_1/zin[1][196] ,
         \modmult_1/zin[1][195] , \modmult_1/zin[1][194] ,
         \modmult_1/zin[1][193] , \modmult_1/zin[1][192] ,
         \modmult_1/zin[1][191] , \modmult_1/zin[1][190] ,
         \modmult_1/zin[1][189] , \modmult_1/zin[1][188] ,
         \modmult_1/zin[1][187] , \modmult_1/zin[1][186] ,
         \modmult_1/zin[1][185] , \modmult_1/zin[1][184] ,
         \modmult_1/zin[1][183] , \modmult_1/zin[1][182] ,
         \modmult_1/zin[1][181] , \modmult_1/zin[1][180] ,
         \modmult_1/zin[1][179] , \modmult_1/zin[1][178] ,
         \modmult_1/zin[1][177] , \modmult_1/zin[1][176] ,
         \modmult_1/zin[1][175] , \modmult_1/zin[1][174] ,
         \modmult_1/zin[1][173] , \modmult_1/zin[1][172] ,
         \modmult_1/zin[1][171] , \modmult_1/zin[1][170] ,
         \modmult_1/zin[1][169] , \modmult_1/zin[1][168] ,
         \modmult_1/zin[1][167] , \modmult_1/zin[1][166] ,
         \modmult_1/zin[1][165] , \modmult_1/zin[1][164] ,
         \modmult_1/zin[1][163] , \modmult_1/zin[1][162] ,
         \modmult_1/zin[1][161] , \modmult_1/zin[1][160] ,
         \modmult_1/zin[1][159] , \modmult_1/zin[1][158] ,
         \modmult_1/zin[1][157] , \modmult_1/zin[1][156] ,
         \modmult_1/zin[1][155] , \modmult_1/zin[1][154] ,
         \modmult_1/zin[1][153] , \modmult_1/zin[1][152] ,
         \modmult_1/zin[1][151] , \modmult_1/zin[1][150] ,
         \modmult_1/zin[1][149] , \modmult_1/zin[1][148] ,
         \modmult_1/zin[1][147] , \modmult_1/zin[1][146] ,
         \modmult_1/zin[1][145] , \modmult_1/zin[1][144] ,
         \modmult_1/zin[1][143] , \modmult_1/zin[1][142] ,
         \modmult_1/zin[1][141] , \modmult_1/zin[1][140] ,
         \modmult_1/zin[1][139] , \modmult_1/zin[1][138] ,
         \modmult_1/zin[1][137] , \modmult_1/zin[1][136] ,
         \modmult_1/zin[1][135] , \modmult_1/zin[1][134] ,
         \modmult_1/zin[1][133] , \modmult_1/zin[1][132] ,
         \modmult_1/zin[1][131] , \modmult_1/zin[1][130] ,
         \modmult_1/zin[1][129] , \modmult_1/zin[1][128] ,
         \modmult_1/zin[1][127] , \modmult_1/zin[1][126] ,
         \modmult_1/zin[1][125] , \modmult_1/zin[1][124] ,
         \modmult_1/zin[1][123] , \modmult_1/zin[1][122] ,
         \modmult_1/zin[1][121] , \modmult_1/zin[1][120] ,
         \modmult_1/zin[1][119] , \modmult_1/zin[1][118] ,
         \modmult_1/zin[1][117] , \modmult_1/zin[1][116] ,
         \modmult_1/zin[1][115] , \modmult_1/zin[1][114] ,
         \modmult_1/zin[1][113] , \modmult_1/zin[1][112] ,
         \modmult_1/zin[1][111] , \modmult_1/zin[1][110] ,
         \modmult_1/zin[1][109] , \modmult_1/zin[1][108] ,
         \modmult_1/zin[1][107] , \modmult_1/zin[1][106] ,
         \modmult_1/zin[1][105] , \modmult_1/zin[1][104] ,
         \modmult_1/zin[1][103] , \modmult_1/zin[1][102] ,
         \modmult_1/zin[1][101] , \modmult_1/zin[1][100] ,
         \modmult_1/zin[1][99] , \modmult_1/zin[1][98] ,
         \modmult_1/zin[1][97] , \modmult_1/zin[1][96] ,
         \modmult_1/zin[1][95] , \modmult_1/zin[1][94] ,
         \modmult_1/zin[1][93] , \modmult_1/zin[1][92] ,
         \modmult_1/zin[1][91] , \modmult_1/zin[1][90] ,
         \modmult_1/zin[1][89] , \modmult_1/zin[1][88] ,
         \modmult_1/zin[1][87] , \modmult_1/zin[1][86] ,
         \modmult_1/zin[1][85] , \modmult_1/zin[1][84] ,
         \modmult_1/zin[1][83] , \modmult_1/zin[1][82] ,
         \modmult_1/zin[1][81] , \modmult_1/zin[1][80] ,
         \modmult_1/zin[1][79] , \modmult_1/zin[1][78] ,
         \modmult_1/zin[1][77] , \modmult_1/zin[1][76] ,
         \modmult_1/zin[1][75] , \modmult_1/zin[1][74] ,
         \modmult_1/zin[1][73] , \modmult_1/zin[1][72] ,
         \modmult_1/zin[1][71] , \modmult_1/zin[1][70] ,
         \modmult_1/zin[1][69] , \modmult_1/zin[1][68] ,
         \modmult_1/zin[1][67] , \modmult_1/zin[1][66] ,
         \modmult_1/zin[1][65] , \modmult_1/zin[1][64] ,
         \modmult_1/zin[1][63] , \modmult_1/zin[1][62] ,
         \modmult_1/zin[1][61] , \modmult_1/zin[1][60] ,
         \modmult_1/zin[1][59] , \modmult_1/zin[1][58] ,
         \modmult_1/zin[1][57] , \modmult_1/zin[1][56] ,
         \modmult_1/zin[1][55] , \modmult_1/zin[1][54] ,
         \modmult_1/zin[1][53] , \modmult_1/zin[1][52] ,
         \modmult_1/zin[1][51] , \modmult_1/zin[1][50] ,
         \modmult_1/zin[1][49] , \modmult_1/zin[1][48] ,
         \modmult_1/zin[1][47] , \modmult_1/zin[1][46] ,
         \modmult_1/zin[1][45] , \modmult_1/zin[1][44] ,
         \modmult_1/zin[1][43] , \modmult_1/zin[1][42] ,
         \modmult_1/zin[1][41] , \modmult_1/zin[1][40] ,
         \modmult_1/zin[1][39] , \modmult_1/zin[1][38] ,
         \modmult_1/zin[1][37] , \modmult_1/zin[1][36] ,
         \modmult_1/zin[1][35] , \modmult_1/zin[1][34] ,
         \modmult_1/zin[1][33] , \modmult_1/zin[1][32] ,
         \modmult_1/zin[1][31] , \modmult_1/zin[1][30] ,
         \modmult_1/zin[1][29] , \modmult_1/zin[1][28] ,
         \modmult_1/zin[1][27] , \modmult_1/zin[1][26] ,
         \modmult_1/zin[1][25] , \modmult_1/zin[1][24] ,
         \modmult_1/zin[1][23] , \modmult_1/zin[1][22] ,
         \modmult_1/zin[1][21] , \modmult_1/zin[1][20] ,
         \modmult_1/zin[1][19] , \modmult_1/zin[1][18] ,
         \modmult_1/zin[1][17] , \modmult_1/zin[1][16] ,
         \modmult_1/zin[1][15] , \modmult_1/zin[1][14] ,
         \modmult_1/zin[1][13] , \modmult_1/zin[1][12] ,
         \modmult_1/zin[1][11] , \modmult_1/zin[1][10] , \modmult_1/zin[1][9] ,
         \modmult_1/zin[1][8] , \modmult_1/zin[1][7] , \modmult_1/zin[1][6] ,
         \modmult_1/zin[1][5] , \modmult_1/zin[1][4] , \modmult_1/zin[1][3] ,
         \modmult_1/zin[1][2] , \modmult_1/zin[1][1] , \modmult_1/zin[1][0] ,
         \modmult_1/zin[0][256] , \modmult_1/zin[0][255] ,
         \modmult_1/zin[0][254] , \modmult_1/zin[0][253] ,
         \modmult_1/zin[0][252] , \modmult_1/zin[0][251] ,
         \modmult_1/zin[0][250] , \modmult_1/zin[0][249] ,
         \modmult_1/zin[0][248] , \modmult_1/zin[0][247] ,
         \modmult_1/zin[0][246] , \modmult_1/zin[0][245] ,
         \modmult_1/zin[0][244] , \modmult_1/zin[0][243] ,
         \modmult_1/zin[0][242] , \modmult_1/zin[0][241] ,
         \modmult_1/zin[0][240] , \modmult_1/zin[0][239] ,
         \modmult_1/zin[0][238] , \modmult_1/zin[0][237] ,
         \modmult_1/zin[0][236] , \modmult_1/zin[0][235] ,
         \modmult_1/zin[0][234] , \modmult_1/zin[0][233] ,
         \modmult_1/zin[0][232] , \modmult_1/zin[0][231] ,
         \modmult_1/zin[0][230] , \modmult_1/zin[0][229] ,
         \modmult_1/zin[0][228] , \modmult_1/zin[0][227] ,
         \modmult_1/zin[0][226] , \modmult_1/zin[0][225] ,
         \modmult_1/zin[0][224] , \modmult_1/zin[0][223] ,
         \modmult_1/zin[0][222] , \modmult_1/zin[0][221] ,
         \modmult_1/zin[0][220] , \modmult_1/zin[0][219] ,
         \modmult_1/zin[0][218] , \modmult_1/zin[0][217] ,
         \modmult_1/zin[0][216] , \modmult_1/zin[0][215] ,
         \modmult_1/zin[0][214] , \modmult_1/zin[0][213] ,
         \modmult_1/zin[0][212] , \modmult_1/zin[0][211] ,
         \modmult_1/zin[0][210] , \modmult_1/zin[0][209] ,
         \modmult_1/zin[0][208] , \modmult_1/zin[0][207] ,
         \modmult_1/zin[0][206] , \modmult_1/zin[0][205] ,
         \modmult_1/zin[0][204] , \modmult_1/zin[0][203] ,
         \modmult_1/zin[0][202] , \modmult_1/zin[0][201] ,
         \modmult_1/zin[0][200] , \modmult_1/zin[0][199] ,
         \modmult_1/zin[0][198] , \modmult_1/zin[0][197] ,
         \modmult_1/zin[0][196] , \modmult_1/zin[0][195] ,
         \modmult_1/zin[0][194] , \modmult_1/zin[0][193] ,
         \modmult_1/zin[0][192] , \modmult_1/zin[0][191] ,
         \modmult_1/zin[0][190] , \modmult_1/zin[0][189] ,
         \modmult_1/zin[0][188] , \modmult_1/zin[0][187] ,
         \modmult_1/zin[0][186] , \modmult_1/zin[0][185] ,
         \modmult_1/zin[0][184] , \modmult_1/zin[0][183] ,
         \modmult_1/zin[0][182] , \modmult_1/zin[0][181] ,
         \modmult_1/zin[0][180] , \modmult_1/zin[0][179] ,
         \modmult_1/zin[0][178] , \modmult_1/zin[0][177] ,
         \modmult_1/zin[0][176] , \modmult_1/zin[0][175] ,
         \modmult_1/zin[0][174] , \modmult_1/zin[0][173] ,
         \modmult_1/zin[0][172] , \modmult_1/zin[0][171] ,
         \modmult_1/zin[0][170] , \modmult_1/zin[0][169] ,
         \modmult_1/zin[0][168] , \modmult_1/zin[0][167] ,
         \modmult_1/zin[0][166] , \modmult_1/zin[0][165] ,
         \modmult_1/zin[0][164] , \modmult_1/zin[0][163] ,
         \modmult_1/zin[0][162] , \modmult_1/zin[0][161] ,
         \modmult_1/zin[0][160] , \modmult_1/zin[0][159] ,
         \modmult_1/zin[0][158] , \modmult_1/zin[0][157] ,
         \modmult_1/zin[0][156] , \modmult_1/zin[0][155] ,
         \modmult_1/zin[0][154] , \modmult_1/zin[0][153] ,
         \modmult_1/zin[0][152] , \modmult_1/zin[0][151] ,
         \modmult_1/zin[0][150] , \modmult_1/zin[0][149] ,
         \modmult_1/zin[0][148] , \modmult_1/zin[0][147] ,
         \modmult_1/zin[0][146] , \modmult_1/zin[0][145] ,
         \modmult_1/zin[0][144] , \modmult_1/zin[0][143] ,
         \modmult_1/zin[0][142] , \modmult_1/zin[0][141] ,
         \modmult_1/zin[0][140] , \modmult_1/zin[0][139] ,
         \modmult_1/zin[0][138] , \modmult_1/zin[0][137] ,
         \modmult_1/zin[0][136] , \modmult_1/zin[0][135] ,
         \modmult_1/zin[0][134] , \modmult_1/zin[0][133] ,
         \modmult_1/zin[0][132] , \modmult_1/zin[0][131] ,
         \modmult_1/zin[0][130] , \modmult_1/zin[0][129] ,
         \modmult_1/zin[0][128] , \modmult_1/zin[0][127] ,
         \modmult_1/zin[0][126] , \modmult_1/zin[0][125] ,
         \modmult_1/zin[0][124] , \modmult_1/zin[0][123] ,
         \modmult_1/zin[0][122] , \modmult_1/zin[0][121] ,
         \modmult_1/zin[0][120] , \modmult_1/zin[0][119] ,
         \modmult_1/zin[0][118] , \modmult_1/zin[0][117] ,
         \modmult_1/zin[0][116] , \modmult_1/zin[0][115] ,
         \modmult_1/zin[0][114] , \modmult_1/zin[0][113] ,
         \modmult_1/zin[0][112] , \modmult_1/zin[0][111] ,
         \modmult_1/zin[0][110] , \modmult_1/zin[0][109] ,
         \modmult_1/zin[0][108] , \modmult_1/zin[0][107] ,
         \modmult_1/zin[0][106] , \modmult_1/zin[0][105] ,
         \modmult_1/zin[0][104] , \modmult_1/zin[0][103] ,
         \modmult_1/zin[0][102] , \modmult_1/zin[0][101] ,
         \modmult_1/zin[0][100] , \modmult_1/zin[0][99] ,
         \modmult_1/zin[0][98] , \modmult_1/zin[0][97] ,
         \modmult_1/zin[0][96] , \modmult_1/zin[0][95] ,
         \modmult_1/zin[0][94] , \modmult_1/zin[0][93] ,
         \modmult_1/zin[0][92] , \modmult_1/zin[0][91] ,
         \modmult_1/zin[0][90] , \modmult_1/zin[0][89] ,
         \modmult_1/zin[0][88] , \modmult_1/zin[0][87] ,
         \modmult_1/zin[0][86] , \modmult_1/zin[0][85] ,
         \modmult_1/zin[0][84] , \modmult_1/zin[0][83] ,
         \modmult_1/zin[0][82] , \modmult_1/zin[0][81] ,
         \modmult_1/zin[0][80] , \modmult_1/zin[0][79] ,
         \modmult_1/zin[0][78] , \modmult_1/zin[0][77] ,
         \modmult_1/zin[0][76] , \modmult_1/zin[0][75] ,
         \modmult_1/zin[0][74] , \modmult_1/zin[0][73] ,
         \modmult_1/zin[0][72] , \modmult_1/zin[0][71] ,
         \modmult_1/zin[0][70] , \modmult_1/zin[0][69] ,
         \modmult_1/zin[0][68] , \modmult_1/zin[0][67] ,
         \modmult_1/zin[0][66] , \modmult_1/zin[0][65] ,
         \modmult_1/zin[0][64] , \modmult_1/zin[0][63] ,
         \modmult_1/zin[0][62] , \modmult_1/zin[0][61] ,
         \modmult_1/zin[0][60] , \modmult_1/zin[0][59] ,
         \modmult_1/zin[0][58] , \modmult_1/zin[0][57] ,
         \modmult_1/zin[0][56] , \modmult_1/zin[0][55] ,
         \modmult_1/zin[0][54] , \modmult_1/zin[0][53] ,
         \modmult_1/zin[0][52] , \modmult_1/zin[0][51] ,
         \modmult_1/zin[0][50] , \modmult_1/zin[0][49] ,
         \modmult_1/zin[0][48] , \modmult_1/zin[0][47] ,
         \modmult_1/zin[0][46] , \modmult_1/zin[0][45] ,
         \modmult_1/zin[0][44] , \modmult_1/zin[0][43] ,
         \modmult_1/zin[0][42] , \modmult_1/zin[0][41] ,
         \modmult_1/zin[0][40] , \modmult_1/zin[0][39] ,
         \modmult_1/zin[0][38] , \modmult_1/zin[0][37] ,
         \modmult_1/zin[0][36] , \modmult_1/zin[0][35] ,
         \modmult_1/zin[0][34] , \modmult_1/zin[0][33] ,
         \modmult_1/zin[0][32] , \modmult_1/zin[0][31] ,
         \modmult_1/zin[0][30] , \modmult_1/zin[0][29] ,
         \modmult_1/zin[0][28] , \modmult_1/zin[0][27] ,
         \modmult_1/zin[0][26] , \modmult_1/zin[0][25] ,
         \modmult_1/zin[0][24] , \modmult_1/zin[0][23] ,
         \modmult_1/zin[0][22] , \modmult_1/zin[0][21] ,
         \modmult_1/zin[0][20] , \modmult_1/zin[0][19] ,
         \modmult_1/zin[0][18] , \modmult_1/zin[0][17] ,
         \modmult_1/zin[0][16] , \modmult_1/zin[0][15] ,
         \modmult_1/zin[0][14] , \modmult_1/zin[0][13] ,
         \modmult_1/zin[0][12] , \modmult_1/zin[0][11] ,
         \modmult_1/zin[0][10] , \modmult_1/zin[0][9] , \modmult_1/zin[0][8] ,
         \modmult_1/zin[0][7] , \modmult_1/zin[0][6] , \modmult_1/zin[0][5] ,
         \modmult_1/zin[0][4] , \modmult_1/zin[0][3] , \modmult_1/zin[0][2] ,
         \modmult_1/zin[0][1] , \modmult_1/zin[0][0] , \modmult_1/zreg[256] ,
         \modmult_1/zreg[255] , \modmult_1/zreg[254] , \modmult_1/zreg[253] ,
         \modmult_1/zreg[252] , \modmult_1/zreg[251] , \modmult_1/zreg[250] ,
         \modmult_1/zreg[249] , \modmult_1/zreg[248] , \modmult_1/zreg[247] ,
         \modmult_1/zreg[246] , \modmult_1/zreg[245] , \modmult_1/zreg[244] ,
         \modmult_1/zreg[243] , \modmult_1/zreg[242] , \modmult_1/zreg[241] ,
         \modmult_1/zreg[240] , \modmult_1/zreg[239] , \modmult_1/zreg[238] ,
         \modmult_1/zreg[237] , \modmult_1/zreg[236] , \modmult_1/zreg[235] ,
         \modmult_1/zreg[234] , \modmult_1/zreg[233] , \modmult_1/zreg[232] ,
         \modmult_1/zreg[231] , \modmult_1/zreg[230] , \modmult_1/zreg[229] ,
         \modmult_1/zreg[228] , \modmult_1/zreg[227] , \modmult_1/zreg[226] ,
         \modmult_1/zreg[225] , \modmult_1/zreg[224] , \modmult_1/zreg[223] ,
         \modmult_1/zreg[222] , \modmult_1/zreg[221] , \modmult_1/zreg[220] ,
         \modmult_1/zreg[219] , \modmult_1/zreg[218] , \modmult_1/zreg[217] ,
         \modmult_1/zreg[216] , \modmult_1/zreg[215] , \modmult_1/zreg[214] ,
         \modmult_1/zreg[213] , \modmult_1/zreg[212] , \modmult_1/zreg[211] ,
         \modmult_1/zreg[210] , \modmult_1/zreg[209] , \modmult_1/zreg[208] ,
         \modmult_1/zreg[207] , \modmult_1/zreg[206] , \modmult_1/zreg[205] ,
         \modmult_1/zreg[204] , \modmult_1/zreg[203] , \modmult_1/zreg[202] ,
         \modmult_1/zreg[201] , \modmult_1/zreg[200] , \modmult_1/zreg[199] ,
         \modmult_1/zreg[198] , \modmult_1/zreg[197] , \modmult_1/zreg[196] ,
         \modmult_1/zreg[195] , \modmult_1/zreg[194] , \modmult_1/zreg[193] ,
         \modmult_1/zreg[192] , \modmult_1/zreg[191] , \modmult_1/zreg[190] ,
         \modmult_1/zreg[189] , \modmult_1/zreg[188] , \modmult_1/zreg[187] ,
         \modmult_1/zreg[186] , \modmult_1/zreg[185] , \modmult_1/zreg[184] ,
         \modmult_1/zreg[183] , \modmult_1/zreg[182] , \modmult_1/zreg[181] ,
         \modmult_1/zreg[180] , \modmult_1/zreg[179] , \modmult_1/zreg[178] ,
         \modmult_1/zreg[177] , \modmult_1/zreg[176] , \modmult_1/zreg[175] ,
         \modmult_1/zreg[174] , \modmult_1/zreg[173] , \modmult_1/zreg[172] ,
         \modmult_1/zreg[171] , \modmult_1/zreg[170] , \modmult_1/zreg[169] ,
         \modmult_1/zreg[168] , \modmult_1/zreg[167] , \modmult_1/zreg[166] ,
         \modmult_1/zreg[165] , \modmult_1/zreg[164] , \modmult_1/zreg[163] ,
         \modmult_1/zreg[162] , \modmult_1/zreg[161] , \modmult_1/zreg[160] ,
         \modmult_1/zreg[159] , \modmult_1/zreg[158] , \modmult_1/zreg[157] ,
         \modmult_1/zreg[156] , \modmult_1/zreg[155] , \modmult_1/zreg[154] ,
         \modmult_1/zreg[153] , \modmult_1/zreg[152] , \modmult_1/zreg[151] ,
         \modmult_1/zreg[150] , \modmult_1/zreg[149] , \modmult_1/zreg[148] ,
         \modmult_1/zreg[147] , \modmult_1/zreg[146] , \modmult_1/zreg[145] ,
         \modmult_1/zreg[144] , \modmult_1/zreg[143] , \modmult_1/zreg[142] ,
         \modmult_1/zreg[141] , \modmult_1/zreg[140] , \modmult_1/zreg[139] ,
         \modmult_1/zreg[138] , \modmult_1/zreg[137] , \modmult_1/zreg[136] ,
         \modmult_1/zreg[135] , \modmult_1/zreg[134] , \modmult_1/zreg[133] ,
         \modmult_1/zreg[132] , \modmult_1/zreg[131] , \modmult_1/zreg[130] ,
         \modmult_1/zreg[129] , \modmult_1/zreg[128] , \modmult_1/zreg[127] ,
         \modmult_1/zreg[126] , \modmult_1/zreg[125] , \modmult_1/zreg[124] ,
         \modmult_1/zreg[123] , \modmult_1/zreg[122] , \modmult_1/zreg[121] ,
         \modmult_1/zreg[120] , \modmult_1/zreg[119] , \modmult_1/zreg[118] ,
         \modmult_1/zreg[117] , \modmult_1/zreg[116] , \modmult_1/zreg[115] ,
         \modmult_1/zreg[114] , \modmult_1/zreg[113] , \modmult_1/zreg[112] ,
         \modmult_1/zreg[111] , \modmult_1/zreg[110] , \modmult_1/zreg[109] ,
         \modmult_1/zreg[108] , \modmult_1/zreg[107] , \modmult_1/zreg[106] ,
         \modmult_1/zreg[105] , \modmult_1/zreg[104] , \modmult_1/zreg[103] ,
         \modmult_1/zreg[102] , \modmult_1/zreg[101] , \modmult_1/zreg[100] ,
         \modmult_1/zreg[99] , \modmult_1/zreg[98] , \modmult_1/zreg[97] ,
         \modmult_1/zreg[96] , \modmult_1/zreg[95] , \modmult_1/zreg[94] ,
         \modmult_1/zreg[93] , \modmult_1/zreg[92] , \modmult_1/zreg[91] ,
         \modmult_1/zreg[90] , \modmult_1/zreg[89] , \modmult_1/zreg[88] ,
         \modmult_1/zreg[87] , \modmult_1/zreg[86] , \modmult_1/zreg[85] ,
         \modmult_1/zreg[84] , \modmult_1/zreg[83] , \modmult_1/zreg[82] ,
         \modmult_1/zreg[81] , \modmult_1/zreg[80] , \modmult_1/zreg[79] ,
         \modmult_1/zreg[78] , \modmult_1/zreg[77] , \modmult_1/zreg[76] ,
         \modmult_1/zreg[75] , \modmult_1/zreg[74] , \modmult_1/zreg[73] ,
         \modmult_1/zreg[72] , \modmult_1/zreg[71] , \modmult_1/zreg[70] ,
         \modmult_1/zreg[69] , \modmult_1/zreg[68] , \modmult_1/zreg[67] ,
         \modmult_1/zreg[66] , \modmult_1/zreg[65] , \modmult_1/zreg[64] ,
         \modmult_1/zreg[63] , \modmult_1/zreg[62] , \modmult_1/zreg[61] ,
         \modmult_1/zreg[60] , \modmult_1/zreg[59] , \modmult_1/zreg[58] ,
         \modmult_1/zreg[57] , \modmult_1/zreg[56] , \modmult_1/zreg[55] ,
         \modmult_1/zreg[54] , \modmult_1/zreg[53] , \modmult_1/zreg[52] ,
         \modmult_1/zreg[51] , \modmult_1/zreg[50] , \modmult_1/zreg[49] ,
         \modmult_1/zreg[48] , \modmult_1/zreg[47] , \modmult_1/zreg[46] ,
         \modmult_1/zreg[45] , \modmult_1/zreg[44] , \modmult_1/zreg[43] ,
         \modmult_1/zreg[42] , \modmult_1/zreg[41] , \modmult_1/zreg[40] ,
         \modmult_1/zreg[39] , \modmult_1/zreg[38] , \modmult_1/zreg[37] ,
         \modmult_1/zreg[36] , \modmult_1/zreg[35] , \modmult_1/zreg[34] ,
         \modmult_1/zreg[33] , \modmult_1/zreg[32] , \modmult_1/zreg[31] ,
         \modmult_1/zreg[30] , \modmult_1/zreg[29] , \modmult_1/zreg[28] ,
         \modmult_1/zreg[27] , \modmult_1/zreg[26] , \modmult_1/zreg[25] ,
         \modmult_1/zreg[24] , \modmult_1/zreg[23] , \modmult_1/zreg[22] ,
         \modmult_1/zreg[21] , \modmult_1/zreg[20] , \modmult_1/zreg[19] ,
         \modmult_1/zreg[18] , \modmult_1/zreg[17] , \modmult_1/zreg[16] ,
         \modmult_1/zreg[15] , \modmult_1/zreg[14] , \modmult_1/zreg[13] ,
         \modmult_1/zreg[12] , \modmult_1/zreg[11] , \modmult_1/zreg[10] ,
         \modmult_1/zreg[9] , \modmult_1/zreg[8] , \modmult_1/zreg[7] ,
         \modmult_1/zreg[6] , \modmult_1/zreg[5] , \modmult_1/zreg[4] ,
         \modmult_1/zreg[3] , \modmult_1/zreg[2] , \modmult_1/zreg[1] ,
         \modmult_1/zreg[0] , \modmult_1/zout[1][256] , n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214;
  wire   [127:0] start_in;
  wire   [127:0] start_reg;
  wire   [255:0] ereg;
  wire   [255:0] o;
  wire   [255:0] creg;
  wire   [255:0] y;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  modmult_step_N256_1 \modmult_1/MODMULT_STEP[1].modmult_step_  ( .xregN_1(
        \modmult_1/xin[254] ), .y(y), .n(n), .zin({1'b0, 
        \modmult_1/zin[1][256] , \modmult_1/zin[1][255] , 
        \modmult_1/zin[1][254] , \modmult_1/zin[1][253] , 
        \modmult_1/zin[1][252] , \modmult_1/zin[1][251] , 
        \modmult_1/zin[1][250] , \modmult_1/zin[1][249] , 
        \modmult_1/zin[1][248] , \modmult_1/zin[1][247] , 
        \modmult_1/zin[1][246] , \modmult_1/zin[1][245] , 
        \modmult_1/zin[1][244] , \modmult_1/zin[1][243] , 
        \modmult_1/zin[1][242] , \modmult_1/zin[1][241] , 
        \modmult_1/zin[1][240] , \modmult_1/zin[1][239] , 
        \modmult_1/zin[1][238] , \modmult_1/zin[1][237] , 
        \modmult_1/zin[1][236] , \modmult_1/zin[1][235] , 
        \modmult_1/zin[1][234] , \modmult_1/zin[1][233] , 
        \modmult_1/zin[1][232] , \modmult_1/zin[1][231] , 
        \modmult_1/zin[1][230] , \modmult_1/zin[1][229] , 
        \modmult_1/zin[1][228] , \modmult_1/zin[1][227] , 
        \modmult_1/zin[1][226] , \modmult_1/zin[1][225] , 
        \modmult_1/zin[1][224] , \modmult_1/zin[1][223] , 
        \modmult_1/zin[1][222] , \modmult_1/zin[1][221] , 
        \modmult_1/zin[1][220] , \modmult_1/zin[1][219] , 
        \modmult_1/zin[1][218] , \modmult_1/zin[1][217] , 
        \modmult_1/zin[1][216] , \modmult_1/zin[1][215] , 
        \modmult_1/zin[1][214] , \modmult_1/zin[1][213] , 
        \modmult_1/zin[1][212] , \modmult_1/zin[1][211] , 
        \modmult_1/zin[1][210] , \modmult_1/zin[1][209] , 
        \modmult_1/zin[1][208] , \modmult_1/zin[1][207] , 
        \modmult_1/zin[1][206] , \modmult_1/zin[1][205] , 
        \modmult_1/zin[1][204] , \modmult_1/zin[1][203] , 
        \modmult_1/zin[1][202] , \modmult_1/zin[1][201] , 
        \modmult_1/zin[1][200] , \modmult_1/zin[1][199] , 
        \modmult_1/zin[1][198] , \modmult_1/zin[1][197] , 
        \modmult_1/zin[1][196] , \modmult_1/zin[1][195] , 
        \modmult_1/zin[1][194] , \modmult_1/zin[1][193] , 
        \modmult_1/zin[1][192] , \modmult_1/zin[1][191] , 
        \modmult_1/zin[1][190] , \modmult_1/zin[1][189] , 
        \modmult_1/zin[1][188] , \modmult_1/zin[1][187] , 
        \modmult_1/zin[1][186] , \modmult_1/zin[1][185] , 
        \modmult_1/zin[1][184] , \modmult_1/zin[1][183] , 
        \modmult_1/zin[1][182] , \modmult_1/zin[1][181] , 
        \modmult_1/zin[1][180] , \modmult_1/zin[1][179] , 
        \modmult_1/zin[1][178] , \modmult_1/zin[1][177] , 
        \modmult_1/zin[1][176] , \modmult_1/zin[1][175] , 
        \modmult_1/zin[1][174] , \modmult_1/zin[1][173] , 
        \modmult_1/zin[1][172] , \modmult_1/zin[1][171] , 
        \modmult_1/zin[1][170] , \modmult_1/zin[1][169] , 
        \modmult_1/zin[1][168] , \modmult_1/zin[1][167] , 
        \modmult_1/zin[1][166] , \modmult_1/zin[1][165] , 
        \modmult_1/zin[1][164] , \modmult_1/zin[1][163] , 
        \modmult_1/zin[1][162] , \modmult_1/zin[1][161] , 
        \modmult_1/zin[1][160] , \modmult_1/zin[1][159] , 
        \modmult_1/zin[1][158] , \modmult_1/zin[1][157] , 
        \modmult_1/zin[1][156] , \modmult_1/zin[1][155] , 
        \modmult_1/zin[1][154] , \modmult_1/zin[1][153] , 
        \modmult_1/zin[1][152] , \modmult_1/zin[1][151] , 
        \modmult_1/zin[1][150] , \modmult_1/zin[1][149] , 
        \modmult_1/zin[1][148] , \modmult_1/zin[1][147] , 
        \modmult_1/zin[1][146] , \modmult_1/zin[1][145] , 
        \modmult_1/zin[1][144] , \modmult_1/zin[1][143] , 
        \modmult_1/zin[1][142] , \modmult_1/zin[1][141] , 
        \modmult_1/zin[1][140] , \modmult_1/zin[1][139] , 
        \modmult_1/zin[1][138] , \modmult_1/zin[1][137] , 
        \modmult_1/zin[1][136] , \modmult_1/zin[1][135] , 
        \modmult_1/zin[1][134] , \modmult_1/zin[1][133] , 
        \modmult_1/zin[1][132] , \modmult_1/zin[1][131] , 
        \modmult_1/zin[1][130] , \modmult_1/zin[1][129] , 
        \modmult_1/zin[1][128] , \modmult_1/zin[1][127] , 
        \modmult_1/zin[1][126] , \modmult_1/zin[1][125] , 
        \modmult_1/zin[1][124] , \modmult_1/zin[1][123] , 
        \modmult_1/zin[1][122] , \modmult_1/zin[1][121] , 
        \modmult_1/zin[1][120] , \modmult_1/zin[1][119] , 
        \modmult_1/zin[1][118] , \modmult_1/zin[1][117] , 
        \modmult_1/zin[1][116] , \modmult_1/zin[1][115] , 
        \modmult_1/zin[1][114] , \modmult_1/zin[1][113] , 
        \modmult_1/zin[1][112] , \modmult_1/zin[1][111] , 
        \modmult_1/zin[1][110] , \modmult_1/zin[1][109] , 
        \modmult_1/zin[1][108] , \modmult_1/zin[1][107] , 
        \modmult_1/zin[1][106] , \modmult_1/zin[1][105] , 
        \modmult_1/zin[1][104] , \modmult_1/zin[1][103] , 
        \modmult_1/zin[1][102] , \modmult_1/zin[1][101] , 
        \modmult_1/zin[1][100] , \modmult_1/zin[1][99] , 
        \modmult_1/zin[1][98] , \modmult_1/zin[1][97] , \modmult_1/zin[1][96] , 
        \modmult_1/zin[1][95] , \modmult_1/zin[1][94] , \modmult_1/zin[1][93] , 
        \modmult_1/zin[1][92] , \modmult_1/zin[1][91] , \modmult_1/zin[1][90] , 
        \modmult_1/zin[1][89] , \modmult_1/zin[1][88] , \modmult_1/zin[1][87] , 
        \modmult_1/zin[1][86] , \modmult_1/zin[1][85] , \modmult_1/zin[1][84] , 
        \modmult_1/zin[1][83] , \modmult_1/zin[1][82] , \modmult_1/zin[1][81] , 
        \modmult_1/zin[1][80] , \modmult_1/zin[1][79] , \modmult_1/zin[1][78] , 
        \modmult_1/zin[1][77] , \modmult_1/zin[1][76] , \modmult_1/zin[1][75] , 
        \modmult_1/zin[1][74] , \modmult_1/zin[1][73] , \modmult_1/zin[1][72] , 
        \modmult_1/zin[1][71] , \modmult_1/zin[1][70] , \modmult_1/zin[1][69] , 
        \modmult_1/zin[1][68] , \modmult_1/zin[1][67] , \modmult_1/zin[1][66] , 
        \modmult_1/zin[1][65] , \modmult_1/zin[1][64] , \modmult_1/zin[1][63] , 
        \modmult_1/zin[1][62] , \modmult_1/zin[1][61] , \modmult_1/zin[1][60] , 
        \modmult_1/zin[1][59] , \modmult_1/zin[1][58] , \modmult_1/zin[1][57] , 
        \modmult_1/zin[1][56] , \modmult_1/zin[1][55] , \modmult_1/zin[1][54] , 
        \modmult_1/zin[1][53] , \modmult_1/zin[1][52] , \modmult_1/zin[1][51] , 
        \modmult_1/zin[1][50] , \modmult_1/zin[1][49] , \modmult_1/zin[1][48] , 
        \modmult_1/zin[1][47] , \modmult_1/zin[1][46] , \modmult_1/zin[1][45] , 
        \modmult_1/zin[1][44] , \modmult_1/zin[1][43] , \modmult_1/zin[1][42] , 
        \modmult_1/zin[1][41] , \modmult_1/zin[1][40] , \modmult_1/zin[1][39] , 
        \modmult_1/zin[1][38] , \modmult_1/zin[1][37] , \modmult_1/zin[1][36] , 
        \modmult_1/zin[1][35] , \modmult_1/zin[1][34] , \modmult_1/zin[1][33] , 
        \modmult_1/zin[1][32] , \modmult_1/zin[1][31] , \modmult_1/zin[1][30] , 
        \modmult_1/zin[1][29] , \modmult_1/zin[1][28] , \modmult_1/zin[1][27] , 
        \modmult_1/zin[1][26] , \modmult_1/zin[1][25] , \modmult_1/zin[1][24] , 
        \modmult_1/zin[1][23] , \modmult_1/zin[1][22] , \modmult_1/zin[1][21] , 
        \modmult_1/zin[1][20] , \modmult_1/zin[1][19] , \modmult_1/zin[1][18] , 
        \modmult_1/zin[1][17] , \modmult_1/zin[1][16] , \modmult_1/zin[1][15] , 
        \modmult_1/zin[1][14] , \modmult_1/zin[1][13] , \modmult_1/zin[1][12] , 
        \modmult_1/zin[1][11] , \modmult_1/zin[1][10] , \modmult_1/zin[1][9] , 
        \modmult_1/zin[1][8] , \modmult_1/zin[1][7] , \modmult_1/zin[1][6] , 
        \modmult_1/zin[1][5] , \modmult_1/zin[1][4] , \modmult_1/zin[1][3] , 
        \modmult_1/zin[1][2] , \modmult_1/zin[1][1] , \modmult_1/zin[1][0] }), 
        .zout({SYNOPSYS_UNCONNECTED__0, \modmult_1/zout[1][256] , o}) );
  modmult_step_N256_0 \modmult_1/MODMULT_STEP[0].modmult_step_  ( .xregN_1(
        \modmult_1/xin[255] ), .y(y), .n(n), .zin({1'b0, 
        \modmult_1/zin[0][256] , \modmult_1/zin[0][255] , 
        \modmult_1/zin[0][254] , \modmult_1/zin[0][253] , 
        \modmult_1/zin[0][252] , \modmult_1/zin[0][251] , 
        \modmult_1/zin[0][250] , \modmult_1/zin[0][249] , 
        \modmult_1/zin[0][248] , \modmult_1/zin[0][247] , 
        \modmult_1/zin[0][246] , \modmult_1/zin[0][245] , 
        \modmult_1/zin[0][244] , \modmult_1/zin[0][243] , 
        \modmult_1/zin[0][242] , \modmult_1/zin[0][241] , 
        \modmult_1/zin[0][240] , \modmult_1/zin[0][239] , 
        \modmult_1/zin[0][238] , \modmult_1/zin[0][237] , 
        \modmult_1/zin[0][236] , \modmult_1/zin[0][235] , 
        \modmult_1/zin[0][234] , \modmult_1/zin[0][233] , 
        \modmult_1/zin[0][232] , \modmult_1/zin[0][231] , 
        \modmult_1/zin[0][230] , \modmult_1/zin[0][229] , 
        \modmult_1/zin[0][228] , \modmult_1/zin[0][227] , 
        \modmult_1/zin[0][226] , \modmult_1/zin[0][225] , 
        \modmult_1/zin[0][224] , \modmult_1/zin[0][223] , 
        \modmult_1/zin[0][222] , \modmult_1/zin[0][221] , 
        \modmult_1/zin[0][220] , \modmult_1/zin[0][219] , 
        \modmult_1/zin[0][218] , \modmult_1/zin[0][217] , 
        \modmult_1/zin[0][216] , \modmult_1/zin[0][215] , 
        \modmult_1/zin[0][214] , \modmult_1/zin[0][213] , 
        \modmult_1/zin[0][212] , \modmult_1/zin[0][211] , 
        \modmult_1/zin[0][210] , \modmult_1/zin[0][209] , 
        \modmult_1/zin[0][208] , \modmult_1/zin[0][207] , 
        \modmult_1/zin[0][206] , \modmult_1/zin[0][205] , 
        \modmult_1/zin[0][204] , \modmult_1/zin[0][203] , 
        \modmult_1/zin[0][202] , \modmult_1/zin[0][201] , 
        \modmult_1/zin[0][200] , \modmult_1/zin[0][199] , 
        \modmult_1/zin[0][198] , \modmult_1/zin[0][197] , 
        \modmult_1/zin[0][196] , \modmult_1/zin[0][195] , 
        \modmult_1/zin[0][194] , \modmult_1/zin[0][193] , 
        \modmult_1/zin[0][192] , \modmult_1/zin[0][191] , 
        \modmult_1/zin[0][190] , \modmult_1/zin[0][189] , 
        \modmult_1/zin[0][188] , \modmult_1/zin[0][187] , 
        \modmult_1/zin[0][186] , \modmult_1/zin[0][185] , 
        \modmult_1/zin[0][184] , \modmult_1/zin[0][183] , 
        \modmult_1/zin[0][182] , \modmult_1/zin[0][181] , 
        \modmult_1/zin[0][180] , \modmult_1/zin[0][179] , 
        \modmult_1/zin[0][178] , \modmult_1/zin[0][177] , 
        \modmult_1/zin[0][176] , \modmult_1/zin[0][175] , 
        \modmult_1/zin[0][174] , \modmult_1/zin[0][173] , 
        \modmult_1/zin[0][172] , \modmult_1/zin[0][171] , 
        \modmult_1/zin[0][170] , \modmult_1/zin[0][169] , 
        \modmult_1/zin[0][168] , \modmult_1/zin[0][167] , 
        \modmult_1/zin[0][166] , \modmult_1/zin[0][165] , 
        \modmult_1/zin[0][164] , \modmult_1/zin[0][163] , 
        \modmult_1/zin[0][162] , \modmult_1/zin[0][161] , 
        \modmult_1/zin[0][160] , \modmult_1/zin[0][159] , 
        \modmult_1/zin[0][158] , \modmult_1/zin[0][157] , 
        \modmult_1/zin[0][156] , \modmult_1/zin[0][155] , 
        \modmult_1/zin[0][154] , \modmult_1/zin[0][153] , 
        \modmult_1/zin[0][152] , \modmult_1/zin[0][151] , 
        \modmult_1/zin[0][150] , \modmult_1/zin[0][149] , 
        \modmult_1/zin[0][148] , \modmult_1/zin[0][147] , 
        \modmult_1/zin[0][146] , \modmult_1/zin[0][145] , 
        \modmult_1/zin[0][144] , \modmult_1/zin[0][143] , 
        \modmult_1/zin[0][142] , \modmult_1/zin[0][141] , 
        \modmult_1/zin[0][140] , \modmult_1/zin[0][139] , 
        \modmult_1/zin[0][138] , \modmult_1/zin[0][137] , 
        \modmult_1/zin[0][136] , \modmult_1/zin[0][135] , 
        \modmult_1/zin[0][134] , \modmult_1/zin[0][133] , 
        \modmult_1/zin[0][132] , \modmult_1/zin[0][131] , 
        \modmult_1/zin[0][130] , \modmult_1/zin[0][129] , 
        \modmult_1/zin[0][128] , \modmult_1/zin[0][127] , 
        \modmult_1/zin[0][126] , \modmult_1/zin[0][125] , 
        \modmult_1/zin[0][124] , \modmult_1/zin[0][123] , 
        \modmult_1/zin[0][122] , \modmult_1/zin[0][121] , 
        \modmult_1/zin[0][120] , \modmult_1/zin[0][119] , 
        \modmult_1/zin[0][118] , \modmult_1/zin[0][117] , 
        \modmult_1/zin[0][116] , \modmult_1/zin[0][115] , 
        \modmult_1/zin[0][114] , \modmult_1/zin[0][113] , 
        \modmult_1/zin[0][112] , \modmult_1/zin[0][111] , 
        \modmult_1/zin[0][110] , \modmult_1/zin[0][109] , 
        \modmult_1/zin[0][108] , \modmult_1/zin[0][107] , 
        \modmult_1/zin[0][106] , \modmult_1/zin[0][105] , 
        \modmult_1/zin[0][104] , \modmult_1/zin[0][103] , 
        \modmult_1/zin[0][102] , \modmult_1/zin[0][101] , 
        \modmult_1/zin[0][100] , \modmult_1/zin[0][99] , 
        \modmult_1/zin[0][98] , \modmult_1/zin[0][97] , \modmult_1/zin[0][96] , 
        \modmult_1/zin[0][95] , \modmult_1/zin[0][94] , \modmult_1/zin[0][93] , 
        \modmult_1/zin[0][92] , \modmult_1/zin[0][91] , \modmult_1/zin[0][90] , 
        \modmult_1/zin[0][89] , \modmult_1/zin[0][88] , \modmult_1/zin[0][87] , 
        \modmult_1/zin[0][86] , \modmult_1/zin[0][85] , \modmult_1/zin[0][84] , 
        \modmult_1/zin[0][83] , \modmult_1/zin[0][82] , \modmult_1/zin[0][81] , 
        \modmult_1/zin[0][80] , \modmult_1/zin[0][79] , \modmult_1/zin[0][78] , 
        \modmult_1/zin[0][77] , \modmult_1/zin[0][76] , \modmult_1/zin[0][75] , 
        \modmult_1/zin[0][74] , \modmult_1/zin[0][73] , \modmult_1/zin[0][72] , 
        \modmult_1/zin[0][71] , \modmult_1/zin[0][70] , \modmult_1/zin[0][69] , 
        \modmult_1/zin[0][68] , \modmult_1/zin[0][67] , \modmult_1/zin[0][66] , 
        \modmult_1/zin[0][65] , \modmult_1/zin[0][64] , \modmult_1/zin[0][63] , 
        \modmult_1/zin[0][62] , \modmult_1/zin[0][61] , \modmult_1/zin[0][60] , 
        \modmult_1/zin[0][59] , \modmult_1/zin[0][58] , \modmult_1/zin[0][57] , 
        \modmult_1/zin[0][56] , \modmult_1/zin[0][55] , \modmult_1/zin[0][54] , 
        \modmult_1/zin[0][53] , \modmult_1/zin[0][52] , \modmult_1/zin[0][51] , 
        \modmult_1/zin[0][50] , \modmult_1/zin[0][49] , \modmult_1/zin[0][48] , 
        \modmult_1/zin[0][47] , \modmult_1/zin[0][46] , \modmult_1/zin[0][45] , 
        \modmult_1/zin[0][44] , \modmult_1/zin[0][43] , \modmult_1/zin[0][42] , 
        \modmult_1/zin[0][41] , \modmult_1/zin[0][40] , \modmult_1/zin[0][39] , 
        \modmult_1/zin[0][38] , \modmult_1/zin[0][37] , \modmult_1/zin[0][36] , 
        \modmult_1/zin[0][35] , \modmult_1/zin[0][34] , \modmult_1/zin[0][33] , 
        \modmult_1/zin[0][32] , \modmult_1/zin[0][31] , \modmult_1/zin[0][30] , 
        \modmult_1/zin[0][29] , \modmult_1/zin[0][28] , \modmult_1/zin[0][27] , 
        \modmult_1/zin[0][26] , \modmult_1/zin[0][25] , \modmult_1/zin[0][24] , 
        \modmult_1/zin[0][23] , \modmult_1/zin[0][22] , \modmult_1/zin[0][21] , 
        \modmult_1/zin[0][20] , \modmult_1/zin[0][19] , \modmult_1/zin[0][18] , 
        \modmult_1/zin[0][17] , \modmult_1/zin[0][16] , \modmult_1/zin[0][15] , 
        \modmult_1/zin[0][14] , \modmult_1/zin[0][13] , \modmult_1/zin[0][12] , 
        \modmult_1/zin[0][11] , \modmult_1/zin[0][10] , \modmult_1/zin[0][9] , 
        \modmult_1/zin[0][8] , \modmult_1/zin[0][7] , \modmult_1/zin[0][6] , 
        \modmult_1/zin[0][5] , \modmult_1/zin[0][4] , \modmult_1/zin[0][3] , 
        \modmult_1/zin[0][2] , \modmult_1/zin[0][1] , \modmult_1/zin[0][0] }), 
        .zout({SYNOPSYS_UNCONNECTED__1, \modmult_1/zin[1][256] , 
        \modmult_1/zin[1][255] , \modmult_1/zin[1][254] , 
        \modmult_1/zin[1][253] , \modmult_1/zin[1][252] , 
        \modmult_1/zin[1][251] , \modmult_1/zin[1][250] , 
        \modmult_1/zin[1][249] , \modmult_1/zin[1][248] , 
        \modmult_1/zin[1][247] , \modmult_1/zin[1][246] , 
        \modmult_1/zin[1][245] , \modmult_1/zin[1][244] , 
        \modmult_1/zin[1][243] , \modmult_1/zin[1][242] , 
        \modmult_1/zin[1][241] , \modmult_1/zin[1][240] , 
        \modmult_1/zin[1][239] , \modmult_1/zin[1][238] , 
        \modmult_1/zin[1][237] , \modmult_1/zin[1][236] , 
        \modmult_1/zin[1][235] , \modmult_1/zin[1][234] , 
        \modmult_1/zin[1][233] , \modmult_1/zin[1][232] , 
        \modmult_1/zin[1][231] , \modmult_1/zin[1][230] , 
        \modmult_1/zin[1][229] , \modmult_1/zin[1][228] , 
        \modmult_1/zin[1][227] , \modmult_1/zin[1][226] , 
        \modmult_1/zin[1][225] , \modmult_1/zin[1][224] , 
        \modmult_1/zin[1][223] , \modmult_1/zin[1][222] , 
        \modmult_1/zin[1][221] , \modmult_1/zin[1][220] , 
        \modmult_1/zin[1][219] , \modmult_1/zin[1][218] , 
        \modmult_1/zin[1][217] , \modmult_1/zin[1][216] , 
        \modmult_1/zin[1][215] , \modmult_1/zin[1][214] , 
        \modmult_1/zin[1][213] , \modmult_1/zin[1][212] , 
        \modmult_1/zin[1][211] , \modmult_1/zin[1][210] , 
        \modmult_1/zin[1][209] , \modmult_1/zin[1][208] , 
        \modmult_1/zin[1][207] , \modmult_1/zin[1][206] , 
        \modmult_1/zin[1][205] , \modmult_1/zin[1][204] , 
        \modmult_1/zin[1][203] , \modmult_1/zin[1][202] , 
        \modmult_1/zin[1][201] , \modmult_1/zin[1][200] , 
        \modmult_1/zin[1][199] , \modmult_1/zin[1][198] , 
        \modmult_1/zin[1][197] , \modmult_1/zin[1][196] , 
        \modmult_1/zin[1][195] , \modmult_1/zin[1][194] , 
        \modmult_1/zin[1][193] , \modmult_1/zin[1][192] , 
        \modmult_1/zin[1][191] , \modmult_1/zin[1][190] , 
        \modmult_1/zin[1][189] , \modmult_1/zin[1][188] , 
        \modmult_1/zin[1][187] , \modmult_1/zin[1][186] , 
        \modmult_1/zin[1][185] , \modmult_1/zin[1][184] , 
        \modmult_1/zin[1][183] , \modmult_1/zin[1][182] , 
        \modmult_1/zin[1][181] , \modmult_1/zin[1][180] , 
        \modmult_1/zin[1][179] , \modmult_1/zin[1][178] , 
        \modmult_1/zin[1][177] , \modmult_1/zin[1][176] , 
        \modmult_1/zin[1][175] , \modmult_1/zin[1][174] , 
        \modmult_1/zin[1][173] , \modmult_1/zin[1][172] , 
        \modmult_1/zin[1][171] , \modmult_1/zin[1][170] , 
        \modmult_1/zin[1][169] , \modmult_1/zin[1][168] , 
        \modmult_1/zin[1][167] , \modmult_1/zin[1][166] , 
        \modmult_1/zin[1][165] , \modmult_1/zin[1][164] , 
        \modmult_1/zin[1][163] , \modmult_1/zin[1][162] , 
        \modmult_1/zin[1][161] , \modmult_1/zin[1][160] , 
        \modmult_1/zin[1][159] , \modmult_1/zin[1][158] , 
        \modmult_1/zin[1][157] , \modmult_1/zin[1][156] , 
        \modmult_1/zin[1][155] , \modmult_1/zin[1][154] , 
        \modmult_1/zin[1][153] , \modmult_1/zin[1][152] , 
        \modmult_1/zin[1][151] , \modmult_1/zin[1][150] , 
        \modmult_1/zin[1][149] , \modmult_1/zin[1][148] , 
        \modmult_1/zin[1][147] , \modmult_1/zin[1][146] , 
        \modmult_1/zin[1][145] , \modmult_1/zin[1][144] , 
        \modmult_1/zin[1][143] , \modmult_1/zin[1][142] , 
        \modmult_1/zin[1][141] , \modmult_1/zin[1][140] , 
        \modmult_1/zin[1][139] , \modmult_1/zin[1][138] , 
        \modmult_1/zin[1][137] , \modmult_1/zin[1][136] , 
        \modmult_1/zin[1][135] , \modmult_1/zin[1][134] , 
        \modmult_1/zin[1][133] , \modmult_1/zin[1][132] , 
        \modmult_1/zin[1][131] , \modmult_1/zin[1][130] , 
        \modmult_1/zin[1][129] , \modmult_1/zin[1][128] , 
        \modmult_1/zin[1][127] , \modmult_1/zin[1][126] , 
        \modmult_1/zin[1][125] , \modmult_1/zin[1][124] , 
        \modmult_1/zin[1][123] , \modmult_1/zin[1][122] , 
        \modmult_1/zin[1][121] , \modmult_1/zin[1][120] , 
        \modmult_1/zin[1][119] , \modmult_1/zin[1][118] , 
        \modmult_1/zin[1][117] , \modmult_1/zin[1][116] , 
        \modmult_1/zin[1][115] , \modmult_1/zin[1][114] , 
        \modmult_1/zin[1][113] , \modmult_1/zin[1][112] , 
        \modmult_1/zin[1][111] , \modmult_1/zin[1][110] , 
        \modmult_1/zin[1][109] , \modmult_1/zin[1][108] , 
        \modmult_1/zin[1][107] , \modmult_1/zin[1][106] , 
        \modmult_1/zin[1][105] , \modmult_1/zin[1][104] , 
        \modmult_1/zin[1][103] , \modmult_1/zin[1][102] , 
        \modmult_1/zin[1][101] , \modmult_1/zin[1][100] , 
        \modmult_1/zin[1][99] , \modmult_1/zin[1][98] , \modmult_1/zin[1][97] , 
        \modmult_1/zin[1][96] , \modmult_1/zin[1][95] , \modmult_1/zin[1][94] , 
        \modmult_1/zin[1][93] , \modmult_1/zin[1][92] , \modmult_1/zin[1][91] , 
        \modmult_1/zin[1][90] , \modmult_1/zin[1][89] , \modmult_1/zin[1][88] , 
        \modmult_1/zin[1][87] , \modmult_1/zin[1][86] , \modmult_1/zin[1][85] , 
        \modmult_1/zin[1][84] , \modmult_1/zin[1][83] , \modmult_1/zin[1][82] , 
        \modmult_1/zin[1][81] , \modmult_1/zin[1][80] , \modmult_1/zin[1][79] , 
        \modmult_1/zin[1][78] , \modmult_1/zin[1][77] , \modmult_1/zin[1][76] , 
        \modmult_1/zin[1][75] , \modmult_1/zin[1][74] , \modmult_1/zin[1][73] , 
        \modmult_1/zin[1][72] , \modmult_1/zin[1][71] , \modmult_1/zin[1][70] , 
        \modmult_1/zin[1][69] , \modmult_1/zin[1][68] , \modmult_1/zin[1][67] , 
        \modmult_1/zin[1][66] , \modmult_1/zin[1][65] , \modmult_1/zin[1][64] , 
        \modmult_1/zin[1][63] , \modmult_1/zin[1][62] , \modmult_1/zin[1][61] , 
        \modmult_1/zin[1][60] , \modmult_1/zin[1][59] , \modmult_1/zin[1][58] , 
        \modmult_1/zin[1][57] , \modmult_1/zin[1][56] , \modmult_1/zin[1][55] , 
        \modmult_1/zin[1][54] , \modmult_1/zin[1][53] , \modmult_1/zin[1][52] , 
        \modmult_1/zin[1][51] , \modmult_1/zin[1][50] , \modmult_1/zin[1][49] , 
        \modmult_1/zin[1][48] , \modmult_1/zin[1][47] , \modmult_1/zin[1][46] , 
        \modmult_1/zin[1][45] , \modmult_1/zin[1][44] , \modmult_1/zin[1][43] , 
        \modmult_1/zin[1][42] , \modmult_1/zin[1][41] , \modmult_1/zin[1][40] , 
        \modmult_1/zin[1][39] , \modmult_1/zin[1][38] , \modmult_1/zin[1][37] , 
        \modmult_1/zin[1][36] , \modmult_1/zin[1][35] , \modmult_1/zin[1][34] , 
        \modmult_1/zin[1][33] , \modmult_1/zin[1][32] , \modmult_1/zin[1][31] , 
        \modmult_1/zin[1][30] , \modmult_1/zin[1][29] , \modmult_1/zin[1][28] , 
        \modmult_1/zin[1][27] , \modmult_1/zin[1][26] , \modmult_1/zin[1][25] , 
        \modmult_1/zin[1][24] , \modmult_1/zin[1][23] , \modmult_1/zin[1][22] , 
        \modmult_1/zin[1][21] , \modmult_1/zin[1][20] , \modmult_1/zin[1][19] , 
        \modmult_1/zin[1][18] , \modmult_1/zin[1][17] , \modmult_1/zin[1][16] , 
        \modmult_1/zin[1][15] , \modmult_1/zin[1][14] , \modmult_1/zin[1][13] , 
        \modmult_1/zin[1][12] , \modmult_1/zin[1][11] , \modmult_1/zin[1][10] , 
        \modmult_1/zin[1][9] , \modmult_1/zin[1][8] , \modmult_1/zin[1][7] , 
        \modmult_1/zin[1][6] , \modmult_1/zin[1][5] , \modmult_1/zin[1][4] , 
        \modmult_1/zin[1][3] , \modmult_1/zin[1][2] , \modmult_1/zin[1][1] , 
        \modmult_1/zin[1][0] }) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .Q(
        start_reg[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .Q(
        start_reg[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .Q(
        start_reg[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .Q(
        start_reg[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .Q(
        start_reg[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .Q(
        start_reg[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .Q(
        start_reg[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .Q(
        start_reg[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .Q(
        start_reg[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .Q(
        start_reg[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .Q(
        start_reg[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .Q(
        start_reg[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .Q(
        start_reg[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .Q(
        start_reg[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .Q(
        start_reg[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .Q(
        start_reg[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .Q(
        start_reg[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .Q(
        start_reg[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .Q(
        start_reg[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .Q(
        start_reg[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .Q(
        start_reg[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .Q(
        start_reg[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .Q(
        start_reg[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .Q(
        start_reg[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .Q(
        start_reg[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .Q(
        start_reg[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .Q(
        start_reg[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .Q(
        start_reg[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .Q(
        start_reg[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .Q(
        start_reg[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .Q(
        start_reg[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .Q(
        start_reg[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .Q(
        start_reg[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .Q(
        start_reg[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .Q(
        start_reg[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .Q(
        start_reg[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .Q(
        start_reg[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .Q(
        start_reg[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .Q(
        start_reg[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .Q(
        start_reg[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .Q(
        start_reg[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .Q(
        start_reg[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .Q(
        start_reg[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .Q(
        start_reg[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .Q(
        start_reg[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .Q(
        start_reg[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .Q(
        start_reg[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .Q(
        start_reg[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .Q(
        start_reg[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .Q(
        start_reg[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .Q(
        start_reg[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .Q(
        start_reg[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .Q(
        start_reg[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .Q(
        start_reg[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .Q(
        start_reg[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .Q(
        start_reg[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .Q(
        start_reg[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .Q(
        start_reg[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .Q(
        start_reg[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .Q(
        start_reg[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .Q(
        start_reg[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .Q(
        start_reg[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .Q(
        start_reg[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .Q(
        start_reg[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .Q(
        start_reg[127]) );
  DFF \modmult_1/zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[0] ) );
  DFF \modmult_1/xreg_reg[2]  ( .D(\modmult_1/xin[0] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[2] ) );
  DFF \modmult_1/zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[1] ) );
  DFF \modmult_1/xreg_reg[3]  ( .D(\modmult_1/xin[1] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[3] ) );
  DFF \modmult_1/zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[2] ) );
  DFF \modmult_1/xreg_reg[4]  ( .D(\modmult_1/xin[2] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[4] ) );
  DFF \modmult_1/zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[3] ) );
  DFF \modmult_1/xreg_reg[5]  ( .D(\modmult_1/xin[3] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[5] ) );
  DFF \modmult_1/zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[4] ) );
  DFF \modmult_1/xreg_reg[6]  ( .D(\modmult_1/xin[4] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[6] ) );
  DFF \modmult_1/zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[5] ) );
  DFF \modmult_1/xreg_reg[7]  ( .D(\modmult_1/xin[5] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[7] ) );
  DFF \modmult_1/zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[6] ) );
  DFF \modmult_1/xreg_reg[8]  ( .D(\modmult_1/xin[6] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[8] ) );
  DFF \modmult_1/zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[7] ) );
  DFF \modmult_1/xreg_reg[9]  ( .D(\modmult_1/xin[7] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[9] ) );
  DFF \modmult_1/zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[8] ) );
  DFF \modmult_1/xreg_reg[10]  ( .D(\modmult_1/xin[8] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[10] ) );
  DFF \modmult_1/zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[9] ) );
  DFF \modmult_1/xreg_reg[11]  ( .D(\modmult_1/xin[9] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[11] ) );
  DFF \modmult_1/zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[10] ) );
  DFF \modmult_1/xreg_reg[12]  ( .D(\modmult_1/xin[10] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[12] ) );
  DFF \modmult_1/zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[11] ) );
  DFF \modmult_1/xreg_reg[13]  ( .D(\modmult_1/xin[11] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[13] ) );
  DFF \modmult_1/zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[12] ) );
  DFF \modmult_1/xreg_reg[14]  ( .D(\modmult_1/xin[12] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[14] ) );
  DFF \modmult_1/zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[13] ) );
  DFF \modmult_1/xreg_reg[15]  ( .D(\modmult_1/xin[13] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[15] ) );
  DFF \modmult_1/zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[14] ) );
  DFF \modmult_1/xreg_reg[16]  ( .D(\modmult_1/xin[14] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[16] ) );
  DFF \modmult_1/zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[15] ) );
  DFF \modmult_1/xreg_reg[17]  ( .D(\modmult_1/xin[15] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[17] ) );
  DFF \modmult_1/zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[16] ) );
  DFF \modmult_1/xreg_reg[18]  ( .D(\modmult_1/xin[16] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[18] ) );
  DFF \modmult_1/zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[17] ) );
  DFF \modmult_1/xreg_reg[19]  ( .D(\modmult_1/xin[17] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[19] ) );
  DFF \modmult_1/zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[18] ) );
  DFF \modmult_1/xreg_reg[20]  ( .D(\modmult_1/xin[18] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[20] ) );
  DFF \modmult_1/zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[19] ) );
  DFF \modmult_1/xreg_reg[21]  ( .D(\modmult_1/xin[19] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[21] ) );
  DFF \modmult_1/zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[20] ) );
  DFF \modmult_1/xreg_reg[22]  ( .D(\modmult_1/xin[20] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[22] ) );
  DFF \modmult_1/zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[21] ) );
  DFF \modmult_1/xreg_reg[23]  ( .D(\modmult_1/xin[21] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[23] ) );
  DFF \modmult_1/zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[22] ) );
  DFF \modmult_1/xreg_reg[24]  ( .D(\modmult_1/xin[22] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[24] ) );
  DFF \modmult_1/zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[23] ) );
  DFF \modmult_1/xreg_reg[25]  ( .D(\modmult_1/xin[23] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[25] ) );
  DFF \modmult_1/zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[24] ) );
  DFF \modmult_1/xreg_reg[26]  ( .D(\modmult_1/xin[24] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[26] ) );
  DFF \modmult_1/zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[25] ) );
  DFF \modmult_1/xreg_reg[27]  ( .D(\modmult_1/xin[25] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[27] ) );
  DFF \modmult_1/zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[26] ) );
  DFF \modmult_1/xreg_reg[28]  ( .D(\modmult_1/xin[26] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[28] ) );
  DFF \modmult_1/zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[27] ) );
  DFF \modmult_1/xreg_reg[29]  ( .D(\modmult_1/xin[27] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[29] ) );
  DFF \modmult_1/zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[28] ) );
  DFF \modmult_1/xreg_reg[30]  ( .D(\modmult_1/xin[28] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[30] ) );
  DFF \modmult_1/zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[29] ) );
  DFF \modmult_1/xreg_reg[31]  ( .D(\modmult_1/xin[29] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[31] ) );
  DFF \modmult_1/zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[30] ) );
  DFF \modmult_1/xreg_reg[32]  ( .D(\modmult_1/xin[30] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[32] ) );
  DFF \modmult_1/zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[31] ) );
  DFF \modmult_1/xreg_reg[33]  ( .D(\modmult_1/xin[31] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[33] ) );
  DFF \modmult_1/zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[32] ) );
  DFF \modmult_1/xreg_reg[34]  ( .D(\modmult_1/xin[32] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[34] ) );
  DFF \modmult_1/zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[33] ) );
  DFF \modmult_1/xreg_reg[35]  ( .D(\modmult_1/xin[33] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[35] ) );
  DFF \modmult_1/zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[34] ) );
  DFF \modmult_1/xreg_reg[36]  ( .D(\modmult_1/xin[34] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[36] ) );
  DFF \modmult_1/zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[35] ) );
  DFF \modmult_1/xreg_reg[37]  ( .D(\modmult_1/xin[35] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[37] ) );
  DFF \modmult_1/zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[36] ) );
  DFF \modmult_1/xreg_reg[38]  ( .D(\modmult_1/xin[36] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[38] ) );
  DFF \modmult_1/zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[37] ) );
  DFF \modmult_1/xreg_reg[39]  ( .D(\modmult_1/xin[37] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[39] ) );
  DFF \modmult_1/zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[38] ) );
  DFF \modmult_1/xreg_reg[40]  ( .D(\modmult_1/xin[38] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[40] ) );
  DFF \modmult_1/zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[39] ) );
  DFF \modmult_1/xreg_reg[41]  ( .D(\modmult_1/xin[39] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[41] ) );
  DFF \modmult_1/zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[40] ) );
  DFF \modmult_1/xreg_reg[42]  ( .D(\modmult_1/xin[40] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[42] ) );
  DFF \modmult_1/zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[41] ) );
  DFF \modmult_1/xreg_reg[43]  ( .D(\modmult_1/xin[41] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[43] ) );
  DFF \modmult_1/zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[42] ) );
  DFF \modmult_1/xreg_reg[44]  ( .D(\modmult_1/xin[42] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[44] ) );
  DFF \modmult_1/zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[43] ) );
  DFF \modmult_1/xreg_reg[45]  ( .D(\modmult_1/xin[43] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[45] ) );
  DFF \modmult_1/zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[44] ) );
  DFF \modmult_1/xreg_reg[46]  ( .D(\modmult_1/xin[44] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[46] ) );
  DFF \modmult_1/zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[45] ) );
  DFF \modmult_1/xreg_reg[47]  ( .D(\modmult_1/xin[45] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[47] ) );
  DFF \modmult_1/zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[46] ) );
  DFF \modmult_1/xreg_reg[48]  ( .D(\modmult_1/xin[46] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[48] ) );
  DFF \modmult_1/zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[47] ) );
  DFF \modmult_1/xreg_reg[49]  ( .D(\modmult_1/xin[47] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[49] ) );
  DFF \modmult_1/zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[48] ) );
  DFF \modmult_1/xreg_reg[50]  ( .D(\modmult_1/xin[48] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[50] ) );
  DFF \modmult_1/zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[49] ) );
  DFF \modmult_1/xreg_reg[51]  ( .D(\modmult_1/xin[49] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[51] ) );
  DFF \modmult_1/zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[50] ) );
  DFF \modmult_1/xreg_reg[52]  ( .D(\modmult_1/xin[50] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[52] ) );
  DFF \modmult_1/zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[51] ) );
  DFF \modmult_1/xreg_reg[53]  ( .D(\modmult_1/xin[51] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[53] ) );
  DFF \modmult_1/zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[52] ) );
  DFF \modmult_1/xreg_reg[54]  ( .D(\modmult_1/xin[52] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[54] ) );
  DFF \modmult_1/zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[53] ) );
  DFF \modmult_1/xreg_reg[55]  ( .D(\modmult_1/xin[53] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[55] ) );
  DFF \modmult_1/zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[54] ) );
  DFF \modmult_1/xreg_reg[56]  ( .D(\modmult_1/xin[54] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[56] ) );
  DFF \modmult_1/zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[55] ) );
  DFF \modmult_1/xreg_reg[57]  ( .D(\modmult_1/xin[55] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[57] ) );
  DFF \modmult_1/zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[56] ) );
  DFF \modmult_1/xreg_reg[58]  ( .D(\modmult_1/xin[56] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[58] ) );
  DFF \modmult_1/zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[57] ) );
  DFF \modmult_1/xreg_reg[59]  ( .D(\modmult_1/xin[57] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[59] ) );
  DFF \modmult_1/zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[58] ) );
  DFF \modmult_1/xreg_reg[60]  ( .D(\modmult_1/xin[58] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[60] ) );
  DFF \modmult_1/zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[59] ) );
  DFF \modmult_1/xreg_reg[61]  ( .D(\modmult_1/xin[59] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[61] ) );
  DFF \modmult_1/zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[60] ) );
  DFF \modmult_1/xreg_reg[62]  ( .D(\modmult_1/xin[60] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[62] ) );
  DFF \modmult_1/zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[61] ) );
  DFF \modmult_1/xreg_reg[63]  ( .D(\modmult_1/xin[61] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[63] ) );
  DFF \modmult_1/zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[62] ) );
  DFF \modmult_1/xreg_reg[64]  ( .D(\modmult_1/xin[62] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[64] ) );
  DFF \modmult_1/zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[63] ) );
  DFF \modmult_1/xreg_reg[65]  ( .D(\modmult_1/xin[63] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[65] ) );
  DFF \modmult_1/zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[64] ) );
  DFF \modmult_1/xreg_reg[66]  ( .D(\modmult_1/xin[64] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[66] ) );
  DFF \modmult_1/zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[65] ) );
  DFF \modmult_1/xreg_reg[67]  ( .D(\modmult_1/xin[65] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[67] ) );
  DFF \modmult_1/zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[66] ) );
  DFF \modmult_1/xreg_reg[68]  ( .D(\modmult_1/xin[66] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[68] ) );
  DFF \modmult_1/zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[67] ) );
  DFF \modmult_1/xreg_reg[69]  ( .D(\modmult_1/xin[67] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[69] ) );
  DFF \modmult_1/zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[68] ) );
  DFF \modmult_1/xreg_reg[70]  ( .D(\modmult_1/xin[68] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[70] ) );
  DFF \modmult_1/zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[69] ) );
  DFF \modmult_1/xreg_reg[71]  ( .D(\modmult_1/xin[69] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[71] ) );
  DFF \modmult_1/zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[70] ) );
  DFF \modmult_1/xreg_reg[72]  ( .D(\modmult_1/xin[70] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[72] ) );
  DFF \modmult_1/zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[71] ) );
  DFF \modmult_1/xreg_reg[73]  ( .D(\modmult_1/xin[71] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[73] ) );
  DFF \modmult_1/zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[72] ) );
  DFF \modmult_1/xreg_reg[74]  ( .D(\modmult_1/xin[72] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[74] ) );
  DFF \modmult_1/zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[73] ) );
  DFF \modmult_1/xreg_reg[75]  ( .D(\modmult_1/xin[73] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[75] ) );
  DFF \modmult_1/zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[74] ) );
  DFF \modmult_1/xreg_reg[76]  ( .D(\modmult_1/xin[74] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[76] ) );
  DFF \modmult_1/zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[75] ) );
  DFF \modmult_1/xreg_reg[77]  ( .D(\modmult_1/xin[75] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[77] ) );
  DFF \modmult_1/zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[76] ) );
  DFF \modmult_1/xreg_reg[78]  ( .D(\modmult_1/xin[76] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[78] ) );
  DFF \modmult_1/zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[77] ) );
  DFF \modmult_1/xreg_reg[79]  ( .D(\modmult_1/xin[77] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[79] ) );
  DFF \modmult_1/zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[78] ) );
  DFF \modmult_1/xreg_reg[80]  ( .D(\modmult_1/xin[78] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[80] ) );
  DFF \modmult_1/zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[79] ) );
  DFF \modmult_1/xreg_reg[81]  ( .D(\modmult_1/xin[79] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[81] ) );
  DFF \modmult_1/zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[80] ) );
  DFF \modmult_1/xreg_reg[82]  ( .D(\modmult_1/xin[80] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[82] ) );
  DFF \modmult_1/zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[81] ) );
  DFF \modmult_1/xreg_reg[83]  ( .D(\modmult_1/xin[81] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[83] ) );
  DFF \modmult_1/zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[82] ) );
  DFF \modmult_1/xreg_reg[84]  ( .D(\modmult_1/xin[82] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[84] ) );
  DFF \modmult_1/zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[83] ) );
  DFF \modmult_1/xreg_reg[85]  ( .D(\modmult_1/xin[83] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[85] ) );
  DFF \modmult_1/zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[84] ) );
  DFF \modmult_1/xreg_reg[86]  ( .D(\modmult_1/xin[84] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[86] ) );
  DFF \modmult_1/zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[85] ) );
  DFF \modmult_1/xreg_reg[87]  ( .D(\modmult_1/xin[85] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[87] ) );
  DFF \modmult_1/zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[86] ) );
  DFF \modmult_1/xreg_reg[88]  ( .D(\modmult_1/xin[86] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[88] ) );
  DFF \modmult_1/zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[87] ) );
  DFF \modmult_1/xreg_reg[89]  ( .D(\modmult_1/xin[87] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[89] ) );
  DFF \modmult_1/zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[88] ) );
  DFF \modmult_1/xreg_reg[90]  ( .D(\modmult_1/xin[88] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[90] ) );
  DFF \modmult_1/zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[89] ) );
  DFF \modmult_1/xreg_reg[91]  ( .D(\modmult_1/xin[89] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[91] ) );
  DFF \modmult_1/zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[90] ) );
  DFF \modmult_1/xreg_reg[92]  ( .D(\modmult_1/xin[90] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[92] ) );
  DFF \modmult_1/zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[91] ) );
  DFF \modmult_1/xreg_reg[93]  ( .D(\modmult_1/xin[91] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[93] ) );
  DFF \modmult_1/zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[92] ) );
  DFF \modmult_1/xreg_reg[94]  ( .D(\modmult_1/xin[92] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[94] ) );
  DFF \modmult_1/zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[93] ) );
  DFF \modmult_1/xreg_reg[95]  ( .D(\modmult_1/xin[93] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[95] ) );
  DFF \modmult_1/zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[94] ) );
  DFF \modmult_1/xreg_reg[96]  ( .D(\modmult_1/xin[94] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[96] ) );
  DFF \modmult_1/zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[95] ) );
  DFF \modmult_1/xreg_reg[97]  ( .D(\modmult_1/xin[95] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[97] ) );
  DFF \modmult_1/zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[96] ) );
  DFF \modmult_1/xreg_reg[98]  ( .D(\modmult_1/xin[96] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[98] ) );
  DFF \modmult_1/zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[97] ) );
  DFF \modmult_1/xreg_reg[99]  ( .D(\modmult_1/xin[97] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[99] ) );
  DFF \modmult_1/zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[98] ) );
  DFF \modmult_1/xreg_reg[100]  ( .D(\modmult_1/xin[98] ), .CLK(clk), .RST(rst), .Q(\modmult_1/xreg[100] ) );
  DFF \modmult_1/zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[99] ) );
  DFF \modmult_1/xreg_reg[101]  ( .D(\modmult_1/xin[99] ), .CLK(clk), .RST(rst), .Q(\modmult_1/xreg[101] ) );
  DFF \modmult_1/zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[100] ) );
  DFF \modmult_1/xreg_reg[102]  ( .D(\modmult_1/xin[100] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[102] ) );
  DFF \modmult_1/zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[101] ) );
  DFF \modmult_1/xreg_reg[103]  ( .D(\modmult_1/xin[101] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[103] ) );
  DFF \modmult_1/zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[102] ) );
  DFF \modmult_1/xreg_reg[104]  ( .D(\modmult_1/xin[102] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[104] ) );
  DFF \modmult_1/zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[103] ) );
  DFF \modmult_1/xreg_reg[105]  ( .D(\modmult_1/xin[103] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[105] ) );
  DFF \modmult_1/zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[104] ) );
  DFF \modmult_1/xreg_reg[106]  ( .D(\modmult_1/xin[104] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[106] ) );
  DFF \modmult_1/zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[105] ) );
  DFF \modmult_1/xreg_reg[107]  ( .D(\modmult_1/xin[105] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[107] ) );
  DFF \modmult_1/zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[106] ) );
  DFF \modmult_1/xreg_reg[108]  ( .D(\modmult_1/xin[106] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[108] ) );
  DFF \modmult_1/zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[107] ) );
  DFF \modmult_1/xreg_reg[109]  ( .D(\modmult_1/xin[107] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[109] ) );
  DFF \modmult_1/zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[108] ) );
  DFF \modmult_1/xreg_reg[110]  ( .D(\modmult_1/xin[108] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[110] ) );
  DFF \modmult_1/zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[109] ) );
  DFF \modmult_1/xreg_reg[111]  ( .D(\modmult_1/xin[109] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[111] ) );
  DFF \modmult_1/zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[110] ) );
  DFF \modmult_1/xreg_reg[112]  ( .D(\modmult_1/xin[110] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[112] ) );
  DFF \modmult_1/zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[111] ) );
  DFF \modmult_1/xreg_reg[113]  ( .D(\modmult_1/xin[111] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[113] ) );
  DFF \modmult_1/zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[112] ) );
  DFF \modmult_1/xreg_reg[114]  ( .D(\modmult_1/xin[112] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[114] ) );
  DFF \modmult_1/zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[113] ) );
  DFF \modmult_1/xreg_reg[115]  ( .D(\modmult_1/xin[113] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[115] ) );
  DFF \modmult_1/zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[114] ) );
  DFF \modmult_1/xreg_reg[116]  ( .D(\modmult_1/xin[114] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[116] ) );
  DFF \modmult_1/zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[115] ) );
  DFF \modmult_1/xreg_reg[117]  ( .D(\modmult_1/xin[115] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[117] ) );
  DFF \modmult_1/zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[116] ) );
  DFF \modmult_1/xreg_reg[118]  ( .D(\modmult_1/xin[116] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[118] ) );
  DFF \modmult_1/zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[117] ) );
  DFF \modmult_1/xreg_reg[119]  ( .D(\modmult_1/xin[117] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[119] ) );
  DFF \modmult_1/zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[118] ) );
  DFF \modmult_1/xreg_reg[120]  ( .D(\modmult_1/xin[118] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[120] ) );
  DFF \modmult_1/zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[119] ) );
  DFF \modmult_1/xreg_reg[121]  ( .D(\modmult_1/xin[119] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[121] ) );
  DFF \modmult_1/zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[120] ) );
  DFF \modmult_1/xreg_reg[122]  ( .D(\modmult_1/xin[120] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[122] ) );
  DFF \modmult_1/zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[121] ) );
  DFF \modmult_1/xreg_reg[123]  ( .D(\modmult_1/xin[121] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[123] ) );
  DFF \modmult_1/zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[122] ) );
  DFF \modmult_1/xreg_reg[124]  ( .D(\modmult_1/xin[122] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[124] ) );
  DFF \modmult_1/zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[123] ) );
  DFF \modmult_1/xreg_reg[125]  ( .D(\modmult_1/xin[123] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[125] ) );
  DFF \modmult_1/zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[124] ) );
  DFF \modmult_1/xreg_reg[126]  ( .D(\modmult_1/xin[124] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[126] ) );
  DFF \modmult_1/zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[125] ) );
  DFF \modmult_1/xreg_reg[127]  ( .D(\modmult_1/xin[125] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[127] ) );
  DFF \modmult_1/zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[126] ) );
  DFF \modmult_1/xreg_reg[128]  ( .D(\modmult_1/xin[126] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[128] ) );
  DFF \modmult_1/zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[127] ) );
  DFF \modmult_1/xreg_reg[129]  ( .D(\modmult_1/xin[127] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[129] ) );
  DFF \modmult_1/zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[128] ) );
  DFF \modmult_1/xreg_reg[130]  ( .D(\modmult_1/xin[128] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[130] ) );
  DFF \modmult_1/zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[129] ) );
  DFF \modmult_1/xreg_reg[131]  ( .D(\modmult_1/xin[129] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[131] ) );
  DFF \modmult_1/zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[130] ) );
  DFF \modmult_1/xreg_reg[132]  ( .D(\modmult_1/xin[130] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[132] ) );
  DFF \modmult_1/zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[131] ) );
  DFF \modmult_1/xreg_reg[133]  ( .D(\modmult_1/xin[131] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[133] ) );
  DFF \modmult_1/zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[132] ) );
  DFF \modmult_1/xreg_reg[134]  ( .D(\modmult_1/xin[132] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[134] ) );
  DFF \modmult_1/zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[133] ) );
  DFF \modmult_1/xreg_reg[135]  ( .D(\modmult_1/xin[133] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[135] ) );
  DFF \modmult_1/zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[134] ) );
  DFF \modmult_1/xreg_reg[136]  ( .D(\modmult_1/xin[134] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[136] ) );
  DFF \modmult_1/zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[135] ) );
  DFF \modmult_1/xreg_reg[137]  ( .D(\modmult_1/xin[135] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[137] ) );
  DFF \modmult_1/zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[136] ) );
  DFF \modmult_1/xreg_reg[138]  ( .D(\modmult_1/xin[136] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[138] ) );
  DFF \modmult_1/zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[137] ) );
  DFF \modmult_1/xreg_reg[139]  ( .D(\modmult_1/xin[137] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[139] ) );
  DFF \modmult_1/zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[138] ) );
  DFF \modmult_1/xreg_reg[140]  ( .D(\modmult_1/xin[138] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[140] ) );
  DFF \modmult_1/zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[139] ) );
  DFF \modmult_1/xreg_reg[141]  ( .D(\modmult_1/xin[139] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[141] ) );
  DFF \modmult_1/zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[140] ) );
  DFF \modmult_1/xreg_reg[142]  ( .D(\modmult_1/xin[140] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[142] ) );
  DFF \modmult_1/zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[141] ) );
  DFF \modmult_1/xreg_reg[143]  ( .D(\modmult_1/xin[141] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[143] ) );
  DFF \modmult_1/zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[142] ) );
  DFF \modmult_1/xreg_reg[144]  ( .D(\modmult_1/xin[142] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[144] ) );
  DFF \modmult_1/zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[143] ) );
  DFF \modmult_1/xreg_reg[145]  ( .D(\modmult_1/xin[143] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[145] ) );
  DFF \modmult_1/zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[144] ) );
  DFF \modmult_1/xreg_reg[146]  ( .D(\modmult_1/xin[144] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[146] ) );
  DFF \modmult_1/zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[145] ) );
  DFF \modmult_1/xreg_reg[147]  ( .D(\modmult_1/xin[145] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[147] ) );
  DFF \modmult_1/zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[146] ) );
  DFF \modmult_1/xreg_reg[148]  ( .D(\modmult_1/xin[146] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[148] ) );
  DFF \modmult_1/zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[147] ) );
  DFF \modmult_1/xreg_reg[149]  ( .D(\modmult_1/xin[147] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[149] ) );
  DFF \modmult_1/zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[148] ) );
  DFF \modmult_1/xreg_reg[150]  ( .D(\modmult_1/xin[148] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[150] ) );
  DFF \modmult_1/zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[149] ) );
  DFF \modmult_1/xreg_reg[151]  ( .D(\modmult_1/xin[149] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[151] ) );
  DFF \modmult_1/zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[150] ) );
  DFF \modmult_1/xreg_reg[152]  ( .D(\modmult_1/xin[150] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[152] ) );
  DFF \modmult_1/zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[151] ) );
  DFF \modmult_1/xreg_reg[153]  ( .D(\modmult_1/xin[151] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[153] ) );
  DFF \modmult_1/zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[152] ) );
  DFF \modmult_1/xreg_reg[154]  ( .D(\modmult_1/xin[152] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[154] ) );
  DFF \modmult_1/zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[153] ) );
  DFF \modmult_1/xreg_reg[155]  ( .D(\modmult_1/xin[153] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[155] ) );
  DFF \modmult_1/zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[154] ) );
  DFF \modmult_1/xreg_reg[156]  ( .D(\modmult_1/xin[154] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[156] ) );
  DFF \modmult_1/zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[155] ) );
  DFF \modmult_1/xreg_reg[157]  ( .D(\modmult_1/xin[155] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[157] ) );
  DFF \modmult_1/zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[156] ) );
  DFF \modmult_1/xreg_reg[158]  ( .D(\modmult_1/xin[156] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[158] ) );
  DFF \modmult_1/zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[157] ) );
  DFF \modmult_1/xreg_reg[159]  ( .D(\modmult_1/xin[157] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[159] ) );
  DFF \modmult_1/zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[158] ) );
  DFF \modmult_1/xreg_reg[160]  ( .D(\modmult_1/xin[158] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[160] ) );
  DFF \modmult_1/zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[159] ) );
  DFF \modmult_1/xreg_reg[161]  ( .D(\modmult_1/xin[159] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[161] ) );
  DFF \modmult_1/zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[160] ) );
  DFF \modmult_1/xreg_reg[162]  ( .D(\modmult_1/xin[160] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[162] ) );
  DFF \modmult_1/zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[161] ) );
  DFF \modmult_1/xreg_reg[163]  ( .D(\modmult_1/xin[161] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[163] ) );
  DFF \modmult_1/zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[162] ) );
  DFF \modmult_1/xreg_reg[164]  ( .D(\modmult_1/xin[162] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[164] ) );
  DFF \modmult_1/zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[163] ) );
  DFF \modmult_1/xreg_reg[165]  ( .D(\modmult_1/xin[163] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[165] ) );
  DFF \modmult_1/zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[164] ) );
  DFF \modmult_1/xreg_reg[166]  ( .D(\modmult_1/xin[164] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[166] ) );
  DFF \modmult_1/zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[165] ) );
  DFF \modmult_1/xreg_reg[167]  ( .D(\modmult_1/xin[165] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[167] ) );
  DFF \modmult_1/zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[166] ) );
  DFF \modmult_1/xreg_reg[168]  ( .D(\modmult_1/xin[166] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[168] ) );
  DFF \modmult_1/zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[167] ) );
  DFF \modmult_1/xreg_reg[169]  ( .D(\modmult_1/xin[167] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[169] ) );
  DFF \modmult_1/zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[168] ) );
  DFF \modmult_1/xreg_reg[170]  ( .D(\modmult_1/xin[168] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[170] ) );
  DFF \modmult_1/zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[169] ) );
  DFF \modmult_1/xreg_reg[171]  ( .D(\modmult_1/xin[169] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[171] ) );
  DFF \modmult_1/zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[170] ) );
  DFF \modmult_1/xreg_reg[172]  ( .D(\modmult_1/xin[170] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[172] ) );
  DFF \modmult_1/zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[171] ) );
  DFF \modmult_1/xreg_reg[173]  ( .D(\modmult_1/xin[171] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[173] ) );
  DFF \modmult_1/zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[172] ) );
  DFF \modmult_1/xreg_reg[174]  ( .D(\modmult_1/xin[172] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[174] ) );
  DFF \modmult_1/zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[173] ) );
  DFF \modmult_1/xreg_reg[175]  ( .D(\modmult_1/xin[173] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[175] ) );
  DFF \modmult_1/zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[174] ) );
  DFF \modmult_1/xreg_reg[176]  ( .D(\modmult_1/xin[174] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[176] ) );
  DFF \modmult_1/zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[175] ) );
  DFF \modmult_1/xreg_reg[177]  ( .D(\modmult_1/xin[175] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[177] ) );
  DFF \modmult_1/zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[176] ) );
  DFF \modmult_1/xreg_reg[178]  ( .D(\modmult_1/xin[176] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[178] ) );
  DFF \modmult_1/zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[177] ) );
  DFF \modmult_1/xreg_reg[179]  ( .D(\modmult_1/xin[177] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[179] ) );
  DFF \modmult_1/zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[178] ) );
  DFF \modmult_1/xreg_reg[180]  ( .D(\modmult_1/xin[178] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[180] ) );
  DFF \modmult_1/zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[179] ) );
  DFF \modmult_1/xreg_reg[181]  ( .D(\modmult_1/xin[179] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[181] ) );
  DFF \modmult_1/zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[180] ) );
  DFF \modmult_1/xreg_reg[182]  ( .D(\modmult_1/xin[180] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[182] ) );
  DFF \modmult_1/zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[181] ) );
  DFF \modmult_1/xreg_reg[183]  ( .D(\modmult_1/xin[181] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[183] ) );
  DFF \modmult_1/zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[182] ) );
  DFF \modmult_1/xreg_reg[184]  ( .D(\modmult_1/xin[182] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[184] ) );
  DFF \modmult_1/zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[183] ) );
  DFF \modmult_1/xreg_reg[185]  ( .D(\modmult_1/xin[183] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[185] ) );
  DFF \modmult_1/zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[184] ) );
  DFF \modmult_1/xreg_reg[186]  ( .D(\modmult_1/xin[184] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[186] ) );
  DFF \modmult_1/zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[185] ) );
  DFF \modmult_1/xreg_reg[187]  ( .D(\modmult_1/xin[185] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[187] ) );
  DFF \modmult_1/zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[186] ) );
  DFF \modmult_1/xreg_reg[188]  ( .D(\modmult_1/xin[186] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[188] ) );
  DFF \modmult_1/zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[187] ) );
  DFF \modmult_1/xreg_reg[189]  ( .D(\modmult_1/xin[187] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[189] ) );
  DFF \modmult_1/zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[188] ) );
  DFF \modmult_1/xreg_reg[190]  ( .D(\modmult_1/xin[188] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[190] ) );
  DFF \modmult_1/zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[189] ) );
  DFF \modmult_1/xreg_reg[191]  ( .D(\modmult_1/xin[189] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[191] ) );
  DFF \modmult_1/zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[190] ) );
  DFF \modmult_1/xreg_reg[192]  ( .D(\modmult_1/xin[190] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[192] ) );
  DFF \modmult_1/zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[191] ) );
  DFF \modmult_1/xreg_reg[193]  ( .D(\modmult_1/xin[191] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[193] ) );
  DFF \modmult_1/zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[192] ) );
  DFF \modmult_1/xreg_reg[194]  ( .D(\modmult_1/xin[192] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[194] ) );
  DFF \modmult_1/zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[193] ) );
  DFF \modmult_1/xreg_reg[195]  ( .D(\modmult_1/xin[193] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[195] ) );
  DFF \modmult_1/zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[194] ) );
  DFF \modmult_1/xreg_reg[196]  ( .D(\modmult_1/xin[194] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[196] ) );
  DFF \modmult_1/zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[195] ) );
  DFF \modmult_1/xreg_reg[197]  ( .D(\modmult_1/xin[195] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[197] ) );
  DFF \modmult_1/zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[196] ) );
  DFF \modmult_1/xreg_reg[198]  ( .D(\modmult_1/xin[196] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[198] ) );
  DFF \modmult_1/zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[197] ) );
  DFF \modmult_1/xreg_reg[199]  ( .D(\modmult_1/xin[197] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[199] ) );
  DFF \modmult_1/zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[198] ) );
  DFF \modmult_1/xreg_reg[200]  ( .D(\modmult_1/xin[198] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[200] ) );
  DFF \modmult_1/zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[199] ) );
  DFF \modmult_1/xreg_reg[201]  ( .D(\modmult_1/xin[199] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[201] ) );
  DFF \modmult_1/zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[200] ) );
  DFF \modmult_1/xreg_reg[202]  ( .D(\modmult_1/xin[200] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[202] ) );
  DFF \modmult_1/zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[201] ) );
  DFF \modmult_1/xreg_reg[203]  ( .D(\modmult_1/xin[201] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[203] ) );
  DFF \modmult_1/zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[202] ) );
  DFF \modmult_1/xreg_reg[204]  ( .D(\modmult_1/xin[202] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[204] ) );
  DFF \modmult_1/zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[203] ) );
  DFF \modmult_1/xreg_reg[205]  ( .D(\modmult_1/xin[203] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[205] ) );
  DFF \modmult_1/zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[204] ) );
  DFF \modmult_1/xreg_reg[206]  ( .D(\modmult_1/xin[204] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[206] ) );
  DFF \modmult_1/zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[205] ) );
  DFF \modmult_1/xreg_reg[207]  ( .D(\modmult_1/xin[205] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[207] ) );
  DFF \modmult_1/zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[206] ) );
  DFF \modmult_1/xreg_reg[208]  ( .D(\modmult_1/xin[206] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[208] ) );
  DFF \modmult_1/zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[207] ) );
  DFF \modmult_1/xreg_reg[209]  ( .D(\modmult_1/xin[207] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[209] ) );
  DFF \modmult_1/zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[208] ) );
  DFF \modmult_1/xreg_reg[210]  ( .D(\modmult_1/xin[208] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[210] ) );
  DFF \modmult_1/zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[209] ) );
  DFF \modmult_1/xreg_reg[211]  ( .D(\modmult_1/xin[209] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[211] ) );
  DFF \modmult_1/zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[210] ) );
  DFF \modmult_1/xreg_reg[212]  ( .D(\modmult_1/xin[210] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[212] ) );
  DFF \modmult_1/zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[211] ) );
  DFF \modmult_1/xreg_reg[213]  ( .D(\modmult_1/xin[211] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[213] ) );
  DFF \modmult_1/zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[212] ) );
  DFF \modmult_1/xreg_reg[214]  ( .D(\modmult_1/xin[212] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[214] ) );
  DFF \modmult_1/zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[213] ) );
  DFF \modmult_1/xreg_reg[215]  ( .D(\modmult_1/xin[213] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[215] ) );
  DFF \modmult_1/zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[214] ) );
  DFF \modmult_1/xreg_reg[216]  ( .D(\modmult_1/xin[214] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[216] ) );
  DFF \modmult_1/zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[215] ) );
  DFF \modmult_1/xreg_reg[217]  ( .D(\modmult_1/xin[215] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[217] ) );
  DFF \modmult_1/zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[216] ) );
  DFF \modmult_1/xreg_reg[218]  ( .D(\modmult_1/xin[216] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[218] ) );
  DFF \modmult_1/zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[217] ) );
  DFF \modmult_1/xreg_reg[219]  ( .D(\modmult_1/xin[217] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[219] ) );
  DFF \modmult_1/zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[218] ) );
  DFF \modmult_1/xreg_reg[220]  ( .D(\modmult_1/xin[218] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[220] ) );
  DFF \modmult_1/zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[219] ) );
  DFF \modmult_1/xreg_reg[221]  ( .D(\modmult_1/xin[219] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[221] ) );
  DFF \modmult_1/zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[220] ) );
  DFF \modmult_1/xreg_reg[222]  ( .D(\modmult_1/xin[220] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[222] ) );
  DFF \modmult_1/zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[221] ) );
  DFF \modmult_1/xreg_reg[223]  ( .D(\modmult_1/xin[221] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[223] ) );
  DFF \modmult_1/zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[222] ) );
  DFF \modmult_1/xreg_reg[224]  ( .D(\modmult_1/xin[222] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[224] ) );
  DFF \modmult_1/zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[223] ) );
  DFF \modmult_1/xreg_reg[225]  ( .D(\modmult_1/xin[223] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[225] ) );
  DFF \modmult_1/zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[224] ) );
  DFF \modmult_1/xreg_reg[226]  ( .D(\modmult_1/xin[224] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[226] ) );
  DFF \modmult_1/zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[225] ) );
  DFF \modmult_1/xreg_reg[227]  ( .D(\modmult_1/xin[225] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[227] ) );
  DFF \modmult_1/zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[226] ) );
  DFF \modmult_1/xreg_reg[228]  ( .D(\modmult_1/xin[226] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[228] ) );
  DFF \modmult_1/zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[227] ) );
  DFF \modmult_1/xreg_reg[229]  ( .D(\modmult_1/xin[227] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[229] ) );
  DFF \modmult_1/zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[228] ) );
  DFF \modmult_1/xreg_reg[230]  ( .D(\modmult_1/xin[228] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[230] ) );
  DFF \modmult_1/zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[229] ) );
  DFF \modmult_1/xreg_reg[231]  ( .D(\modmult_1/xin[229] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[231] ) );
  DFF \modmult_1/zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[230] ) );
  DFF \modmult_1/xreg_reg[232]  ( .D(\modmult_1/xin[230] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[232] ) );
  DFF \modmult_1/zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[231] ) );
  DFF \modmult_1/xreg_reg[233]  ( .D(\modmult_1/xin[231] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[233] ) );
  DFF \modmult_1/zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[232] ) );
  DFF \modmult_1/xreg_reg[234]  ( .D(\modmult_1/xin[232] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[234] ) );
  DFF \modmult_1/zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[233] ) );
  DFF \modmult_1/xreg_reg[235]  ( .D(\modmult_1/xin[233] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[235] ) );
  DFF \modmult_1/zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[234] ) );
  DFF \modmult_1/xreg_reg[236]  ( .D(\modmult_1/xin[234] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[236] ) );
  DFF \modmult_1/zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[235] ) );
  DFF \modmult_1/xreg_reg[237]  ( .D(\modmult_1/xin[235] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[237] ) );
  DFF \modmult_1/zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[236] ) );
  DFF \modmult_1/xreg_reg[238]  ( .D(\modmult_1/xin[236] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[238] ) );
  DFF \modmult_1/zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[237] ) );
  DFF \modmult_1/xreg_reg[239]  ( .D(\modmult_1/xin[237] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[239] ) );
  DFF \modmult_1/zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[238] ) );
  DFF \modmult_1/xreg_reg[240]  ( .D(\modmult_1/xin[238] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[240] ) );
  DFF \modmult_1/zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[239] ) );
  DFF \modmult_1/xreg_reg[241]  ( .D(\modmult_1/xin[239] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[241] ) );
  DFF \modmult_1/zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[240] ) );
  DFF \modmult_1/xreg_reg[242]  ( .D(\modmult_1/xin[240] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[242] ) );
  DFF \modmult_1/zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[241] ) );
  DFF \modmult_1/xreg_reg[243]  ( .D(\modmult_1/xin[241] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[243] ) );
  DFF \modmult_1/zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[242] ) );
  DFF \modmult_1/xreg_reg[244]  ( .D(\modmult_1/xin[242] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[244] ) );
  DFF \modmult_1/zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[243] ) );
  DFF \modmult_1/xreg_reg[245]  ( .D(\modmult_1/xin[243] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[245] ) );
  DFF \modmult_1/zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[244] ) );
  DFF \modmult_1/xreg_reg[246]  ( .D(\modmult_1/xin[244] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[246] ) );
  DFF \modmult_1/zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[245] ) );
  DFF \modmult_1/xreg_reg[247]  ( .D(\modmult_1/xin[245] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[247] ) );
  DFF \modmult_1/zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[246] ) );
  DFF \modmult_1/xreg_reg[248]  ( .D(\modmult_1/xin[246] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[248] ) );
  DFF \modmult_1/zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[247] ) );
  DFF \modmult_1/xreg_reg[249]  ( .D(\modmult_1/xin[247] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[249] ) );
  DFF \modmult_1/zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[248] ) );
  DFF \modmult_1/xreg_reg[250]  ( .D(\modmult_1/xin[248] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[250] ) );
  DFF \modmult_1/zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[249] ) );
  DFF \modmult_1/xreg_reg[251]  ( .D(\modmult_1/xin[249] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[251] ) );
  DFF \modmult_1/zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[250] ) );
  DFF \modmult_1/xreg_reg[252]  ( .D(\modmult_1/xin[250] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[252] ) );
  DFF \modmult_1/zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[251] ) );
  DFF \modmult_1/xreg_reg[253]  ( .D(\modmult_1/xin[251] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[253] ) );
  DFF \modmult_1/zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[252] ) );
  DFF \modmult_1/xreg_reg[254]  ( .D(\modmult_1/xin[252] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[254] ) );
  DFF \modmult_1/zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[253] ) );
  DFF \modmult_1/xreg_reg[255]  ( .D(\modmult_1/xin[253] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/xreg[255] ) );
  DFF \modmult_1/zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[254] ) );
  DFF \modmult_1/zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[255] ) );
  DFF \modmult_1/zreg_reg[256]  ( .D(\modmult_1/zout[1][256] ), .CLK(clk), 
        .RST(rst), .Q(\modmult_1/zreg[256] ) );
  DFF mul_pow_reg ( .D(n2314), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n2313), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n2312), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n2311), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n2310), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n2309), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n2308), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n2307), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n2306), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n2305), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n2304), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n2303), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n2302), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n2301), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n2300), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n2299), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n2298), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n2297), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n2296), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n2295), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n2294), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n2293), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n2292), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n2291), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n2290), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n2289), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n2288), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n2287), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n2286), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n2285), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n2284), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n2283), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n2282), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n2281), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n2280), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n2279), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n2278), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n2277), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n2276), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n2275), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n2274), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n2273), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n2272), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n2271), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n2270), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n2269), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n2268), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n2267), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n2266), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n2265), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n2264), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n2263), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n2262), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n2261), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n2260), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n2259), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n2258), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n2257), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n2256), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n2255), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n2254), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n2253), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n2252), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n2251), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n2250), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n2249), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n2248), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n2247), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n2246), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n2245), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n2244), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n2243), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n2242), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n2241), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n2240), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n2239), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n2238), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n2237), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n2236), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n2235), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n2234), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n2233), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n2232), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n2231), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n2230), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n2229), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n2228), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n2227), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n2226), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n2225), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n2224), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n2223), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n2222), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n2221), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n2220), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n2219), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n2218), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n2217), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n2216), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n2215), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n2214), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n2213), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n2212), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n2211), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n2210), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n2209), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n2208), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n2207), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n2206), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n2205), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n2204), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n2203), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n2202), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n2201), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n2200), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n2199), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n2198), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n2197), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n2196), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n2195), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n2194), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n2193), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n2192), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n2191), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n2190), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n2189), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n2188), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n2187), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n2186), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n2185), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n2184), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n2183), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n2182), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n2181), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n2180), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n2179), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n2178), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n2177), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n2176), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n2175), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n2174), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n2173), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n2172), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n2171), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n2170), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n2169), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n2168), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n2167), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n2166), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n2165), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n2164), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n2163), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n2162), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n2161), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n2160), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n2159), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n2158), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n2157), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n2156), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n2155), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n2154), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n2153), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n2152), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n2151), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n2150), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n2149), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n2148), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n2147), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n2146), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n2145), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n2144), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n2143), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n2142), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n2141), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n2140), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n2139), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n2138), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n2137), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n2136), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n2135), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n2134), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n2133), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n2132), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n2131), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n2130), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n2129), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n2128), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n2127), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n2126), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n2125), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n2124), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n2123), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n2122), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n2121), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n2120), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n2119), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n2118), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n2117), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n2116), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n2115), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n2114), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n2113), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n2112), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n2111), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n2110), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n2109), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n2108), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n2107), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n2106), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n2105), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n2104), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n2103), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n2102), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n2101), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n2100), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n2099), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n2098), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n2097), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n2096), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n2095), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n2094), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n2093), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n2092), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n2091), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n2090), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n2089), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n2088), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n2087), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n2086), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n2085), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n2084), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n2083), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n2082), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n2081), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n2080), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n2079), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n2078), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n2077), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n2076), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n2075), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n2074), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n2073), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n2072), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n2071), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n2070), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n2069), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n2068), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n2067), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n2066), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n2065), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n2064), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n2063), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n2062), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n2061), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n2060), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n2059), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n2058), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF first_one_reg ( .D(n2057), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n2056), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n2055), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n2054), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n2053), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n2052), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n2051), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n2050), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n2049), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n2048), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n2047), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n2046), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n2045), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n2044), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n2043), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n2042), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n2041), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n2040), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n2039), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n2038), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n2037), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n2036), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n2035), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n2034), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n2033), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n2032), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n2031), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n2030), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n2029), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n2028), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n2027), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n2026), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n2025), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n2024), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n2023), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n2022), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n2021), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n2020), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n2019), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n2018), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n2017), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n2016), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n2015), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n2014), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n2013), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n2012), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n2011), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n2010), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n2009), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n2008), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n2007), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n2006), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n2005), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n2004), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n2003), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n2002), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n2001), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n2000), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n1999), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n1998), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n1997), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n1996), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n1995), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n1994), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n1993), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n1992), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n1991), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n1990), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n1989), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n1988), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n1987), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n1986), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n1985), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n1984), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n1983), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n1982), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n1981), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n1980), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n1979), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n1978), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n1977), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n1976), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n1975), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n1974), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n1973), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n1972), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n1971), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n1970), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n1969), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n1968), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n1967), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n1966), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n1965), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n1964), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n1963), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n1962), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n1961), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n1960), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n1959), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n1958), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n1957), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n1956), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n1955), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n1954), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n1953), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n1952), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n1951), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n1950), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n1949), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n1948), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n1947), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n1946), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n1945), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n1944), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n1943), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n1942), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n1941), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n1940), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n1939), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n1938), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n1937), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n1936), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n1935), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n1934), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n1933), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n1932), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n1931), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n1930), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n1929), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n1928), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n1927), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n1926), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n1925), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n1924), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n1923), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n1922), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n1921), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n1920), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n1919), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n1918), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n1917), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n1916), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n1915), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n1914), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n1913), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n1912), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n1911), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n1910), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n1909), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n1908), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n1907), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n1906), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n1905), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n1904), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n1903), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n1902), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n1901), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n1900), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n1899), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n1898), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n1897), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n1896), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n1895), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n1894), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n1893), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n1892), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n1891), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n1890), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n1889), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n1888), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n1887), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n1886), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n1885), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n1884), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n1883), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n1882), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n1881), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n1880), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n1879), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n1878), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n1877), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n1876), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n1875), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n1874), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n1873), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n1872), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n1871), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n1870), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n1869), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n1868), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n1867), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n1866), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n1865), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n1864), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n1863), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n1862), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n1861), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n1860), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n1859), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n1858), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n1857), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n1856), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n1855), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n1854), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n1853), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n1852), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n1851), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n1850), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n1849), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n1848), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n1847), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n1846), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n1845), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n1844), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n1843), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n1842), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n1841), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n1840), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n1839), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n1838), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n1837), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n1836), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n1835), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n1834), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n1833), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n1832), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n1831), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n1830), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n1829), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n1828), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n1827), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n1826), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n1825), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n1824), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n1823), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n1822), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n1821), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n1820), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n1819), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n1818), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n1817), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n1816), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n1815), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n1814), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n1813), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n1812), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n1811), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n1810), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n1809), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n1808), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n1807), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n1806), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n1805), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n1804), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n1803), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n1802), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n1801), .CLK(clk), .RST(rst), .Q(creg[255]) );
  IV U5522 ( .A(n6157), .Z(n4366) );
  IV U5523 ( .A(n7188), .Z(n4367) );
  IV U5524 ( .A(init), .Z(n4368) );
  NANDN U5526 ( .A(n4368), .B(ereg[255]), .Z(n4369) );
  AND U5527 ( .A(e[255]), .B(n4368), .Z(n7193) );
  ANDN U5528 ( .B(n4369), .A(n7193), .Z(n7188) );
  NANDN U5529 ( .A(n4367), .B(creg[0]), .Z(n4371) );
  NANDN U5530 ( .A(n7188), .B(o[0]), .Z(n4370) );
  NAND U5531 ( .A(n4371), .B(n4370), .Z(c[0]) );
  NANDN U5532 ( .A(n4367), .B(creg[100]), .Z(n4373) );
  NANDN U5533 ( .A(n7188), .B(o[100]), .Z(n4372) );
  NAND U5534 ( .A(n4373), .B(n4372), .Z(c[100]) );
  NANDN U5535 ( .A(n4367), .B(creg[101]), .Z(n4375) );
  NANDN U5536 ( .A(n7188), .B(o[101]), .Z(n4374) );
  NAND U5537 ( .A(n4375), .B(n4374), .Z(c[101]) );
  NANDN U5538 ( .A(n4367), .B(creg[102]), .Z(n4377) );
  NANDN U5539 ( .A(n7188), .B(o[102]), .Z(n4376) );
  NAND U5540 ( .A(n4377), .B(n4376), .Z(c[102]) );
  NANDN U5541 ( .A(n4367), .B(creg[103]), .Z(n4379) );
  NANDN U5542 ( .A(n7188), .B(o[103]), .Z(n4378) );
  NAND U5543 ( .A(n4379), .B(n4378), .Z(c[103]) );
  NANDN U5544 ( .A(n4367), .B(creg[104]), .Z(n4381) );
  NANDN U5545 ( .A(n7188), .B(o[104]), .Z(n4380) );
  NAND U5546 ( .A(n4381), .B(n4380), .Z(c[104]) );
  NANDN U5547 ( .A(n4367), .B(creg[105]), .Z(n4383) );
  NANDN U5548 ( .A(n7188), .B(o[105]), .Z(n4382) );
  NAND U5549 ( .A(n4383), .B(n4382), .Z(c[105]) );
  NANDN U5550 ( .A(n4367), .B(creg[106]), .Z(n4385) );
  NANDN U5551 ( .A(n7188), .B(o[106]), .Z(n4384) );
  NAND U5552 ( .A(n4385), .B(n4384), .Z(c[106]) );
  NANDN U5553 ( .A(n4367), .B(creg[107]), .Z(n4387) );
  NANDN U5554 ( .A(n7188), .B(o[107]), .Z(n4386) );
  NAND U5555 ( .A(n4387), .B(n4386), .Z(c[107]) );
  NANDN U5556 ( .A(n4367), .B(creg[108]), .Z(n4389) );
  NANDN U5557 ( .A(n7188), .B(o[108]), .Z(n4388) );
  NAND U5558 ( .A(n4389), .B(n4388), .Z(c[108]) );
  NANDN U5559 ( .A(n4367), .B(creg[109]), .Z(n4391) );
  NANDN U5560 ( .A(n7188), .B(o[109]), .Z(n4390) );
  NAND U5561 ( .A(n4391), .B(n4390), .Z(c[109]) );
  NANDN U5562 ( .A(n4367), .B(creg[10]), .Z(n4393) );
  NANDN U5563 ( .A(n7188), .B(o[10]), .Z(n4392) );
  NAND U5564 ( .A(n4393), .B(n4392), .Z(c[10]) );
  NANDN U5565 ( .A(n4367), .B(creg[110]), .Z(n4395) );
  NANDN U5566 ( .A(n7188), .B(o[110]), .Z(n4394) );
  NAND U5567 ( .A(n4395), .B(n4394), .Z(c[110]) );
  NANDN U5568 ( .A(n4367), .B(creg[111]), .Z(n4397) );
  NANDN U5569 ( .A(n7188), .B(o[111]), .Z(n4396) );
  NAND U5570 ( .A(n4397), .B(n4396), .Z(c[111]) );
  NANDN U5571 ( .A(n4367), .B(creg[112]), .Z(n4399) );
  NANDN U5572 ( .A(n7188), .B(o[112]), .Z(n4398) );
  NAND U5573 ( .A(n4399), .B(n4398), .Z(c[112]) );
  NANDN U5574 ( .A(n4367), .B(creg[113]), .Z(n4401) );
  NANDN U5575 ( .A(n7188), .B(o[113]), .Z(n4400) );
  NAND U5576 ( .A(n4401), .B(n4400), .Z(c[113]) );
  NANDN U5577 ( .A(n4367), .B(creg[114]), .Z(n4403) );
  NANDN U5578 ( .A(n7188), .B(o[114]), .Z(n4402) );
  NAND U5579 ( .A(n4403), .B(n4402), .Z(c[114]) );
  NANDN U5580 ( .A(n4367), .B(creg[115]), .Z(n4405) );
  NANDN U5581 ( .A(n7188), .B(o[115]), .Z(n4404) );
  NAND U5582 ( .A(n4405), .B(n4404), .Z(c[115]) );
  NANDN U5583 ( .A(n4367), .B(creg[116]), .Z(n4407) );
  NANDN U5584 ( .A(n7188), .B(o[116]), .Z(n4406) );
  NAND U5585 ( .A(n4407), .B(n4406), .Z(c[116]) );
  NANDN U5586 ( .A(n4367), .B(creg[117]), .Z(n4409) );
  NANDN U5587 ( .A(n7188), .B(o[117]), .Z(n4408) );
  NAND U5588 ( .A(n4409), .B(n4408), .Z(c[117]) );
  NANDN U5589 ( .A(n4367), .B(creg[118]), .Z(n4411) );
  NANDN U5590 ( .A(n7188), .B(o[118]), .Z(n4410) );
  NAND U5591 ( .A(n4411), .B(n4410), .Z(c[118]) );
  NANDN U5592 ( .A(n4367), .B(creg[119]), .Z(n4413) );
  NANDN U5593 ( .A(n7188), .B(o[119]), .Z(n4412) );
  NAND U5594 ( .A(n4413), .B(n4412), .Z(c[119]) );
  NANDN U5595 ( .A(n4367), .B(creg[11]), .Z(n4415) );
  NANDN U5596 ( .A(n7188), .B(o[11]), .Z(n4414) );
  NAND U5597 ( .A(n4415), .B(n4414), .Z(c[11]) );
  NANDN U5598 ( .A(n4367), .B(creg[120]), .Z(n4417) );
  NANDN U5599 ( .A(n7188), .B(o[120]), .Z(n4416) );
  NAND U5600 ( .A(n4417), .B(n4416), .Z(c[120]) );
  NANDN U5601 ( .A(n4367), .B(creg[121]), .Z(n4419) );
  NANDN U5602 ( .A(n7188), .B(o[121]), .Z(n4418) );
  NAND U5603 ( .A(n4419), .B(n4418), .Z(c[121]) );
  NANDN U5604 ( .A(n4367), .B(creg[122]), .Z(n4421) );
  NANDN U5605 ( .A(n7188), .B(o[122]), .Z(n4420) );
  NAND U5606 ( .A(n4421), .B(n4420), .Z(c[122]) );
  NANDN U5607 ( .A(n4367), .B(creg[123]), .Z(n4423) );
  NANDN U5608 ( .A(n7188), .B(o[123]), .Z(n4422) );
  NAND U5609 ( .A(n4423), .B(n4422), .Z(c[123]) );
  NANDN U5610 ( .A(n4367), .B(creg[124]), .Z(n4425) );
  NANDN U5611 ( .A(n7188), .B(o[124]), .Z(n4424) );
  NAND U5612 ( .A(n4425), .B(n4424), .Z(c[124]) );
  NANDN U5613 ( .A(n4367), .B(creg[125]), .Z(n4427) );
  NANDN U5614 ( .A(n7188), .B(o[125]), .Z(n4426) );
  NAND U5615 ( .A(n4427), .B(n4426), .Z(c[125]) );
  NANDN U5616 ( .A(n4367), .B(creg[126]), .Z(n4429) );
  NANDN U5617 ( .A(n7188), .B(o[126]), .Z(n4428) );
  NAND U5618 ( .A(n4429), .B(n4428), .Z(c[126]) );
  NANDN U5619 ( .A(n4367), .B(creg[127]), .Z(n4431) );
  NANDN U5620 ( .A(n7188), .B(o[127]), .Z(n4430) );
  NAND U5621 ( .A(n4431), .B(n4430), .Z(c[127]) );
  NANDN U5622 ( .A(n4367), .B(creg[128]), .Z(n4433) );
  NANDN U5623 ( .A(n7188), .B(o[128]), .Z(n4432) );
  NAND U5624 ( .A(n4433), .B(n4432), .Z(c[128]) );
  NANDN U5625 ( .A(n4367), .B(creg[129]), .Z(n4435) );
  NANDN U5626 ( .A(n7188), .B(o[129]), .Z(n4434) );
  NAND U5627 ( .A(n4435), .B(n4434), .Z(c[129]) );
  NANDN U5628 ( .A(n4367), .B(creg[12]), .Z(n4437) );
  NANDN U5629 ( .A(n7188), .B(o[12]), .Z(n4436) );
  NAND U5630 ( .A(n4437), .B(n4436), .Z(c[12]) );
  NANDN U5631 ( .A(n4367), .B(creg[130]), .Z(n4439) );
  NANDN U5632 ( .A(n7188), .B(o[130]), .Z(n4438) );
  NAND U5633 ( .A(n4439), .B(n4438), .Z(c[130]) );
  NANDN U5634 ( .A(n4367), .B(creg[131]), .Z(n4441) );
  NANDN U5635 ( .A(n7188), .B(o[131]), .Z(n4440) );
  NAND U5636 ( .A(n4441), .B(n4440), .Z(c[131]) );
  NANDN U5637 ( .A(n4367), .B(creg[132]), .Z(n4443) );
  NANDN U5638 ( .A(n7188), .B(o[132]), .Z(n4442) );
  NAND U5639 ( .A(n4443), .B(n4442), .Z(c[132]) );
  NANDN U5640 ( .A(n4367), .B(creg[133]), .Z(n4445) );
  NANDN U5641 ( .A(n7188), .B(o[133]), .Z(n4444) );
  NAND U5642 ( .A(n4445), .B(n4444), .Z(c[133]) );
  NANDN U5643 ( .A(n4367), .B(creg[134]), .Z(n4447) );
  NANDN U5644 ( .A(n7188), .B(o[134]), .Z(n4446) );
  NAND U5645 ( .A(n4447), .B(n4446), .Z(c[134]) );
  NANDN U5646 ( .A(n4367), .B(creg[135]), .Z(n4449) );
  NANDN U5647 ( .A(n7188), .B(o[135]), .Z(n4448) );
  NAND U5648 ( .A(n4449), .B(n4448), .Z(c[135]) );
  NANDN U5649 ( .A(n4367), .B(creg[136]), .Z(n4451) );
  NANDN U5650 ( .A(n7188), .B(o[136]), .Z(n4450) );
  NAND U5651 ( .A(n4451), .B(n4450), .Z(c[136]) );
  NANDN U5652 ( .A(n4367), .B(creg[137]), .Z(n4453) );
  NANDN U5653 ( .A(n7188), .B(o[137]), .Z(n4452) );
  NAND U5654 ( .A(n4453), .B(n4452), .Z(c[137]) );
  NANDN U5655 ( .A(n4367), .B(creg[138]), .Z(n4455) );
  NANDN U5656 ( .A(n7188), .B(o[138]), .Z(n4454) );
  NAND U5657 ( .A(n4455), .B(n4454), .Z(c[138]) );
  NANDN U5658 ( .A(n4367), .B(creg[139]), .Z(n4457) );
  NANDN U5659 ( .A(n7188), .B(o[139]), .Z(n4456) );
  NAND U5660 ( .A(n4457), .B(n4456), .Z(c[139]) );
  NANDN U5661 ( .A(n4367), .B(creg[13]), .Z(n4459) );
  NANDN U5662 ( .A(n7188), .B(o[13]), .Z(n4458) );
  NAND U5663 ( .A(n4459), .B(n4458), .Z(c[13]) );
  NANDN U5664 ( .A(n4367), .B(creg[140]), .Z(n4461) );
  NANDN U5665 ( .A(n7188), .B(o[140]), .Z(n4460) );
  NAND U5666 ( .A(n4461), .B(n4460), .Z(c[140]) );
  NANDN U5667 ( .A(n4367), .B(creg[141]), .Z(n4463) );
  NANDN U5668 ( .A(n7188), .B(o[141]), .Z(n4462) );
  NAND U5669 ( .A(n4463), .B(n4462), .Z(c[141]) );
  NANDN U5670 ( .A(n4367), .B(creg[142]), .Z(n4465) );
  NANDN U5671 ( .A(n7188), .B(o[142]), .Z(n4464) );
  NAND U5672 ( .A(n4465), .B(n4464), .Z(c[142]) );
  NANDN U5673 ( .A(n4367), .B(creg[143]), .Z(n4467) );
  NANDN U5674 ( .A(n7188), .B(o[143]), .Z(n4466) );
  NAND U5675 ( .A(n4467), .B(n4466), .Z(c[143]) );
  NANDN U5676 ( .A(n4367), .B(creg[144]), .Z(n4469) );
  NANDN U5677 ( .A(n7188), .B(o[144]), .Z(n4468) );
  NAND U5678 ( .A(n4469), .B(n4468), .Z(c[144]) );
  NANDN U5679 ( .A(n4367), .B(creg[145]), .Z(n4471) );
  NANDN U5680 ( .A(n7188), .B(o[145]), .Z(n4470) );
  NAND U5681 ( .A(n4471), .B(n4470), .Z(c[145]) );
  NANDN U5682 ( .A(n4367), .B(creg[146]), .Z(n4473) );
  NANDN U5683 ( .A(n7188), .B(o[146]), .Z(n4472) );
  NAND U5684 ( .A(n4473), .B(n4472), .Z(c[146]) );
  NANDN U5685 ( .A(n4367), .B(creg[147]), .Z(n4475) );
  NANDN U5686 ( .A(n7188), .B(o[147]), .Z(n4474) );
  NAND U5687 ( .A(n4475), .B(n4474), .Z(c[147]) );
  NANDN U5688 ( .A(n4367), .B(creg[148]), .Z(n4477) );
  NANDN U5689 ( .A(n7188), .B(o[148]), .Z(n4476) );
  NAND U5690 ( .A(n4477), .B(n4476), .Z(c[148]) );
  NANDN U5691 ( .A(n4367), .B(creg[149]), .Z(n4479) );
  NANDN U5692 ( .A(n7188), .B(o[149]), .Z(n4478) );
  NAND U5693 ( .A(n4479), .B(n4478), .Z(c[149]) );
  NANDN U5694 ( .A(n4367), .B(creg[14]), .Z(n4481) );
  NANDN U5695 ( .A(n7188), .B(o[14]), .Z(n4480) );
  NAND U5696 ( .A(n4481), .B(n4480), .Z(c[14]) );
  NANDN U5697 ( .A(n4367), .B(creg[150]), .Z(n4483) );
  NANDN U5698 ( .A(n7188), .B(o[150]), .Z(n4482) );
  NAND U5699 ( .A(n4483), .B(n4482), .Z(c[150]) );
  NANDN U5700 ( .A(n4367), .B(creg[151]), .Z(n4485) );
  NANDN U5701 ( .A(n7188), .B(o[151]), .Z(n4484) );
  NAND U5702 ( .A(n4485), .B(n4484), .Z(c[151]) );
  NANDN U5703 ( .A(n4367), .B(creg[152]), .Z(n4487) );
  NANDN U5704 ( .A(n7188), .B(o[152]), .Z(n4486) );
  NAND U5705 ( .A(n4487), .B(n4486), .Z(c[152]) );
  NANDN U5706 ( .A(n4367), .B(creg[153]), .Z(n4489) );
  NANDN U5707 ( .A(n7188), .B(o[153]), .Z(n4488) );
  NAND U5708 ( .A(n4489), .B(n4488), .Z(c[153]) );
  NANDN U5709 ( .A(n4367), .B(creg[154]), .Z(n4491) );
  NANDN U5710 ( .A(n7188), .B(o[154]), .Z(n4490) );
  NAND U5711 ( .A(n4491), .B(n4490), .Z(c[154]) );
  NANDN U5712 ( .A(n4367), .B(creg[155]), .Z(n4493) );
  NANDN U5713 ( .A(n7188), .B(o[155]), .Z(n4492) );
  NAND U5714 ( .A(n4493), .B(n4492), .Z(c[155]) );
  NANDN U5715 ( .A(n4367), .B(creg[156]), .Z(n4495) );
  NANDN U5716 ( .A(n7188), .B(o[156]), .Z(n4494) );
  NAND U5717 ( .A(n4495), .B(n4494), .Z(c[156]) );
  NANDN U5718 ( .A(n4367), .B(creg[157]), .Z(n4497) );
  NANDN U5719 ( .A(n7188), .B(o[157]), .Z(n4496) );
  NAND U5720 ( .A(n4497), .B(n4496), .Z(c[157]) );
  NANDN U5721 ( .A(n4367), .B(creg[158]), .Z(n4499) );
  NANDN U5722 ( .A(n7188), .B(o[158]), .Z(n4498) );
  NAND U5723 ( .A(n4499), .B(n4498), .Z(c[158]) );
  NANDN U5724 ( .A(n4367), .B(creg[159]), .Z(n4501) );
  NANDN U5725 ( .A(n7188), .B(o[159]), .Z(n4500) );
  NAND U5726 ( .A(n4501), .B(n4500), .Z(c[159]) );
  NANDN U5727 ( .A(n4367), .B(creg[15]), .Z(n4503) );
  NANDN U5728 ( .A(n7188), .B(o[15]), .Z(n4502) );
  NAND U5729 ( .A(n4503), .B(n4502), .Z(c[15]) );
  NANDN U5730 ( .A(n4367), .B(creg[160]), .Z(n4505) );
  NANDN U5731 ( .A(n7188), .B(o[160]), .Z(n4504) );
  NAND U5732 ( .A(n4505), .B(n4504), .Z(c[160]) );
  NANDN U5733 ( .A(n4367), .B(creg[161]), .Z(n4507) );
  NANDN U5734 ( .A(n7188), .B(o[161]), .Z(n4506) );
  NAND U5735 ( .A(n4507), .B(n4506), .Z(c[161]) );
  NANDN U5736 ( .A(n4367), .B(creg[162]), .Z(n4509) );
  NANDN U5737 ( .A(n7188), .B(o[162]), .Z(n4508) );
  NAND U5738 ( .A(n4509), .B(n4508), .Z(c[162]) );
  NANDN U5739 ( .A(n4367), .B(creg[163]), .Z(n4511) );
  NANDN U5740 ( .A(n7188), .B(o[163]), .Z(n4510) );
  NAND U5741 ( .A(n4511), .B(n4510), .Z(c[163]) );
  NANDN U5742 ( .A(n4367), .B(creg[164]), .Z(n4513) );
  NANDN U5743 ( .A(n7188), .B(o[164]), .Z(n4512) );
  NAND U5744 ( .A(n4513), .B(n4512), .Z(c[164]) );
  NANDN U5745 ( .A(n4367), .B(creg[165]), .Z(n4515) );
  NANDN U5746 ( .A(n7188), .B(o[165]), .Z(n4514) );
  NAND U5747 ( .A(n4515), .B(n4514), .Z(c[165]) );
  NANDN U5748 ( .A(n4367), .B(creg[166]), .Z(n4517) );
  NANDN U5749 ( .A(n7188), .B(o[166]), .Z(n4516) );
  NAND U5750 ( .A(n4517), .B(n4516), .Z(c[166]) );
  NANDN U5751 ( .A(n4367), .B(creg[167]), .Z(n4519) );
  NANDN U5752 ( .A(n7188), .B(o[167]), .Z(n4518) );
  NAND U5753 ( .A(n4519), .B(n4518), .Z(c[167]) );
  NANDN U5754 ( .A(n4367), .B(creg[168]), .Z(n4521) );
  NANDN U5755 ( .A(n7188), .B(o[168]), .Z(n4520) );
  NAND U5756 ( .A(n4521), .B(n4520), .Z(c[168]) );
  NANDN U5757 ( .A(n4367), .B(creg[169]), .Z(n4523) );
  NANDN U5758 ( .A(n7188), .B(o[169]), .Z(n4522) );
  NAND U5759 ( .A(n4523), .B(n4522), .Z(c[169]) );
  NANDN U5760 ( .A(n4367), .B(creg[16]), .Z(n4525) );
  NANDN U5761 ( .A(n7188), .B(o[16]), .Z(n4524) );
  NAND U5762 ( .A(n4525), .B(n4524), .Z(c[16]) );
  NANDN U5763 ( .A(n4367), .B(creg[170]), .Z(n4527) );
  NANDN U5764 ( .A(n7188), .B(o[170]), .Z(n4526) );
  NAND U5765 ( .A(n4527), .B(n4526), .Z(c[170]) );
  NANDN U5766 ( .A(n4367), .B(creg[171]), .Z(n4529) );
  NANDN U5767 ( .A(n7188), .B(o[171]), .Z(n4528) );
  NAND U5768 ( .A(n4529), .B(n4528), .Z(c[171]) );
  NANDN U5769 ( .A(n4367), .B(creg[172]), .Z(n4531) );
  NANDN U5770 ( .A(n7188), .B(o[172]), .Z(n4530) );
  NAND U5771 ( .A(n4531), .B(n4530), .Z(c[172]) );
  NANDN U5772 ( .A(n4367), .B(creg[173]), .Z(n4533) );
  NANDN U5773 ( .A(n7188), .B(o[173]), .Z(n4532) );
  NAND U5774 ( .A(n4533), .B(n4532), .Z(c[173]) );
  NANDN U5775 ( .A(n4367), .B(creg[174]), .Z(n4535) );
  NANDN U5776 ( .A(n7188), .B(o[174]), .Z(n4534) );
  NAND U5777 ( .A(n4535), .B(n4534), .Z(c[174]) );
  NANDN U5778 ( .A(n4367), .B(creg[175]), .Z(n4537) );
  NANDN U5779 ( .A(n7188), .B(o[175]), .Z(n4536) );
  NAND U5780 ( .A(n4537), .B(n4536), .Z(c[175]) );
  NANDN U5781 ( .A(n4367), .B(creg[176]), .Z(n4539) );
  NANDN U5782 ( .A(n7188), .B(o[176]), .Z(n4538) );
  NAND U5783 ( .A(n4539), .B(n4538), .Z(c[176]) );
  NANDN U5784 ( .A(n4367), .B(creg[177]), .Z(n4541) );
  NANDN U5785 ( .A(n7188), .B(o[177]), .Z(n4540) );
  NAND U5786 ( .A(n4541), .B(n4540), .Z(c[177]) );
  NANDN U5787 ( .A(n4367), .B(creg[178]), .Z(n4543) );
  NANDN U5788 ( .A(n7188), .B(o[178]), .Z(n4542) );
  NAND U5789 ( .A(n4543), .B(n4542), .Z(c[178]) );
  NANDN U5790 ( .A(n4367), .B(creg[179]), .Z(n4545) );
  NANDN U5791 ( .A(n7188), .B(o[179]), .Z(n4544) );
  NAND U5792 ( .A(n4545), .B(n4544), .Z(c[179]) );
  NANDN U5793 ( .A(n4367), .B(creg[17]), .Z(n4547) );
  NANDN U5794 ( .A(n7188), .B(o[17]), .Z(n4546) );
  NAND U5795 ( .A(n4547), .B(n4546), .Z(c[17]) );
  NANDN U5796 ( .A(n4367), .B(creg[180]), .Z(n4549) );
  NANDN U5797 ( .A(n7188), .B(o[180]), .Z(n4548) );
  NAND U5798 ( .A(n4549), .B(n4548), .Z(c[180]) );
  NANDN U5799 ( .A(n4367), .B(creg[181]), .Z(n4551) );
  NANDN U5800 ( .A(n7188), .B(o[181]), .Z(n4550) );
  NAND U5801 ( .A(n4551), .B(n4550), .Z(c[181]) );
  NANDN U5802 ( .A(n4367), .B(creg[182]), .Z(n4553) );
  NANDN U5803 ( .A(n7188), .B(o[182]), .Z(n4552) );
  NAND U5804 ( .A(n4553), .B(n4552), .Z(c[182]) );
  NANDN U5805 ( .A(n4367), .B(creg[183]), .Z(n4555) );
  NANDN U5806 ( .A(n7188), .B(o[183]), .Z(n4554) );
  NAND U5807 ( .A(n4555), .B(n4554), .Z(c[183]) );
  NANDN U5808 ( .A(n4367), .B(creg[184]), .Z(n4557) );
  NANDN U5809 ( .A(n7188), .B(o[184]), .Z(n4556) );
  NAND U5810 ( .A(n4557), .B(n4556), .Z(c[184]) );
  NANDN U5811 ( .A(n4367), .B(creg[185]), .Z(n4559) );
  NANDN U5812 ( .A(n7188), .B(o[185]), .Z(n4558) );
  NAND U5813 ( .A(n4559), .B(n4558), .Z(c[185]) );
  NANDN U5814 ( .A(n4367), .B(creg[186]), .Z(n4561) );
  NANDN U5815 ( .A(n7188), .B(o[186]), .Z(n4560) );
  NAND U5816 ( .A(n4561), .B(n4560), .Z(c[186]) );
  NANDN U5817 ( .A(n4367), .B(creg[187]), .Z(n4563) );
  NANDN U5818 ( .A(n7188), .B(o[187]), .Z(n4562) );
  NAND U5819 ( .A(n4563), .B(n4562), .Z(c[187]) );
  NANDN U5820 ( .A(n4367), .B(creg[188]), .Z(n4565) );
  NANDN U5821 ( .A(n7188), .B(o[188]), .Z(n4564) );
  NAND U5822 ( .A(n4565), .B(n4564), .Z(c[188]) );
  NANDN U5823 ( .A(n4367), .B(creg[189]), .Z(n4567) );
  NANDN U5824 ( .A(n7188), .B(o[189]), .Z(n4566) );
  NAND U5825 ( .A(n4567), .B(n4566), .Z(c[189]) );
  NANDN U5826 ( .A(n4367), .B(creg[18]), .Z(n4569) );
  NANDN U5827 ( .A(n7188), .B(o[18]), .Z(n4568) );
  NAND U5828 ( .A(n4569), .B(n4568), .Z(c[18]) );
  NANDN U5829 ( .A(n4367), .B(creg[190]), .Z(n4571) );
  NANDN U5830 ( .A(n7188), .B(o[190]), .Z(n4570) );
  NAND U5831 ( .A(n4571), .B(n4570), .Z(c[190]) );
  NANDN U5832 ( .A(n4367), .B(creg[191]), .Z(n4573) );
  NANDN U5833 ( .A(n7188), .B(o[191]), .Z(n4572) );
  NAND U5834 ( .A(n4573), .B(n4572), .Z(c[191]) );
  NANDN U5835 ( .A(n4367), .B(creg[192]), .Z(n4575) );
  NANDN U5836 ( .A(n7188), .B(o[192]), .Z(n4574) );
  NAND U5837 ( .A(n4575), .B(n4574), .Z(c[192]) );
  NANDN U5838 ( .A(n4367), .B(creg[193]), .Z(n4577) );
  NANDN U5839 ( .A(n7188), .B(o[193]), .Z(n4576) );
  NAND U5840 ( .A(n4577), .B(n4576), .Z(c[193]) );
  NANDN U5841 ( .A(n4367), .B(creg[194]), .Z(n4579) );
  NANDN U5842 ( .A(n7188), .B(o[194]), .Z(n4578) );
  NAND U5843 ( .A(n4579), .B(n4578), .Z(c[194]) );
  NANDN U5844 ( .A(n4367), .B(creg[195]), .Z(n4581) );
  NANDN U5845 ( .A(n7188), .B(o[195]), .Z(n4580) );
  NAND U5846 ( .A(n4581), .B(n4580), .Z(c[195]) );
  NANDN U5847 ( .A(n4367), .B(creg[196]), .Z(n4583) );
  NANDN U5848 ( .A(n7188), .B(o[196]), .Z(n4582) );
  NAND U5849 ( .A(n4583), .B(n4582), .Z(c[196]) );
  NANDN U5850 ( .A(n4367), .B(creg[197]), .Z(n4585) );
  NANDN U5851 ( .A(n7188), .B(o[197]), .Z(n4584) );
  NAND U5852 ( .A(n4585), .B(n4584), .Z(c[197]) );
  NANDN U5853 ( .A(n4367), .B(creg[198]), .Z(n4587) );
  NANDN U5854 ( .A(n7188), .B(o[198]), .Z(n4586) );
  NAND U5855 ( .A(n4587), .B(n4586), .Z(c[198]) );
  NANDN U5856 ( .A(n4367), .B(creg[199]), .Z(n4589) );
  NANDN U5857 ( .A(n7188), .B(o[199]), .Z(n4588) );
  NAND U5858 ( .A(n4589), .B(n4588), .Z(c[199]) );
  NANDN U5859 ( .A(n4367), .B(creg[19]), .Z(n4591) );
  NANDN U5860 ( .A(n7188), .B(o[19]), .Z(n4590) );
  NAND U5861 ( .A(n4591), .B(n4590), .Z(c[19]) );
  NANDN U5862 ( .A(n4367), .B(creg[1]), .Z(n4593) );
  NANDN U5863 ( .A(n7188), .B(o[1]), .Z(n4592) );
  NAND U5864 ( .A(n4593), .B(n4592), .Z(c[1]) );
  NANDN U5865 ( .A(n4367), .B(creg[200]), .Z(n4595) );
  NANDN U5866 ( .A(n7188), .B(o[200]), .Z(n4594) );
  NAND U5867 ( .A(n4595), .B(n4594), .Z(c[200]) );
  NANDN U5868 ( .A(n4367), .B(creg[201]), .Z(n4597) );
  NANDN U5869 ( .A(n7188), .B(o[201]), .Z(n4596) );
  NAND U5870 ( .A(n4597), .B(n4596), .Z(c[201]) );
  NANDN U5871 ( .A(n4367), .B(creg[202]), .Z(n4599) );
  NANDN U5872 ( .A(n7188), .B(o[202]), .Z(n4598) );
  NAND U5873 ( .A(n4599), .B(n4598), .Z(c[202]) );
  NANDN U5874 ( .A(n4367), .B(creg[203]), .Z(n4601) );
  NANDN U5875 ( .A(n7188), .B(o[203]), .Z(n4600) );
  NAND U5876 ( .A(n4601), .B(n4600), .Z(c[203]) );
  NANDN U5877 ( .A(n4367), .B(creg[204]), .Z(n4603) );
  NANDN U5878 ( .A(n7188), .B(o[204]), .Z(n4602) );
  NAND U5879 ( .A(n4603), .B(n4602), .Z(c[204]) );
  NANDN U5880 ( .A(n4367), .B(creg[205]), .Z(n4605) );
  NANDN U5881 ( .A(n7188), .B(o[205]), .Z(n4604) );
  NAND U5882 ( .A(n4605), .B(n4604), .Z(c[205]) );
  NANDN U5883 ( .A(n4367), .B(creg[206]), .Z(n4607) );
  NANDN U5884 ( .A(n7188), .B(o[206]), .Z(n4606) );
  NAND U5885 ( .A(n4607), .B(n4606), .Z(c[206]) );
  NANDN U5886 ( .A(n4367), .B(creg[207]), .Z(n4609) );
  NANDN U5887 ( .A(n7188), .B(o[207]), .Z(n4608) );
  NAND U5888 ( .A(n4609), .B(n4608), .Z(c[207]) );
  NANDN U5889 ( .A(n4367), .B(creg[208]), .Z(n4611) );
  NANDN U5890 ( .A(n7188), .B(o[208]), .Z(n4610) );
  NAND U5891 ( .A(n4611), .B(n4610), .Z(c[208]) );
  NANDN U5892 ( .A(n4367), .B(creg[209]), .Z(n4613) );
  NANDN U5893 ( .A(n7188), .B(o[209]), .Z(n4612) );
  NAND U5894 ( .A(n4613), .B(n4612), .Z(c[209]) );
  NANDN U5895 ( .A(n4367), .B(creg[20]), .Z(n4615) );
  NANDN U5896 ( .A(n7188), .B(o[20]), .Z(n4614) );
  NAND U5897 ( .A(n4615), .B(n4614), .Z(c[20]) );
  NANDN U5898 ( .A(n4367), .B(creg[210]), .Z(n4617) );
  NANDN U5899 ( .A(n7188), .B(o[210]), .Z(n4616) );
  NAND U5900 ( .A(n4617), .B(n4616), .Z(c[210]) );
  NANDN U5901 ( .A(n4367), .B(creg[211]), .Z(n4619) );
  NANDN U5902 ( .A(n7188), .B(o[211]), .Z(n4618) );
  NAND U5903 ( .A(n4619), .B(n4618), .Z(c[211]) );
  NANDN U5904 ( .A(n4367), .B(creg[212]), .Z(n4621) );
  NANDN U5905 ( .A(n7188), .B(o[212]), .Z(n4620) );
  NAND U5906 ( .A(n4621), .B(n4620), .Z(c[212]) );
  NANDN U5907 ( .A(n4367), .B(creg[213]), .Z(n4623) );
  NANDN U5908 ( .A(n7188), .B(o[213]), .Z(n4622) );
  NAND U5909 ( .A(n4623), .B(n4622), .Z(c[213]) );
  NANDN U5910 ( .A(n4367), .B(creg[214]), .Z(n4625) );
  NANDN U5911 ( .A(n7188), .B(o[214]), .Z(n4624) );
  NAND U5912 ( .A(n4625), .B(n4624), .Z(c[214]) );
  NANDN U5913 ( .A(n4367), .B(creg[215]), .Z(n4627) );
  NANDN U5914 ( .A(n7188), .B(o[215]), .Z(n4626) );
  NAND U5915 ( .A(n4627), .B(n4626), .Z(c[215]) );
  NANDN U5916 ( .A(n4367), .B(creg[216]), .Z(n4629) );
  NANDN U5917 ( .A(n7188), .B(o[216]), .Z(n4628) );
  NAND U5918 ( .A(n4629), .B(n4628), .Z(c[216]) );
  NANDN U5919 ( .A(n4367), .B(creg[217]), .Z(n4631) );
  NANDN U5920 ( .A(n7188), .B(o[217]), .Z(n4630) );
  NAND U5921 ( .A(n4631), .B(n4630), .Z(c[217]) );
  NANDN U5922 ( .A(n4367), .B(creg[218]), .Z(n4633) );
  NANDN U5923 ( .A(n7188), .B(o[218]), .Z(n4632) );
  NAND U5924 ( .A(n4633), .B(n4632), .Z(c[218]) );
  NANDN U5925 ( .A(n4367), .B(creg[219]), .Z(n4635) );
  NANDN U5926 ( .A(n7188), .B(o[219]), .Z(n4634) );
  NAND U5927 ( .A(n4635), .B(n4634), .Z(c[219]) );
  NANDN U5928 ( .A(n4367), .B(creg[21]), .Z(n4637) );
  NANDN U5929 ( .A(n7188), .B(o[21]), .Z(n4636) );
  NAND U5930 ( .A(n4637), .B(n4636), .Z(c[21]) );
  NANDN U5931 ( .A(n4367), .B(creg[220]), .Z(n4639) );
  NANDN U5932 ( .A(n7188), .B(o[220]), .Z(n4638) );
  NAND U5933 ( .A(n4639), .B(n4638), .Z(c[220]) );
  NANDN U5934 ( .A(n4367), .B(creg[221]), .Z(n4641) );
  NANDN U5935 ( .A(n7188), .B(o[221]), .Z(n4640) );
  NAND U5936 ( .A(n4641), .B(n4640), .Z(c[221]) );
  NANDN U5937 ( .A(n4367), .B(creg[222]), .Z(n4643) );
  NANDN U5938 ( .A(n7188), .B(o[222]), .Z(n4642) );
  NAND U5939 ( .A(n4643), .B(n4642), .Z(c[222]) );
  NANDN U5940 ( .A(n4367), .B(creg[223]), .Z(n4645) );
  NANDN U5941 ( .A(n7188), .B(o[223]), .Z(n4644) );
  NAND U5942 ( .A(n4645), .B(n4644), .Z(c[223]) );
  NANDN U5943 ( .A(n4367), .B(creg[224]), .Z(n4647) );
  NANDN U5944 ( .A(n7188), .B(o[224]), .Z(n4646) );
  NAND U5945 ( .A(n4647), .B(n4646), .Z(c[224]) );
  NANDN U5946 ( .A(n4367), .B(creg[225]), .Z(n4649) );
  NANDN U5947 ( .A(n7188), .B(o[225]), .Z(n4648) );
  NAND U5948 ( .A(n4649), .B(n4648), .Z(c[225]) );
  NANDN U5949 ( .A(n4367), .B(creg[226]), .Z(n4651) );
  NANDN U5950 ( .A(n7188), .B(o[226]), .Z(n4650) );
  NAND U5951 ( .A(n4651), .B(n4650), .Z(c[226]) );
  NANDN U5952 ( .A(n4367), .B(creg[227]), .Z(n4653) );
  NANDN U5953 ( .A(n7188), .B(o[227]), .Z(n4652) );
  NAND U5954 ( .A(n4653), .B(n4652), .Z(c[227]) );
  NANDN U5955 ( .A(n4367), .B(creg[228]), .Z(n4655) );
  NANDN U5956 ( .A(n7188), .B(o[228]), .Z(n4654) );
  NAND U5957 ( .A(n4655), .B(n4654), .Z(c[228]) );
  NANDN U5958 ( .A(n4367), .B(creg[229]), .Z(n4657) );
  NANDN U5959 ( .A(n7188), .B(o[229]), .Z(n4656) );
  NAND U5960 ( .A(n4657), .B(n4656), .Z(c[229]) );
  NANDN U5961 ( .A(n4367), .B(creg[22]), .Z(n4659) );
  NANDN U5962 ( .A(n7188), .B(o[22]), .Z(n4658) );
  NAND U5963 ( .A(n4659), .B(n4658), .Z(c[22]) );
  NANDN U5964 ( .A(n4367), .B(creg[230]), .Z(n4661) );
  NANDN U5965 ( .A(n7188), .B(o[230]), .Z(n4660) );
  NAND U5966 ( .A(n4661), .B(n4660), .Z(c[230]) );
  NANDN U5967 ( .A(n4367), .B(creg[231]), .Z(n4663) );
  NANDN U5968 ( .A(n7188), .B(o[231]), .Z(n4662) );
  NAND U5969 ( .A(n4663), .B(n4662), .Z(c[231]) );
  NANDN U5970 ( .A(n4367), .B(creg[232]), .Z(n4665) );
  NANDN U5971 ( .A(n7188), .B(o[232]), .Z(n4664) );
  NAND U5972 ( .A(n4665), .B(n4664), .Z(c[232]) );
  NANDN U5973 ( .A(n4367), .B(creg[233]), .Z(n4667) );
  NANDN U5974 ( .A(n7188), .B(o[233]), .Z(n4666) );
  NAND U5975 ( .A(n4667), .B(n4666), .Z(c[233]) );
  NANDN U5976 ( .A(n4367), .B(creg[234]), .Z(n4669) );
  NANDN U5977 ( .A(n7188), .B(o[234]), .Z(n4668) );
  NAND U5978 ( .A(n4669), .B(n4668), .Z(c[234]) );
  NANDN U5979 ( .A(n4367), .B(creg[235]), .Z(n4671) );
  NANDN U5980 ( .A(n7188), .B(o[235]), .Z(n4670) );
  NAND U5981 ( .A(n4671), .B(n4670), .Z(c[235]) );
  NANDN U5982 ( .A(n4367), .B(creg[236]), .Z(n4673) );
  NANDN U5983 ( .A(n7188), .B(o[236]), .Z(n4672) );
  NAND U5984 ( .A(n4673), .B(n4672), .Z(c[236]) );
  NANDN U5985 ( .A(n4367), .B(creg[237]), .Z(n4675) );
  NANDN U5986 ( .A(n7188), .B(o[237]), .Z(n4674) );
  NAND U5987 ( .A(n4675), .B(n4674), .Z(c[237]) );
  NANDN U5988 ( .A(n4367), .B(creg[238]), .Z(n4677) );
  NANDN U5989 ( .A(n7188), .B(o[238]), .Z(n4676) );
  NAND U5990 ( .A(n4677), .B(n4676), .Z(c[238]) );
  NANDN U5991 ( .A(n4367), .B(creg[239]), .Z(n4679) );
  NANDN U5992 ( .A(n7188), .B(o[239]), .Z(n4678) );
  NAND U5993 ( .A(n4679), .B(n4678), .Z(c[239]) );
  NANDN U5994 ( .A(n4367), .B(creg[23]), .Z(n4681) );
  NANDN U5995 ( .A(n7188), .B(o[23]), .Z(n4680) );
  NAND U5996 ( .A(n4681), .B(n4680), .Z(c[23]) );
  NANDN U5997 ( .A(n4367), .B(creg[240]), .Z(n4683) );
  NANDN U5998 ( .A(n7188), .B(o[240]), .Z(n4682) );
  NAND U5999 ( .A(n4683), .B(n4682), .Z(c[240]) );
  NANDN U6000 ( .A(n4367), .B(creg[241]), .Z(n4685) );
  NANDN U6001 ( .A(n7188), .B(o[241]), .Z(n4684) );
  NAND U6002 ( .A(n4685), .B(n4684), .Z(c[241]) );
  NANDN U6003 ( .A(n4367), .B(creg[242]), .Z(n4687) );
  NANDN U6004 ( .A(n7188), .B(o[242]), .Z(n4686) );
  NAND U6005 ( .A(n4687), .B(n4686), .Z(c[242]) );
  NANDN U6006 ( .A(n4367), .B(creg[243]), .Z(n4689) );
  NANDN U6007 ( .A(n7188), .B(o[243]), .Z(n4688) );
  NAND U6008 ( .A(n4689), .B(n4688), .Z(c[243]) );
  NANDN U6009 ( .A(n4367), .B(creg[244]), .Z(n4691) );
  NANDN U6010 ( .A(n7188), .B(o[244]), .Z(n4690) );
  NAND U6011 ( .A(n4691), .B(n4690), .Z(c[244]) );
  NANDN U6012 ( .A(n4367), .B(creg[245]), .Z(n4693) );
  NANDN U6013 ( .A(n7188), .B(o[245]), .Z(n4692) );
  NAND U6014 ( .A(n4693), .B(n4692), .Z(c[245]) );
  NANDN U6015 ( .A(n4367), .B(creg[246]), .Z(n4695) );
  NANDN U6016 ( .A(n7188), .B(o[246]), .Z(n4694) );
  NAND U6017 ( .A(n4695), .B(n4694), .Z(c[246]) );
  NANDN U6018 ( .A(n4367), .B(creg[247]), .Z(n4697) );
  NANDN U6019 ( .A(n7188), .B(o[247]), .Z(n4696) );
  NAND U6020 ( .A(n4697), .B(n4696), .Z(c[247]) );
  NANDN U6021 ( .A(n4367), .B(creg[248]), .Z(n4699) );
  NANDN U6022 ( .A(n7188), .B(o[248]), .Z(n4698) );
  NAND U6023 ( .A(n4699), .B(n4698), .Z(c[248]) );
  NANDN U6024 ( .A(n4367), .B(creg[249]), .Z(n4701) );
  NANDN U6025 ( .A(n7188), .B(o[249]), .Z(n4700) );
  NAND U6026 ( .A(n4701), .B(n4700), .Z(c[249]) );
  NANDN U6027 ( .A(n4367), .B(creg[24]), .Z(n4703) );
  NANDN U6028 ( .A(n7188), .B(o[24]), .Z(n4702) );
  NAND U6029 ( .A(n4703), .B(n4702), .Z(c[24]) );
  NANDN U6030 ( .A(n4367), .B(creg[250]), .Z(n4705) );
  NANDN U6031 ( .A(n7188), .B(o[250]), .Z(n4704) );
  NAND U6032 ( .A(n4705), .B(n4704), .Z(c[250]) );
  NANDN U6033 ( .A(n4367), .B(creg[251]), .Z(n4707) );
  NANDN U6034 ( .A(n7188), .B(o[251]), .Z(n4706) );
  NAND U6035 ( .A(n4707), .B(n4706), .Z(c[251]) );
  NANDN U6036 ( .A(n4367), .B(creg[252]), .Z(n4709) );
  NANDN U6037 ( .A(n7188), .B(o[252]), .Z(n4708) );
  NAND U6038 ( .A(n4709), .B(n4708), .Z(c[252]) );
  NANDN U6039 ( .A(n4367), .B(creg[253]), .Z(n4711) );
  NANDN U6040 ( .A(n7188), .B(o[253]), .Z(n4710) );
  NAND U6041 ( .A(n4711), .B(n4710), .Z(c[253]) );
  NANDN U6042 ( .A(n4367), .B(creg[254]), .Z(n4713) );
  NANDN U6043 ( .A(n7188), .B(o[254]), .Z(n4712) );
  NAND U6044 ( .A(n4713), .B(n4712), .Z(c[254]) );
  NANDN U6045 ( .A(n4367), .B(creg[255]), .Z(n4715) );
  NANDN U6046 ( .A(n7188), .B(o[255]), .Z(n4714) );
  NAND U6047 ( .A(n4715), .B(n4714), .Z(c[255]) );
  NANDN U6048 ( .A(n4367), .B(creg[25]), .Z(n4717) );
  NANDN U6049 ( .A(n7188), .B(o[25]), .Z(n4716) );
  NAND U6050 ( .A(n4717), .B(n4716), .Z(c[25]) );
  NANDN U6051 ( .A(n4367), .B(creg[26]), .Z(n4719) );
  NANDN U6052 ( .A(n7188), .B(o[26]), .Z(n4718) );
  NAND U6053 ( .A(n4719), .B(n4718), .Z(c[26]) );
  NANDN U6054 ( .A(n4367), .B(creg[27]), .Z(n4721) );
  NANDN U6055 ( .A(n7188), .B(o[27]), .Z(n4720) );
  NAND U6056 ( .A(n4721), .B(n4720), .Z(c[27]) );
  NANDN U6057 ( .A(n4367), .B(creg[28]), .Z(n4723) );
  NANDN U6058 ( .A(n7188), .B(o[28]), .Z(n4722) );
  NAND U6059 ( .A(n4723), .B(n4722), .Z(c[28]) );
  NANDN U6060 ( .A(n4367), .B(creg[29]), .Z(n4725) );
  NANDN U6061 ( .A(n7188), .B(o[29]), .Z(n4724) );
  NAND U6062 ( .A(n4725), .B(n4724), .Z(c[29]) );
  NANDN U6063 ( .A(n4367), .B(creg[2]), .Z(n4727) );
  NANDN U6064 ( .A(n7188), .B(o[2]), .Z(n4726) );
  NAND U6065 ( .A(n4727), .B(n4726), .Z(c[2]) );
  NANDN U6066 ( .A(n4367), .B(creg[30]), .Z(n4729) );
  NANDN U6067 ( .A(n7188), .B(o[30]), .Z(n4728) );
  NAND U6068 ( .A(n4729), .B(n4728), .Z(c[30]) );
  NANDN U6069 ( .A(n4367), .B(creg[31]), .Z(n4731) );
  NANDN U6070 ( .A(n7188), .B(o[31]), .Z(n4730) );
  NAND U6071 ( .A(n4731), .B(n4730), .Z(c[31]) );
  NANDN U6072 ( .A(n4367), .B(creg[32]), .Z(n4733) );
  NANDN U6073 ( .A(n7188), .B(o[32]), .Z(n4732) );
  NAND U6074 ( .A(n4733), .B(n4732), .Z(c[32]) );
  NANDN U6075 ( .A(n4367), .B(creg[33]), .Z(n4735) );
  NANDN U6076 ( .A(n7188), .B(o[33]), .Z(n4734) );
  NAND U6077 ( .A(n4735), .B(n4734), .Z(c[33]) );
  NANDN U6078 ( .A(n4367), .B(creg[34]), .Z(n4737) );
  NANDN U6079 ( .A(n7188), .B(o[34]), .Z(n4736) );
  NAND U6080 ( .A(n4737), .B(n4736), .Z(c[34]) );
  NANDN U6081 ( .A(n4367), .B(creg[35]), .Z(n4739) );
  NANDN U6082 ( .A(n7188), .B(o[35]), .Z(n4738) );
  NAND U6083 ( .A(n4739), .B(n4738), .Z(c[35]) );
  NANDN U6084 ( .A(n4367), .B(creg[36]), .Z(n4741) );
  NANDN U6085 ( .A(n7188), .B(o[36]), .Z(n4740) );
  NAND U6086 ( .A(n4741), .B(n4740), .Z(c[36]) );
  NANDN U6087 ( .A(n4367), .B(creg[37]), .Z(n4743) );
  NANDN U6088 ( .A(n7188), .B(o[37]), .Z(n4742) );
  NAND U6089 ( .A(n4743), .B(n4742), .Z(c[37]) );
  NANDN U6090 ( .A(n4367), .B(creg[38]), .Z(n4745) );
  NANDN U6091 ( .A(n7188), .B(o[38]), .Z(n4744) );
  NAND U6092 ( .A(n4745), .B(n4744), .Z(c[38]) );
  NANDN U6093 ( .A(n4367), .B(creg[39]), .Z(n4747) );
  NANDN U6094 ( .A(n7188), .B(o[39]), .Z(n4746) );
  NAND U6095 ( .A(n4747), .B(n4746), .Z(c[39]) );
  NANDN U6096 ( .A(n4367), .B(creg[3]), .Z(n4749) );
  NANDN U6097 ( .A(n7188), .B(o[3]), .Z(n4748) );
  NAND U6098 ( .A(n4749), .B(n4748), .Z(c[3]) );
  NANDN U6099 ( .A(n4367), .B(creg[40]), .Z(n4751) );
  NANDN U6100 ( .A(n7188), .B(o[40]), .Z(n4750) );
  NAND U6101 ( .A(n4751), .B(n4750), .Z(c[40]) );
  NANDN U6102 ( .A(n4367), .B(creg[41]), .Z(n4753) );
  NANDN U6103 ( .A(n7188), .B(o[41]), .Z(n4752) );
  NAND U6104 ( .A(n4753), .B(n4752), .Z(c[41]) );
  NANDN U6105 ( .A(n4367), .B(creg[42]), .Z(n4755) );
  NANDN U6106 ( .A(n7188), .B(o[42]), .Z(n4754) );
  NAND U6107 ( .A(n4755), .B(n4754), .Z(c[42]) );
  NANDN U6108 ( .A(n4367), .B(creg[43]), .Z(n4757) );
  NANDN U6109 ( .A(n7188), .B(o[43]), .Z(n4756) );
  NAND U6110 ( .A(n4757), .B(n4756), .Z(c[43]) );
  NANDN U6111 ( .A(n4367), .B(creg[44]), .Z(n4759) );
  NANDN U6112 ( .A(n7188), .B(o[44]), .Z(n4758) );
  NAND U6113 ( .A(n4759), .B(n4758), .Z(c[44]) );
  NANDN U6114 ( .A(n4367), .B(creg[45]), .Z(n4761) );
  NANDN U6115 ( .A(n7188), .B(o[45]), .Z(n4760) );
  NAND U6116 ( .A(n4761), .B(n4760), .Z(c[45]) );
  NANDN U6117 ( .A(n4367), .B(creg[46]), .Z(n4763) );
  NANDN U6118 ( .A(n7188), .B(o[46]), .Z(n4762) );
  NAND U6119 ( .A(n4763), .B(n4762), .Z(c[46]) );
  NANDN U6120 ( .A(n4367), .B(creg[47]), .Z(n4765) );
  NANDN U6121 ( .A(n7188), .B(o[47]), .Z(n4764) );
  NAND U6122 ( .A(n4765), .B(n4764), .Z(c[47]) );
  NANDN U6123 ( .A(n4367), .B(creg[48]), .Z(n4767) );
  NANDN U6124 ( .A(n7188), .B(o[48]), .Z(n4766) );
  NAND U6125 ( .A(n4767), .B(n4766), .Z(c[48]) );
  NANDN U6126 ( .A(n4367), .B(creg[49]), .Z(n4769) );
  NANDN U6127 ( .A(n7188), .B(o[49]), .Z(n4768) );
  NAND U6128 ( .A(n4769), .B(n4768), .Z(c[49]) );
  NANDN U6129 ( .A(n4367), .B(creg[4]), .Z(n4771) );
  NANDN U6130 ( .A(n7188), .B(o[4]), .Z(n4770) );
  NAND U6131 ( .A(n4771), .B(n4770), .Z(c[4]) );
  NANDN U6132 ( .A(n4367), .B(creg[50]), .Z(n4773) );
  NANDN U6133 ( .A(n7188), .B(o[50]), .Z(n4772) );
  NAND U6134 ( .A(n4773), .B(n4772), .Z(c[50]) );
  NANDN U6135 ( .A(n4367), .B(creg[51]), .Z(n4775) );
  NANDN U6136 ( .A(n7188), .B(o[51]), .Z(n4774) );
  NAND U6137 ( .A(n4775), .B(n4774), .Z(c[51]) );
  NANDN U6138 ( .A(n4367), .B(creg[52]), .Z(n4777) );
  NANDN U6139 ( .A(n7188), .B(o[52]), .Z(n4776) );
  NAND U6140 ( .A(n4777), .B(n4776), .Z(c[52]) );
  NANDN U6141 ( .A(n4367), .B(creg[53]), .Z(n4779) );
  NANDN U6142 ( .A(n7188), .B(o[53]), .Z(n4778) );
  NAND U6143 ( .A(n4779), .B(n4778), .Z(c[53]) );
  NANDN U6144 ( .A(n4367), .B(creg[54]), .Z(n4781) );
  NANDN U6145 ( .A(n7188), .B(o[54]), .Z(n4780) );
  NAND U6146 ( .A(n4781), .B(n4780), .Z(c[54]) );
  NANDN U6147 ( .A(n4367), .B(creg[55]), .Z(n4783) );
  NANDN U6148 ( .A(n7188), .B(o[55]), .Z(n4782) );
  NAND U6149 ( .A(n4783), .B(n4782), .Z(c[55]) );
  NANDN U6150 ( .A(n4367), .B(creg[56]), .Z(n4785) );
  NANDN U6151 ( .A(n7188), .B(o[56]), .Z(n4784) );
  NAND U6152 ( .A(n4785), .B(n4784), .Z(c[56]) );
  NANDN U6153 ( .A(n4367), .B(creg[57]), .Z(n4787) );
  NANDN U6154 ( .A(n7188), .B(o[57]), .Z(n4786) );
  NAND U6155 ( .A(n4787), .B(n4786), .Z(c[57]) );
  NANDN U6156 ( .A(n4367), .B(creg[58]), .Z(n4789) );
  NANDN U6157 ( .A(n7188), .B(o[58]), .Z(n4788) );
  NAND U6158 ( .A(n4789), .B(n4788), .Z(c[58]) );
  NANDN U6159 ( .A(n4367), .B(creg[59]), .Z(n4791) );
  NANDN U6160 ( .A(n7188), .B(o[59]), .Z(n4790) );
  NAND U6161 ( .A(n4791), .B(n4790), .Z(c[59]) );
  NANDN U6162 ( .A(n4367), .B(creg[5]), .Z(n4793) );
  NANDN U6163 ( .A(n7188), .B(o[5]), .Z(n4792) );
  NAND U6164 ( .A(n4793), .B(n4792), .Z(c[5]) );
  NANDN U6165 ( .A(n4367), .B(creg[60]), .Z(n4795) );
  NANDN U6166 ( .A(n7188), .B(o[60]), .Z(n4794) );
  NAND U6167 ( .A(n4795), .B(n4794), .Z(c[60]) );
  NANDN U6168 ( .A(n4367), .B(creg[61]), .Z(n4797) );
  NANDN U6169 ( .A(n7188), .B(o[61]), .Z(n4796) );
  NAND U6170 ( .A(n4797), .B(n4796), .Z(c[61]) );
  NANDN U6171 ( .A(n4367), .B(creg[62]), .Z(n4799) );
  NANDN U6172 ( .A(n7188), .B(o[62]), .Z(n4798) );
  NAND U6173 ( .A(n4799), .B(n4798), .Z(c[62]) );
  NANDN U6174 ( .A(n4367), .B(creg[63]), .Z(n4801) );
  NANDN U6175 ( .A(n7188), .B(o[63]), .Z(n4800) );
  NAND U6176 ( .A(n4801), .B(n4800), .Z(c[63]) );
  NANDN U6177 ( .A(n4367), .B(creg[64]), .Z(n4803) );
  NANDN U6178 ( .A(n7188), .B(o[64]), .Z(n4802) );
  NAND U6179 ( .A(n4803), .B(n4802), .Z(c[64]) );
  NANDN U6180 ( .A(n4367), .B(creg[65]), .Z(n4805) );
  NANDN U6181 ( .A(n7188), .B(o[65]), .Z(n4804) );
  NAND U6182 ( .A(n4805), .B(n4804), .Z(c[65]) );
  NANDN U6183 ( .A(n4367), .B(creg[66]), .Z(n4807) );
  NANDN U6184 ( .A(n7188), .B(o[66]), .Z(n4806) );
  NAND U6185 ( .A(n4807), .B(n4806), .Z(c[66]) );
  NANDN U6186 ( .A(n4367), .B(creg[67]), .Z(n4809) );
  NANDN U6187 ( .A(n7188), .B(o[67]), .Z(n4808) );
  NAND U6188 ( .A(n4809), .B(n4808), .Z(c[67]) );
  NANDN U6189 ( .A(n4367), .B(creg[68]), .Z(n4811) );
  NANDN U6190 ( .A(n7188), .B(o[68]), .Z(n4810) );
  NAND U6191 ( .A(n4811), .B(n4810), .Z(c[68]) );
  NANDN U6192 ( .A(n4367), .B(creg[69]), .Z(n4813) );
  NANDN U6193 ( .A(n7188), .B(o[69]), .Z(n4812) );
  NAND U6194 ( .A(n4813), .B(n4812), .Z(c[69]) );
  NANDN U6195 ( .A(n4367), .B(creg[6]), .Z(n4815) );
  NANDN U6196 ( .A(n7188), .B(o[6]), .Z(n4814) );
  NAND U6197 ( .A(n4815), .B(n4814), .Z(c[6]) );
  NANDN U6198 ( .A(n4367), .B(creg[70]), .Z(n4817) );
  NANDN U6199 ( .A(n7188), .B(o[70]), .Z(n4816) );
  NAND U6200 ( .A(n4817), .B(n4816), .Z(c[70]) );
  NANDN U6201 ( .A(n4367), .B(creg[71]), .Z(n4819) );
  NANDN U6202 ( .A(n7188), .B(o[71]), .Z(n4818) );
  NAND U6203 ( .A(n4819), .B(n4818), .Z(c[71]) );
  NANDN U6204 ( .A(n4367), .B(creg[72]), .Z(n4821) );
  NANDN U6205 ( .A(n7188), .B(o[72]), .Z(n4820) );
  NAND U6206 ( .A(n4821), .B(n4820), .Z(c[72]) );
  NANDN U6207 ( .A(n4367), .B(creg[73]), .Z(n4823) );
  NANDN U6208 ( .A(n7188), .B(o[73]), .Z(n4822) );
  NAND U6209 ( .A(n4823), .B(n4822), .Z(c[73]) );
  NANDN U6210 ( .A(n4367), .B(creg[74]), .Z(n4825) );
  NANDN U6211 ( .A(n7188), .B(o[74]), .Z(n4824) );
  NAND U6212 ( .A(n4825), .B(n4824), .Z(c[74]) );
  NANDN U6213 ( .A(n4367), .B(creg[75]), .Z(n4827) );
  NANDN U6214 ( .A(n7188), .B(o[75]), .Z(n4826) );
  NAND U6215 ( .A(n4827), .B(n4826), .Z(c[75]) );
  NANDN U6216 ( .A(n4367), .B(creg[76]), .Z(n4829) );
  NANDN U6217 ( .A(n7188), .B(o[76]), .Z(n4828) );
  NAND U6218 ( .A(n4829), .B(n4828), .Z(c[76]) );
  NANDN U6219 ( .A(n4367), .B(creg[77]), .Z(n4831) );
  NANDN U6220 ( .A(n7188), .B(o[77]), .Z(n4830) );
  NAND U6221 ( .A(n4831), .B(n4830), .Z(c[77]) );
  NANDN U6222 ( .A(n4367), .B(creg[78]), .Z(n4833) );
  NANDN U6223 ( .A(n7188), .B(o[78]), .Z(n4832) );
  NAND U6224 ( .A(n4833), .B(n4832), .Z(c[78]) );
  NANDN U6225 ( .A(n4367), .B(creg[79]), .Z(n4835) );
  NANDN U6226 ( .A(n7188), .B(o[79]), .Z(n4834) );
  NAND U6227 ( .A(n4835), .B(n4834), .Z(c[79]) );
  NANDN U6228 ( .A(n4367), .B(creg[7]), .Z(n4837) );
  NANDN U6229 ( .A(n7188), .B(o[7]), .Z(n4836) );
  NAND U6230 ( .A(n4837), .B(n4836), .Z(c[7]) );
  NANDN U6231 ( .A(n4367), .B(creg[80]), .Z(n4839) );
  NANDN U6232 ( .A(n7188), .B(o[80]), .Z(n4838) );
  NAND U6233 ( .A(n4839), .B(n4838), .Z(c[80]) );
  NANDN U6234 ( .A(n4367), .B(creg[81]), .Z(n4841) );
  NANDN U6235 ( .A(n7188), .B(o[81]), .Z(n4840) );
  NAND U6236 ( .A(n4841), .B(n4840), .Z(c[81]) );
  NANDN U6237 ( .A(n4367), .B(creg[82]), .Z(n4843) );
  NANDN U6238 ( .A(n7188), .B(o[82]), .Z(n4842) );
  NAND U6239 ( .A(n4843), .B(n4842), .Z(c[82]) );
  NANDN U6240 ( .A(n4367), .B(creg[83]), .Z(n4845) );
  NANDN U6241 ( .A(n7188), .B(o[83]), .Z(n4844) );
  NAND U6242 ( .A(n4845), .B(n4844), .Z(c[83]) );
  NANDN U6243 ( .A(n4367), .B(creg[84]), .Z(n4847) );
  NANDN U6244 ( .A(n7188), .B(o[84]), .Z(n4846) );
  NAND U6245 ( .A(n4847), .B(n4846), .Z(c[84]) );
  NANDN U6246 ( .A(n4367), .B(creg[85]), .Z(n4849) );
  NANDN U6247 ( .A(n7188), .B(o[85]), .Z(n4848) );
  NAND U6248 ( .A(n4849), .B(n4848), .Z(c[85]) );
  NANDN U6249 ( .A(n4367), .B(creg[86]), .Z(n4851) );
  NANDN U6250 ( .A(n7188), .B(o[86]), .Z(n4850) );
  NAND U6251 ( .A(n4851), .B(n4850), .Z(c[86]) );
  NANDN U6252 ( .A(n4367), .B(creg[87]), .Z(n4853) );
  NANDN U6253 ( .A(n7188), .B(o[87]), .Z(n4852) );
  NAND U6254 ( .A(n4853), .B(n4852), .Z(c[87]) );
  NANDN U6255 ( .A(n4367), .B(creg[88]), .Z(n4855) );
  NANDN U6256 ( .A(n7188), .B(o[88]), .Z(n4854) );
  NAND U6257 ( .A(n4855), .B(n4854), .Z(c[88]) );
  NANDN U6258 ( .A(n4367), .B(creg[89]), .Z(n4857) );
  NANDN U6259 ( .A(n7188), .B(o[89]), .Z(n4856) );
  NAND U6260 ( .A(n4857), .B(n4856), .Z(c[89]) );
  NANDN U6261 ( .A(n4367), .B(creg[8]), .Z(n4859) );
  NANDN U6262 ( .A(n7188), .B(o[8]), .Z(n4858) );
  NAND U6263 ( .A(n4859), .B(n4858), .Z(c[8]) );
  NANDN U6264 ( .A(n4367), .B(creg[90]), .Z(n4861) );
  NANDN U6265 ( .A(n7188), .B(o[90]), .Z(n4860) );
  NAND U6266 ( .A(n4861), .B(n4860), .Z(c[90]) );
  NANDN U6267 ( .A(n4367), .B(creg[91]), .Z(n4863) );
  NANDN U6268 ( .A(n7188), .B(o[91]), .Z(n4862) );
  NAND U6269 ( .A(n4863), .B(n4862), .Z(c[91]) );
  NANDN U6270 ( .A(n4367), .B(creg[92]), .Z(n4865) );
  NANDN U6271 ( .A(n7188), .B(o[92]), .Z(n4864) );
  NAND U6272 ( .A(n4865), .B(n4864), .Z(c[92]) );
  NANDN U6273 ( .A(n4367), .B(creg[93]), .Z(n4867) );
  NANDN U6274 ( .A(n7188), .B(o[93]), .Z(n4866) );
  NAND U6275 ( .A(n4867), .B(n4866), .Z(c[93]) );
  NANDN U6276 ( .A(n4367), .B(creg[94]), .Z(n4869) );
  NANDN U6277 ( .A(n7188), .B(o[94]), .Z(n4868) );
  NAND U6278 ( .A(n4869), .B(n4868), .Z(c[94]) );
  NANDN U6279 ( .A(n4367), .B(creg[95]), .Z(n4871) );
  NANDN U6280 ( .A(n7188), .B(o[95]), .Z(n4870) );
  NAND U6281 ( .A(n4871), .B(n4870), .Z(c[95]) );
  NANDN U6282 ( .A(n4367), .B(creg[96]), .Z(n4873) );
  NANDN U6283 ( .A(n7188), .B(o[96]), .Z(n4872) );
  NAND U6284 ( .A(n4873), .B(n4872), .Z(c[96]) );
  NANDN U6285 ( .A(n4367), .B(creg[97]), .Z(n4875) );
  NANDN U6286 ( .A(n7188), .B(o[97]), .Z(n4874) );
  NAND U6287 ( .A(n4875), .B(n4874), .Z(c[97]) );
  NANDN U6288 ( .A(n4367), .B(creg[98]), .Z(n4877) );
  NANDN U6289 ( .A(n7188), .B(o[98]), .Z(n4876) );
  NAND U6290 ( .A(n4877), .B(n4876), .Z(c[98]) );
  NANDN U6291 ( .A(n4367), .B(creg[99]), .Z(n4879) );
  NANDN U6292 ( .A(n7188), .B(o[99]), .Z(n4878) );
  NAND U6293 ( .A(n4879), .B(n4878), .Z(c[99]) );
  NANDN U6294 ( .A(n4367), .B(creg[9]), .Z(n4881) );
  NANDN U6295 ( .A(n7188), .B(o[9]), .Z(n4880) );
  NAND U6296 ( .A(n4881), .B(n4880), .Z(c[9]) );
  AND U6297 ( .A(m[0]), .B(n4368), .Z(n7187) );
  NANDN U6298 ( .A(n4368), .B(start_reg[0]), .Z(n5643) );
  NANDN U6299 ( .A(n5643), .B(creg[0]), .Z(n4882) );
  NANDN U6300 ( .A(n7187), .B(n4882), .Z(\modmult_1/xin[0] ) );
  OR U6301 ( .A(start_reg[0]), .B(n4368), .Z(start_in[0]) );
  NANDN U6302 ( .A(n5643), .B(creg[100]), .Z(n4883) );
  AND U6303 ( .A(m[100]), .B(n4368), .Z(n6785) );
  ANDN U6304 ( .B(n4883), .A(n6785), .Z(n4885) );
  NANDN U6305 ( .A(start_in[0]), .B(\modmult_1/xreg[100] ), .Z(n4884) );
  NAND U6306 ( .A(n4885), .B(n4884), .Z(\modmult_1/xin[100] ) );
  AND U6307 ( .A(m[101]), .B(n4368), .Z(n6781) );
  NANDN U6308 ( .A(start_in[0]), .B(\modmult_1/xreg[101] ), .Z(n4887) );
  NANDN U6309 ( .A(n5643), .B(creg[101]), .Z(n4886) );
  AND U6310 ( .A(n4887), .B(n4886), .Z(n4888) );
  NANDN U6311 ( .A(n6781), .B(n4888), .Z(\modmult_1/xin[101] ) );
  AND U6312 ( .A(m[102]), .B(n4368), .Z(n6777) );
  NANDN U6313 ( .A(start_in[0]), .B(\modmult_1/xreg[102] ), .Z(n4890) );
  NANDN U6314 ( .A(n5643), .B(creg[102]), .Z(n4889) );
  AND U6315 ( .A(n4890), .B(n4889), .Z(n4891) );
  NANDN U6316 ( .A(n6777), .B(n4891), .Z(\modmult_1/xin[102] ) );
  AND U6317 ( .A(m[103]), .B(n4368), .Z(n6773) );
  NANDN U6318 ( .A(start_in[0]), .B(\modmult_1/xreg[103] ), .Z(n4893) );
  NANDN U6319 ( .A(n5643), .B(creg[103]), .Z(n4892) );
  AND U6320 ( .A(n4893), .B(n4892), .Z(n4894) );
  NANDN U6321 ( .A(n6773), .B(n4894), .Z(\modmult_1/xin[103] ) );
  AND U6322 ( .A(m[104]), .B(n4368), .Z(n6769) );
  NANDN U6323 ( .A(start_in[0]), .B(\modmult_1/xreg[104] ), .Z(n4896) );
  NANDN U6324 ( .A(n5643), .B(creg[104]), .Z(n4895) );
  AND U6325 ( .A(n4896), .B(n4895), .Z(n4897) );
  NANDN U6326 ( .A(n6769), .B(n4897), .Z(\modmult_1/xin[104] ) );
  AND U6327 ( .A(m[105]), .B(n4368), .Z(n6765) );
  NANDN U6328 ( .A(start_in[0]), .B(\modmult_1/xreg[105] ), .Z(n4899) );
  NANDN U6329 ( .A(n5643), .B(creg[105]), .Z(n4898) );
  AND U6330 ( .A(n4899), .B(n4898), .Z(n4900) );
  NANDN U6331 ( .A(n6765), .B(n4900), .Z(\modmult_1/xin[105] ) );
  AND U6332 ( .A(m[106]), .B(n4368), .Z(n6761) );
  NANDN U6333 ( .A(start_in[0]), .B(\modmult_1/xreg[106] ), .Z(n4902) );
  NANDN U6334 ( .A(n5643), .B(creg[106]), .Z(n4901) );
  AND U6335 ( .A(n4902), .B(n4901), .Z(n4903) );
  NANDN U6336 ( .A(n6761), .B(n4903), .Z(\modmult_1/xin[106] ) );
  AND U6337 ( .A(m[107]), .B(n4368), .Z(n6757) );
  NANDN U6338 ( .A(start_in[0]), .B(\modmult_1/xreg[107] ), .Z(n4905) );
  NANDN U6339 ( .A(n5643), .B(creg[107]), .Z(n4904) );
  AND U6340 ( .A(n4905), .B(n4904), .Z(n4906) );
  NANDN U6341 ( .A(n6757), .B(n4906), .Z(\modmult_1/xin[107] ) );
  AND U6342 ( .A(m[108]), .B(n4368), .Z(n6753) );
  NANDN U6343 ( .A(start_in[0]), .B(\modmult_1/xreg[108] ), .Z(n4908) );
  NANDN U6344 ( .A(n5643), .B(creg[108]), .Z(n4907) );
  AND U6345 ( .A(n4908), .B(n4907), .Z(n4909) );
  NANDN U6346 ( .A(n6753), .B(n4909), .Z(\modmult_1/xin[108] ) );
  AND U6347 ( .A(m[109]), .B(n4368), .Z(n6749) );
  NANDN U6348 ( .A(start_in[0]), .B(\modmult_1/xreg[109] ), .Z(n4911) );
  NANDN U6349 ( .A(n5643), .B(creg[109]), .Z(n4910) );
  AND U6350 ( .A(n4911), .B(n4910), .Z(n4912) );
  NANDN U6351 ( .A(n6749), .B(n4912), .Z(\modmult_1/xin[109] ) );
  AND U6352 ( .A(m[10]), .B(n4368), .Z(n7145) );
  NANDN U6353 ( .A(start_in[0]), .B(\modmult_1/xreg[10] ), .Z(n4914) );
  NANDN U6354 ( .A(n5643), .B(creg[10]), .Z(n4913) );
  AND U6355 ( .A(n4914), .B(n4913), .Z(n4915) );
  NANDN U6356 ( .A(n7145), .B(n4915), .Z(\modmult_1/xin[10] ) );
  AND U6357 ( .A(m[110]), .B(n4368), .Z(n6745) );
  NANDN U6358 ( .A(start_in[0]), .B(\modmult_1/xreg[110] ), .Z(n4917) );
  NANDN U6359 ( .A(n5643), .B(creg[110]), .Z(n4916) );
  AND U6360 ( .A(n4917), .B(n4916), .Z(n4918) );
  NANDN U6361 ( .A(n6745), .B(n4918), .Z(\modmult_1/xin[110] ) );
  AND U6362 ( .A(m[111]), .B(n4368), .Z(n6741) );
  NANDN U6363 ( .A(start_in[0]), .B(\modmult_1/xreg[111] ), .Z(n4920) );
  NANDN U6364 ( .A(n5643), .B(creg[111]), .Z(n4919) );
  AND U6365 ( .A(n4920), .B(n4919), .Z(n4921) );
  NANDN U6366 ( .A(n6741), .B(n4921), .Z(\modmult_1/xin[111] ) );
  AND U6367 ( .A(m[112]), .B(n4368), .Z(n6737) );
  NANDN U6368 ( .A(start_in[0]), .B(\modmult_1/xreg[112] ), .Z(n4923) );
  NANDN U6369 ( .A(n5643), .B(creg[112]), .Z(n4922) );
  AND U6370 ( .A(n4923), .B(n4922), .Z(n4924) );
  NANDN U6371 ( .A(n6737), .B(n4924), .Z(\modmult_1/xin[112] ) );
  AND U6372 ( .A(m[113]), .B(n4368), .Z(n6733) );
  NANDN U6373 ( .A(start_in[0]), .B(\modmult_1/xreg[113] ), .Z(n4926) );
  NANDN U6374 ( .A(n5643), .B(creg[113]), .Z(n4925) );
  AND U6375 ( .A(n4926), .B(n4925), .Z(n4927) );
  NANDN U6376 ( .A(n6733), .B(n4927), .Z(\modmult_1/xin[113] ) );
  AND U6377 ( .A(m[114]), .B(n4368), .Z(n6729) );
  NANDN U6378 ( .A(start_in[0]), .B(\modmult_1/xreg[114] ), .Z(n4929) );
  NANDN U6379 ( .A(n5643), .B(creg[114]), .Z(n4928) );
  AND U6380 ( .A(n4929), .B(n4928), .Z(n4930) );
  NANDN U6381 ( .A(n6729), .B(n4930), .Z(\modmult_1/xin[114] ) );
  AND U6382 ( .A(m[115]), .B(n4368), .Z(n6725) );
  NANDN U6383 ( .A(start_in[0]), .B(\modmult_1/xreg[115] ), .Z(n4932) );
  NANDN U6384 ( .A(n5643), .B(creg[115]), .Z(n4931) );
  AND U6385 ( .A(n4932), .B(n4931), .Z(n4933) );
  NANDN U6386 ( .A(n6725), .B(n4933), .Z(\modmult_1/xin[115] ) );
  AND U6387 ( .A(m[116]), .B(n4368), .Z(n6721) );
  NANDN U6388 ( .A(start_in[0]), .B(\modmult_1/xreg[116] ), .Z(n4935) );
  NANDN U6389 ( .A(n5643), .B(creg[116]), .Z(n4934) );
  AND U6390 ( .A(n4935), .B(n4934), .Z(n4936) );
  NANDN U6391 ( .A(n6721), .B(n4936), .Z(\modmult_1/xin[116] ) );
  AND U6392 ( .A(m[117]), .B(n4368), .Z(n6717) );
  NANDN U6393 ( .A(start_in[0]), .B(\modmult_1/xreg[117] ), .Z(n4938) );
  NANDN U6394 ( .A(n5643), .B(creg[117]), .Z(n4937) );
  AND U6395 ( .A(n4938), .B(n4937), .Z(n4939) );
  NANDN U6396 ( .A(n6717), .B(n4939), .Z(\modmult_1/xin[117] ) );
  AND U6397 ( .A(m[118]), .B(n4368), .Z(n6713) );
  NANDN U6398 ( .A(start_in[0]), .B(\modmult_1/xreg[118] ), .Z(n4941) );
  NANDN U6399 ( .A(n5643), .B(creg[118]), .Z(n4940) );
  AND U6400 ( .A(n4941), .B(n4940), .Z(n4942) );
  NANDN U6401 ( .A(n6713), .B(n4942), .Z(\modmult_1/xin[118] ) );
  AND U6402 ( .A(m[119]), .B(n4368), .Z(n6709) );
  NANDN U6403 ( .A(start_in[0]), .B(\modmult_1/xreg[119] ), .Z(n4944) );
  NANDN U6404 ( .A(n5643), .B(creg[119]), .Z(n4943) );
  AND U6405 ( .A(n4944), .B(n4943), .Z(n4945) );
  NANDN U6406 ( .A(n6709), .B(n4945), .Z(\modmult_1/xin[119] ) );
  AND U6407 ( .A(m[11]), .B(n4368), .Z(n7141) );
  NANDN U6408 ( .A(start_in[0]), .B(\modmult_1/xreg[11] ), .Z(n4947) );
  NANDN U6409 ( .A(n5643), .B(creg[11]), .Z(n4946) );
  AND U6410 ( .A(n4947), .B(n4946), .Z(n4948) );
  NANDN U6411 ( .A(n7141), .B(n4948), .Z(\modmult_1/xin[11] ) );
  AND U6412 ( .A(m[120]), .B(n4368), .Z(n6705) );
  NANDN U6413 ( .A(start_in[0]), .B(\modmult_1/xreg[120] ), .Z(n4950) );
  NANDN U6414 ( .A(n5643), .B(creg[120]), .Z(n4949) );
  AND U6415 ( .A(n4950), .B(n4949), .Z(n4951) );
  NANDN U6416 ( .A(n6705), .B(n4951), .Z(\modmult_1/xin[120] ) );
  AND U6417 ( .A(m[121]), .B(n4368), .Z(n6701) );
  NANDN U6418 ( .A(start_in[0]), .B(\modmult_1/xreg[121] ), .Z(n4953) );
  NANDN U6419 ( .A(n5643), .B(creg[121]), .Z(n4952) );
  AND U6420 ( .A(n4953), .B(n4952), .Z(n4954) );
  NANDN U6421 ( .A(n6701), .B(n4954), .Z(\modmult_1/xin[121] ) );
  AND U6422 ( .A(m[122]), .B(n4368), .Z(n6697) );
  NANDN U6423 ( .A(start_in[0]), .B(\modmult_1/xreg[122] ), .Z(n4956) );
  NANDN U6424 ( .A(n5643), .B(creg[122]), .Z(n4955) );
  AND U6425 ( .A(n4956), .B(n4955), .Z(n4957) );
  NANDN U6426 ( .A(n6697), .B(n4957), .Z(\modmult_1/xin[122] ) );
  AND U6427 ( .A(m[123]), .B(n4368), .Z(n6693) );
  NANDN U6428 ( .A(start_in[0]), .B(\modmult_1/xreg[123] ), .Z(n4959) );
  NANDN U6429 ( .A(n5643), .B(creg[123]), .Z(n4958) );
  AND U6430 ( .A(n4959), .B(n4958), .Z(n4960) );
  NANDN U6431 ( .A(n6693), .B(n4960), .Z(\modmult_1/xin[123] ) );
  AND U6432 ( .A(m[124]), .B(n4368), .Z(n6689) );
  NANDN U6433 ( .A(start_in[0]), .B(\modmult_1/xreg[124] ), .Z(n4962) );
  NANDN U6434 ( .A(n5643), .B(creg[124]), .Z(n4961) );
  AND U6435 ( .A(n4962), .B(n4961), .Z(n4963) );
  NANDN U6436 ( .A(n6689), .B(n4963), .Z(\modmult_1/xin[124] ) );
  AND U6437 ( .A(m[125]), .B(n4368), .Z(n6685) );
  NANDN U6438 ( .A(start_in[0]), .B(\modmult_1/xreg[125] ), .Z(n4965) );
  NANDN U6439 ( .A(n5643), .B(creg[125]), .Z(n4964) );
  AND U6440 ( .A(n4965), .B(n4964), .Z(n4966) );
  NANDN U6441 ( .A(n6685), .B(n4966), .Z(\modmult_1/xin[125] ) );
  AND U6442 ( .A(m[126]), .B(n4368), .Z(n6681) );
  NANDN U6443 ( .A(start_in[0]), .B(\modmult_1/xreg[126] ), .Z(n4968) );
  NANDN U6444 ( .A(n5643), .B(creg[126]), .Z(n4967) );
  AND U6445 ( .A(n4968), .B(n4967), .Z(n4969) );
  NANDN U6446 ( .A(n6681), .B(n4969), .Z(\modmult_1/xin[126] ) );
  AND U6447 ( .A(m[127]), .B(n4368), .Z(n6677) );
  NANDN U6448 ( .A(start_in[0]), .B(\modmult_1/xreg[127] ), .Z(n4971) );
  NANDN U6449 ( .A(n5643), .B(creg[127]), .Z(n4970) );
  AND U6450 ( .A(n4971), .B(n4970), .Z(n4972) );
  NANDN U6451 ( .A(n6677), .B(n4972), .Z(\modmult_1/xin[127] ) );
  AND U6452 ( .A(m[128]), .B(n4368), .Z(n6673) );
  NANDN U6453 ( .A(start_in[0]), .B(\modmult_1/xreg[128] ), .Z(n4974) );
  NANDN U6454 ( .A(n5643), .B(creg[128]), .Z(n4973) );
  AND U6455 ( .A(n4974), .B(n4973), .Z(n4975) );
  NANDN U6456 ( .A(n6673), .B(n4975), .Z(\modmult_1/xin[128] ) );
  AND U6457 ( .A(m[129]), .B(n4368), .Z(n6669) );
  NANDN U6458 ( .A(start_in[0]), .B(\modmult_1/xreg[129] ), .Z(n4977) );
  NANDN U6459 ( .A(n5643), .B(creg[129]), .Z(n4976) );
  AND U6460 ( .A(n4977), .B(n4976), .Z(n4978) );
  NANDN U6461 ( .A(n6669), .B(n4978), .Z(\modmult_1/xin[129] ) );
  AND U6462 ( .A(m[12]), .B(n4368), .Z(n7137) );
  NANDN U6463 ( .A(start_in[0]), .B(\modmult_1/xreg[12] ), .Z(n4980) );
  NANDN U6464 ( .A(n5643), .B(creg[12]), .Z(n4979) );
  AND U6465 ( .A(n4980), .B(n4979), .Z(n4981) );
  NANDN U6466 ( .A(n7137), .B(n4981), .Z(\modmult_1/xin[12] ) );
  AND U6467 ( .A(m[130]), .B(n4368), .Z(n6665) );
  NANDN U6468 ( .A(start_in[0]), .B(\modmult_1/xreg[130] ), .Z(n4983) );
  NANDN U6469 ( .A(n5643), .B(creg[130]), .Z(n4982) );
  AND U6470 ( .A(n4983), .B(n4982), .Z(n4984) );
  NANDN U6471 ( .A(n6665), .B(n4984), .Z(\modmult_1/xin[130] ) );
  AND U6472 ( .A(m[131]), .B(n4368), .Z(n6661) );
  NANDN U6473 ( .A(start_in[0]), .B(\modmult_1/xreg[131] ), .Z(n4986) );
  NANDN U6474 ( .A(n5643), .B(creg[131]), .Z(n4985) );
  AND U6475 ( .A(n4986), .B(n4985), .Z(n4987) );
  NANDN U6476 ( .A(n6661), .B(n4987), .Z(\modmult_1/xin[131] ) );
  AND U6477 ( .A(m[132]), .B(n4368), .Z(n6657) );
  NANDN U6478 ( .A(start_in[0]), .B(\modmult_1/xreg[132] ), .Z(n4989) );
  NANDN U6479 ( .A(n5643), .B(creg[132]), .Z(n4988) );
  AND U6480 ( .A(n4989), .B(n4988), .Z(n4990) );
  NANDN U6481 ( .A(n6657), .B(n4990), .Z(\modmult_1/xin[132] ) );
  AND U6482 ( .A(m[133]), .B(n4368), .Z(n6653) );
  NANDN U6483 ( .A(start_in[0]), .B(\modmult_1/xreg[133] ), .Z(n4992) );
  NANDN U6484 ( .A(n5643), .B(creg[133]), .Z(n4991) );
  AND U6485 ( .A(n4992), .B(n4991), .Z(n4993) );
  NANDN U6486 ( .A(n6653), .B(n4993), .Z(\modmult_1/xin[133] ) );
  AND U6487 ( .A(m[134]), .B(n4368), .Z(n6649) );
  NANDN U6488 ( .A(start_in[0]), .B(\modmult_1/xreg[134] ), .Z(n4995) );
  NANDN U6489 ( .A(n5643), .B(creg[134]), .Z(n4994) );
  AND U6490 ( .A(n4995), .B(n4994), .Z(n4996) );
  NANDN U6491 ( .A(n6649), .B(n4996), .Z(\modmult_1/xin[134] ) );
  AND U6492 ( .A(m[135]), .B(n4368), .Z(n6645) );
  NANDN U6493 ( .A(start_in[0]), .B(\modmult_1/xreg[135] ), .Z(n4998) );
  NANDN U6494 ( .A(n5643), .B(creg[135]), .Z(n4997) );
  AND U6495 ( .A(n4998), .B(n4997), .Z(n4999) );
  NANDN U6496 ( .A(n6645), .B(n4999), .Z(\modmult_1/xin[135] ) );
  AND U6497 ( .A(m[136]), .B(n4368), .Z(n6641) );
  NANDN U6498 ( .A(start_in[0]), .B(\modmult_1/xreg[136] ), .Z(n5001) );
  NANDN U6499 ( .A(n5643), .B(creg[136]), .Z(n5000) );
  AND U6500 ( .A(n5001), .B(n5000), .Z(n5002) );
  NANDN U6501 ( .A(n6641), .B(n5002), .Z(\modmult_1/xin[136] ) );
  AND U6502 ( .A(m[137]), .B(n4368), .Z(n6637) );
  NANDN U6503 ( .A(start_in[0]), .B(\modmult_1/xreg[137] ), .Z(n5004) );
  NANDN U6504 ( .A(n5643), .B(creg[137]), .Z(n5003) );
  AND U6505 ( .A(n5004), .B(n5003), .Z(n5005) );
  NANDN U6506 ( .A(n6637), .B(n5005), .Z(\modmult_1/xin[137] ) );
  AND U6507 ( .A(m[138]), .B(n4368), .Z(n6633) );
  NANDN U6508 ( .A(start_in[0]), .B(\modmult_1/xreg[138] ), .Z(n5007) );
  NANDN U6509 ( .A(n5643), .B(creg[138]), .Z(n5006) );
  AND U6510 ( .A(n5007), .B(n5006), .Z(n5008) );
  NANDN U6511 ( .A(n6633), .B(n5008), .Z(\modmult_1/xin[138] ) );
  AND U6512 ( .A(m[139]), .B(n4368), .Z(n6629) );
  NANDN U6513 ( .A(start_in[0]), .B(\modmult_1/xreg[139] ), .Z(n5010) );
  NANDN U6514 ( .A(n5643), .B(creg[139]), .Z(n5009) );
  AND U6515 ( .A(n5010), .B(n5009), .Z(n5011) );
  NANDN U6516 ( .A(n6629), .B(n5011), .Z(\modmult_1/xin[139] ) );
  AND U6517 ( .A(m[13]), .B(n4368), .Z(n7133) );
  NANDN U6518 ( .A(start_in[0]), .B(\modmult_1/xreg[13] ), .Z(n5013) );
  NANDN U6519 ( .A(n5643), .B(creg[13]), .Z(n5012) );
  AND U6520 ( .A(n5013), .B(n5012), .Z(n5014) );
  NANDN U6521 ( .A(n7133), .B(n5014), .Z(\modmult_1/xin[13] ) );
  AND U6522 ( .A(m[140]), .B(n4368), .Z(n6625) );
  NANDN U6523 ( .A(start_in[0]), .B(\modmult_1/xreg[140] ), .Z(n5016) );
  NANDN U6524 ( .A(n5643), .B(creg[140]), .Z(n5015) );
  AND U6525 ( .A(n5016), .B(n5015), .Z(n5017) );
  NANDN U6526 ( .A(n6625), .B(n5017), .Z(\modmult_1/xin[140] ) );
  AND U6527 ( .A(m[141]), .B(n4368), .Z(n6621) );
  NANDN U6528 ( .A(start_in[0]), .B(\modmult_1/xreg[141] ), .Z(n5019) );
  NANDN U6529 ( .A(n5643), .B(creg[141]), .Z(n5018) );
  AND U6530 ( .A(n5019), .B(n5018), .Z(n5020) );
  NANDN U6531 ( .A(n6621), .B(n5020), .Z(\modmult_1/xin[141] ) );
  AND U6532 ( .A(m[142]), .B(n4368), .Z(n6617) );
  NANDN U6533 ( .A(start_in[0]), .B(\modmult_1/xreg[142] ), .Z(n5022) );
  NANDN U6534 ( .A(n5643), .B(creg[142]), .Z(n5021) );
  AND U6535 ( .A(n5022), .B(n5021), .Z(n5023) );
  NANDN U6536 ( .A(n6617), .B(n5023), .Z(\modmult_1/xin[142] ) );
  AND U6537 ( .A(m[143]), .B(n4368), .Z(n6613) );
  NANDN U6538 ( .A(start_in[0]), .B(\modmult_1/xreg[143] ), .Z(n5025) );
  NANDN U6539 ( .A(n5643), .B(creg[143]), .Z(n5024) );
  AND U6540 ( .A(n5025), .B(n5024), .Z(n5026) );
  NANDN U6541 ( .A(n6613), .B(n5026), .Z(\modmult_1/xin[143] ) );
  AND U6542 ( .A(m[144]), .B(n4368), .Z(n6609) );
  NANDN U6543 ( .A(start_in[0]), .B(\modmult_1/xreg[144] ), .Z(n5028) );
  NANDN U6544 ( .A(n5643), .B(creg[144]), .Z(n5027) );
  AND U6545 ( .A(n5028), .B(n5027), .Z(n5029) );
  NANDN U6546 ( .A(n6609), .B(n5029), .Z(\modmult_1/xin[144] ) );
  AND U6547 ( .A(m[145]), .B(n4368), .Z(n6605) );
  NANDN U6548 ( .A(start_in[0]), .B(\modmult_1/xreg[145] ), .Z(n5031) );
  NANDN U6549 ( .A(n5643), .B(creg[145]), .Z(n5030) );
  AND U6550 ( .A(n5031), .B(n5030), .Z(n5032) );
  NANDN U6551 ( .A(n6605), .B(n5032), .Z(\modmult_1/xin[145] ) );
  AND U6552 ( .A(m[146]), .B(n4368), .Z(n6601) );
  NANDN U6553 ( .A(start_in[0]), .B(\modmult_1/xreg[146] ), .Z(n5034) );
  NANDN U6554 ( .A(n5643), .B(creg[146]), .Z(n5033) );
  AND U6555 ( .A(n5034), .B(n5033), .Z(n5035) );
  NANDN U6556 ( .A(n6601), .B(n5035), .Z(\modmult_1/xin[146] ) );
  AND U6557 ( .A(m[147]), .B(n4368), .Z(n6597) );
  NANDN U6558 ( .A(start_in[0]), .B(\modmult_1/xreg[147] ), .Z(n5037) );
  NANDN U6559 ( .A(n5643), .B(creg[147]), .Z(n5036) );
  AND U6560 ( .A(n5037), .B(n5036), .Z(n5038) );
  NANDN U6561 ( .A(n6597), .B(n5038), .Z(\modmult_1/xin[147] ) );
  AND U6562 ( .A(m[148]), .B(n4368), .Z(n6593) );
  NANDN U6563 ( .A(start_in[0]), .B(\modmult_1/xreg[148] ), .Z(n5040) );
  NANDN U6564 ( .A(n5643), .B(creg[148]), .Z(n5039) );
  AND U6565 ( .A(n5040), .B(n5039), .Z(n5041) );
  NANDN U6566 ( .A(n6593), .B(n5041), .Z(\modmult_1/xin[148] ) );
  AND U6567 ( .A(m[149]), .B(n4368), .Z(n6589) );
  NANDN U6568 ( .A(start_in[0]), .B(\modmult_1/xreg[149] ), .Z(n5043) );
  NANDN U6569 ( .A(n5643), .B(creg[149]), .Z(n5042) );
  AND U6570 ( .A(n5043), .B(n5042), .Z(n5044) );
  NANDN U6571 ( .A(n6589), .B(n5044), .Z(\modmult_1/xin[149] ) );
  AND U6572 ( .A(m[14]), .B(n4368), .Z(n7129) );
  NANDN U6573 ( .A(start_in[0]), .B(\modmult_1/xreg[14] ), .Z(n5046) );
  NANDN U6574 ( .A(n5643), .B(creg[14]), .Z(n5045) );
  AND U6575 ( .A(n5046), .B(n5045), .Z(n5047) );
  NANDN U6576 ( .A(n7129), .B(n5047), .Z(\modmult_1/xin[14] ) );
  AND U6577 ( .A(m[150]), .B(n4368), .Z(n6585) );
  NANDN U6578 ( .A(start_in[0]), .B(\modmult_1/xreg[150] ), .Z(n5049) );
  NANDN U6579 ( .A(n5643), .B(creg[150]), .Z(n5048) );
  AND U6580 ( .A(n5049), .B(n5048), .Z(n5050) );
  NANDN U6581 ( .A(n6585), .B(n5050), .Z(\modmult_1/xin[150] ) );
  AND U6582 ( .A(m[151]), .B(n4368), .Z(n6581) );
  NANDN U6583 ( .A(start_in[0]), .B(\modmult_1/xreg[151] ), .Z(n5052) );
  NANDN U6584 ( .A(n5643), .B(creg[151]), .Z(n5051) );
  AND U6585 ( .A(n5052), .B(n5051), .Z(n5053) );
  NANDN U6586 ( .A(n6581), .B(n5053), .Z(\modmult_1/xin[151] ) );
  AND U6587 ( .A(m[152]), .B(n4368), .Z(n6577) );
  NANDN U6588 ( .A(start_in[0]), .B(\modmult_1/xreg[152] ), .Z(n5055) );
  NANDN U6589 ( .A(n5643), .B(creg[152]), .Z(n5054) );
  AND U6590 ( .A(n5055), .B(n5054), .Z(n5056) );
  NANDN U6591 ( .A(n6577), .B(n5056), .Z(\modmult_1/xin[152] ) );
  AND U6592 ( .A(m[153]), .B(n4368), .Z(n6573) );
  NANDN U6593 ( .A(start_in[0]), .B(\modmult_1/xreg[153] ), .Z(n5058) );
  NANDN U6594 ( .A(n5643), .B(creg[153]), .Z(n5057) );
  AND U6595 ( .A(n5058), .B(n5057), .Z(n5059) );
  NANDN U6596 ( .A(n6573), .B(n5059), .Z(\modmult_1/xin[153] ) );
  AND U6597 ( .A(m[154]), .B(n4368), .Z(n6569) );
  NANDN U6598 ( .A(start_in[0]), .B(\modmult_1/xreg[154] ), .Z(n5061) );
  NANDN U6599 ( .A(n5643), .B(creg[154]), .Z(n5060) );
  AND U6600 ( .A(n5061), .B(n5060), .Z(n5062) );
  NANDN U6601 ( .A(n6569), .B(n5062), .Z(\modmult_1/xin[154] ) );
  AND U6602 ( .A(m[155]), .B(n4368), .Z(n6565) );
  NANDN U6603 ( .A(start_in[0]), .B(\modmult_1/xreg[155] ), .Z(n5064) );
  NANDN U6604 ( .A(n5643), .B(creg[155]), .Z(n5063) );
  AND U6605 ( .A(n5064), .B(n5063), .Z(n5065) );
  NANDN U6606 ( .A(n6565), .B(n5065), .Z(\modmult_1/xin[155] ) );
  AND U6607 ( .A(m[156]), .B(n4368), .Z(n6561) );
  NANDN U6608 ( .A(start_in[0]), .B(\modmult_1/xreg[156] ), .Z(n5067) );
  NANDN U6609 ( .A(n5643), .B(creg[156]), .Z(n5066) );
  AND U6610 ( .A(n5067), .B(n5066), .Z(n5068) );
  NANDN U6611 ( .A(n6561), .B(n5068), .Z(\modmult_1/xin[156] ) );
  AND U6612 ( .A(m[157]), .B(n4368), .Z(n6557) );
  NANDN U6613 ( .A(start_in[0]), .B(\modmult_1/xreg[157] ), .Z(n5070) );
  NANDN U6614 ( .A(n5643), .B(creg[157]), .Z(n5069) );
  AND U6615 ( .A(n5070), .B(n5069), .Z(n5071) );
  NANDN U6616 ( .A(n6557), .B(n5071), .Z(\modmult_1/xin[157] ) );
  AND U6617 ( .A(m[158]), .B(n4368), .Z(n6553) );
  NANDN U6618 ( .A(start_in[0]), .B(\modmult_1/xreg[158] ), .Z(n5073) );
  NANDN U6619 ( .A(n5643), .B(creg[158]), .Z(n5072) );
  AND U6620 ( .A(n5073), .B(n5072), .Z(n5074) );
  NANDN U6621 ( .A(n6553), .B(n5074), .Z(\modmult_1/xin[158] ) );
  AND U6622 ( .A(m[159]), .B(n4368), .Z(n6549) );
  NANDN U6623 ( .A(start_in[0]), .B(\modmult_1/xreg[159] ), .Z(n5076) );
  NANDN U6624 ( .A(n5643), .B(creg[159]), .Z(n5075) );
  AND U6625 ( .A(n5076), .B(n5075), .Z(n5077) );
  NANDN U6626 ( .A(n6549), .B(n5077), .Z(\modmult_1/xin[159] ) );
  AND U6627 ( .A(m[15]), .B(n4368), .Z(n7125) );
  NANDN U6628 ( .A(start_in[0]), .B(\modmult_1/xreg[15] ), .Z(n5079) );
  NANDN U6629 ( .A(n5643), .B(creg[15]), .Z(n5078) );
  AND U6630 ( .A(n5079), .B(n5078), .Z(n5080) );
  NANDN U6631 ( .A(n7125), .B(n5080), .Z(\modmult_1/xin[15] ) );
  AND U6632 ( .A(m[160]), .B(n4368), .Z(n6545) );
  NANDN U6633 ( .A(start_in[0]), .B(\modmult_1/xreg[160] ), .Z(n5082) );
  NANDN U6634 ( .A(n5643), .B(creg[160]), .Z(n5081) );
  AND U6635 ( .A(n5082), .B(n5081), .Z(n5083) );
  NANDN U6636 ( .A(n6545), .B(n5083), .Z(\modmult_1/xin[160] ) );
  AND U6637 ( .A(m[161]), .B(n4368), .Z(n6541) );
  NANDN U6638 ( .A(start_in[0]), .B(\modmult_1/xreg[161] ), .Z(n5085) );
  NANDN U6639 ( .A(n5643), .B(creg[161]), .Z(n5084) );
  AND U6640 ( .A(n5085), .B(n5084), .Z(n5086) );
  NANDN U6641 ( .A(n6541), .B(n5086), .Z(\modmult_1/xin[161] ) );
  AND U6642 ( .A(m[162]), .B(n4368), .Z(n6537) );
  NANDN U6643 ( .A(start_in[0]), .B(\modmult_1/xreg[162] ), .Z(n5088) );
  NANDN U6644 ( .A(n5643), .B(creg[162]), .Z(n5087) );
  AND U6645 ( .A(n5088), .B(n5087), .Z(n5089) );
  NANDN U6646 ( .A(n6537), .B(n5089), .Z(\modmult_1/xin[162] ) );
  AND U6647 ( .A(m[163]), .B(n4368), .Z(n6533) );
  NANDN U6648 ( .A(start_in[0]), .B(\modmult_1/xreg[163] ), .Z(n5091) );
  NANDN U6649 ( .A(n5643), .B(creg[163]), .Z(n5090) );
  AND U6650 ( .A(n5091), .B(n5090), .Z(n5092) );
  NANDN U6651 ( .A(n6533), .B(n5092), .Z(\modmult_1/xin[163] ) );
  AND U6652 ( .A(m[164]), .B(n4368), .Z(n6529) );
  NANDN U6653 ( .A(start_in[0]), .B(\modmult_1/xreg[164] ), .Z(n5094) );
  NANDN U6654 ( .A(n5643), .B(creg[164]), .Z(n5093) );
  AND U6655 ( .A(n5094), .B(n5093), .Z(n5095) );
  NANDN U6656 ( .A(n6529), .B(n5095), .Z(\modmult_1/xin[164] ) );
  AND U6657 ( .A(m[165]), .B(n4368), .Z(n6525) );
  NANDN U6658 ( .A(start_in[0]), .B(\modmult_1/xreg[165] ), .Z(n5097) );
  NANDN U6659 ( .A(n5643), .B(creg[165]), .Z(n5096) );
  AND U6660 ( .A(n5097), .B(n5096), .Z(n5098) );
  NANDN U6661 ( .A(n6525), .B(n5098), .Z(\modmult_1/xin[165] ) );
  AND U6662 ( .A(m[166]), .B(n4368), .Z(n6521) );
  NANDN U6663 ( .A(start_in[0]), .B(\modmult_1/xreg[166] ), .Z(n5100) );
  NANDN U6664 ( .A(n5643), .B(creg[166]), .Z(n5099) );
  AND U6665 ( .A(n5100), .B(n5099), .Z(n5101) );
  NANDN U6666 ( .A(n6521), .B(n5101), .Z(\modmult_1/xin[166] ) );
  AND U6667 ( .A(m[167]), .B(n4368), .Z(n6517) );
  NANDN U6668 ( .A(start_in[0]), .B(\modmult_1/xreg[167] ), .Z(n5103) );
  NANDN U6669 ( .A(n5643), .B(creg[167]), .Z(n5102) );
  AND U6670 ( .A(n5103), .B(n5102), .Z(n5104) );
  NANDN U6671 ( .A(n6517), .B(n5104), .Z(\modmult_1/xin[167] ) );
  AND U6672 ( .A(m[168]), .B(n4368), .Z(n6513) );
  NANDN U6673 ( .A(start_in[0]), .B(\modmult_1/xreg[168] ), .Z(n5106) );
  NANDN U6674 ( .A(n5643), .B(creg[168]), .Z(n5105) );
  AND U6675 ( .A(n5106), .B(n5105), .Z(n5107) );
  NANDN U6676 ( .A(n6513), .B(n5107), .Z(\modmult_1/xin[168] ) );
  AND U6677 ( .A(m[169]), .B(n4368), .Z(n6509) );
  NANDN U6678 ( .A(start_in[0]), .B(\modmult_1/xreg[169] ), .Z(n5109) );
  NANDN U6679 ( .A(n5643), .B(creg[169]), .Z(n5108) );
  AND U6680 ( .A(n5109), .B(n5108), .Z(n5110) );
  NANDN U6681 ( .A(n6509), .B(n5110), .Z(\modmult_1/xin[169] ) );
  AND U6682 ( .A(m[16]), .B(n4368), .Z(n7121) );
  NANDN U6683 ( .A(start_in[0]), .B(\modmult_1/xreg[16] ), .Z(n5112) );
  NANDN U6684 ( .A(n5643), .B(creg[16]), .Z(n5111) );
  AND U6685 ( .A(n5112), .B(n5111), .Z(n5113) );
  NANDN U6686 ( .A(n7121), .B(n5113), .Z(\modmult_1/xin[16] ) );
  AND U6687 ( .A(m[170]), .B(n4368), .Z(n6505) );
  NANDN U6688 ( .A(start_in[0]), .B(\modmult_1/xreg[170] ), .Z(n5115) );
  NANDN U6689 ( .A(n5643), .B(creg[170]), .Z(n5114) );
  AND U6690 ( .A(n5115), .B(n5114), .Z(n5116) );
  NANDN U6691 ( .A(n6505), .B(n5116), .Z(\modmult_1/xin[170] ) );
  AND U6692 ( .A(m[171]), .B(n4368), .Z(n6501) );
  NANDN U6693 ( .A(start_in[0]), .B(\modmult_1/xreg[171] ), .Z(n5118) );
  NANDN U6694 ( .A(n5643), .B(creg[171]), .Z(n5117) );
  AND U6695 ( .A(n5118), .B(n5117), .Z(n5119) );
  NANDN U6696 ( .A(n6501), .B(n5119), .Z(\modmult_1/xin[171] ) );
  AND U6697 ( .A(m[172]), .B(n4368), .Z(n6497) );
  NANDN U6698 ( .A(start_in[0]), .B(\modmult_1/xreg[172] ), .Z(n5121) );
  NANDN U6699 ( .A(n5643), .B(creg[172]), .Z(n5120) );
  AND U6700 ( .A(n5121), .B(n5120), .Z(n5122) );
  NANDN U6701 ( .A(n6497), .B(n5122), .Z(\modmult_1/xin[172] ) );
  AND U6702 ( .A(m[173]), .B(n4368), .Z(n6493) );
  NANDN U6703 ( .A(start_in[0]), .B(\modmult_1/xreg[173] ), .Z(n5124) );
  NANDN U6704 ( .A(n5643), .B(creg[173]), .Z(n5123) );
  AND U6705 ( .A(n5124), .B(n5123), .Z(n5125) );
  NANDN U6706 ( .A(n6493), .B(n5125), .Z(\modmult_1/xin[173] ) );
  AND U6707 ( .A(m[174]), .B(n4368), .Z(n6489) );
  NANDN U6708 ( .A(start_in[0]), .B(\modmult_1/xreg[174] ), .Z(n5127) );
  NANDN U6709 ( .A(n5643), .B(creg[174]), .Z(n5126) );
  AND U6710 ( .A(n5127), .B(n5126), .Z(n5128) );
  NANDN U6711 ( .A(n6489), .B(n5128), .Z(\modmult_1/xin[174] ) );
  AND U6712 ( .A(m[175]), .B(n4368), .Z(n6485) );
  NANDN U6713 ( .A(start_in[0]), .B(\modmult_1/xreg[175] ), .Z(n5130) );
  NANDN U6714 ( .A(n5643), .B(creg[175]), .Z(n5129) );
  AND U6715 ( .A(n5130), .B(n5129), .Z(n5131) );
  NANDN U6716 ( .A(n6485), .B(n5131), .Z(\modmult_1/xin[175] ) );
  AND U6717 ( .A(m[176]), .B(n4368), .Z(n6481) );
  NANDN U6718 ( .A(start_in[0]), .B(\modmult_1/xreg[176] ), .Z(n5133) );
  NANDN U6719 ( .A(n5643), .B(creg[176]), .Z(n5132) );
  AND U6720 ( .A(n5133), .B(n5132), .Z(n5134) );
  NANDN U6721 ( .A(n6481), .B(n5134), .Z(\modmult_1/xin[176] ) );
  AND U6722 ( .A(m[177]), .B(n4368), .Z(n6477) );
  NANDN U6723 ( .A(start_in[0]), .B(\modmult_1/xreg[177] ), .Z(n5136) );
  NANDN U6724 ( .A(n5643), .B(creg[177]), .Z(n5135) );
  AND U6725 ( .A(n5136), .B(n5135), .Z(n5137) );
  NANDN U6726 ( .A(n6477), .B(n5137), .Z(\modmult_1/xin[177] ) );
  AND U6727 ( .A(m[178]), .B(n4368), .Z(n6473) );
  NANDN U6728 ( .A(start_in[0]), .B(\modmult_1/xreg[178] ), .Z(n5139) );
  NANDN U6729 ( .A(n5643), .B(creg[178]), .Z(n5138) );
  AND U6730 ( .A(n5139), .B(n5138), .Z(n5140) );
  NANDN U6731 ( .A(n6473), .B(n5140), .Z(\modmult_1/xin[178] ) );
  AND U6732 ( .A(m[179]), .B(n4368), .Z(n6469) );
  NANDN U6733 ( .A(start_in[0]), .B(\modmult_1/xreg[179] ), .Z(n5142) );
  NANDN U6734 ( .A(n5643), .B(creg[179]), .Z(n5141) );
  AND U6735 ( .A(n5142), .B(n5141), .Z(n5143) );
  NANDN U6736 ( .A(n6469), .B(n5143), .Z(\modmult_1/xin[179] ) );
  AND U6737 ( .A(m[17]), .B(n4368), .Z(n7117) );
  NANDN U6738 ( .A(start_in[0]), .B(\modmult_1/xreg[17] ), .Z(n5145) );
  NANDN U6739 ( .A(n5643), .B(creg[17]), .Z(n5144) );
  AND U6740 ( .A(n5145), .B(n5144), .Z(n5146) );
  NANDN U6741 ( .A(n7117), .B(n5146), .Z(\modmult_1/xin[17] ) );
  AND U6742 ( .A(m[180]), .B(n4368), .Z(n6465) );
  NANDN U6743 ( .A(start_in[0]), .B(\modmult_1/xreg[180] ), .Z(n5148) );
  NANDN U6744 ( .A(n5643), .B(creg[180]), .Z(n5147) );
  AND U6745 ( .A(n5148), .B(n5147), .Z(n5149) );
  NANDN U6746 ( .A(n6465), .B(n5149), .Z(\modmult_1/xin[180] ) );
  AND U6747 ( .A(m[181]), .B(n4368), .Z(n6461) );
  NANDN U6748 ( .A(start_in[0]), .B(\modmult_1/xreg[181] ), .Z(n5151) );
  NANDN U6749 ( .A(n5643), .B(creg[181]), .Z(n5150) );
  AND U6750 ( .A(n5151), .B(n5150), .Z(n5152) );
  NANDN U6751 ( .A(n6461), .B(n5152), .Z(\modmult_1/xin[181] ) );
  AND U6752 ( .A(m[182]), .B(n4368), .Z(n6457) );
  NANDN U6753 ( .A(start_in[0]), .B(\modmult_1/xreg[182] ), .Z(n5154) );
  NANDN U6754 ( .A(n5643), .B(creg[182]), .Z(n5153) );
  AND U6755 ( .A(n5154), .B(n5153), .Z(n5155) );
  NANDN U6756 ( .A(n6457), .B(n5155), .Z(\modmult_1/xin[182] ) );
  AND U6757 ( .A(m[183]), .B(n4368), .Z(n6453) );
  NANDN U6758 ( .A(start_in[0]), .B(\modmult_1/xreg[183] ), .Z(n5157) );
  NANDN U6759 ( .A(n5643), .B(creg[183]), .Z(n5156) );
  AND U6760 ( .A(n5157), .B(n5156), .Z(n5158) );
  NANDN U6761 ( .A(n6453), .B(n5158), .Z(\modmult_1/xin[183] ) );
  AND U6762 ( .A(m[184]), .B(n4368), .Z(n6449) );
  NANDN U6763 ( .A(start_in[0]), .B(\modmult_1/xreg[184] ), .Z(n5160) );
  NANDN U6764 ( .A(n5643), .B(creg[184]), .Z(n5159) );
  AND U6765 ( .A(n5160), .B(n5159), .Z(n5161) );
  NANDN U6766 ( .A(n6449), .B(n5161), .Z(\modmult_1/xin[184] ) );
  AND U6767 ( .A(m[185]), .B(n4368), .Z(n6445) );
  NANDN U6768 ( .A(start_in[0]), .B(\modmult_1/xreg[185] ), .Z(n5163) );
  NANDN U6769 ( .A(n5643), .B(creg[185]), .Z(n5162) );
  AND U6770 ( .A(n5163), .B(n5162), .Z(n5164) );
  NANDN U6771 ( .A(n6445), .B(n5164), .Z(\modmult_1/xin[185] ) );
  AND U6772 ( .A(m[186]), .B(n4368), .Z(n6441) );
  NANDN U6773 ( .A(start_in[0]), .B(\modmult_1/xreg[186] ), .Z(n5166) );
  NANDN U6774 ( .A(n5643), .B(creg[186]), .Z(n5165) );
  AND U6775 ( .A(n5166), .B(n5165), .Z(n5167) );
  NANDN U6776 ( .A(n6441), .B(n5167), .Z(\modmult_1/xin[186] ) );
  AND U6777 ( .A(m[187]), .B(n4368), .Z(n6437) );
  NANDN U6778 ( .A(start_in[0]), .B(\modmult_1/xreg[187] ), .Z(n5169) );
  NANDN U6779 ( .A(n5643), .B(creg[187]), .Z(n5168) );
  AND U6780 ( .A(n5169), .B(n5168), .Z(n5170) );
  NANDN U6781 ( .A(n6437), .B(n5170), .Z(\modmult_1/xin[187] ) );
  AND U6782 ( .A(m[188]), .B(n4368), .Z(n6433) );
  NANDN U6783 ( .A(start_in[0]), .B(\modmult_1/xreg[188] ), .Z(n5172) );
  NANDN U6784 ( .A(n5643), .B(creg[188]), .Z(n5171) );
  AND U6785 ( .A(n5172), .B(n5171), .Z(n5173) );
  NANDN U6786 ( .A(n6433), .B(n5173), .Z(\modmult_1/xin[188] ) );
  AND U6787 ( .A(m[189]), .B(n4368), .Z(n6429) );
  NANDN U6788 ( .A(start_in[0]), .B(\modmult_1/xreg[189] ), .Z(n5175) );
  NANDN U6789 ( .A(n5643), .B(creg[189]), .Z(n5174) );
  AND U6790 ( .A(n5175), .B(n5174), .Z(n5176) );
  NANDN U6791 ( .A(n6429), .B(n5176), .Z(\modmult_1/xin[189] ) );
  AND U6792 ( .A(m[18]), .B(n4368), .Z(n7113) );
  NANDN U6793 ( .A(start_in[0]), .B(\modmult_1/xreg[18] ), .Z(n5178) );
  NANDN U6794 ( .A(n5643), .B(creg[18]), .Z(n5177) );
  AND U6795 ( .A(n5178), .B(n5177), .Z(n5179) );
  NANDN U6796 ( .A(n7113), .B(n5179), .Z(\modmult_1/xin[18] ) );
  AND U6797 ( .A(m[190]), .B(n4368), .Z(n6425) );
  NANDN U6798 ( .A(start_in[0]), .B(\modmult_1/xreg[190] ), .Z(n5181) );
  NANDN U6799 ( .A(n5643), .B(creg[190]), .Z(n5180) );
  AND U6800 ( .A(n5181), .B(n5180), .Z(n5182) );
  NANDN U6801 ( .A(n6425), .B(n5182), .Z(\modmult_1/xin[190] ) );
  AND U6802 ( .A(m[191]), .B(n4368), .Z(n6421) );
  NANDN U6803 ( .A(start_in[0]), .B(\modmult_1/xreg[191] ), .Z(n5184) );
  NANDN U6804 ( .A(n5643), .B(creg[191]), .Z(n5183) );
  AND U6805 ( .A(n5184), .B(n5183), .Z(n5185) );
  NANDN U6806 ( .A(n6421), .B(n5185), .Z(\modmult_1/xin[191] ) );
  AND U6807 ( .A(m[192]), .B(n4368), .Z(n6417) );
  NANDN U6808 ( .A(start_in[0]), .B(\modmult_1/xreg[192] ), .Z(n5187) );
  NANDN U6809 ( .A(n5643), .B(creg[192]), .Z(n5186) );
  AND U6810 ( .A(n5187), .B(n5186), .Z(n5188) );
  NANDN U6811 ( .A(n6417), .B(n5188), .Z(\modmult_1/xin[192] ) );
  AND U6812 ( .A(m[193]), .B(n4368), .Z(n6413) );
  NANDN U6813 ( .A(start_in[0]), .B(\modmult_1/xreg[193] ), .Z(n5190) );
  NANDN U6814 ( .A(n5643), .B(creg[193]), .Z(n5189) );
  AND U6815 ( .A(n5190), .B(n5189), .Z(n5191) );
  NANDN U6816 ( .A(n6413), .B(n5191), .Z(\modmult_1/xin[193] ) );
  AND U6817 ( .A(m[194]), .B(n4368), .Z(n6409) );
  NANDN U6818 ( .A(start_in[0]), .B(\modmult_1/xreg[194] ), .Z(n5193) );
  NANDN U6819 ( .A(n5643), .B(creg[194]), .Z(n5192) );
  AND U6820 ( .A(n5193), .B(n5192), .Z(n5194) );
  NANDN U6821 ( .A(n6409), .B(n5194), .Z(\modmult_1/xin[194] ) );
  AND U6822 ( .A(m[195]), .B(n4368), .Z(n6405) );
  NANDN U6823 ( .A(start_in[0]), .B(\modmult_1/xreg[195] ), .Z(n5196) );
  NANDN U6824 ( .A(n5643), .B(creg[195]), .Z(n5195) );
  AND U6825 ( .A(n5196), .B(n5195), .Z(n5197) );
  NANDN U6826 ( .A(n6405), .B(n5197), .Z(\modmult_1/xin[195] ) );
  AND U6827 ( .A(m[196]), .B(n4368), .Z(n6401) );
  NANDN U6828 ( .A(start_in[0]), .B(\modmult_1/xreg[196] ), .Z(n5199) );
  NANDN U6829 ( .A(n5643), .B(creg[196]), .Z(n5198) );
  AND U6830 ( .A(n5199), .B(n5198), .Z(n5200) );
  NANDN U6831 ( .A(n6401), .B(n5200), .Z(\modmult_1/xin[196] ) );
  AND U6832 ( .A(m[197]), .B(n4368), .Z(n6397) );
  NANDN U6833 ( .A(start_in[0]), .B(\modmult_1/xreg[197] ), .Z(n5202) );
  NANDN U6834 ( .A(n5643), .B(creg[197]), .Z(n5201) );
  AND U6835 ( .A(n5202), .B(n5201), .Z(n5203) );
  NANDN U6836 ( .A(n6397), .B(n5203), .Z(\modmult_1/xin[197] ) );
  AND U6837 ( .A(m[198]), .B(n4368), .Z(n6393) );
  NANDN U6838 ( .A(start_in[0]), .B(\modmult_1/xreg[198] ), .Z(n5205) );
  NANDN U6839 ( .A(n5643), .B(creg[198]), .Z(n5204) );
  AND U6840 ( .A(n5205), .B(n5204), .Z(n5206) );
  NANDN U6841 ( .A(n6393), .B(n5206), .Z(\modmult_1/xin[198] ) );
  AND U6842 ( .A(m[199]), .B(n4368), .Z(n6389) );
  NANDN U6843 ( .A(start_in[0]), .B(\modmult_1/xreg[199] ), .Z(n5208) );
  NANDN U6844 ( .A(n5643), .B(creg[199]), .Z(n5207) );
  AND U6845 ( .A(n5208), .B(n5207), .Z(n5209) );
  NANDN U6846 ( .A(n6389), .B(n5209), .Z(\modmult_1/xin[199] ) );
  AND U6847 ( .A(m[19]), .B(n4368), .Z(n7109) );
  NANDN U6848 ( .A(start_in[0]), .B(\modmult_1/xreg[19] ), .Z(n5211) );
  NANDN U6849 ( .A(n5643), .B(creg[19]), .Z(n5210) );
  AND U6850 ( .A(n5211), .B(n5210), .Z(n5212) );
  NANDN U6851 ( .A(n7109), .B(n5212), .Z(\modmult_1/xin[19] ) );
  AND U6852 ( .A(m[1]), .B(n4368), .Z(n7181) );
  NANDN U6853 ( .A(n5643), .B(creg[1]), .Z(n5213) );
  NANDN U6854 ( .A(n7181), .B(n5213), .Z(\modmult_1/xin[1] ) );
  AND U6855 ( .A(m[200]), .B(n4368), .Z(n6385) );
  NANDN U6856 ( .A(start_in[0]), .B(\modmult_1/xreg[200] ), .Z(n5215) );
  NANDN U6857 ( .A(n5643), .B(creg[200]), .Z(n5214) );
  AND U6858 ( .A(n5215), .B(n5214), .Z(n5216) );
  NANDN U6859 ( .A(n6385), .B(n5216), .Z(\modmult_1/xin[200] ) );
  AND U6860 ( .A(m[201]), .B(n4368), .Z(n6381) );
  NANDN U6861 ( .A(start_in[0]), .B(\modmult_1/xreg[201] ), .Z(n5218) );
  NANDN U6862 ( .A(n5643), .B(creg[201]), .Z(n5217) );
  AND U6863 ( .A(n5218), .B(n5217), .Z(n5219) );
  NANDN U6864 ( .A(n6381), .B(n5219), .Z(\modmult_1/xin[201] ) );
  AND U6865 ( .A(m[202]), .B(n4368), .Z(n6377) );
  NANDN U6866 ( .A(start_in[0]), .B(\modmult_1/xreg[202] ), .Z(n5221) );
  NANDN U6867 ( .A(n5643), .B(creg[202]), .Z(n5220) );
  AND U6868 ( .A(n5221), .B(n5220), .Z(n5222) );
  NANDN U6869 ( .A(n6377), .B(n5222), .Z(\modmult_1/xin[202] ) );
  AND U6870 ( .A(m[203]), .B(n4368), .Z(n6373) );
  NANDN U6871 ( .A(start_in[0]), .B(\modmult_1/xreg[203] ), .Z(n5224) );
  NANDN U6872 ( .A(n5643), .B(creg[203]), .Z(n5223) );
  AND U6873 ( .A(n5224), .B(n5223), .Z(n5225) );
  NANDN U6874 ( .A(n6373), .B(n5225), .Z(\modmult_1/xin[203] ) );
  AND U6875 ( .A(m[204]), .B(n4368), .Z(n6369) );
  NANDN U6876 ( .A(start_in[0]), .B(\modmult_1/xreg[204] ), .Z(n5227) );
  NANDN U6877 ( .A(n5643), .B(creg[204]), .Z(n5226) );
  AND U6878 ( .A(n5227), .B(n5226), .Z(n5228) );
  NANDN U6879 ( .A(n6369), .B(n5228), .Z(\modmult_1/xin[204] ) );
  AND U6880 ( .A(m[205]), .B(n4368), .Z(n6365) );
  NANDN U6881 ( .A(start_in[0]), .B(\modmult_1/xreg[205] ), .Z(n5230) );
  NANDN U6882 ( .A(n5643), .B(creg[205]), .Z(n5229) );
  AND U6883 ( .A(n5230), .B(n5229), .Z(n5231) );
  NANDN U6884 ( .A(n6365), .B(n5231), .Z(\modmult_1/xin[205] ) );
  AND U6885 ( .A(m[206]), .B(n4368), .Z(n6361) );
  NANDN U6886 ( .A(start_in[0]), .B(\modmult_1/xreg[206] ), .Z(n5233) );
  NANDN U6887 ( .A(n5643), .B(creg[206]), .Z(n5232) );
  AND U6888 ( .A(n5233), .B(n5232), .Z(n5234) );
  NANDN U6889 ( .A(n6361), .B(n5234), .Z(\modmult_1/xin[206] ) );
  AND U6890 ( .A(m[207]), .B(n4368), .Z(n6357) );
  NANDN U6891 ( .A(start_in[0]), .B(\modmult_1/xreg[207] ), .Z(n5236) );
  NANDN U6892 ( .A(n5643), .B(creg[207]), .Z(n5235) );
  AND U6893 ( .A(n5236), .B(n5235), .Z(n5237) );
  NANDN U6894 ( .A(n6357), .B(n5237), .Z(\modmult_1/xin[207] ) );
  AND U6895 ( .A(m[208]), .B(n4368), .Z(n6353) );
  NANDN U6896 ( .A(start_in[0]), .B(\modmult_1/xreg[208] ), .Z(n5239) );
  NANDN U6897 ( .A(n5643), .B(creg[208]), .Z(n5238) );
  AND U6898 ( .A(n5239), .B(n5238), .Z(n5240) );
  NANDN U6899 ( .A(n6353), .B(n5240), .Z(\modmult_1/xin[208] ) );
  AND U6900 ( .A(m[209]), .B(n4368), .Z(n6349) );
  NANDN U6901 ( .A(start_in[0]), .B(\modmult_1/xreg[209] ), .Z(n5242) );
  NANDN U6902 ( .A(n5643), .B(creg[209]), .Z(n5241) );
  AND U6903 ( .A(n5242), .B(n5241), .Z(n5243) );
  NANDN U6904 ( .A(n6349), .B(n5243), .Z(\modmult_1/xin[209] ) );
  AND U6905 ( .A(m[20]), .B(n4368), .Z(n7105) );
  NANDN U6906 ( .A(start_in[0]), .B(\modmult_1/xreg[20] ), .Z(n5245) );
  NANDN U6907 ( .A(n5643), .B(creg[20]), .Z(n5244) );
  AND U6908 ( .A(n5245), .B(n5244), .Z(n5246) );
  NANDN U6909 ( .A(n7105), .B(n5246), .Z(\modmult_1/xin[20] ) );
  AND U6910 ( .A(m[210]), .B(n4368), .Z(n6345) );
  NANDN U6911 ( .A(start_in[0]), .B(\modmult_1/xreg[210] ), .Z(n5248) );
  NANDN U6912 ( .A(n5643), .B(creg[210]), .Z(n5247) );
  AND U6913 ( .A(n5248), .B(n5247), .Z(n5249) );
  NANDN U6914 ( .A(n6345), .B(n5249), .Z(\modmult_1/xin[210] ) );
  AND U6915 ( .A(m[211]), .B(n4368), .Z(n6341) );
  NANDN U6916 ( .A(start_in[0]), .B(\modmult_1/xreg[211] ), .Z(n5251) );
  NANDN U6917 ( .A(n5643), .B(creg[211]), .Z(n5250) );
  AND U6918 ( .A(n5251), .B(n5250), .Z(n5252) );
  NANDN U6919 ( .A(n6341), .B(n5252), .Z(\modmult_1/xin[211] ) );
  AND U6920 ( .A(m[212]), .B(n4368), .Z(n6337) );
  NANDN U6921 ( .A(start_in[0]), .B(\modmult_1/xreg[212] ), .Z(n5254) );
  NANDN U6922 ( .A(n5643), .B(creg[212]), .Z(n5253) );
  AND U6923 ( .A(n5254), .B(n5253), .Z(n5255) );
  NANDN U6924 ( .A(n6337), .B(n5255), .Z(\modmult_1/xin[212] ) );
  AND U6925 ( .A(m[213]), .B(n4368), .Z(n6333) );
  NANDN U6926 ( .A(start_in[0]), .B(\modmult_1/xreg[213] ), .Z(n5257) );
  NANDN U6927 ( .A(n5643), .B(creg[213]), .Z(n5256) );
  AND U6928 ( .A(n5257), .B(n5256), .Z(n5258) );
  NANDN U6929 ( .A(n6333), .B(n5258), .Z(\modmult_1/xin[213] ) );
  AND U6930 ( .A(m[214]), .B(n4368), .Z(n6329) );
  NANDN U6931 ( .A(start_in[0]), .B(\modmult_1/xreg[214] ), .Z(n5260) );
  NANDN U6932 ( .A(n5643), .B(creg[214]), .Z(n5259) );
  AND U6933 ( .A(n5260), .B(n5259), .Z(n5261) );
  NANDN U6934 ( .A(n6329), .B(n5261), .Z(\modmult_1/xin[214] ) );
  AND U6935 ( .A(m[215]), .B(n4368), .Z(n6325) );
  NANDN U6936 ( .A(start_in[0]), .B(\modmult_1/xreg[215] ), .Z(n5263) );
  NANDN U6937 ( .A(n5643), .B(creg[215]), .Z(n5262) );
  AND U6938 ( .A(n5263), .B(n5262), .Z(n5264) );
  NANDN U6939 ( .A(n6325), .B(n5264), .Z(\modmult_1/xin[215] ) );
  AND U6940 ( .A(m[216]), .B(n4368), .Z(n6321) );
  NANDN U6941 ( .A(start_in[0]), .B(\modmult_1/xreg[216] ), .Z(n5266) );
  NANDN U6942 ( .A(n5643), .B(creg[216]), .Z(n5265) );
  AND U6943 ( .A(n5266), .B(n5265), .Z(n5267) );
  NANDN U6944 ( .A(n6321), .B(n5267), .Z(\modmult_1/xin[216] ) );
  AND U6945 ( .A(m[217]), .B(n4368), .Z(n6317) );
  NANDN U6946 ( .A(start_in[0]), .B(\modmult_1/xreg[217] ), .Z(n5269) );
  NANDN U6947 ( .A(n5643), .B(creg[217]), .Z(n5268) );
  AND U6948 ( .A(n5269), .B(n5268), .Z(n5270) );
  NANDN U6949 ( .A(n6317), .B(n5270), .Z(\modmult_1/xin[217] ) );
  AND U6950 ( .A(m[218]), .B(n4368), .Z(n6313) );
  NANDN U6951 ( .A(start_in[0]), .B(\modmult_1/xreg[218] ), .Z(n5272) );
  NANDN U6952 ( .A(n5643), .B(creg[218]), .Z(n5271) );
  AND U6953 ( .A(n5272), .B(n5271), .Z(n5273) );
  NANDN U6954 ( .A(n6313), .B(n5273), .Z(\modmult_1/xin[218] ) );
  AND U6955 ( .A(m[219]), .B(n4368), .Z(n6309) );
  NANDN U6956 ( .A(start_in[0]), .B(\modmult_1/xreg[219] ), .Z(n5275) );
  NANDN U6957 ( .A(n5643), .B(creg[219]), .Z(n5274) );
  AND U6958 ( .A(n5275), .B(n5274), .Z(n5276) );
  NANDN U6959 ( .A(n6309), .B(n5276), .Z(\modmult_1/xin[219] ) );
  AND U6960 ( .A(m[21]), .B(n4368), .Z(n7101) );
  NANDN U6961 ( .A(start_in[0]), .B(\modmult_1/xreg[21] ), .Z(n5278) );
  NANDN U6962 ( .A(n5643), .B(creg[21]), .Z(n5277) );
  AND U6963 ( .A(n5278), .B(n5277), .Z(n5279) );
  NANDN U6964 ( .A(n7101), .B(n5279), .Z(\modmult_1/xin[21] ) );
  AND U6965 ( .A(m[220]), .B(n4368), .Z(n6305) );
  NANDN U6966 ( .A(start_in[0]), .B(\modmult_1/xreg[220] ), .Z(n5281) );
  NANDN U6967 ( .A(n5643), .B(creg[220]), .Z(n5280) );
  AND U6968 ( .A(n5281), .B(n5280), .Z(n5282) );
  NANDN U6969 ( .A(n6305), .B(n5282), .Z(\modmult_1/xin[220] ) );
  AND U6970 ( .A(m[221]), .B(n4368), .Z(n6301) );
  NANDN U6971 ( .A(start_in[0]), .B(\modmult_1/xreg[221] ), .Z(n5284) );
  NANDN U6972 ( .A(n5643), .B(creg[221]), .Z(n5283) );
  AND U6973 ( .A(n5284), .B(n5283), .Z(n5285) );
  NANDN U6974 ( .A(n6301), .B(n5285), .Z(\modmult_1/xin[221] ) );
  AND U6975 ( .A(m[222]), .B(n4368), .Z(n6297) );
  NANDN U6976 ( .A(start_in[0]), .B(\modmult_1/xreg[222] ), .Z(n5287) );
  NANDN U6977 ( .A(n5643), .B(creg[222]), .Z(n5286) );
  AND U6978 ( .A(n5287), .B(n5286), .Z(n5288) );
  NANDN U6979 ( .A(n6297), .B(n5288), .Z(\modmult_1/xin[222] ) );
  AND U6980 ( .A(m[223]), .B(n4368), .Z(n6293) );
  NANDN U6981 ( .A(start_in[0]), .B(\modmult_1/xreg[223] ), .Z(n5290) );
  NANDN U6982 ( .A(n5643), .B(creg[223]), .Z(n5289) );
  AND U6983 ( .A(n5290), .B(n5289), .Z(n5291) );
  NANDN U6984 ( .A(n6293), .B(n5291), .Z(\modmult_1/xin[223] ) );
  AND U6985 ( .A(m[224]), .B(n4368), .Z(n6289) );
  NANDN U6986 ( .A(start_in[0]), .B(\modmult_1/xreg[224] ), .Z(n5293) );
  NANDN U6987 ( .A(n5643), .B(creg[224]), .Z(n5292) );
  AND U6988 ( .A(n5293), .B(n5292), .Z(n5294) );
  NANDN U6989 ( .A(n6289), .B(n5294), .Z(\modmult_1/xin[224] ) );
  AND U6990 ( .A(m[225]), .B(n4368), .Z(n6285) );
  NANDN U6991 ( .A(start_in[0]), .B(\modmult_1/xreg[225] ), .Z(n5296) );
  NANDN U6992 ( .A(n5643), .B(creg[225]), .Z(n5295) );
  AND U6993 ( .A(n5296), .B(n5295), .Z(n5297) );
  NANDN U6994 ( .A(n6285), .B(n5297), .Z(\modmult_1/xin[225] ) );
  AND U6995 ( .A(m[226]), .B(n4368), .Z(n6281) );
  NANDN U6996 ( .A(start_in[0]), .B(\modmult_1/xreg[226] ), .Z(n5299) );
  NANDN U6997 ( .A(n5643), .B(creg[226]), .Z(n5298) );
  AND U6998 ( .A(n5299), .B(n5298), .Z(n5300) );
  NANDN U6999 ( .A(n6281), .B(n5300), .Z(\modmult_1/xin[226] ) );
  AND U7000 ( .A(m[227]), .B(n4368), .Z(n6277) );
  NANDN U7001 ( .A(start_in[0]), .B(\modmult_1/xreg[227] ), .Z(n5302) );
  NANDN U7002 ( .A(n5643), .B(creg[227]), .Z(n5301) );
  AND U7003 ( .A(n5302), .B(n5301), .Z(n5303) );
  NANDN U7004 ( .A(n6277), .B(n5303), .Z(\modmult_1/xin[227] ) );
  AND U7005 ( .A(m[228]), .B(n4368), .Z(n6273) );
  NANDN U7006 ( .A(start_in[0]), .B(\modmult_1/xreg[228] ), .Z(n5305) );
  NANDN U7007 ( .A(n5643), .B(creg[228]), .Z(n5304) );
  AND U7008 ( .A(n5305), .B(n5304), .Z(n5306) );
  NANDN U7009 ( .A(n6273), .B(n5306), .Z(\modmult_1/xin[228] ) );
  AND U7010 ( .A(m[229]), .B(n4368), .Z(n6269) );
  NANDN U7011 ( .A(start_in[0]), .B(\modmult_1/xreg[229] ), .Z(n5308) );
  NANDN U7012 ( .A(n5643), .B(creg[229]), .Z(n5307) );
  AND U7013 ( .A(n5308), .B(n5307), .Z(n5309) );
  NANDN U7014 ( .A(n6269), .B(n5309), .Z(\modmult_1/xin[229] ) );
  AND U7015 ( .A(m[22]), .B(n4368), .Z(n7097) );
  NANDN U7016 ( .A(start_in[0]), .B(\modmult_1/xreg[22] ), .Z(n5311) );
  NANDN U7017 ( .A(n5643), .B(creg[22]), .Z(n5310) );
  AND U7018 ( .A(n5311), .B(n5310), .Z(n5312) );
  NANDN U7019 ( .A(n7097), .B(n5312), .Z(\modmult_1/xin[22] ) );
  AND U7020 ( .A(m[230]), .B(n4368), .Z(n6265) );
  NANDN U7021 ( .A(start_in[0]), .B(\modmult_1/xreg[230] ), .Z(n5314) );
  NANDN U7022 ( .A(n5643), .B(creg[230]), .Z(n5313) );
  AND U7023 ( .A(n5314), .B(n5313), .Z(n5315) );
  NANDN U7024 ( .A(n6265), .B(n5315), .Z(\modmult_1/xin[230] ) );
  AND U7025 ( .A(m[231]), .B(n4368), .Z(n6261) );
  NANDN U7026 ( .A(start_in[0]), .B(\modmult_1/xreg[231] ), .Z(n5317) );
  NANDN U7027 ( .A(n5643), .B(creg[231]), .Z(n5316) );
  AND U7028 ( .A(n5317), .B(n5316), .Z(n5318) );
  NANDN U7029 ( .A(n6261), .B(n5318), .Z(\modmult_1/xin[231] ) );
  AND U7030 ( .A(m[232]), .B(n4368), .Z(n6257) );
  NANDN U7031 ( .A(start_in[0]), .B(\modmult_1/xreg[232] ), .Z(n5320) );
  NANDN U7032 ( .A(n5643), .B(creg[232]), .Z(n5319) );
  AND U7033 ( .A(n5320), .B(n5319), .Z(n5321) );
  NANDN U7034 ( .A(n6257), .B(n5321), .Z(\modmult_1/xin[232] ) );
  AND U7035 ( .A(m[233]), .B(n4368), .Z(n6253) );
  NANDN U7036 ( .A(start_in[0]), .B(\modmult_1/xreg[233] ), .Z(n5323) );
  NANDN U7037 ( .A(n5643), .B(creg[233]), .Z(n5322) );
  AND U7038 ( .A(n5323), .B(n5322), .Z(n5324) );
  NANDN U7039 ( .A(n6253), .B(n5324), .Z(\modmult_1/xin[233] ) );
  AND U7040 ( .A(m[234]), .B(n4368), .Z(n6249) );
  NANDN U7041 ( .A(start_in[0]), .B(\modmult_1/xreg[234] ), .Z(n5326) );
  NANDN U7042 ( .A(n5643), .B(creg[234]), .Z(n5325) );
  AND U7043 ( .A(n5326), .B(n5325), .Z(n5327) );
  NANDN U7044 ( .A(n6249), .B(n5327), .Z(\modmult_1/xin[234] ) );
  AND U7045 ( .A(m[235]), .B(n4368), .Z(n6245) );
  NANDN U7046 ( .A(start_in[0]), .B(\modmult_1/xreg[235] ), .Z(n5329) );
  NANDN U7047 ( .A(n5643), .B(creg[235]), .Z(n5328) );
  AND U7048 ( .A(n5329), .B(n5328), .Z(n5330) );
  NANDN U7049 ( .A(n6245), .B(n5330), .Z(\modmult_1/xin[235] ) );
  AND U7050 ( .A(m[236]), .B(n4368), .Z(n6241) );
  NANDN U7051 ( .A(start_in[0]), .B(\modmult_1/xreg[236] ), .Z(n5332) );
  NANDN U7052 ( .A(n5643), .B(creg[236]), .Z(n5331) );
  AND U7053 ( .A(n5332), .B(n5331), .Z(n5333) );
  NANDN U7054 ( .A(n6241), .B(n5333), .Z(\modmult_1/xin[236] ) );
  AND U7055 ( .A(m[237]), .B(n4368), .Z(n6237) );
  NANDN U7056 ( .A(start_in[0]), .B(\modmult_1/xreg[237] ), .Z(n5335) );
  NANDN U7057 ( .A(n5643), .B(creg[237]), .Z(n5334) );
  AND U7058 ( .A(n5335), .B(n5334), .Z(n5336) );
  NANDN U7059 ( .A(n6237), .B(n5336), .Z(\modmult_1/xin[237] ) );
  AND U7060 ( .A(m[238]), .B(n4368), .Z(n6233) );
  NANDN U7061 ( .A(start_in[0]), .B(\modmult_1/xreg[238] ), .Z(n5338) );
  NANDN U7062 ( .A(n5643), .B(creg[238]), .Z(n5337) );
  AND U7063 ( .A(n5338), .B(n5337), .Z(n5339) );
  NANDN U7064 ( .A(n6233), .B(n5339), .Z(\modmult_1/xin[238] ) );
  AND U7065 ( .A(m[239]), .B(n4368), .Z(n6229) );
  NANDN U7066 ( .A(start_in[0]), .B(\modmult_1/xreg[239] ), .Z(n5341) );
  NANDN U7067 ( .A(n5643), .B(creg[239]), .Z(n5340) );
  AND U7068 ( .A(n5341), .B(n5340), .Z(n5342) );
  NANDN U7069 ( .A(n6229), .B(n5342), .Z(\modmult_1/xin[239] ) );
  AND U7070 ( .A(m[23]), .B(n4368), .Z(n7093) );
  NANDN U7071 ( .A(start_in[0]), .B(\modmult_1/xreg[23] ), .Z(n5344) );
  NANDN U7072 ( .A(n5643), .B(creg[23]), .Z(n5343) );
  AND U7073 ( .A(n5344), .B(n5343), .Z(n5345) );
  NANDN U7074 ( .A(n7093), .B(n5345), .Z(\modmult_1/xin[23] ) );
  AND U7075 ( .A(m[240]), .B(n4368), .Z(n6225) );
  NANDN U7076 ( .A(start_in[0]), .B(\modmult_1/xreg[240] ), .Z(n5347) );
  NANDN U7077 ( .A(n5643), .B(creg[240]), .Z(n5346) );
  AND U7078 ( .A(n5347), .B(n5346), .Z(n5348) );
  NANDN U7079 ( .A(n6225), .B(n5348), .Z(\modmult_1/xin[240] ) );
  AND U7080 ( .A(m[241]), .B(n4368), .Z(n6221) );
  NANDN U7081 ( .A(start_in[0]), .B(\modmult_1/xreg[241] ), .Z(n5350) );
  NANDN U7082 ( .A(n5643), .B(creg[241]), .Z(n5349) );
  AND U7083 ( .A(n5350), .B(n5349), .Z(n5351) );
  NANDN U7084 ( .A(n6221), .B(n5351), .Z(\modmult_1/xin[241] ) );
  AND U7085 ( .A(m[242]), .B(n4368), .Z(n6217) );
  NANDN U7086 ( .A(start_in[0]), .B(\modmult_1/xreg[242] ), .Z(n5353) );
  NANDN U7087 ( .A(n5643), .B(creg[242]), .Z(n5352) );
  AND U7088 ( .A(n5353), .B(n5352), .Z(n5354) );
  NANDN U7089 ( .A(n6217), .B(n5354), .Z(\modmult_1/xin[242] ) );
  AND U7090 ( .A(m[243]), .B(n4368), .Z(n6213) );
  NANDN U7091 ( .A(start_in[0]), .B(\modmult_1/xreg[243] ), .Z(n5356) );
  NANDN U7092 ( .A(n5643), .B(creg[243]), .Z(n5355) );
  AND U7093 ( .A(n5356), .B(n5355), .Z(n5357) );
  NANDN U7094 ( .A(n6213), .B(n5357), .Z(\modmult_1/xin[243] ) );
  AND U7095 ( .A(m[244]), .B(n4368), .Z(n6209) );
  NANDN U7096 ( .A(start_in[0]), .B(\modmult_1/xreg[244] ), .Z(n5359) );
  NANDN U7097 ( .A(n5643), .B(creg[244]), .Z(n5358) );
  AND U7098 ( .A(n5359), .B(n5358), .Z(n5360) );
  NANDN U7099 ( .A(n6209), .B(n5360), .Z(\modmult_1/xin[244] ) );
  AND U7100 ( .A(m[245]), .B(n4368), .Z(n6205) );
  NANDN U7101 ( .A(start_in[0]), .B(\modmult_1/xreg[245] ), .Z(n5362) );
  NANDN U7102 ( .A(n5643), .B(creg[245]), .Z(n5361) );
  AND U7103 ( .A(n5362), .B(n5361), .Z(n5363) );
  NANDN U7104 ( .A(n6205), .B(n5363), .Z(\modmult_1/xin[245] ) );
  AND U7105 ( .A(m[246]), .B(n4368), .Z(n6201) );
  NANDN U7106 ( .A(start_in[0]), .B(\modmult_1/xreg[246] ), .Z(n5365) );
  NANDN U7107 ( .A(n5643), .B(creg[246]), .Z(n5364) );
  AND U7108 ( .A(n5365), .B(n5364), .Z(n5366) );
  NANDN U7109 ( .A(n6201), .B(n5366), .Z(\modmult_1/xin[246] ) );
  AND U7110 ( .A(m[247]), .B(n4368), .Z(n6197) );
  NANDN U7111 ( .A(start_in[0]), .B(\modmult_1/xreg[247] ), .Z(n5368) );
  NANDN U7112 ( .A(n5643), .B(creg[247]), .Z(n5367) );
  AND U7113 ( .A(n5368), .B(n5367), .Z(n5369) );
  NANDN U7114 ( .A(n6197), .B(n5369), .Z(\modmult_1/xin[247] ) );
  AND U7115 ( .A(m[248]), .B(n4368), .Z(n6193) );
  NANDN U7116 ( .A(start_in[0]), .B(\modmult_1/xreg[248] ), .Z(n5371) );
  NANDN U7117 ( .A(n5643), .B(creg[248]), .Z(n5370) );
  AND U7118 ( .A(n5371), .B(n5370), .Z(n5372) );
  NANDN U7119 ( .A(n6193), .B(n5372), .Z(\modmult_1/xin[248] ) );
  AND U7120 ( .A(m[249]), .B(n4368), .Z(n6189) );
  NANDN U7121 ( .A(start_in[0]), .B(\modmult_1/xreg[249] ), .Z(n5374) );
  NANDN U7122 ( .A(n5643), .B(creg[249]), .Z(n5373) );
  AND U7123 ( .A(n5374), .B(n5373), .Z(n5375) );
  NANDN U7124 ( .A(n6189), .B(n5375), .Z(\modmult_1/xin[249] ) );
  AND U7125 ( .A(m[24]), .B(n4368), .Z(n7089) );
  NANDN U7126 ( .A(start_in[0]), .B(\modmult_1/xreg[24] ), .Z(n5377) );
  NANDN U7127 ( .A(n5643), .B(creg[24]), .Z(n5376) );
  AND U7128 ( .A(n5377), .B(n5376), .Z(n5378) );
  NANDN U7129 ( .A(n7089), .B(n5378), .Z(\modmult_1/xin[24] ) );
  AND U7130 ( .A(m[250]), .B(n4368), .Z(n6185) );
  NANDN U7131 ( .A(start_in[0]), .B(\modmult_1/xreg[250] ), .Z(n5380) );
  NANDN U7132 ( .A(n5643), .B(creg[250]), .Z(n5379) );
  AND U7133 ( .A(n5380), .B(n5379), .Z(n5381) );
  NANDN U7134 ( .A(n6185), .B(n5381), .Z(\modmult_1/xin[250] ) );
  AND U7135 ( .A(m[251]), .B(n4368), .Z(n6181) );
  NANDN U7136 ( .A(start_in[0]), .B(\modmult_1/xreg[251] ), .Z(n5383) );
  NANDN U7137 ( .A(n5643), .B(creg[251]), .Z(n5382) );
  AND U7138 ( .A(n5383), .B(n5382), .Z(n5384) );
  NANDN U7139 ( .A(n6181), .B(n5384), .Z(\modmult_1/xin[251] ) );
  AND U7140 ( .A(m[252]), .B(n4368), .Z(n6177) );
  NANDN U7141 ( .A(start_in[0]), .B(\modmult_1/xreg[252] ), .Z(n5386) );
  NANDN U7142 ( .A(n5643), .B(creg[252]), .Z(n5385) );
  AND U7143 ( .A(n5386), .B(n5385), .Z(n5387) );
  NANDN U7144 ( .A(n6177), .B(n5387), .Z(\modmult_1/xin[252] ) );
  AND U7145 ( .A(m[253]), .B(n4368), .Z(n6173) );
  NANDN U7146 ( .A(start_in[0]), .B(\modmult_1/xreg[253] ), .Z(n5389) );
  NANDN U7147 ( .A(n5643), .B(creg[253]), .Z(n5388) );
  AND U7148 ( .A(n5389), .B(n5388), .Z(n5390) );
  NANDN U7149 ( .A(n6173), .B(n5390), .Z(\modmult_1/xin[253] ) );
  AND U7150 ( .A(m[254]), .B(n4368), .Z(n6169) );
  NANDN U7151 ( .A(start_in[0]), .B(\modmult_1/xreg[254] ), .Z(n5392) );
  NANDN U7152 ( .A(n5643), .B(creg[254]), .Z(n5391) );
  AND U7153 ( .A(n5392), .B(n5391), .Z(n5393) );
  NANDN U7154 ( .A(n6169), .B(n5393), .Z(\modmult_1/xin[254] ) );
  AND U7155 ( .A(m[255]), .B(n4368), .Z(n6162) );
  NANDN U7156 ( .A(start_in[0]), .B(\modmult_1/xreg[255] ), .Z(n5395) );
  NANDN U7157 ( .A(n5643), .B(creg[255]), .Z(n5394) );
  AND U7158 ( .A(n5395), .B(n5394), .Z(n5396) );
  NANDN U7159 ( .A(n6162), .B(n5396), .Z(\modmult_1/xin[255] ) );
  AND U7160 ( .A(m[25]), .B(n4368), .Z(n7085) );
  NANDN U7161 ( .A(start_in[0]), .B(\modmult_1/xreg[25] ), .Z(n5398) );
  NANDN U7162 ( .A(n5643), .B(creg[25]), .Z(n5397) );
  AND U7163 ( .A(n5398), .B(n5397), .Z(n5399) );
  NANDN U7164 ( .A(n7085), .B(n5399), .Z(\modmult_1/xin[25] ) );
  AND U7165 ( .A(m[26]), .B(n4368), .Z(n7081) );
  NANDN U7166 ( .A(start_in[0]), .B(\modmult_1/xreg[26] ), .Z(n5401) );
  NANDN U7167 ( .A(n5643), .B(creg[26]), .Z(n5400) );
  AND U7168 ( .A(n5401), .B(n5400), .Z(n5402) );
  NANDN U7169 ( .A(n7081), .B(n5402), .Z(\modmult_1/xin[26] ) );
  AND U7170 ( .A(m[27]), .B(n4368), .Z(n7077) );
  NANDN U7171 ( .A(start_in[0]), .B(\modmult_1/xreg[27] ), .Z(n5404) );
  NANDN U7172 ( .A(n5643), .B(creg[27]), .Z(n5403) );
  AND U7173 ( .A(n5404), .B(n5403), .Z(n5405) );
  NANDN U7174 ( .A(n7077), .B(n5405), .Z(\modmult_1/xin[27] ) );
  AND U7175 ( .A(m[28]), .B(n4368), .Z(n7073) );
  NANDN U7176 ( .A(start_in[0]), .B(\modmult_1/xreg[28] ), .Z(n5407) );
  NANDN U7177 ( .A(n5643), .B(creg[28]), .Z(n5406) );
  AND U7178 ( .A(n5407), .B(n5406), .Z(n5408) );
  NANDN U7179 ( .A(n7073), .B(n5408), .Z(\modmult_1/xin[28] ) );
  AND U7180 ( .A(m[29]), .B(n4368), .Z(n7069) );
  NANDN U7181 ( .A(start_in[0]), .B(\modmult_1/xreg[29] ), .Z(n5410) );
  NANDN U7182 ( .A(n5643), .B(creg[29]), .Z(n5409) );
  AND U7183 ( .A(n5410), .B(n5409), .Z(n5411) );
  NANDN U7184 ( .A(n7069), .B(n5411), .Z(\modmult_1/xin[29] ) );
  AND U7185 ( .A(m[2]), .B(n4368), .Z(n7177) );
  NANDN U7186 ( .A(start_in[0]), .B(\modmult_1/xreg[2] ), .Z(n5413) );
  NANDN U7187 ( .A(n5643), .B(creg[2]), .Z(n5412) );
  AND U7188 ( .A(n5413), .B(n5412), .Z(n5414) );
  NANDN U7189 ( .A(n7177), .B(n5414), .Z(\modmult_1/xin[2] ) );
  AND U7190 ( .A(m[30]), .B(n4368), .Z(n7065) );
  NANDN U7191 ( .A(start_in[0]), .B(\modmult_1/xreg[30] ), .Z(n5416) );
  NANDN U7192 ( .A(n5643), .B(creg[30]), .Z(n5415) );
  AND U7193 ( .A(n5416), .B(n5415), .Z(n5417) );
  NANDN U7194 ( .A(n7065), .B(n5417), .Z(\modmult_1/xin[30] ) );
  AND U7195 ( .A(m[31]), .B(n4368), .Z(n7061) );
  NANDN U7196 ( .A(start_in[0]), .B(\modmult_1/xreg[31] ), .Z(n5419) );
  NANDN U7197 ( .A(n5643), .B(creg[31]), .Z(n5418) );
  AND U7198 ( .A(n5419), .B(n5418), .Z(n5420) );
  NANDN U7199 ( .A(n7061), .B(n5420), .Z(\modmult_1/xin[31] ) );
  AND U7200 ( .A(m[32]), .B(n4368), .Z(n7057) );
  NANDN U7201 ( .A(start_in[0]), .B(\modmult_1/xreg[32] ), .Z(n5422) );
  NANDN U7202 ( .A(n5643), .B(creg[32]), .Z(n5421) );
  AND U7203 ( .A(n5422), .B(n5421), .Z(n5423) );
  NANDN U7204 ( .A(n7057), .B(n5423), .Z(\modmult_1/xin[32] ) );
  AND U7205 ( .A(m[33]), .B(n4368), .Z(n7053) );
  NANDN U7206 ( .A(start_in[0]), .B(\modmult_1/xreg[33] ), .Z(n5425) );
  NANDN U7207 ( .A(n5643), .B(creg[33]), .Z(n5424) );
  AND U7208 ( .A(n5425), .B(n5424), .Z(n5426) );
  NANDN U7209 ( .A(n7053), .B(n5426), .Z(\modmult_1/xin[33] ) );
  AND U7210 ( .A(m[34]), .B(n4368), .Z(n7049) );
  NANDN U7211 ( .A(start_in[0]), .B(\modmult_1/xreg[34] ), .Z(n5428) );
  NANDN U7212 ( .A(n5643), .B(creg[34]), .Z(n5427) );
  AND U7213 ( .A(n5428), .B(n5427), .Z(n5429) );
  NANDN U7214 ( .A(n7049), .B(n5429), .Z(\modmult_1/xin[34] ) );
  AND U7215 ( .A(m[35]), .B(n4368), .Z(n7045) );
  NANDN U7216 ( .A(start_in[0]), .B(\modmult_1/xreg[35] ), .Z(n5431) );
  NANDN U7217 ( .A(n5643), .B(creg[35]), .Z(n5430) );
  AND U7218 ( .A(n5431), .B(n5430), .Z(n5432) );
  NANDN U7219 ( .A(n7045), .B(n5432), .Z(\modmult_1/xin[35] ) );
  AND U7220 ( .A(m[36]), .B(n4368), .Z(n7041) );
  NANDN U7221 ( .A(start_in[0]), .B(\modmult_1/xreg[36] ), .Z(n5434) );
  NANDN U7222 ( .A(n5643), .B(creg[36]), .Z(n5433) );
  AND U7223 ( .A(n5434), .B(n5433), .Z(n5435) );
  NANDN U7224 ( .A(n7041), .B(n5435), .Z(\modmult_1/xin[36] ) );
  AND U7225 ( .A(m[37]), .B(n4368), .Z(n7037) );
  NANDN U7226 ( .A(start_in[0]), .B(\modmult_1/xreg[37] ), .Z(n5437) );
  NANDN U7227 ( .A(n5643), .B(creg[37]), .Z(n5436) );
  AND U7228 ( .A(n5437), .B(n5436), .Z(n5438) );
  NANDN U7229 ( .A(n7037), .B(n5438), .Z(\modmult_1/xin[37] ) );
  AND U7230 ( .A(m[38]), .B(n4368), .Z(n7033) );
  NANDN U7231 ( .A(start_in[0]), .B(\modmult_1/xreg[38] ), .Z(n5440) );
  NANDN U7232 ( .A(n5643), .B(creg[38]), .Z(n5439) );
  AND U7233 ( .A(n5440), .B(n5439), .Z(n5441) );
  NANDN U7234 ( .A(n7033), .B(n5441), .Z(\modmult_1/xin[38] ) );
  AND U7235 ( .A(m[39]), .B(n4368), .Z(n7029) );
  NANDN U7236 ( .A(start_in[0]), .B(\modmult_1/xreg[39] ), .Z(n5443) );
  NANDN U7237 ( .A(n5643), .B(creg[39]), .Z(n5442) );
  AND U7238 ( .A(n5443), .B(n5442), .Z(n5444) );
  NANDN U7239 ( .A(n7029), .B(n5444), .Z(\modmult_1/xin[39] ) );
  AND U7240 ( .A(m[3]), .B(n4368), .Z(n7173) );
  NANDN U7241 ( .A(start_in[0]), .B(\modmult_1/xreg[3] ), .Z(n5446) );
  NANDN U7242 ( .A(n5643), .B(creg[3]), .Z(n5445) );
  AND U7243 ( .A(n5446), .B(n5445), .Z(n5447) );
  NANDN U7244 ( .A(n7173), .B(n5447), .Z(\modmult_1/xin[3] ) );
  AND U7245 ( .A(m[40]), .B(n4368), .Z(n7025) );
  NANDN U7246 ( .A(start_in[0]), .B(\modmult_1/xreg[40] ), .Z(n5449) );
  NANDN U7247 ( .A(n5643), .B(creg[40]), .Z(n5448) );
  AND U7248 ( .A(n5449), .B(n5448), .Z(n5450) );
  NANDN U7249 ( .A(n7025), .B(n5450), .Z(\modmult_1/xin[40] ) );
  AND U7250 ( .A(m[41]), .B(n4368), .Z(n7021) );
  NANDN U7251 ( .A(start_in[0]), .B(\modmult_1/xreg[41] ), .Z(n5452) );
  NANDN U7252 ( .A(n5643), .B(creg[41]), .Z(n5451) );
  AND U7253 ( .A(n5452), .B(n5451), .Z(n5453) );
  NANDN U7254 ( .A(n7021), .B(n5453), .Z(\modmult_1/xin[41] ) );
  AND U7255 ( .A(m[42]), .B(n4368), .Z(n7017) );
  NANDN U7256 ( .A(start_in[0]), .B(\modmult_1/xreg[42] ), .Z(n5455) );
  NANDN U7257 ( .A(n5643), .B(creg[42]), .Z(n5454) );
  AND U7258 ( .A(n5455), .B(n5454), .Z(n5456) );
  NANDN U7259 ( .A(n7017), .B(n5456), .Z(\modmult_1/xin[42] ) );
  AND U7260 ( .A(m[43]), .B(n4368), .Z(n7013) );
  NANDN U7261 ( .A(start_in[0]), .B(\modmult_1/xreg[43] ), .Z(n5458) );
  NANDN U7262 ( .A(n5643), .B(creg[43]), .Z(n5457) );
  AND U7263 ( .A(n5458), .B(n5457), .Z(n5459) );
  NANDN U7264 ( .A(n7013), .B(n5459), .Z(\modmult_1/xin[43] ) );
  AND U7265 ( .A(m[44]), .B(n4368), .Z(n7009) );
  NANDN U7266 ( .A(start_in[0]), .B(\modmult_1/xreg[44] ), .Z(n5461) );
  NANDN U7267 ( .A(n5643), .B(creg[44]), .Z(n5460) );
  AND U7268 ( .A(n5461), .B(n5460), .Z(n5462) );
  NANDN U7269 ( .A(n7009), .B(n5462), .Z(\modmult_1/xin[44] ) );
  AND U7270 ( .A(m[45]), .B(n4368), .Z(n7005) );
  NANDN U7271 ( .A(start_in[0]), .B(\modmult_1/xreg[45] ), .Z(n5464) );
  NANDN U7272 ( .A(n5643), .B(creg[45]), .Z(n5463) );
  AND U7273 ( .A(n5464), .B(n5463), .Z(n5465) );
  NANDN U7274 ( .A(n7005), .B(n5465), .Z(\modmult_1/xin[45] ) );
  AND U7275 ( .A(m[46]), .B(n4368), .Z(n7001) );
  NANDN U7276 ( .A(start_in[0]), .B(\modmult_1/xreg[46] ), .Z(n5467) );
  NANDN U7277 ( .A(n5643), .B(creg[46]), .Z(n5466) );
  AND U7278 ( .A(n5467), .B(n5466), .Z(n5468) );
  NANDN U7279 ( .A(n7001), .B(n5468), .Z(\modmult_1/xin[46] ) );
  AND U7280 ( .A(m[47]), .B(n4368), .Z(n6997) );
  NANDN U7281 ( .A(start_in[0]), .B(\modmult_1/xreg[47] ), .Z(n5470) );
  NANDN U7282 ( .A(n5643), .B(creg[47]), .Z(n5469) );
  AND U7283 ( .A(n5470), .B(n5469), .Z(n5471) );
  NANDN U7284 ( .A(n6997), .B(n5471), .Z(\modmult_1/xin[47] ) );
  AND U7285 ( .A(m[48]), .B(n4368), .Z(n6993) );
  NANDN U7286 ( .A(start_in[0]), .B(\modmult_1/xreg[48] ), .Z(n5473) );
  NANDN U7287 ( .A(n5643), .B(creg[48]), .Z(n5472) );
  AND U7288 ( .A(n5473), .B(n5472), .Z(n5474) );
  NANDN U7289 ( .A(n6993), .B(n5474), .Z(\modmult_1/xin[48] ) );
  AND U7290 ( .A(m[49]), .B(n4368), .Z(n6989) );
  NANDN U7291 ( .A(start_in[0]), .B(\modmult_1/xreg[49] ), .Z(n5476) );
  NANDN U7292 ( .A(n5643), .B(creg[49]), .Z(n5475) );
  AND U7293 ( .A(n5476), .B(n5475), .Z(n5477) );
  NANDN U7294 ( .A(n6989), .B(n5477), .Z(\modmult_1/xin[49] ) );
  AND U7295 ( .A(m[4]), .B(n4368), .Z(n7169) );
  NANDN U7296 ( .A(start_in[0]), .B(\modmult_1/xreg[4] ), .Z(n5479) );
  NANDN U7297 ( .A(n5643), .B(creg[4]), .Z(n5478) );
  AND U7298 ( .A(n5479), .B(n5478), .Z(n5480) );
  NANDN U7299 ( .A(n7169), .B(n5480), .Z(\modmult_1/xin[4] ) );
  AND U7300 ( .A(m[50]), .B(n4368), .Z(n6985) );
  NANDN U7301 ( .A(start_in[0]), .B(\modmult_1/xreg[50] ), .Z(n5482) );
  NANDN U7302 ( .A(n5643), .B(creg[50]), .Z(n5481) );
  AND U7303 ( .A(n5482), .B(n5481), .Z(n5483) );
  NANDN U7304 ( .A(n6985), .B(n5483), .Z(\modmult_1/xin[50] ) );
  AND U7305 ( .A(m[51]), .B(n4368), .Z(n6981) );
  NANDN U7306 ( .A(start_in[0]), .B(\modmult_1/xreg[51] ), .Z(n5485) );
  NANDN U7307 ( .A(n5643), .B(creg[51]), .Z(n5484) );
  AND U7308 ( .A(n5485), .B(n5484), .Z(n5486) );
  NANDN U7309 ( .A(n6981), .B(n5486), .Z(\modmult_1/xin[51] ) );
  AND U7310 ( .A(m[52]), .B(n4368), .Z(n6977) );
  NANDN U7311 ( .A(start_in[0]), .B(\modmult_1/xreg[52] ), .Z(n5488) );
  NANDN U7312 ( .A(n5643), .B(creg[52]), .Z(n5487) );
  AND U7313 ( .A(n5488), .B(n5487), .Z(n5489) );
  NANDN U7314 ( .A(n6977), .B(n5489), .Z(\modmult_1/xin[52] ) );
  AND U7315 ( .A(m[53]), .B(n4368), .Z(n6973) );
  NANDN U7316 ( .A(start_in[0]), .B(\modmult_1/xreg[53] ), .Z(n5491) );
  NANDN U7317 ( .A(n5643), .B(creg[53]), .Z(n5490) );
  AND U7318 ( .A(n5491), .B(n5490), .Z(n5492) );
  NANDN U7319 ( .A(n6973), .B(n5492), .Z(\modmult_1/xin[53] ) );
  AND U7320 ( .A(m[54]), .B(n4368), .Z(n6969) );
  NANDN U7321 ( .A(start_in[0]), .B(\modmult_1/xreg[54] ), .Z(n5494) );
  NANDN U7322 ( .A(n5643), .B(creg[54]), .Z(n5493) );
  AND U7323 ( .A(n5494), .B(n5493), .Z(n5495) );
  NANDN U7324 ( .A(n6969), .B(n5495), .Z(\modmult_1/xin[54] ) );
  AND U7325 ( .A(m[55]), .B(n4368), .Z(n6965) );
  NANDN U7326 ( .A(start_in[0]), .B(\modmult_1/xreg[55] ), .Z(n5497) );
  NANDN U7327 ( .A(n5643), .B(creg[55]), .Z(n5496) );
  AND U7328 ( .A(n5497), .B(n5496), .Z(n5498) );
  NANDN U7329 ( .A(n6965), .B(n5498), .Z(\modmult_1/xin[55] ) );
  AND U7330 ( .A(m[56]), .B(n4368), .Z(n6961) );
  NANDN U7331 ( .A(start_in[0]), .B(\modmult_1/xreg[56] ), .Z(n5500) );
  NANDN U7332 ( .A(n5643), .B(creg[56]), .Z(n5499) );
  AND U7333 ( .A(n5500), .B(n5499), .Z(n5501) );
  NANDN U7334 ( .A(n6961), .B(n5501), .Z(\modmult_1/xin[56] ) );
  AND U7335 ( .A(m[57]), .B(n4368), .Z(n6957) );
  NANDN U7336 ( .A(start_in[0]), .B(\modmult_1/xreg[57] ), .Z(n5503) );
  NANDN U7337 ( .A(n5643), .B(creg[57]), .Z(n5502) );
  AND U7338 ( .A(n5503), .B(n5502), .Z(n5504) );
  NANDN U7339 ( .A(n6957), .B(n5504), .Z(\modmult_1/xin[57] ) );
  AND U7340 ( .A(m[58]), .B(n4368), .Z(n6953) );
  NANDN U7341 ( .A(start_in[0]), .B(\modmult_1/xreg[58] ), .Z(n5506) );
  NANDN U7342 ( .A(n5643), .B(creg[58]), .Z(n5505) );
  AND U7343 ( .A(n5506), .B(n5505), .Z(n5507) );
  NANDN U7344 ( .A(n6953), .B(n5507), .Z(\modmult_1/xin[58] ) );
  AND U7345 ( .A(m[59]), .B(n4368), .Z(n6949) );
  NANDN U7346 ( .A(start_in[0]), .B(\modmult_1/xreg[59] ), .Z(n5509) );
  NANDN U7347 ( .A(n5643), .B(creg[59]), .Z(n5508) );
  AND U7348 ( .A(n5509), .B(n5508), .Z(n5510) );
  NANDN U7349 ( .A(n6949), .B(n5510), .Z(\modmult_1/xin[59] ) );
  AND U7350 ( .A(m[5]), .B(n4368), .Z(n7165) );
  NANDN U7351 ( .A(start_in[0]), .B(\modmult_1/xreg[5] ), .Z(n5512) );
  NANDN U7352 ( .A(n5643), .B(creg[5]), .Z(n5511) );
  AND U7353 ( .A(n5512), .B(n5511), .Z(n5513) );
  NANDN U7354 ( .A(n7165), .B(n5513), .Z(\modmult_1/xin[5] ) );
  AND U7355 ( .A(m[60]), .B(n4368), .Z(n6945) );
  NANDN U7356 ( .A(start_in[0]), .B(\modmult_1/xreg[60] ), .Z(n5515) );
  NANDN U7357 ( .A(n5643), .B(creg[60]), .Z(n5514) );
  AND U7358 ( .A(n5515), .B(n5514), .Z(n5516) );
  NANDN U7359 ( .A(n6945), .B(n5516), .Z(\modmult_1/xin[60] ) );
  AND U7360 ( .A(m[61]), .B(n4368), .Z(n6941) );
  NANDN U7361 ( .A(start_in[0]), .B(\modmult_1/xreg[61] ), .Z(n5518) );
  NANDN U7362 ( .A(n5643), .B(creg[61]), .Z(n5517) );
  AND U7363 ( .A(n5518), .B(n5517), .Z(n5519) );
  NANDN U7364 ( .A(n6941), .B(n5519), .Z(\modmult_1/xin[61] ) );
  AND U7365 ( .A(m[62]), .B(n4368), .Z(n6937) );
  NANDN U7366 ( .A(start_in[0]), .B(\modmult_1/xreg[62] ), .Z(n5521) );
  NANDN U7367 ( .A(n5643), .B(creg[62]), .Z(n5520) );
  AND U7368 ( .A(n5521), .B(n5520), .Z(n5522) );
  NANDN U7369 ( .A(n6937), .B(n5522), .Z(\modmult_1/xin[62] ) );
  AND U7370 ( .A(m[63]), .B(n4368), .Z(n6933) );
  NANDN U7371 ( .A(start_in[0]), .B(\modmult_1/xreg[63] ), .Z(n5524) );
  NANDN U7372 ( .A(n5643), .B(creg[63]), .Z(n5523) );
  AND U7373 ( .A(n5524), .B(n5523), .Z(n5525) );
  NANDN U7374 ( .A(n6933), .B(n5525), .Z(\modmult_1/xin[63] ) );
  AND U7375 ( .A(m[64]), .B(n4368), .Z(n6929) );
  NANDN U7376 ( .A(start_in[0]), .B(\modmult_1/xreg[64] ), .Z(n5527) );
  NANDN U7377 ( .A(n5643), .B(creg[64]), .Z(n5526) );
  AND U7378 ( .A(n5527), .B(n5526), .Z(n5528) );
  NANDN U7379 ( .A(n6929), .B(n5528), .Z(\modmult_1/xin[64] ) );
  AND U7380 ( .A(m[65]), .B(n4368), .Z(n6925) );
  NANDN U7381 ( .A(start_in[0]), .B(\modmult_1/xreg[65] ), .Z(n5530) );
  NANDN U7382 ( .A(n5643), .B(creg[65]), .Z(n5529) );
  AND U7383 ( .A(n5530), .B(n5529), .Z(n5531) );
  NANDN U7384 ( .A(n6925), .B(n5531), .Z(\modmult_1/xin[65] ) );
  AND U7385 ( .A(m[66]), .B(n4368), .Z(n6921) );
  NANDN U7386 ( .A(start_in[0]), .B(\modmult_1/xreg[66] ), .Z(n5533) );
  NANDN U7387 ( .A(n5643), .B(creg[66]), .Z(n5532) );
  AND U7388 ( .A(n5533), .B(n5532), .Z(n5534) );
  NANDN U7389 ( .A(n6921), .B(n5534), .Z(\modmult_1/xin[66] ) );
  AND U7390 ( .A(m[67]), .B(n4368), .Z(n6917) );
  NANDN U7391 ( .A(start_in[0]), .B(\modmult_1/xreg[67] ), .Z(n5536) );
  NANDN U7392 ( .A(n5643), .B(creg[67]), .Z(n5535) );
  AND U7393 ( .A(n5536), .B(n5535), .Z(n5537) );
  NANDN U7394 ( .A(n6917), .B(n5537), .Z(\modmult_1/xin[67] ) );
  AND U7395 ( .A(m[68]), .B(n4368), .Z(n6913) );
  NANDN U7396 ( .A(start_in[0]), .B(\modmult_1/xreg[68] ), .Z(n5539) );
  NANDN U7397 ( .A(n5643), .B(creg[68]), .Z(n5538) );
  AND U7398 ( .A(n5539), .B(n5538), .Z(n5540) );
  NANDN U7399 ( .A(n6913), .B(n5540), .Z(\modmult_1/xin[68] ) );
  AND U7400 ( .A(m[69]), .B(n4368), .Z(n6909) );
  NANDN U7401 ( .A(start_in[0]), .B(\modmult_1/xreg[69] ), .Z(n5542) );
  NANDN U7402 ( .A(n5643), .B(creg[69]), .Z(n5541) );
  AND U7403 ( .A(n5542), .B(n5541), .Z(n5543) );
  NANDN U7404 ( .A(n6909), .B(n5543), .Z(\modmult_1/xin[69] ) );
  AND U7405 ( .A(m[6]), .B(n4368), .Z(n7161) );
  NANDN U7406 ( .A(start_in[0]), .B(\modmult_1/xreg[6] ), .Z(n5545) );
  NANDN U7407 ( .A(n5643), .B(creg[6]), .Z(n5544) );
  AND U7408 ( .A(n5545), .B(n5544), .Z(n5546) );
  NANDN U7409 ( .A(n7161), .B(n5546), .Z(\modmult_1/xin[6] ) );
  AND U7410 ( .A(m[70]), .B(n4368), .Z(n6905) );
  NANDN U7411 ( .A(start_in[0]), .B(\modmult_1/xreg[70] ), .Z(n5548) );
  NANDN U7412 ( .A(n5643), .B(creg[70]), .Z(n5547) );
  AND U7413 ( .A(n5548), .B(n5547), .Z(n5549) );
  NANDN U7414 ( .A(n6905), .B(n5549), .Z(\modmult_1/xin[70] ) );
  AND U7415 ( .A(m[71]), .B(n4368), .Z(n6901) );
  NANDN U7416 ( .A(start_in[0]), .B(\modmult_1/xreg[71] ), .Z(n5551) );
  NANDN U7417 ( .A(n5643), .B(creg[71]), .Z(n5550) );
  AND U7418 ( .A(n5551), .B(n5550), .Z(n5552) );
  NANDN U7419 ( .A(n6901), .B(n5552), .Z(\modmult_1/xin[71] ) );
  AND U7420 ( .A(m[72]), .B(n4368), .Z(n6897) );
  NANDN U7421 ( .A(start_in[0]), .B(\modmult_1/xreg[72] ), .Z(n5554) );
  NANDN U7422 ( .A(n5643), .B(creg[72]), .Z(n5553) );
  AND U7423 ( .A(n5554), .B(n5553), .Z(n5555) );
  NANDN U7424 ( .A(n6897), .B(n5555), .Z(\modmult_1/xin[72] ) );
  AND U7425 ( .A(m[73]), .B(n4368), .Z(n6893) );
  NANDN U7426 ( .A(start_in[0]), .B(\modmult_1/xreg[73] ), .Z(n5557) );
  NANDN U7427 ( .A(n5643), .B(creg[73]), .Z(n5556) );
  AND U7428 ( .A(n5557), .B(n5556), .Z(n5558) );
  NANDN U7429 ( .A(n6893), .B(n5558), .Z(\modmult_1/xin[73] ) );
  AND U7430 ( .A(m[74]), .B(n4368), .Z(n6889) );
  NANDN U7431 ( .A(start_in[0]), .B(\modmult_1/xreg[74] ), .Z(n5560) );
  NANDN U7432 ( .A(n5643), .B(creg[74]), .Z(n5559) );
  AND U7433 ( .A(n5560), .B(n5559), .Z(n5561) );
  NANDN U7434 ( .A(n6889), .B(n5561), .Z(\modmult_1/xin[74] ) );
  AND U7435 ( .A(m[75]), .B(n4368), .Z(n6885) );
  NANDN U7436 ( .A(start_in[0]), .B(\modmult_1/xreg[75] ), .Z(n5563) );
  NANDN U7437 ( .A(n5643), .B(creg[75]), .Z(n5562) );
  AND U7438 ( .A(n5563), .B(n5562), .Z(n5564) );
  NANDN U7439 ( .A(n6885), .B(n5564), .Z(\modmult_1/xin[75] ) );
  AND U7440 ( .A(m[76]), .B(n4368), .Z(n6881) );
  NANDN U7441 ( .A(start_in[0]), .B(\modmult_1/xreg[76] ), .Z(n5566) );
  NANDN U7442 ( .A(n5643), .B(creg[76]), .Z(n5565) );
  AND U7443 ( .A(n5566), .B(n5565), .Z(n5567) );
  NANDN U7444 ( .A(n6881), .B(n5567), .Z(\modmult_1/xin[76] ) );
  AND U7445 ( .A(m[77]), .B(n4368), .Z(n6877) );
  NANDN U7446 ( .A(start_in[0]), .B(\modmult_1/xreg[77] ), .Z(n5569) );
  NANDN U7447 ( .A(n5643), .B(creg[77]), .Z(n5568) );
  AND U7448 ( .A(n5569), .B(n5568), .Z(n5570) );
  NANDN U7449 ( .A(n6877), .B(n5570), .Z(\modmult_1/xin[77] ) );
  AND U7450 ( .A(m[78]), .B(n4368), .Z(n6873) );
  NANDN U7451 ( .A(start_in[0]), .B(\modmult_1/xreg[78] ), .Z(n5572) );
  NANDN U7452 ( .A(n5643), .B(creg[78]), .Z(n5571) );
  AND U7453 ( .A(n5572), .B(n5571), .Z(n5573) );
  NANDN U7454 ( .A(n6873), .B(n5573), .Z(\modmult_1/xin[78] ) );
  AND U7455 ( .A(m[79]), .B(n4368), .Z(n6869) );
  NANDN U7456 ( .A(start_in[0]), .B(\modmult_1/xreg[79] ), .Z(n5575) );
  NANDN U7457 ( .A(n5643), .B(creg[79]), .Z(n5574) );
  AND U7458 ( .A(n5575), .B(n5574), .Z(n5576) );
  NANDN U7459 ( .A(n6869), .B(n5576), .Z(\modmult_1/xin[79] ) );
  AND U7460 ( .A(m[7]), .B(n4368), .Z(n7157) );
  NANDN U7461 ( .A(start_in[0]), .B(\modmult_1/xreg[7] ), .Z(n5578) );
  NANDN U7462 ( .A(n5643), .B(creg[7]), .Z(n5577) );
  AND U7463 ( .A(n5578), .B(n5577), .Z(n5579) );
  NANDN U7464 ( .A(n7157), .B(n5579), .Z(\modmult_1/xin[7] ) );
  AND U7465 ( .A(m[80]), .B(n4368), .Z(n6865) );
  NANDN U7466 ( .A(start_in[0]), .B(\modmult_1/xreg[80] ), .Z(n5581) );
  NANDN U7467 ( .A(n5643), .B(creg[80]), .Z(n5580) );
  AND U7468 ( .A(n5581), .B(n5580), .Z(n5582) );
  NANDN U7469 ( .A(n6865), .B(n5582), .Z(\modmult_1/xin[80] ) );
  AND U7470 ( .A(m[81]), .B(n4368), .Z(n6861) );
  NANDN U7471 ( .A(start_in[0]), .B(\modmult_1/xreg[81] ), .Z(n5584) );
  NANDN U7472 ( .A(n5643), .B(creg[81]), .Z(n5583) );
  AND U7473 ( .A(n5584), .B(n5583), .Z(n5585) );
  NANDN U7474 ( .A(n6861), .B(n5585), .Z(\modmult_1/xin[81] ) );
  AND U7475 ( .A(m[82]), .B(n4368), .Z(n6857) );
  NANDN U7476 ( .A(start_in[0]), .B(\modmult_1/xreg[82] ), .Z(n5587) );
  NANDN U7477 ( .A(n5643), .B(creg[82]), .Z(n5586) );
  AND U7478 ( .A(n5587), .B(n5586), .Z(n5588) );
  NANDN U7479 ( .A(n6857), .B(n5588), .Z(\modmult_1/xin[82] ) );
  AND U7480 ( .A(m[83]), .B(n4368), .Z(n6853) );
  NANDN U7481 ( .A(start_in[0]), .B(\modmult_1/xreg[83] ), .Z(n5590) );
  NANDN U7482 ( .A(n5643), .B(creg[83]), .Z(n5589) );
  AND U7483 ( .A(n5590), .B(n5589), .Z(n5591) );
  NANDN U7484 ( .A(n6853), .B(n5591), .Z(\modmult_1/xin[83] ) );
  AND U7485 ( .A(m[84]), .B(n4368), .Z(n6849) );
  NANDN U7486 ( .A(start_in[0]), .B(\modmult_1/xreg[84] ), .Z(n5593) );
  NANDN U7487 ( .A(n5643), .B(creg[84]), .Z(n5592) );
  AND U7488 ( .A(n5593), .B(n5592), .Z(n5594) );
  NANDN U7489 ( .A(n6849), .B(n5594), .Z(\modmult_1/xin[84] ) );
  AND U7490 ( .A(m[85]), .B(n4368), .Z(n6845) );
  NANDN U7491 ( .A(start_in[0]), .B(\modmult_1/xreg[85] ), .Z(n5596) );
  NANDN U7492 ( .A(n5643), .B(creg[85]), .Z(n5595) );
  AND U7493 ( .A(n5596), .B(n5595), .Z(n5597) );
  NANDN U7494 ( .A(n6845), .B(n5597), .Z(\modmult_1/xin[85] ) );
  AND U7495 ( .A(m[86]), .B(n4368), .Z(n6841) );
  NANDN U7496 ( .A(start_in[0]), .B(\modmult_1/xreg[86] ), .Z(n5599) );
  NANDN U7497 ( .A(n5643), .B(creg[86]), .Z(n5598) );
  AND U7498 ( .A(n5599), .B(n5598), .Z(n5600) );
  NANDN U7499 ( .A(n6841), .B(n5600), .Z(\modmult_1/xin[86] ) );
  AND U7500 ( .A(m[87]), .B(n4368), .Z(n6837) );
  NANDN U7501 ( .A(start_in[0]), .B(\modmult_1/xreg[87] ), .Z(n5602) );
  NANDN U7502 ( .A(n5643), .B(creg[87]), .Z(n5601) );
  AND U7503 ( .A(n5602), .B(n5601), .Z(n5603) );
  NANDN U7504 ( .A(n6837), .B(n5603), .Z(\modmult_1/xin[87] ) );
  AND U7505 ( .A(m[88]), .B(n4368), .Z(n6833) );
  NANDN U7506 ( .A(start_in[0]), .B(\modmult_1/xreg[88] ), .Z(n5605) );
  NANDN U7507 ( .A(n5643), .B(creg[88]), .Z(n5604) );
  AND U7508 ( .A(n5605), .B(n5604), .Z(n5606) );
  NANDN U7509 ( .A(n6833), .B(n5606), .Z(\modmult_1/xin[88] ) );
  AND U7510 ( .A(m[89]), .B(n4368), .Z(n6829) );
  NANDN U7511 ( .A(start_in[0]), .B(\modmult_1/xreg[89] ), .Z(n5608) );
  NANDN U7512 ( .A(n5643), .B(creg[89]), .Z(n5607) );
  AND U7513 ( .A(n5608), .B(n5607), .Z(n5609) );
  NANDN U7514 ( .A(n6829), .B(n5609), .Z(\modmult_1/xin[89] ) );
  AND U7515 ( .A(m[8]), .B(n4368), .Z(n7153) );
  NANDN U7516 ( .A(start_in[0]), .B(\modmult_1/xreg[8] ), .Z(n5611) );
  NANDN U7517 ( .A(n5643), .B(creg[8]), .Z(n5610) );
  AND U7518 ( .A(n5611), .B(n5610), .Z(n5612) );
  NANDN U7519 ( .A(n7153), .B(n5612), .Z(\modmult_1/xin[8] ) );
  AND U7520 ( .A(m[90]), .B(n4368), .Z(n6825) );
  NANDN U7521 ( .A(start_in[0]), .B(\modmult_1/xreg[90] ), .Z(n5614) );
  NANDN U7522 ( .A(n5643), .B(creg[90]), .Z(n5613) );
  AND U7523 ( .A(n5614), .B(n5613), .Z(n5615) );
  NANDN U7524 ( .A(n6825), .B(n5615), .Z(\modmult_1/xin[90] ) );
  AND U7525 ( .A(m[91]), .B(n4368), .Z(n6821) );
  NANDN U7526 ( .A(start_in[0]), .B(\modmult_1/xreg[91] ), .Z(n5617) );
  NANDN U7527 ( .A(n5643), .B(creg[91]), .Z(n5616) );
  AND U7528 ( .A(n5617), .B(n5616), .Z(n5618) );
  NANDN U7529 ( .A(n6821), .B(n5618), .Z(\modmult_1/xin[91] ) );
  AND U7530 ( .A(m[92]), .B(n4368), .Z(n6817) );
  NANDN U7531 ( .A(start_in[0]), .B(\modmult_1/xreg[92] ), .Z(n5620) );
  NANDN U7532 ( .A(n5643), .B(creg[92]), .Z(n5619) );
  AND U7533 ( .A(n5620), .B(n5619), .Z(n5621) );
  NANDN U7534 ( .A(n6817), .B(n5621), .Z(\modmult_1/xin[92] ) );
  AND U7535 ( .A(m[93]), .B(n4368), .Z(n6813) );
  NANDN U7536 ( .A(start_in[0]), .B(\modmult_1/xreg[93] ), .Z(n5623) );
  NANDN U7537 ( .A(n5643), .B(creg[93]), .Z(n5622) );
  AND U7538 ( .A(n5623), .B(n5622), .Z(n5624) );
  NANDN U7539 ( .A(n6813), .B(n5624), .Z(\modmult_1/xin[93] ) );
  AND U7540 ( .A(m[94]), .B(n4368), .Z(n6809) );
  NANDN U7541 ( .A(start_in[0]), .B(\modmult_1/xreg[94] ), .Z(n5626) );
  NANDN U7542 ( .A(n5643), .B(creg[94]), .Z(n5625) );
  AND U7543 ( .A(n5626), .B(n5625), .Z(n5627) );
  NANDN U7544 ( .A(n6809), .B(n5627), .Z(\modmult_1/xin[94] ) );
  AND U7545 ( .A(m[95]), .B(n4368), .Z(n6805) );
  NANDN U7546 ( .A(start_in[0]), .B(\modmult_1/xreg[95] ), .Z(n5629) );
  NANDN U7547 ( .A(n5643), .B(creg[95]), .Z(n5628) );
  AND U7548 ( .A(n5629), .B(n5628), .Z(n5630) );
  NANDN U7549 ( .A(n6805), .B(n5630), .Z(\modmult_1/xin[95] ) );
  AND U7550 ( .A(m[96]), .B(n4368), .Z(n6801) );
  NANDN U7551 ( .A(start_in[0]), .B(\modmult_1/xreg[96] ), .Z(n5632) );
  NANDN U7552 ( .A(n5643), .B(creg[96]), .Z(n5631) );
  AND U7553 ( .A(n5632), .B(n5631), .Z(n5633) );
  NANDN U7554 ( .A(n6801), .B(n5633), .Z(\modmult_1/xin[96] ) );
  AND U7555 ( .A(m[97]), .B(n4368), .Z(n6797) );
  NANDN U7556 ( .A(start_in[0]), .B(\modmult_1/xreg[97] ), .Z(n5635) );
  NANDN U7557 ( .A(n5643), .B(creg[97]), .Z(n5634) );
  AND U7558 ( .A(n5635), .B(n5634), .Z(n5636) );
  NANDN U7559 ( .A(n6797), .B(n5636), .Z(\modmult_1/xin[97] ) );
  AND U7560 ( .A(m[98]), .B(n4368), .Z(n6793) );
  NANDN U7561 ( .A(start_in[0]), .B(\modmult_1/xreg[98] ), .Z(n5638) );
  NANDN U7562 ( .A(n5643), .B(creg[98]), .Z(n5637) );
  AND U7563 ( .A(n5638), .B(n5637), .Z(n5639) );
  NANDN U7564 ( .A(n6793), .B(n5639), .Z(\modmult_1/xin[98] ) );
  AND U7565 ( .A(m[99]), .B(n4368), .Z(n6789) );
  NANDN U7566 ( .A(start_in[0]), .B(\modmult_1/xreg[99] ), .Z(n5641) );
  NANDN U7567 ( .A(n5643), .B(creg[99]), .Z(n5640) );
  AND U7568 ( .A(n5641), .B(n5640), .Z(n5642) );
  NANDN U7569 ( .A(n6789), .B(n5642), .Z(\modmult_1/xin[99] ) );
  AND U7570 ( .A(m[9]), .B(n4368), .Z(n7149) );
  NANDN U7571 ( .A(start_in[0]), .B(\modmult_1/xreg[9] ), .Z(n5645) );
  NANDN U7572 ( .A(n5643), .B(creg[9]), .Z(n5644) );
  AND U7573 ( .A(n5645), .B(n5644), .Z(n5646) );
  NANDN U7574 ( .A(n7149), .B(n5646), .Z(\modmult_1/xin[9] ) );
  ANDN U7575 ( .B(\modmult_1/zreg[0] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][0] ) );
  ANDN U7576 ( .B(\modmult_1/zreg[100] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][100] ) );
  ANDN U7577 ( .B(\modmult_1/zreg[101] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][101] ) );
  ANDN U7578 ( .B(\modmult_1/zreg[102] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][102] ) );
  ANDN U7579 ( .B(\modmult_1/zreg[103] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][103] ) );
  ANDN U7580 ( .B(\modmult_1/zreg[104] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][104] ) );
  ANDN U7581 ( .B(\modmult_1/zreg[105] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][105] ) );
  ANDN U7582 ( .B(\modmult_1/zreg[106] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][106] ) );
  ANDN U7583 ( .B(\modmult_1/zreg[107] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][107] ) );
  ANDN U7584 ( .B(\modmult_1/zreg[108] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][108] ) );
  ANDN U7585 ( .B(\modmult_1/zreg[109] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][109] ) );
  ANDN U7586 ( .B(\modmult_1/zreg[10] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][10] ) );
  ANDN U7587 ( .B(\modmult_1/zreg[110] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][110] ) );
  ANDN U7588 ( .B(\modmult_1/zreg[111] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][111] ) );
  ANDN U7589 ( .B(\modmult_1/zreg[112] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][112] ) );
  ANDN U7590 ( .B(\modmult_1/zreg[113] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][113] ) );
  ANDN U7591 ( .B(\modmult_1/zreg[114] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][114] ) );
  ANDN U7592 ( .B(\modmult_1/zreg[115] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][115] ) );
  ANDN U7593 ( .B(\modmult_1/zreg[116] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][116] ) );
  ANDN U7594 ( .B(\modmult_1/zreg[117] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][117] ) );
  ANDN U7595 ( .B(\modmult_1/zreg[118] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][118] ) );
  ANDN U7596 ( .B(\modmult_1/zreg[119] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][119] ) );
  ANDN U7597 ( .B(\modmult_1/zreg[11] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][11] ) );
  ANDN U7598 ( .B(\modmult_1/zreg[120] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][120] ) );
  ANDN U7599 ( .B(\modmult_1/zreg[121] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][121] ) );
  ANDN U7600 ( .B(\modmult_1/zreg[122] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][122] ) );
  ANDN U7601 ( .B(\modmult_1/zreg[123] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][123] ) );
  ANDN U7602 ( .B(\modmult_1/zreg[124] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][124] ) );
  ANDN U7603 ( .B(\modmult_1/zreg[125] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][125] ) );
  ANDN U7604 ( .B(\modmult_1/zreg[126] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][126] ) );
  ANDN U7605 ( .B(\modmult_1/zreg[127] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][127] ) );
  ANDN U7606 ( .B(\modmult_1/zreg[128] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][128] ) );
  ANDN U7607 ( .B(\modmult_1/zreg[129] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][129] ) );
  ANDN U7608 ( .B(\modmult_1/zreg[12] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][12] ) );
  ANDN U7609 ( .B(\modmult_1/zreg[130] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][130] ) );
  ANDN U7610 ( .B(\modmult_1/zreg[131] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][131] ) );
  ANDN U7611 ( .B(\modmult_1/zreg[132] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][132] ) );
  ANDN U7612 ( .B(\modmult_1/zreg[133] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][133] ) );
  ANDN U7613 ( .B(\modmult_1/zreg[134] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][134] ) );
  ANDN U7614 ( .B(\modmult_1/zreg[135] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][135] ) );
  ANDN U7615 ( .B(\modmult_1/zreg[136] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][136] ) );
  ANDN U7616 ( .B(\modmult_1/zreg[137] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][137] ) );
  ANDN U7617 ( .B(\modmult_1/zreg[138] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][138] ) );
  ANDN U7618 ( .B(\modmult_1/zreg[139] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][139] ) );
  ANDN U7619 ( .B(\modmult_1/zreg[13] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][13] ) );
  ANDN U7620 ( .B(\modmult_1/zreg[140] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][140] ) );
  ANDN U7621 ( .B(\modmult_1/zreg[141] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][141] ) );
  ANDN U7622 ( .B(\modmult_1/zreg[142] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][142] ) );
  ANDN U7623 ( .B(\modmult_1/zreg[143] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][143] ) );
  ANDN U7624 ( .B(\modmult_1/zreg[144] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][144] ) );
  ANDN U7625 ( .B(\modmult_1/zreg[145] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][145] ) );
  ANDN U7626 ( .B(\modmult_1/zreg[146] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][146] ) );
  ANDN U7627 ( .B(\modmult_1/zreg[147] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][147] ) );
  ANDN U7628 ( .B(\modmult_1/zreg[148] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][148] ) );
  ANDN U7629 ( .B(\modmult_1/zreg[149] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][149] ) );
  ANDN U7630 ( .B(\modmult_1/zreg[14] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][14] ) );
  ANDN U7631 ( .B(\modmult_1/zreg[150] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][150] ) );
  ANDN U7632 ( .B(\modmult_1/zreg[151] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][151] ) );
  ANDN U7633 ( .B(\modmult_1/zreg[152] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][152] ) );
  ANDN U7634 ( .B(\modmult_1/zreg[153] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][153] ) );
  ANDN U7635 ( .B(\modmult_1/zreg[154] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][154] ) );
  ANDN U7636 ( .B(\modmult_1/zreg[155] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][155] ) );
  ANDN U7637 ( .B(\modmult_1/zreg[156] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][156] ) );
  ANDN U7638 ( .B(\modmult_1/zreg[157] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][157] ) );
  ANDN U7639 ( .B(\modmult_1/zreg[158] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][158] ) );
  ANDN U7640 ( .B(\modmult_1/zreg[159] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][159] ) );
  ANDN U7641 ( .B(\modmult_1/zreg[15] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][15] ) );
  ANDN U7642 ( .B(\modmult_1/zreg[160] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][160] ) );
  ANDN U7643 ( .B(\modmult_1/zreg[161] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][161] ) );
  ANDN U7644 ( .B(\modmult_1/zreg[162] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][162] ) );
  ANDN U7645 ( .B(\modmult_1/zreg[163] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][163] ) );
  ANDN U7646 ( .B(\modmult_1/zreg[164] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][164] ) );
  ANDN U7647 ( .B(\modmult_1/zreg[165] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][165] ) );
  ANDN U7648 ( .B(\modmult_1/zreg[166] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][166] ) );
  ANDN U7649 ( .B(\modmult_1/zreg[167] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][167] ) );
  ANDN U7650 ( .B(\modmult_1/zreg[168] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][168] ) );
  ANDN U7651 ( .B(\modmult_1/zreg[169] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][169] ) );
  ANDN U7652 ( .B(\modmult_1/zreg[16] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][16] ) );
  ANDN U7653 ( .B(\modmult_1/zreg[170] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][170] ) );
  ANDN U7654 ( .B(\modmult_1/zreg[171] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][171] ) );
  ANDN U7655 ( .B(\modmult_1/zreg[172] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][172] ) );
  ANDN U7656 ( .B(\modmult_1/zreg[173] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][173] ) );
  ANDN U7657 ( .B(\modmult_1/zreg[174] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][174] ) );
  ANDN U7658 ( .B(\modmult_1/zreg[175] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][175] ) );
  ANDN U7659 ( .B(\modmult_1/zreg[176] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][176] ) );
  ANDN U7660 ( .B(\modmult_1/zreg[177] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][177] ) );
  ANDN U7661 ( .B(\modmult_1/zreg[178] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][178] ) );
  ANDN U7662 ( .B(\modmult_1/zreg[179] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][179] ) );
  ANDN U7663 ( .B(\modmult_1/zreg[17] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][17] ) );
  ANDN U7664 ( .B(\modmult_1/zreg[180] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][180] ) );
  ANDN U7665 ( .B(\modmult_1/zreg[181] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][181] ) );
  ANDN U7666 ( .B(\modmult_1/zreg[182] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][182] ) );
  ANDN U7667 ( .B(\modmult_1/zreg[183] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][183] ) );
  ANDN U7668 ( .B(\modmult_1/zreg[184] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][184] ) );
  ANDN U7669 ( .B(\modmult_1/zreg[185] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][185] ) );
  ANDN U7670 ( .B(\modmult_1/zreg[186] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][186] ) );
  ANDN U7671 ( .B(\modmult_1/zreg[187] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][187] ) );
  ANDN U7672 ( .B(\modmult_1/zreg[188] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][188] ) );
  ANDN U7673 ( .B(\modmult_1/zreg[189] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][189] ) );
  ANDN U7674 ( .B(\modmult_1/zreg[18] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][18] ) );
  ANDN U7675 ( .B(\modmult_1/zreg[190] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][190] ) );
  ANDN U7676 ( .B(\modmult_1/zreg[191] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][191] ) );
  ANDN U7677 ( .B(\modmult_1/zreg[192] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][192] ) );
  ANDN U7678 ( .B(\modmult_1/zreg[193] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][193] ) );
  ANDN U7679 ( .B(\modmult_1/zreg[194] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][194] ) );
  ANDN U7680 ( .B(\modmult_1/zreg[195] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][195] ) );
  ANDN U7681 ( .B(\modmult_1/zreg[196] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][196] ) );
  ANDN U7682 ( .B(\modmult_1/zreg[197] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][197] ) );
  ANDN U7683 ( .B(\modmult_1/zreg[198] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][198] ) );
  ANDN U7684 ( .B(\modmult_1/zreg[199] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][199] ) );
  ANDN U7685 ( .B(\modmult_1/zreg[19] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][19] ) );
  ANDN U7686 ( .B(\modmult_1/zreg[1] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][1] ) );
  ANDN U7687 ( .B(\modmult_1/zreg[200] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][200] ) );
  ANDN U7688 ( .B(\modmult_1/zreg[201] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][201] ) );
  ANDN U7689 ( .B(\modmult_1/zreg[202] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][202] ) );
  ANDN U7690 ( .B(\modmult_1/zreg[203] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][203] ) );
  ANDN U7691 ( .B(\modmult_1/zreg[204] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][204] ) );
  ANDN U7692 ( .B(\modmult_1/zreg[205] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][205] ) );
  ANDN U7693 ( .B(\modmult_1/zreg[206] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][206] ) );
  ANDN U7694 ( .B(\modmult_1/zreg[207] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][207] ) );
  ANDN U7695 ( .B(\modmult_1/zreg[208] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][208] ) );
  ANDN U7696 ( .B(\modmult_1/zreg[209] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][209] ) );
  ANDN U7697 ( .B(\modmult_1/zreg[20] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][20] ) );
  ANDN U7698 ( .B(\modmult_1/zreg[210] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][210] ) );
  ANDN U7699 ( .B(\modmult_1/zreg[211] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][211] ) );
  ANDN U7700 ( .B(\modmult_1/zreg[212] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][212] ) );
  ANDN U7701 ( .B(\modmult_1/zreg[213] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][213] ) );
  ANDN U7702 ( .B(\modmult_1/zreg[214] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][214] ) );
  ANDN U7703 ( .B(\modmult_1/zreg[215] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][215] ) );
  ANDN U7704 ( .B(\modmult_1/zreg[216] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][216] ) );
  ANDN U7705 ( .B(\modmult_1/zreg[217] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][217] ) );
  ANDN U7706 ( .B(\modmult_1/zreg[218] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][218] ) );
  ANDN U7707 ( .B(\modmult_1/zreg[219] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][219] ) );
  ANDN U7708 ( .B(\modmult_1/zreg[21] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][21] ) );
  ANDN U7709 ( .B(\modmult_1/zreg[220] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][220] ) );
  ANDN U7710 ( .B(\modmult_1/zreg[221] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][221] ) );
  ANDN U7711 ( .B(\modmult_1/zreg[222] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][222] ) );
  ANDN U7712 ( .B(\modmult_1/zreg[223] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][223] ) );
  ANDN U7713 ( .B(\modmult_1/zreg[224] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][224] ) );
  ANDN U7714 ( .B(\modmult_1/zreg[225] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][225] ) );
  ANDN U7715 ( .B(\modmult_1/zreg[226] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][226] ) );
  ANDN U7716 ( .B(\modmult_1/zreg[227] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][227] ) );
  ANDN U7717 ( .B(\modmult_1/zreg[228] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][228] ) );
  ANDN U7718 ( .B(\modmult_1/zreg[229] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][229] ) );
  ANDN U7719 ( .B(\modmult_1/zreg[22] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][22] ) );
  ANDN U7720 ( .B(\modmult_1/zreg[230] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][230] ) );
  ANDN U7721 ( .B(\modmult_1/zreg[231] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][231] ) );
  ANDN U7722 ( .B(\modmult_1/zreg[232] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][232] ) );
  ANDN U7723 ( .B(\modmult_1/zreg[233] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][233] ) );
  ANDN U7724 ( .B(\modmult_1/zreg[234] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][234] ) );
  ANDN U7725 ( .B(\modmult_1/zreg[235] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][235] ) );
  ANDN U7726 ( .B(\modmult_1/zreg[236] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][236] ) );
  ANDN U7727 ( .B(\modmult_1/zreg[237] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][237] ) );
  ANDN U7728 ( .B(\modmult_1/zreg[238] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][238] ) );
  ANDN U7729 ( .B(\modmult_1/zreg[239] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][239] ) );
  ANDN U7730 ( .B(\modmult_1/zreg[23] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][23] ) );
  ANDN U7731 ( .B(\modmult_1/zreg[240] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][240] ) );
  ANDN U7732 ( .B(\modmult_1/zreg[241] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][241] ) );
  ANDN U7733 ( .B(\modmult_1/zreg[242] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][242] ) );
  ANDN U7734 ( .B(\modmult_1/zreg[243] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][243] ) );
  ANDN U7735 ( .B(\modmult_1/zreg[244] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][244] ) );
  ANDN U7736 ( .B(\modmult_1/zreg[245] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][245] ) );
  ANDN U7737 ( .B(\modmult_1/zreg[246] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][246] ) );
  ANDN U7738 ( .B(\modmult_1/zreg[247] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][247] ) );
  ANDN U7739 ( .B(\modmult_1/zreg[248] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][248] ) );
  ANDN U7740 ( .B(\modmult_1/zreg[249] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][249] ) );
  ANDN U7741 ( .B(\modmult_1/zreg[24] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][24] ) );
  ANDN U7742 ( .B(\modmult_1/zreg[250] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][250] ) );
  ANDN U7743 ( .B(\modmult_1/zreg[251] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][251] ) );
  ANDN U7744 ( .B(\modmult_1/zreg[252] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][252] ) );
  ANDN U7745 ( .B(\modmult_1/zreg[253] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][253] ) );
  ANDN U7746 ( .B(\modmult_1/zreg[254] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][254] ) );
  ANDN U7747 ( .B(\modmult_1/zreg[255] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][255] ) );
  ANDN U7748 ( .B(\modmult_1/zreg[256] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][256] ) );
  ANDN U7749 ( .B(\modmult_1/zreg[25] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][25] ) );
  ANDN U7750 ( .B(\modmult_1/zreg[26] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][26] ) );
  ANDN U7751 ( .B(\modmult_1/zreg[27] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][27] ) );
  ANDN U7752 ( .B(\modmult_1/zreg[28] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][28] ) );
  ANDN U7753 ( .B(\modmult_1/zreg[29] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][29] ) );
  ANDN U7754 ( .B(\modmult_1/zreg[2] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][2] ) );
  ANDN U7755 ( .B(\modmult_1/zreg[30] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][30] ) );
  ANDN U7756 ( .B(\modmult_1/zreg[31] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][31] ) );
  ANDN U7757 ( .B(\modmult_1/zreg[32] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][32] ) );
  ANDN U7758 ( .B(\modmult_1/zreg[33] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][33] ) );
  ANDN U7759 ( .B(\modmult_1/zreg[34] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][34] ) );
  ANDN U7760 ( .B(\modmult_1/zreg[35] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][35] ) );
  ANDN U7761 ( .B(\modmult_1/zreg[36] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][36] ) );
  ANDN U7762 ( .B(\modmult_1/zreg[37] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][37] ) );
  ANDN U7763 ( .B(\modmult_1/zreg[38] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][38] ) );
  ANDN U7764 ( .B(\modmult_1/zreg[39] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][39] ) );
  ANDN U7765 ( .B(\modmult_1/zreg[3] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][3] ) );
  ANDN U7766 ( .B(\modmult_1/zreg[40] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][40] ) );
  ANDN U7767 ( .B(\modmult_1/zreg[41] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][41] ) );
  ANDN U7768 ( .B(\modmult_1/zreg[42] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][42] ) );
  ANDN U7769 ( .B(\modmult_1/zreg[43] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][43] ) );
  ANDN U7770 ( .B(\modmult_1/zreg[44] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][44] ) );
  ANDN U7771 ( .B(\modmult_1/zreg[45] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][45] ) );
  ANDN U7772 ( .B(\modmult_1/zreg[46] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][46] ) );
  ANDN U7773 ( .B(\modmult_1/zreg[47] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][47] ) );
  ANDN U7774 ( .B(\modmult_1/zreg[48] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][48] ) );
  ANDN U7775 ( .B(\modmult_1/zreg[49] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][49] ) );
  ANDN U7776 ( .B(\modmult_1/zreg[4] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][4] ) );
  ANDN U7777 ( .B(\modmult_1/zreg[50] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][50] ) );
  ANDN U7778 ( .B(\modmult_1/zreg[51] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][51] ) );
  ANDN U7779 ( .B(\modmult_1/zreg[52] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][52] ) );
  ANDN U7780 ( .B(\modmult_1/zreg[53] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][53] ) );
  ANDN U7781 ( .B(\modmult_1/zreg[54] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][54] ) );
  ANDN U7782 ( .B(\modmult_1/zreg[55] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][55] ) );
  ANDN U7783 ( .B(\modmult_1/zreg[56] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][56] ) );
  ANDN U7784 ( .B(\modmult_1/zreg[57] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][57] ) );
  ANDN U7785 ( .B(\modmult_1/zreg[58] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][58] ) );
  ANDN U7786 ( .B(\modmult_1/zreg[59] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][59] ) );
  ANDN U7787 ( .B(\modmult_1/zreg[5] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][5] ) );
  ANDN U7788 ( .B(\modmult_1/zreg[60] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][60] ) );
  ANDN U7789 ( .B(\modmult_1/zreg[61] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][61] ) );
  ANDN U7790 ( .B(\modmult_1/zreg[62] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][62] ) );
  ANDN U7791 ( .B(\modmult_1/zreg[63] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][63] ) );
  ANDN U7792 ( .B(\modmult_1/zreg[64] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][64] ) );
  ANDN U7793 ( .B(\modmult_1/zreg[65] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][65] ) );
  ANDN U7794 ( .B(\modmult_1/zreg[66] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][66] ) );
  ANDN U7795 ( .B(\modmult_1/zreg[67] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][67] ) );
  ANDN U7796 ( .B(\modmult_1/zreg[68] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][68] ) );
  ANDN U7797 ( .B(\modmult_1/zreg[69] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][69] ) );
  ANDN U7798 ( .B(\modmult_1/zreg[6] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][6] ) );
  ANDN U7799 ( .B(\modmult_1/zreg[70] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][70] ) );
  ANDN U7800 ( .B(\modmult_1/zreg[71] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][71] ) );
  ANDN U7801 ( .B(\modmult_1/zreg[72] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][72] ) );
  ANDN U7802 ( .B(\modmult_1/zreg[73] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][73] ) );
  ANDN U7803 ( .B(\modmult_1/zreg[74] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][74] ) );
  ANDN U7804 ( .B(\modmult_1/zreg[75] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][75] ) );
  ANDN U7805 ( .B(\modmult_1/zreg[76] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][76] ) );
  ANDN U7806 ( .B(\modmult_1/zreg[77] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][77] ) );
  ANDN U7807 ( .B(\modmult_1/zreg[78] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][78] ) );
  ANDN U7808 ( .B(\modmult_1/zreg[79] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][79] ) );
  ANDN U7809 ( .B(\modmult_1/zreg[7] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][7] ) );
  ANDN U7810 ( .B(\modmult_1/zreg[80] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][80] ) );
  ANDN U7811 ( .B(\modmult_1/zreg[81] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][81] ) );
  ANDN U7812 ( .B(\modmult_1/zreg[82] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][82] ) );
  ANDN U7813 ( .B(\modmult_1/zreg[83] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][83] ) );
  ANDN U7814 ( .B(\modmult_1/zreg[84] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][84] ) );
  ANDN U7815 ( .B(\modmult_1/zreg[85] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][85] ) );
  ANDN U7816 ( .B(\modmult_1/zreg[86] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][86] ) );
  ANDN U7817 ( .B(\modmult_1/zreg[87] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][87] ) );
  ANDN U7818 ( .B(\modmult_1/zreg[88] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][88] ) );
  ANDN U7819 ( .B(\modmult_1/zreg[89] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][89] ) );
  ANDN U7820 ( .B(\modmult_1/zreg[8] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][8] ) );
  ANDN U7821 ( .B(\modmult_1/zreg[90] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][90] ) );
  ANDN U7822 ( .B(\modmult_1/zreg[91] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][91] ) );
  ANDN U7823 ( .B(\modmult_1/zreg[92] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][92] ) );
  ANDN U7824 ( .B(\modmult_1/zreg[93] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][93] ) );
  ANDN U7825 ( .B(\modmult_1/zreg[94] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][94] ) );
  ANDN U7826 ( .B(\modmult_1/zreg[95] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][95] ) );
  ANDN U7827 ( .B(\modmult_1/zreg[96] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][96] ) );
  ANDN U7828 ( .B(\modmult_1/zreg[97] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][97] ) );
  ANDN U7829 ( .B(\modmult_1/zreg[98] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][98] ) );
  ANDN U7830 ( .B(\modmult_1/zreg[99] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][99] ) );
  ANDN U7831 ( .B(\modmult_1/zreg[9] ), .A(start_in[0]), .Z(
        \modmult_1/zin[0][9] ) );
  ANDN U7832 ( .B(start_reg[100]), .A(n4368), .Z(start_in[100]) );
  ANDN U7833 ( .B(start_reg[101]), .A(n4368), .Z(start_in[101]) );
  ANDN U7834 ( .B(start_reg[102]), .A(n4368), .Z(start_in[102]) );
  ANDN U7835 ( .B(start_reg[103]), .A(n4368), .Z(start_in[103]) );
  ANDN U7836 ( .B(start_reg[104]), .A(n4368), .Z(start_in[104]) );
  ANDN U7837 ( .B(start_reg[105]), .A(n4368), .Z(start_in[105]) );
  ANDN U7838 ( .B(start_reg[106]), .A(n4368), .Z(start_in[106]) );
  ANDN U7839 ( .B(start_reg[107]), .A(n4368), .Z(start_in[107]) );
  ANDN U7840 ( .B(start_reg[108]), .A(n4368), .Z(start_in[108]) );
  ANDN U7841 ( .B(start_reg[109]), .A(n4368), .Z(start_in[109]) );
  ANDN U7842 ( .B(start_reg[10]), .A(n4368), .Z(start_in[10]) );
  ANDN U7843 ( .B(start_reg[110]), .A(n4368), .Z(start_in[110]) );
  ANDN U7844 ( .B(start_reg[111]), .A(n4368), .Z(start_in[111]) );
  ANDN U7845 ( .B(start_reg[112]), .A(n4368), .Z(start_in[112]) );
  ANDN U7846 ( .B(start_reg[113]), .A(n4368), .Z(start_in[113]) );
  ANDN U7847 ( .B(start_reg[114]), .A(n4368), .Z(start_in[114]) );
  ANDN U7848 ( .B(start_reg[115]), .A(n4368), .Z(start_in[115]) );
  ANDN U7849 ( .B(start_reg[116]), .A(n4368), .Z(start_in[116]) );
  ANDN U7850 ( .B(start_reg[117]), .A(n4368), .Z(start_in[117]) );
  ANDN U7851 ( .B(start_reg[118]), .A(n4368), .Z(start_in[118]) );
  ANDN U7852 ( .B(start_reg[119]), .A(n4368), .Z(start_in[119]) );
  ANDN U7853 ( .B(start_reg[11]), .A(n4368), .Z(start_in[11]) );
  ANDN U7854 ( .B(start_reg[120]), .A(n4368), .Z(start_in[120]) );
  ANDN U7855 ( .B(start_reg[121]), .A(n4368), .Z(start_in[121]) );
  ANDN U7856 ( .B(start_reg[122]), .A(n4368), .Z(start_in[122]) );
  ANDN U7857 ( .B(start_reg[123]), .A(n4368), .Z(start_in[123]) );
  ANDN U7858 ( .B(start_reg[124]), .A(n4368), .Z(start_in[124]) );
  ANDN U7859 ( .B(start_reg[125]), .A(n4368), .Z(start_in[125]) );
  ANDN U7860 ( .B(start_reg[126]), .A(n4368), .Z(start_in[126]) );
  ANDN U7861 ( .B(start_reg[12]), .A(n4368), .Z(start_in[12]) );
  ANDN U7862 ( .B(start_reg[13]), .A(n4368), .Z(start_in[13]) );
  ANDN U7863 ( .B(start_reg[14]), .A(n4368), .Z(start_in[14]) );
  ANDN U7864 ( .B(start_reg[15]), .A(n4368), .Z(start_in[15]) );
  ANDN U7865 ( .B(start_reg[16]), .A(n4368), .Z(start_in[16]) );
  ANDN U7866 ( .B(start_reg[17]), .A(n4368), .Z(start_in[17]) );
  ANDN U7867 ( .B(start_reg[18]), .A(n4368), .Z(start_in[18]) );
  ANDN U7868 ( .B(start_reg[19]), .A(n4368), .Z(start_in[19]) );
  ANDN U7869 ( .B(start_reg[1]), .A(n4368), .Z(start_in[1]) );
  ANDN U7870 ( .B(start_reg[20]), .A(n4368), .Z(start_in[20]) );
  ANDN U7871 ( .B(start_reg[21]), .A(n4368), .Z(start_in[21]) );
  ANDN U7872 ( .B(start_reg[22]), .A(n4368), .Z(start_in[22]) );
  ANDN U7873 ( .B(start_reg[23]), .A(n4368), .Z(start_in[23]) );
  ANDN U7874 ( .B(start_reg[24]), .A(n4368), .Z(start_in[24]) );
  ANDN U7875 ( .B(start_reg[25]), .A(n4368), .Z(start_in[25]) );
  ANDN U7876 ( .B(start_reg[26]), .A(n4368), .Z(start_in[26]) );
  ANDN U7877 ( .B(start_reg[27]), .A(n4368), .Z(start_in[27]) );
  ANDN U7878 ( .B(start_reg[28]), .A(n4368), .Z(start_in[28]) );
  ANDN U7879 ( .B(start_reg[29]), .A(n4368), .Z(start_in[29]) );
  ANDN U7880 ( .B(start_reg[2]), .A(n4368), .Z(start_in[2]) );
  ANDN U7881 ( .B(start_reg[30]), .A(n4368), .Z(start_in[30]) );
  ANDN U7882 ( .B(start_reg[31]), .A(n4368), .Z(start_in[31]) );
  ANDN U7883 ( .B(start_reg[32]), .A(n4368), .Z(start_in[32]) );
  ANDN U7884 ( .B(start_reg[33]), .A(n4368), .Z(start_in[33]) );
  ANDN U7885 ( .B(start_reg[34]), .A(n4368), .Z(start_in[34]) );
  ANDN U7886 ( .B(start_reg[35]), .A(n4368), .Z(start_in[35]) );
  ANDN U7887 ( .B(start_reg[36]), .A(n4368), .Z(start_in[36]) );
  ANDN U7888 ( .B(start_reg[37]), .A(n4368), .Z(start_in[37]) );
  ANDN U7889 ( .B(start_reg[38]), .A(n4368), .Z(start_in[38]) );
  ANDN U7890 ( .B(start_reg[39]), .A(n4368), .Z(start_in[39]) );
  ANDN U7891 ( .B(start_reg[3]), .A(n4368), .Z(start_in[3]) );
  ANDN U7892 ( .B(start_reg[40]), .A(n4368), .Z(start_in[40]) );
  ANDN U7893 ( .B(start_reg[41]), .A(n4368), .Z(start_in[41]) );
  ANDN U7894 ( .B(start_reg[42]), .A(n4368), .Z(start_in[42]) );
  ANDN U7895 ( .B(start_reg[43]), .A(n4368), .Z(start_in[43]) );
  ANDN U7896 ( .B(start_reg[44]), .A(n4368), .Z(start_in[44]) );
  ANDN U7897 ( .B(start_reg[45]), .A(n4368), .Z(start_in[45]) );
  ANDN U7898 ( .B(start_reg[46]), .A(n4368), .Z(start_in[46]) );
  ANDN U7899 ( .B(start_reg[47]), .A(n4368), .Z(start_in[47]) );
  ANDN U7900 ( .B(start_reg[48]), .A(n4368), .Z(start_in[48]) );
  ANDN U7901 ( .B(start_reg[49]), .A(n4368), .Z(start_in[49]) );
  ANDN U7902 ( .B(start_reg[4]), .A(n4368), .Z(start_in[4]) );
  ANDN U7903 ( .B(start_reg[50]), .A(n4368), .Z(start_in[50]) );
  ANDN U7904 ( .B(start_reg[51]), .A(n4368), .Z(start_in[51]) );
  ANDN U7905 ( .B(start_reg[52]), .A(n4368), .Z(start_in[52]) );
  ANDN U7906 ( .B(start_reg[53]), .A(n4368), .Z(start_in[53]) );
  ANDN U7907 ( .B(start_reg[54]), .A(n4368), .Z(start_in[54]) );
  ANDN U7908 ( .B(start_reg[55]), .A(n4368), .Z(start_in[55]) );
  ANDN U7909 ( .B(start_reg[56]), .A(n4368), .Z(start_in[56]) );
  ANDN U7910 ( .B(start_reg[57]), .A(n4368), .Z(start_in[57]) );
  ANDN U7911 ( .B(start_reg[58]), .A(n4368), .Z(start_in[58]) );
  ANDN U7912 ( .B(start_reg[59]), .A(n4368), .Z(start_in[59]) );
  ANDN U7913 ( .B(start_reg[5]), .A(n4368), .Z(start_in[5]) );
  ANDN U7914 ( .B(start_reg[60]), .A(n4368), .Z(start_in[60]) );
  ANDN U7915 ( .B(start_reg[61]), .A(n4368), .Z(start_in[61]) );
  ANDN U7916 ( .B(start_reg[62]), .A(n4368), .Z(start_in[62]) );
  ANDN U7917 ( .B(start_reg[63]), .A(n4368), .Z(start_in[63]) );
  ANDN U7918 ( .B(start_reg[64]), .A(n4368), .Z(start_in[64]) );
  ANDN U7919 ( .B(start_reg[65]), .A(n4368), .Z(start_in[65]) );
  ANDN U7920 ( .B(start_reg[66]), .A(n4368), .Z(start_in[66]) );
  ANDN U7921 ( .B(start_reg[67]), .A(n4368), .Z(start_in[67]) );
  ANDN U7922 ( .B(start_reg[68]), .A(n4368), .Z(start_in[68]) );
  ANDN U7923 ( .B(start_reg[69]), .A(n4368), .Z(start_in[69]) );
  ANDN U7924 ( .B(start_reg[6]), .A(n4368), .Z(start_in[6]) );
  ANDN U7925 ( .B(start_reg[70]), .A(n4368), .Z(start_in[70]) );
  ANDN U7926 ( .B(start_reg[71]), .A(n4368), .Z(start_in[71]) );
  ANDN U7927 ( .B(start_reg[72]), .A(n4368), .Z(start_in[72]) );
  ANDN U7928 ( .B(start_reg[73]), .A(n4368), .Z(start_in[73]) );
  ANDN U7929 ( .B(start_reg[74]), .A(n4368), .Z(start_in[74]) );
  ANDN U7930 ( .B(start_reg[75]), .A(n4368), .Z(start_in[75]) );
  ANDN U7931 ( .B(start_reg[76]), .A(n4368), .Z(start_in[76]) );
  ANDN U7932 ( .B(start_reg[77]), .A(n4368), .Z(start_in[77]) );
  ANDN U7933 ( .B(start_reg[78]), .A(n4368), .Z(start_in[78]) );
  ANDN U7934 ( .B(start_reg[79]), .A(n4368), .Z(start_in[79]) );
  ANDN U7935 ( .B(start_reg[7]), .A(n4368), .Z(start_in[7]) );
  ANDN U7936 ( .B(start_reg[80]), .A(n4368), .Z(start_in[80]) );
  ANDN U7937 ( .B(start_reg[81]), .A(n4368), .Z(start_in[81]) );
  ANDN U7938 ( .B(start_reg[82]), .A(n4368), .Z(start_in[82]) );
  ANDN U7939 ( .B(start_reg[83]), .A(n4368), .Z(start_in[83]) );
  ANDN U7940 ( .B(start_reg[84]), .A(n4368), .Z(start_in[84]) );
  ANDN U7941 ( .B(start_reg[85]), .A(n4368), .Z(start_in[85]) );
  ANDN U7942 ( .B(start_reg[86]), .A(n4368), .Z(start_in[86]) );
  ANDN U7943 ( .B(start_reg[87]), .A(n4368), .Z(start_in[87]) );
  ANDN U7944 ( .B(start_reg[88]), .A(n4368), .Z(start_in[88]) );
  ANDN U7945 ( .B(start_reg[89]), .A(n4368), .Z(start_in[89]) );
  ANDN U7946 ( .B(start_reg[8]), .A(n4368), .Z(start_in[8]) );
  ANDN U7947 ( .B(start_reg[90]), .A(n4368), .Z(start_in[90]) );
  ANDN U7948 ( .B(start_reg[91]), .A(n4368), .Z(start_in[91]) );
  ANDN U7949 ( .B(start_reg[92]), .A(n4368), .Z(start_in[92]) );
  ANDN U7950 ( .B(start_reg[93]), .A(n4368), .Z(start_in[93]) );
  ANDN U7951 ( .B(start_reg[94]), .A(n4368), .Z(start_in[94]) );
  ANDN U7952 ( .B(start_reg[95]), .A(n4368), .Z(start_in[95]) );
  ANDN U7953 ( .B(start_reg[96]), .A(n4368), .Z(start_in[96]) );
  ANDN U7954 ( .B(start_reg[97]), .A(n4368), .Z(start_in[97]) );
  ANDN U7955 ( .B(start_reg[98]), .A(n4368), .Z(start_in[98]) );
  ANDN U7956 ( .B(start_reg[99]), .A(n4368), .Z(start_in[99]) );
  ANDN U7957 ( .B(start_reg[9]), .A(n4368), .Z(start_in[9]) );
  NOR U7958 ( .A(n4368), .B(mul_pow), .Z(n6157) );
  NANDN U7959 ( .A(n4366), .B(creg[0]), .Z(n5648) );
  NANDN U7960 ( .A(n6157), .B(m[0]), .Z(n5647) );
  NAND U7961 ( .A(n5648), .B(n5647), .Z(y[0]) );
  NANDN U7962 ( .A(n4366), .B(creg[100]), .Z(n5650) );
  NANDN U7963 ( .A(n6157), .B(m[100]), .Z(n5649) );
  NAND U7964 ( .A(n5650), .B(n5649), .Z(y[100]) );
  NANDN U7965 ( .A(n4366), .B(creg[101]), .Z(n5652) );
  NANDN U7966 ( .A(n6157), .B(m[101]), .Z(n5651) );
  NAND U7967 ( .A(n5652), .B(n5651), .Z(y[101]) );
  NANDN U7968 ( .A(n4366), .B(creg[102]), .Z(n5654) );
  NANDN U7969 ( .A(n6157), .B(m[102]), .Z(n5653) );
  NAND U7970 ( .A(n5654), .B(n5653), .Z(y[102]) );
  NANDN U7971 ( .A(n4366), .B(creg[103]), .Z(n5656) );
  NANDN U7972 ( .A(n6157), .B(m[103]), .Z(n5655) );
  NAND U7973 ( .A(n5656), .B(n5655), .Z(y[103]) );
  NANDN U7974 ( .A(n4366), .B(creg[104]), .Z(n5658) );
  NANDN U7975 ( .A(n6157), .B(m[104]), .Z(n5657) );
  NAND U7976 ( .A(n5658), .B(n5657), .Z(y[104]) );
  NANDN U7977 ( .A(n4366), .B(creg[105]), .Z(n5660) );
  NANDN U7978 ( .A(n6157), .B(m[105]), .Z(n5659) );
  NAND U7979 ( .A(n5660), .B(n5659), .Z(y[105]) );
  NANDN U7980 ( .A(n4366), .B(creg[106]), .Z(n5662) );
  NANDN U7981 ( .A(n6157), .B(m[106]), .Z(n5661) );
  NAND U7982 ( .A(n5662), .B(n5661), .Z(y[106]) );
  NANDN U7983 ( .A(n4366), .B(creg[107]), .Z(n5664) );
  NANDN U7984 ( .A(n6157), .B(m[107]), .Z(n5663) );
  NAND U7985 ( .A(n5664), .B(n5663), .Z(y[107]) );
  NANDN U7986 ( .A(n4366), .B(creg[108]), .Z(n5666) );
  NANDN U7987 ( .A(n6157), .B(m[108]), .Z(n5665) );
  NAND U7988 ( .A(n5666), .B(n5665), .Z(y[108]) );
  NANDN U7989 ( .A(n4366), .B(creg[109]), .Z(n5668) );
  NANDN U7990 ( .A(n6157), .B(m[109]), .Z(n5667) );
  NAND U7991 ( .A(n5668), .B(n5667), .Z(y[109]) );
  NANDN U7992 ( .A(n4366), .B(creg[10]), .Z(n5670) );
  NANDN U7993 ( .A(n6157), .B(m[10]), .Z(n5669) );
  NAND U7994 ( .A(n5670), .B(n5669), .Z(y[10]) );
  NANDN U7995 ( .A(n4366), .B(creg[110]), .Z(n5672) );
  NANDN U7996 ( .A(n6157), .B(m[110]), .Z(n5671) );
  NAND U7997 ( .A(n5672), .B(n5671), .Z(y[110]) );
  NANDN U7998 ( .A(n4366), .B(creg[111]), .Z(n5674) );
  NANDN U7999 ( .A(n6157), .B(m[111]), .Z(n5673) );
  NAND U8000 ( .A(n5674), .B(n5673), .Z(y[111]) );
  NANDN U8001 ( .A(n4366), .B(creg[112]), .Z(n5676) );
  NANDN U8002 ( .A(n6157), .B(m[112]), .Z(n5675) );
  NAND U8003 ( .A(n5676), .B(n5675), .Z(y[112]) );
  NANDN U8004 ( .A(n4366), .B(creg[113]), .Z(n5678) );
  NANDN U8005 ( .A(n6157), .B(m[113]), .Z(n5677) );
  NAND U8006 ( .A(n5678), .B(n5677), .Z(y[113]) );
  NANDN U8007 ( .A(n4366), .B(creg[114]), .Z(n5680) );
  NANDN U8008 ( .A(n6157), .B(m[114]), .Z(n5679) );
  NAND U8009 ( .A(n5680), .B(n5679), .Z(y[114]) );
  NANDN U8010 ( .A(n4366), .B(creg[115]), .Z(n5682) );
  NANDN U8011 ( .A(n6157), .B(m[115]), .Z(n5681) );
  NAND U8012 ( .A(n5682), .B(n5681), .Z(y[115]) );
  NANDN U8013 ( .A(n4366), .B(creg[116]), .Z(n5684) );
  NANDN U8014 ( .A(n6157), .B(m[116]), .Z(n5683) );
  NAND U8015 ( .A(n5684), .B(n5683), .Z(y[116]) );
  NANDN U8016 ( .A(n4366), .B(creg[117]), .Z(n5686) );
  NANDN U8017 ( .A(n6157), .B(m[117]), .Z(n5685) );
  NAND U8018 ( .A(n5686), .B(n5685), .Z(y[117]) );
  NANDN U8019 ( .A(n4366), .B(creg[118]), .Z(n5688) );
  NANDN U8020 ( .A(n6157), .B(m[118]), .Z(n5687) );
  NAND U8021 ( .A(n5688), .B(n5687), .Z(y[118]) );
  NANDN U8022 ( .A(n4366), .B(creg[119]), .Z(n5690) );
  NANDN U8023 ( .A(n6157), .B(m[119]), .Z(n5689) );
  NAND U8024 ( .A(n5690), .B(n5689), .Z(y[119]) );
  NANDN U8025 ( .A(n4366), .B(creg[11]), .Z(n5692) );
  NANDN U8026 ( .A(n6157), .B(m[11]), .Z(n5691) );
  NAND U8027 ( .A(n5692), .B(n5691), .Z(y[11]) );
  NANDN U8028 ( .A(n4366), .B(creg[120]), .Z(n5694) );
  NANDN U8029 ( .A(n6157), .B(m[120]), .Z(n5693) );
  NAND U8030 ( .A(n5694), .B(n5693), .Z(y[120]) );
  NANDN U8031 ( .A(n4366), .B(creg[121]), .Z(n5696) );
  NANDN U8032 ( .A(n6157), .B(m[121]), .Z(n5695) );
  NAND U8033 ( .A(n5696), .B(n5695), .Z(y[121]) );
  NANDN U8034 ( .A(n4366), .B(creg[122]), .Z(n5698) );
  NANDN U8035 ( .A(n6157), .B(m[122]), .Z(n5697) );
  NAND U8036 ( .A(n5698), .B(n5697), .Z(y[122]) );
  NANDN U8037 ( .A(n4366), .B(creg[123]), .Z(n5700) );
  NANDN U8038 ( .A(n6157), .B(m[123]), .Z(n5699) );
  NAND U8039 ( .A(n5700), .B(n5699), .Z(y[123]) );
  NANDN U8040 ( .A(n4366), .B(creg[124]), .Z(n5702) );
  NANDN U8041 ( .A(n6157), .B(m[124]), .Z(n5701) );
  NAND U8042 ( .A(n5702), .B(n5701), .Z(y[124]) );
  NANDN U8043 ( .A(n4366), .B(creg[125]), .Z(n5704) );
  NANDN U8044 ( .A(n6157), .B(m[125]), .Z(n5703) );
  NAND U8045 ( .A(n5704), .B(n5703), .Z(y[125]) );
  NANDN U8046 ( .A(n4366), .B(creg[126]), .Z(n5706) );
  NANDN U8047 ( .A(n6157), .B(m[126]), .Z(n5705) );
  NAND U8048 ( .A(n5706), .B(n5705), .Z(y[126]) );
  NANDN U8049 ( .A(n4366), .B(creg[127]), .Z(n5708) );
  NANDN U8050 ( .A(n6157), .B(m[127]), .Z(n5707) );
  NAND U8051 ( .A(n5708), .B(n5707), .Z(y[127]) );
  NANDN U8052 ( .A(n4366), .B(creg[128]), .Z(n5710) );
  NANDN U8053 ( .A(n6157), .B(m[128]), .Z(n5709) );
  NAND U8054 ( .A(n5710), .B(n5709), .Z(y[128]) );
  NANDN U8055 ( .A(n4366), .B(creg[129]), .Z(n5712) );
  NANDN U8056 ( .A(n6157), .B(m[129]), .Z(n5711) );
  NAND U8057 ( .A(n5712), .B(n5711), .Z(y[129]) );
  NANDN U8058 ( .A(n4366), .B(creg[12]), .Z(n5714) );
  NANDN U8059 ( .A(n6157), .B(m[12]), .Z(n5713) );
  NAND U8060 ( .A(n5714), .B(n5713), .Z(y[12]) );
  NANDN U8061 ( .A(n4366), .B(creg[130]), .Z(n5716) );
  NANDN U8062 ( .A(n6157), .B(m[130]), .Z(n5715) );
  NAND U8063 ( .A(n5716), .B(n5715), .Z(y[130]) );
  NANDN U8064 ( .A(n4366), .B(creg[131]), .Z(n5718) );
  NANDN U8065 ( .A(n6157), .B(m[131]), .Z(n5717) );
  NAND U8066 ( .A(n5718), .B(n5717), .Z(y[131]) );
  NANDN U8067 ( .A(n4366), .B(creg[132]), .Z(n5720) );
  NANDN U8068 ( .A(n6157), .B(m[132]), .Z(n5719) );
  NAND U8069 ( .A(n5720), .B(n5719), .Z(y[132]) );
  NANDN U8070 ( .A(n4366), .B(creg[133]), .Z(n5722) );
  NANDN U8071 ( .A(n6157), .B(m[133]), .Z(n5721) );
  NAND U8072 ( .A(n5722), .B(n5721), .Z(y[133]) );
  NANDN U8073 ( .A(n4366), .B(creg[134]), .Z(n5724) );
  NANDN U8074 ( .A(n6157), .B(m[134]), .Z(n5723) );
  NAND U8075 ( .A(n5724), .B(n5723), .Z(y[134]) );
  NANDN U8076 ( .A(n4366), .B(creg[135]), .Z(n5726) );
  NANDN U8077 ( .A(n6157), .B(m[135]), .Z(n5725) );
  NAND U8078 ( .A(n5726), .B(n5725), .Z(y[135]) );
  NANDN U8079 ( .A(n4366), .B(creg[136]), .Z(n5728) );
  NANDN U8080 ( .A(n6157), .B(m[136]), .Z(n5727) );
  NAND U8081 ( .A(n5728), .B(n5727), .Z(y[136]) );
  NANDN U8082 ( .A(n4366), .B(creg[137]), .Z(n5730) );
  NANDN U8083 ( .A(n6157), .B(m[137]), .Z(n5729) );
  NAND U8084 ( .A(n5730), .B(n5729), .Z(y[137]) );
  NANDN U8085 ( .A(n4366), .B(creg[138]), .Z(n5732) );
  NANDN U8086 ( .A(n6157), .B(m[138]), .Z(n5731) );
  NAND U8087 ( .A(n5732), .B(n5731), .Z(y[138]) );
  NANDN U8088 ( .A(n4366), .B(creg[139]), .Z(n5734) );
  NANDN U8089 ( .A(n6157), .B(m[139]), .Z(n5733) );
  NAND U8090 ( .A(n5734), .B(n5733), .Z(y[139]) );
  NANDN U8091 ( .A(n4366), .B(creg[13]), .Z(n5736) );
  NANDN U8092 ( .A(n6157), .B(m[13]), .Z(n5735) );
  NAND U8093 ( .A(n5736), .B(n5735), .Z(y[13]) );
  NANDN U8094 ( .A(n4366), .B(creg[140]), .Z(n5738) );
  NANDN U8095 ( .A(n6157), .B(m[140]), .Z(n5737) );
  NAND U8096 ( .A(n5738), .B(n5737), .Z(y[140]) );
  NANDN U8097 ( .A(n4366), .B(creg[141]), .Z(n5740) );
  NANDN U8098 ( .A(n6157), .B(m[141]), .Z(n5739) );
  NAND U8099 ( .A(n5740), .B(n5739), .Z(y[141]) );
  NANDN U8100 ( .A(n4366), .B(creg[142]), .Z(n5742) );
  NANDN U8101 ( .A(n6157), .B(m[142]), .Z(n5741) );
  NAND U8102 ( .A(n5742), .B(n5741), .Z(y[142]) );
  NANDN U8103 ( .A(n4366), .B(creg[143]), .Z(n5744) );
  NANDN U8104 ( .A(n6157), .B(m[143]), .Z(n5743) );
  NAND U8105 ( .A(n5744), .B(n5743), .Z(y[143]) );
  NANDN U8106 ( .A(n4366), .B(creg[144]), .Z(n5746) );
  NANDN U8107 ( .A(n6157), .B(m[144]), .Z(n5745) );
  NAND U8108 ( .A(n5746), .B(n5745), .Z(y[144]) );
  NANDN U8109 ( .A(n4366), .B(creg[145]), .Z(n5748) );
  NANDN U8110 ( .A(n6157), .B(m[145]), .Z(n5747) );
  NAND U8111 ( .A(n5748), .B(n5747), .Z(y[145]) );
  NANDN U8112 ( .A(n4366), .B(creg[146]), .Z(n5750) );
  NANDN U8113 ( .A(n6157), .B(m[146]), .Z(n5749) );
  NAND U8114 ( .A(n5750), .B(n5749), .Z(y[146]) );
  NANDN U8115 ( .A(n4366), .B(creg[147]), .Z(n5752) );
  NANDN U8116 ( .A(n6157), .B(m[147]), .Z(n5751) );
  NAND U8117 ( .A(n5752), .B(n5751), .Z(y[147]) );
  NANDN U8118 ( .A(n4366), .B(creg[148]), .Z(n5754) );
  NANDN U8119 ( .A(n6157), .B(m[148]), .Z(n5753) );
  NAND U8120 ( .A(n5754), .B(n5753), .Z(y[148]) );
  NANDN U8121 ( .A(n4366), .B(creg[149]), .Z(n5756) );
  NANDN U8122 ( .A(n6157), .B(m[149]), .Z(n5755) );
  NAND U8123 ( .A(n5756), .B(n5755), .Z(y[149]) );
  NANDN U8124 ( .A(n4366), .B(creg[14]), .Z(n5758) );
  NANDN U8125 ( .A(n6157), .B(m[14]), .Z(n5757) );
  NAND U8126 ( .A(n5758), .B(n5757), .Z(y[14]) );
  NANDN U8127 ( .A(n4366), .B(creg[150]), .Z(n5760) );
  NANDN U8128 ( .A(n6157), .B(m[150]), .Z(n5759) );
  NAND U8129 ( .A(n5760), .B(n5759), .Z(y[150]) );
  NANDN U8130 ( .A(n4366), .B(creg[151]), .Z(n5762) );
  NANDN U8131 ( .A(n6157), .B(m[151]), .Z(n5761) );
  NAND U8132 ( .A(n5762), .B(n5761), .Z(y[151]) );
  NANDN U8133 ( .A(n4366), .B(creg[152]), .Z(n5764) );
  NANDN U8134 ( .A(n6157), .B(m[152]), .Z(n5763) );
  NAND U8135 ( .A(n5764), .B(n5763), .Z(y[152]) );
  NANDN U8136 ( .A(n4366), .B(creg[153]), .Z(n5766) );
  NANDN U8137 ( .A(n6157), .B(m[153]), .Z(n5765) );
  NAND U8138 ( .A(n5766), .B(n5765), .Z(y[153]) );
  NANDN U8139 ( .A(n4366), .B(creg[154]), .Z(n5768) );
  NANDN U8140 ( .A(n6157), .B(m[154]), .Z(n5767) );
  NAND U8141 ( .A(n5768), .B(n5767), .Z(y[154]) );
  NANDN U8142 ( .A(n4366), .B(creg[155]), .Z(n5770) );
  NANDN U8143 ( .A(n6157), .B(m[155]), .Z(n5769) );
  NAND U8144 ( .A(n5770), .B(n5769), .Z(y[155]) );
  NANDN U8145 ( .A(n4366), .B(creg[156]), .Z(n5772) );
  NANDN U8146 ( .A(n6157), .B(m[156]), .Z(n5771) );
  NAND U8147 ( .A(n5772), .B(n5771), .Z(y[156]) );
  NANDN U8148 ( .A(n4366), .B(creg[157]), .Z(n5774) );
  NANDN U8149 ( .A(n6157), .B(m[157]), .Z(n5773) );
  NAND U8150 ( .A(n5774), .B(n5773), .Z(y[157]) );
  NANDN U8151 ( .A(n4366), .B(creg[158]), .Z(n5776) );
  NANDN U8152 ( .A(n6157), .B(m[158]), .Z(n5775) );
  NAND U8153 ( .A(n5776), .B(n5775), .Z(y[158]) );
  NANDN U8154 ( .A(n4366), .B(creg[159]), .Z(n5778) );
  NANDN U8155 ( .A(n6157), .B(m[159]), .Z(n5777) );
  NAND U8156 ( .A(n5778), .B(n5777), .Z(y[159]) );
  NANDN U8157 ( .A(n4366), .B(creg[15]), .Z(n5780) );
  NANDN U8158 ( .A(n6157), .B(m[15]), .Z(n5779) );
  NAND U8159 ( .A(n5780), .B(n5779), .Z(y[15]) );
  NANDN U8160 ( .A(n4366), .B(creg[160]), .Z(n5782) );
  NANDN U8161 ( .A(n6157), .B(m[160]), .Z(n5781) );
  NAND U8162 ( .A(n5782), .B(n5781), .Z(y[160]) );
  NANDN U8163 ( .A(n4366), .B(creg[161]), .Z(n5784) );
  NANDN U8164 ( .A(n6157), .B(m[161]), .Z(n5783) );
  NAND U8165 ( .A(n5784), .B(n5783), .Z(y[161]) );
  NANDN U8166 ( .A(n4366), .B(creg[162]), .Z(n5786) );
  NANDN U8167 ( .A(n6157), .B(m[162]), .Z(n5785) );
  NAND U8168 ( .A(n5786), .B(n5785), .Z(y[162]) );
  NANDN U8169 ( .A(n4366), .B(creg[163]), .Z(n5788) );
  NANDN U8170 ( .A(n6157), .B(m[163]), .Z(n5787) );
  NAND U8171 ( .A(n5788), .B(n5787), .Z(y[163]) );
  NANDN U8172 ( .A(n4366), .B(creg[164]), .Z(n5790) );
  NANDN U8173 ( .A(n6157), .B(m[164]), .Z(n5789) );
  NAND U8174 ( .A(n5790), .B(n5789), .Z(y[164]) );
  NANDN U8175 ( .A(n4366), .B(creg[165]), .Z(n5792) );
  NANDN U8176 ( .A(n6157), .B(m[165]), .Z(n5791) );
  NAND U8177 ( .A(n5792), .B(n5791), .Z(y[165]) );
  NANDN U8178 ( .A(n4366), .B(creg[166]), .Z(n5794) );
  NANDN U8179 ( .A(n6157), .B(m[166]), .Z(n5793) );
  NAND U8180 ( .A(n5794), .B(n5793), .Z(y[166]) );
  NANDN U8181 ( .A(n4366), .B(creg[167]), .Z(n5796) );
  NANDN U8182 ( .A(n6157), .B(m[167]), .Z(n5795) );
  NAND U8183 ( .A(n5796), .B(n5795), .Z(y[167]) );
  NANDN U8184 ( .A(n4366), .B(creg[168]), .Z(n5798) );
  NANDN U8185 ( .A(n6157), .B(m[168]), .Z(n5797) );
  NAND U8186 ( .A(n5798), .B(n5797), .Z(y[168]) );
  NANDN U8187 ( .A(n4366), .B(creg[169]), .Z(n5800) );
  NANDN U8188 ( .A(n6157), .B(m[169]), .Z(n5799) );
  NAND U8189 ( .A(n5800), .B(n5799), .Z(y[169]) );
  NANDN U8190 ( .A(n4366), .B(creg[16]), .Z(n5802) );
  NANDN U8191 ( .A(n6157), .B(m[16]), .Z(n5801) );
  NAND U8192 ( .A(n5802), .B(n5801), .Z(y[16]) );
  NANDN U8193 ( .A(n4366), .B(creg[170]), .Z(n5804) );
  NANDN U8194 ( .A(n6157), .B(m[170]), .Z(n5803) );
  NAND U8195 ( .A(n5804), .B(n5803), .Z(y[170]) );
  NANDN U8196 ( .A(n4366), .B(creg[171]), .Z(n5806) );
  NANDN U8197 ( .A(n6157), .B(m[171]), .Z(n5805) );
  NAND U8198 ( .A(n5806), .B(n5805), .Z(y[171]) );
  NANDN U8199 ( .A(n4366), .B(creg[172]), .Z(n5808) );
  NANDN U8200 ( .A(n6157), .B(m[172]), .Z(n5807) );
  NAND U8201 ( .A(n5808), .B(n5807), .Z(y[172]) );
  NANDN U8202 ( .A(n4366), .B(creg[173]), .Z(n5810) );
  NANDN U8203 ( .A(n6157), .B(m[173]), .Z(n5809) );
  NAND U8204 ( .A(n5810), .B(n5809), .Z(y[173]) );
  NANDN U8205 ( .A(n4366), .B(creg[174]), .Z(n5812) );
  NANDN U8206 ( .A(n6157), .B(m[174]), .Z(n5811) );
  NAND U8207 ( .A(n5812), .B(n5811), .Z(y[174]) );
  NANDN U8208 ( .A(n4366), .B(creg[175]), .Z(n5814) );
  NANDN U8209 ( .A(n6157), .B(m[175]), .Z(n5813) );
  NAND U8210 ( .A(n5814), .B(n5813), .Z(y[175]) );
  NANDN U8211 ( .A(n4366), .B(creg[176]), .Z(n5816) );
  NANDN U8212 ( .A(n6157), .B(m[176]), .Z(n5815) );
  NAND U8213 ( .A(n5816), .B(n5815), .Z(y[176]) );
  NANDN U8214 ( .A(n4366), .B(creg[177]), .Z(n5818) );
  NANDN U8215 ( .A(n6157), .B(m[177]), .Z(n5817) );
  NAND U8216 ( .A(n5818), .B(n5817), .Z(y[177]) );
  NANDN U8217 ( .A(n4366), .B(creg[178]), .Z(n5820) );
  NANDN U8218 ( .A(n6157), .B(m[178]), .Z(n5819) );
  NAND U8219 ( .A(n5820), .B(n5819), .Z(y[178]) );
  NANDN U8220 ( .A(n4366), .B(creg[179]), .Z(n5822) );
  NANDN U8221 ( .A(n6157), .B(m[179]), .Z(n5821) );
  NAND U8222 ( .A(n5822), .B(n5821), .Z(y[179]) );
  NANDN U8223 ( .A(n4366), .B(creg[17]), .Z(n5824) );
  NANDN U8224 ( .A(n6157), .B(m[17]), .Z(n5823) );
  NAND U8225 ( .A(n5824), .B(n5823), .Z(y[17]) );
  NANDN U8226 ( .A(n4366), .B(creg[180]), .Z(n5826) );
  NANDN U8227 ( .A(n6157), .B(m[180]), .Z(n5825) );
  NAND U8228 ( .A(n5826), .B(n5825), .Z(y[180]) );
  NANDN U8229 ( .A(n4366), .B(creg[181]), .Z(n5828) );
  NANDN U8230 ( .A(n6157), .B(m[181]), .Z(n5827) );
  NAND U8231 ( .A(n5828), .B(n5827), .Z(y[181]) );
  NANDN U8232 ( .A(n4366), .B(creg[182]), .Z(n5830) );
  NANDN U8233 ( .A(n6157), .B(m[182]), .Z(n5829) );
  NAND U8234 ( .A(n5830), .B(n5829), .Z(y[182]) );
  NANDN U8235 ( .A(n4366), .B(creg[183]), .Z(n5832) );
  NANDN U8236 ( .A(n6157), .B(m[183]), .Z(n5831) );
  NAND U8237 ( .A(n5832), .B(n5831), .Z(y[183]) );
  NANDN U8238 ( .A(n4366), .B(creg[184]), .Z(n5834) );
  NANDN U8239 ( .A(n6157), .B(m[184]), .Z(n5833) );
  NAND U8240 ( .A(n5834), .B(n5833), .Z(y[184]) );
  NANDN U8241 ( .A(n4366), .B(creg[185]), .Z(n5836) );
  NANDN U8242 ( .A(n6157), .B(m[185]), .Z(n5835) );
  NAND U8243 ( .A(n5836), .B(n5835), .Z(y[185]) );
  NANDN U8244 ( .A(n4366), .B(creg[186]), .Z(n5838) );
  NANDN U8245 ( .A(n6157), .B(m[186]), .Z(n5837) );
  NAND U8246 ( .A(n5838), .B(n5837), .Z(y[186]) );
  NANDN U8247 ( .A(n4366), .B(creg[187]), .Z(n5840) );
  NANDN U8248 ( .A(n6157), .B(m[187]), .Z(n5839) );
  NAND U8249 ( .A(n5840), .B(n5839), .Z(y[187]) );
  NANDN U8250 ( .A(n4366), .B(creg[188]), .Z(n5842) );
  NANDN U8251 ( .A(n6157), .B(m[188]), .Z(n5841) );
  NAND U8252 ( .A(n5842), .B(n5841), .Z(y[188]) );
  NANDN U8253 ( .A(n4366), .B(creg[189]), .Z(n5844) );
  NANDN U8254 ( .A(n6157), .B(m[189]), .Z(n5843) );
  NAND U8255 ( .A(n5844), .B(n5843), .Z(y[189]) );
  NANDN U8256 ( .A(n4366), .B(creg[18]), .Z(n5846) );
  NANDN U8257 ( .A(n6157), .B(m[18]), .Z(n5845) );
  NAND U8258 ( .A(n5846), .B(n5845), .Z(y[18]) );
  NANDN U8259 ( .A(n4366), .B(creg[190]), .Z(n5848) );
  NANDN U8260 ( .A(n6157), .B(m[190]), .Z(n5847) );
  NAND U8261 ( .A(n5848), .B(n5847), .Z(y[190]) );
  NANDN U8262 ( .A(n4366), .B(creg[191]), .Z(n5850) );
  NANDN U8263 ( .A(n6157), .B(m[191]), .Z(n5849) );
  NAND U8264 ( .A(n5850), .B(n5849), .Z(y[191]) );
  NANDN U8265 ( .A(n4366), .B(creg[192]), .Z(n5852) );
  NANDN U8266 ( .A(n6157), .B(m[192]), .Z(n5851) );
  NAND U8267 ( .A(n5852), .B(n5851), .Z(y[192]) );
  NANDN U8268 ( .A(n4366), .B(creg[193]), .Z(n5854) );
  NANDN U8269 ( .A(n6157), .B(m[193]), .Z(n5853) );
  NAND U8270 ( .A(n5854), .B(n5853), .Z(y[193]) );
  NANDN U8271 ( .A(n4366), .B(creg[194]), .Z(n5856) );
  NANDN U8272 ( .A(n6157), .B(m[194]), .Z(n5855) );
  NAND U8273 ( .A(n5856), .B(n5855), .Z(y[194]) );
  NANDN U8274 ( .A(n4366), .B(creg[195]), .Z(n5858) );
  NANDN U8275 ( .A(n6157), .B(m[195]), .Z(n5857) );
  NAND U8276 ( .A(n5858), .B(n5857), .Z(y[195]) );
  NANDN U8277 ( .A(n4366), .B(creg[196]), .Z(n5860) );
  NANDN U8278 ( .A(n6157), .B(m[196]), .Z(n5859) );
  NAND U8279 ( .A(n5860), .B(n5859), .Z(y[196]) );
  NANDN U8280 ( .A(n4366), .B(creg[197]), .Z(n5862) );
  NANDN U8281 ( .A(n6157), .B(m[197]), .Z(n5861) );
  NAND U8282 ( .A(n5862), .B(n5861), .Z(y[197]) );
  NANDN U8283 ( .A(n4366), .B(creg[198]), .Z(n5864) );
  NANDN U8284 ( .A(n6157), .B(m[198]), .Z(n5863) );
  NAND U8285 ( .A(n5864), .B(n5863), .Z(y[198]) );
  NANDN U8286 ( .A(n4366), .B(creg[199]), .Z(n5866) );
  NANDN U8287 ( .A(n6157), .B(m[199]), .Z(n5865) );
  NAND U8288 ( .A(n5866), .B(n5865), .Z(y[199]) );
  NANDN U8289 ( .A(n4366), .B(creg[19]), .Z(n5868) );
  NANDN U8290 ( .A(n6157), .B(m[19]), .Z(n5867) );
  NAND U8291 ( .A(n5868), .B(n5867), .Z(y[19]) );
  NANDN U8292 ( .A(n4366), .B(creg[1]), .Z(n5870) );
  NANDN U8293 ( .A(n6157), .B(m[1]), .Z(n5869) );
  NAND U8294 ( .A(n5870), .B(n5869), .Z(y[1]) );
  NANDN U8295 ( .A(n4366), .B(creg[200]), .Z(n5872) );
  NANDN U8296 ( .A(n6157), .B(m[200]), .Z(n5871) );
  NAND U8297 ( .A(n5872), .B(n5871), .Z(y[200]) );
  NANDN U8298 ( .A(n4366), .B(creg[201]), .Z(n5874) );
  NANDN U8299 ( .A(n6157), .B(m[201]), .Z(n5873) );
  NAND U8300 ( .A(n5874), .B(n5873), .Z(y[201]) );
  NANDN U8301 ( .A(n4366), .B(creg[202]), .Z(n5876) );
  NANDN U8302 ( .A(n6157), .B(m[202]), .Z(n5875) );
  NAND U8303 ( .A(n5876), .B(n5875), .Z(y[202]) );
  NANDN U8304 ( .A(n4366), .B(creg[203]), .Z(n5878) );
  NANDN U8305 ( .A(n6157), .B(m[203]), .Z(n5877) );
  NAND U8306 ( .A(n5878), .B(n5877), .Z(y[203]) );
  NANDN U8307 ( .A(n4366), .B(creg[204]), .Z(n5880) );
  NANDN U8308 ( .A(n6157), .B(m[204]), .Z(n5879) );
  NAND U8309 ( .A(n5880), .B(n5879), .Z(y[204]) );
  NANDN U8310 ( .A(n4366), .B(creg[205]), .Z(n5882) );
  NANDN U8311 ( .A(n6157), .B(m[205]), .Z(n5881) );
  NAND U8312 ( .A(n5882), .B(n5881), .Z(y[205]) );
  NANDN U8313 ( .A(n4366), .B(creg[206]), .Z(n5884) );
  NANDN U8314 ( .A(n6157), .B(m[206]), .Z(n5883) );
  NAND U8315 ( .A(n5884), .B(n5883), .Z(y[206]) );
  NANDN U8316 ( .A(n4366), .B(creg[207]), .Z(n5886) );
  NANDN U8317 ( .A(n6157), .B(m[207]), .Z(n5885) );
  NAND U8318 ( .A(n5886), .B(n5885), .Z(y[207]) );
  NANDN U8319 ( .A(n4366), .B(creg[208]), .Z(n5888) );
  NANDN U8320 ( .A(n6157), .B(m[208]), .Z(n5887) );
  NAND U8321 ( .A(n5888), .B(n5887), .Z(y[208]) );
  NANDN U8322 ( .A(n4366), .B(creg[209]), .Z(n5890) );
  NANDN U8323 ( .A(n6157), .B(m[209]), .Z(n5889) );
  NAND U8324 ( .A(n5890), .B(n5889), .Z(y[209]) );
  NANDN U8325 ( .A(n4366), .B(creg[20]), .Z(n5892) );
  NANDN U8326 ( .A(n6157), .B(m[20]), .Z(n5891) );
  NAND U8327 ( .A(n5892), .B(n5891), .Z(y[20]) );
  NANDN U8328 ( .A(n4366), .B(creg[210]), .Z(n5894) );
  NANDN U8329 ( .A(n6157), .B(m[210]), .Z(n5893) );
  NAND U8330 ( .A(n5894), .B(n5893), .Z(y[210]) );
  NANDN U8331 ( .A(n4366), .B(creg[211]), .Z(n5896) );
  NANDN U8332 ( .A(n6157), .B(m[211]), .Z(n5895) );
  NAND U8333 ( .A(n5896), .B(n5895), .Z(y[211]) );
  NANDN U8334 ( .A(n4366), .B(creg[212]), .Z(n5898) );
  NANDN U8335 ( .A(n6157), .B(m[212]), .Z(n5897) );
  NAND U8336 ( .A(n5898), .B(n5897), .Z(y[212]) );
  NANDN U8337 ( .A(n4366), .B(creg[213]), .Z(n5900) );
  NANDN U8338 ( .A(n6157), .B(m[213]), .Z(n5899) );
  NAND U8339 ( .A(n5900), .B(n5899), .Z(y[213]) );
  NANDN U8340 ( .A(n4366), .B(creg[214]), .Z(n5902) );
  NANDN U8341 ( .A(n6157), .B(m[214]), .Z(n5901) );
  NAND U8342 ( .A(n5902), .B(n5901), .Z(y[214]) );
  NANDN U8343 ( .A(n4366), .B(creg[215]), .Z(n5904) );
  NANDN U8344 ( .A(n6157), .B(m[215]), .Z(n5903) );
  NAND U8345 ( .A(n5904), .B(n5903), .Z(y[215]) );
  NANDN U8346 ( .A(n4366), .B(creg[216]), .Z(n5906) );
  NANDN U8347 ( .A(n6157), .B(m[216]), .Z(n5905) );
  NAND U8348 ( .A(n5906), .B(n5905), .Z(y[216]) );
  NANDN U8349 ( .A(n4366), .B(creg[217]), .Z(n5908) );
  NANDN U8350 ( .A(n6157), .B(m[217]), .Z(n5907) );
  NAND U8351 ( .A(n5908), .B(n5907), .Z(y[217]) );
  NANDN U8352 ( .A(n4366), .B(creg[218]), .Z(n5910) );
  NANDN U8353 ( .A(n6157), .B(m[218]), .Z(n5909) );
  NAND U8354 ( .A(n5910), .B(n5909), .Z(y[218]) );
  NANDN U8355 ( .A(n4366), .B(creg[219]), .Z(n5912) );
  NANDN U8356 ( .A(n6157), .B(m[219]), .Z(n5911) );
  NAND U8357 ( .A(n5912), .B(n5911), .Z(y[219]) );
  NANDN U8358 ( .A(n4366), .B(creg[21]), .Z(n5914) );
  NANDN U8359 ( .A(n6157), .B(m[21]), .Z(n5913) );
  NAND U8360 ( .A(n5914), .B(n5913), .Z(y[21]) );
  NANDN U8361 ( .A(n4366), .B(creg[220]), .Z(n5916) );
  NANDN U8362 ( .A(n6157), .B(m[220]), .Z(n5915) );
  NAND U8363 ( .A(n5916), .B(n5915), .Z(y[220]) );
  NANDN U8364 ( .A(n4366), .B(creg[221]), .Z(n5918) );
  NANDN U8365 ( .A(n6157), .B(m[221]), .Z(n5917) );
  NAND U8366 ( .A(n5918), .B(n5917), .Z(y[221]) );
  NANDN U8367 ( .A(n4366), .B(creg[222]), .Z(n5920) );
  NANDN U8368 ( .A(n6157), .B(m[222]), .Z(n5919) );
  NAND U8369 ( .A(n5920), .B(n5919), .Z(y[222]) );
  NANDN U8370 ( .A(n4366), .B(creg[223]), .Z(n5922) );
  NANDN U8371 ( .A(n6157), .B(m[223]), .Z(n5921) );
  NAND U8372 ( .A(n5922), .B(n5921), .Z(y[223]) );
  NANDN U8373 ( .A(n4366), .B(creg[224]), .Z(n5924) );
  NANDN U8374 ( .A(n6157), .B(m[224]), .Z(n5923) );
  NAND U8375 ( .A(n5924), .B(n5923), .Z(y[224]) );
  NANDN U8376 ( .A(n4366), .B(creg[225]), .Z(n5926) );
  NANDN U8377 ( .A(n6157), .B(m[225]), .Z(n5925) );
  NAND U8378 ( .A(n5926), .B(n5925), .Z(y[225]) );
  NANDN U8379 ( .A(n4366), .B(creg[226]), .Z(n5928) );
  NANDN U8380 ( .A(n6157), .B(m[226]), .Z(n5927) );
  NAND U8381 ( .A(n5928), .B(n5927), .Z(y[226]) );
  NANDN U8382 ( .A(n4366), .B(creg[227]), .Z(n5930) );
  NANDN U8383 ( .A(n6157), .B(m[227]), .Z(n5929) );
  NAND U8384 ( .A(n5930), .B(n5929), .Z(y[227]) );
  NANDN U8385 ( .A(n4366), .B(creg[228]), .Z(n5932) );
  NANDN U8386 ( .A(n6157), .B(m[228]), .Z(n5931) );
  NAND U8387 ( .A(n5932), .B(n5931), .Z(y[228]) );
  NANDN U8388 ( .A(n4366), .B(creg[229]), .Z(n5934) );
  NANDN U8389 ( .A(n6157), .B(m[229]), .Z(n5933) );
  NAND U8390 ( .A(n5934), .B(n5933), .Z(y[229]) );
  NANDN U8391 ( .A(n4366), .B(creg[22]), .Z(n5936) );
  NANDN U8392 ( .A(n6157), .B(m[22]), .Z(n5935) );
  NAND U8393 ( .A(n5936), .B(n5935), .Z(y[22]) );
  NANDN U8394 ( .A(n4366), .B(creg[230]), .Z(n5938) );
  NANDN U8395 ( .A(n6157), .B(m[230]), .Z(n5937) );
  NAND U8396 ( .A(n5938), .B(n5937), .Z(y[230]) );
  NANDN U8397 ( .A(n4366), .B(creg[231]), .Z(n5940) );
  NANDN U8398 ( .A(n6157), .B(m[231]), .Z(n5939) );
  NAND U8399 ( .A(n5940), .B(n5939), .Z(y[231]) );
  NANDN U8400 ( .A(n4366), .B(creg[232]), .Z(n5942) );
  NANDN U8401 ( .A(n6157), .B(m[232]), .Z(n5941) );
  NAND U8402 ( .A(n5942), .B(n5941), .Z(y[232]) );
  NANDN U8403 ( .A(n4366), .B(creg[233]), .Z(n5944) );
  NANDN U8404 ( .A(n6157), .B(m[233]), .Z(n5943) );
  NAND U8405 ( .A(n5944), .B(n5943), .Z(y[233]) );
  NANDN U8406 ( .A(n4366), .B(creg[234]), .Z(n5946) );
  NANDN U8407 ( .A(n6157), .B(m[234]), .Z(n5945) );
  NAND U8408 ( .A(n5946), .B(n5945), .Z(y[234]) );
  NANDN U8409 ( .A(n4366), .B(creg[235]), .Z(n5948) );
  NANDN U8410 ( .A(n6157), .B(m[235]), .Z(n5947) );
  NAND U8411 ( .A(n5948), .B(n5947), .Z(y[235]) );
  NANDN U8412 ( .A(n4366), .B(creg[236]), .Z(n5950) );
  NANDN U8413 ( .A(n6157), .B(m[236]), .Z(n5949) );
  NAND U8414 ( .A(n5950), .B(n5949), .Z(y[236]) );
  NANDN U8415 ( .A(n4366), .B(creg[237]), .Z(n5952) );
  NANDN U8416 ( .A(n6157), .B(m[237]), .Z(n5951) );
  NAND U8417 ( .A(n5952), .B(n5951), .Z(y[237]) );
  NANDN U8418 ( .A(n4366), .B(creg[238]), .Z(n5954) );
  NANDN U8419 ( .A(n6157), .B(m[238]), .Z(n5953) );
  NAND U8420 ( .A(n5954), .B(n5953), .Z(y[238]) );
  NANDN U8421 ( .A(n4366), .B(creg[239]), .Z(n5956) );
  NANDN U8422 ( .A(n6157), .B(m[239]), .Z(n5955) );
  NAND U8423 ( .A(n5956), .B(n5955), .Z(y[239]) );
  NANDN U8424 ( .A(n4366), .B(creg[23]), .Z(n5958) );
  NANDN U8425 ( .A(n6157), .B(m[23]), .Z(n5957) );
  NAND U8426 ( .A(n5958), .B(n5957), .Z(y[23]) );
  NANDN U8427 ( .A(n4366), .B(creg[240]), .Z(n5960) );
  NANDN U8428 ( .A(n6157), .B(m[240]), .Z(n5959) );
  NAND U8429 ( .A(n5960), .B(n5959), .Z(y[240]) );
  NANDN U8430 ( .A(n4366), .B(creg[241]), .Z(n5962) );
  NANDN U8431 ( .A(n6157), .B(m[241]), .Z(n5961) );
  NAND U8432 ( .A(n5962), .B(n5961), .Z(y[241]) );
  NANDN U8433 ( .A(n4366), .B(creg[242]), .Z(n5964) );
  NANDN U8434 ( .A(n6157), .B(m[242]), .Z(n5963) );
  NAND U8435 ( .A(n5964), .B(n5963), .Z(y[242]) );
  NANDN U8436 ( .A(n4366), .B(creg[243]), .Z(n5966) );
  NANDN U8437 ( .A(n6157), .B(m[243]), .Z(n5965) );
  NAND U8438 ( .A(n5966), .B(n5965), .Z(y[243]) );
  NANDN U8439 ( .A(n4366), .B(creg[244]), .Z(n5968) );
  NANDN U8440 ( .A(n6157), .B(m[244]), .Z(n5967) );
  NAND U8441 ( .A(n5968), .B(n5967), .Z(y[244]) );
  NANDN U8442 ( .A(n4366), .B(creg[245]), .Z(n5970) );
  NANDN U8443 ( .A(n6157), .B(m[245]), .Z(n5969) );
  NAND U8444 ( .A(n5970), .B(n5969), .Z(y[245]) );
  NANDN U8445 ( .A(n4366), .B(creg[246]), .Z(n5972) );
  NANDN U8446 ( .A(n6157), .B(m[246]), .Z(n5971) );
  NAND U8447 ( .A(n5972), .B(n5971), .Z(y[246]) );
  NANDN U8448 ( .A(n4366), .B(creg[247]), .Z(n5974) );
  NANDN U8449 ( .A(n6157), .B(m[247]), .Z(n5973) );
  NAND U8450 ( .A(n5974), .B(n5973), .Z(y[247]) );
  NANDN U8451 ( .A(n4366), .B(creg[248]), .Z(n5976) );
  NANDN U8452 ( .A(n6157), .B(m[248]), .Z(n5975) );
  NAND U8453 ( .A(n5976), .B(n5975), .Z(y[248]) );
  NANDN U8454 ( .A(n4366), .B(creg[249]), .Z(n5978) );
  NANDN U8455 ( .A(n6157), .B(m[249]), .Z(n5977) );
  NAND U8456 ( .A(n5978), .B(n5977), .Z(y[249]) );
  NANDN U8457 ( .A(n4366), .B(creg[24]), .Z(n5980) );
  NANDN U8458 ( .A(n6157), .B(m[24]), .Z(n5979) );
  NAND U8459 ( .A(n5980), .B(n5979), .Z(y[24]) );
  NANDN U8460 ( .A(n4366), .B(creg[250]), .Z(n5982) );
  NANDN U8461 ( .A(n6157), .B(m[250]), .Z(n5981) );
  NAND U8462 ( .A(n5982), .B(n5981), .Z(y[250]) );
  NANDN U8463 ( .A(n4366), .B(creg[251]), .Z(n5984) );
  NANDN U8464 ( .A(n6157), .B(m[251]), .Z(n5983) );
  NAND U8465 ( .A(n5984), .B(n5983), .Z(y[251]) );
  NANDN U8466 ( .A(n4366), .B(creg[252]), .Z(n5986) );
  NANDN U8467 ( .A(n6157), .B(m[252]), .Z(n5985) );
  NAND U8468 ( .A(n5986), .B(n5985), .Z(y[252]) );
  NANDN U8469 ( .A(n4366), .B(creg[253]), .Z(n5988) );
  NANDN U8470 ( .A(n6157), .B(m[253]), .Z(n5987) );
  NAND U8471 ( .A(n5988), .B(n5987), .Z(y[253]) );
  NANDN U8472 ( .A(n4366), .B(creg[254]), .Z(n5990) );
  NANDN U8473 ( .A(n6157), .B(m[254]), .Z(n5989) );
  NAND U8474 ( .A(n5990), .B(n5989), .Z(y[254]) );
  NANDN U8475 ( .A(n4366), .B(creg[255]), .Z(n5992) );
  NANDN U8476 ( .A(n6157), .B(m[255]), .Z(n5991) );
  NAND U8477 ( .A(n5992), .B(n5991), .Z(y[255]) );
  NANDN U8478 ( .A(n4366), .B(creg[25]), .Z(n5994) );
  NANDN U8479 ( .A(n6157), .B(m[25]), .Z(n5993) );
  NAND U8480 ( .A(n5994), .B(n5993), .Z(y[25]) );
  NANDN U8481 ( .A(n4366), .B(creg[26]), .Z(n5996) );
  NANDN U8482 ( .A(n6157), .B(m[26]), .Z(n5995) );
  NAND U8483 ( .A(n5996), .B(n5995), .Z(y[26]) );
  NANDN U8484 ( .A(n4366), .B(creg[27]), .Z(n5998) );
  NANDN U8485 ( .A(n6157), .B(m[27]), .Z(n5997) );
  NAND U8486 ( .A(n5998), .B(n5997), .Z(y[27]) );
  NANDN U8487 ( .A(n4366), .B(creg[28]), .Z(n6000) );
  NANDN U8488 ( .A(n6157), .B(m[28]), .Z(n5999) );
  NAND U8489 ( .A(n6000), .B(n5999), .Z(y[28]) );
  NANDN U8490 ( .A(n4366), .B(creg[29]), .Z(n6002) );
  NANDN U8491 ( .A(n6157), .B(m[29]), .Z(n6001) );
  NAND U8492 ( .A(n6002), .B(n6001), .Z(y[29]) );
  NANDN U8493 ( .A(n4366), .B(creg[2]), .Z(n6004) );
  NANDN U8494 ( .A(n6157), .B(m[2]), .Z(n6003) );
  NAND U8495 ( .A(n6004), .B(n6003), .Z(y[2]) );
  NANDN U8496 ( .A(n4366), .B(creg[30]), .Z(n6006) );
  NANDN U8497 ( .A(n6157), .B(m[30]), .Z(n6005) );
  NAND U8498 ( .A(n6006), .B(n6005), .Z(y[30]) );
  NANDN U8499 ( .A(n4366), .B(creg[31]), .Z(n6008) );
  NANDN U8500 ( .A(n6157), .B(m[31]), .Z(n6007) );
  NAND U8501 ( .A(n6008), .B(n6007), .Z(y[31]) );
  NANDN U8502 ( .A(n4366), .B(creg[32]), .Z(n6010) );
  NANDN U8503 ( .A(n6157), .B(m[32]), .Z(n6009) );
  NAND U8504 ( .A(n6010), .B(n6009), .Z(y[32]) );
  NANDN U8505 ( .A(n4366), .B(creg[33]), .Z(n6012) );
  NANDN U8506 ( .A(n6157), .B(m[33]), .Z(n6011) );
  NAND U8507 ( .A(n6012), .B(n6011), .Z(y[33]) );
  NANDN U8508 ( .A(n4366), .B(creg[34]), .Z(n6014) );
  NANDN U8509 ( .A(n6157), .B(m[34]), .Z(n6013) );
  NAND U8510 ( .A(n6014), .B(n6013), .Z(y[34]) );
  NANDN U8511 ( .A(n4366), .B(creg[35]), .Z(n6016) );
  NANDN U8512 ( .A(n6157), .B(m[35]), .Z(n6015) );
  NAND U8513 ( .A(n6016), .B(n6015), .Z(y[35]) );
  NANDN U8514 ( .A(n4366), .B(creg[36]), .Z(n6018) );
  NANDN U8515 ( .A(n6157), .B(m[36]), .Z(n6017) );
  NAND U8516 ( .A(n6018), .B(n6017), .Z(y[36]) );
  NANDN U8517 ( .A(n4366), .B(creg[37]), .Z(n6020) );
  NANDN U8518 ( .A(n6157), .B(m[37]), .Z(n6019) );
  NAND U8519 ( .A(n6020), .B(n6019), .Z(y[37]) );
  NANDN U8520 ( .A(n4366), .B(creg[38]), .Z(n6022) );
  NANDN U8521 ( .A(n6157), .B(m[38]), .Z(n6021) );
  NAND U8522 ( .A(n6022), .B(n6021), .Z(y[38]) );
  NANDN U8523 ( .A(n4366), .B(creg[39]), .Z(n6024) );
  NANDN U8524 ( .A(n6157), .B(m[39]), .Z(n6023) );
  NAND U8525 ( .A(n6024), .B(n6023), .Z(y[39]) );
  NANDN U8526 ( .A(n4366), .B(creg[3]), .Z(n6026) );
  NANDN U8527 ( .A(n6157), .B(m[3]), .Z(n6025) );
  NAND U8528 ( .A(n6026), .B(n6025), .Z(y[3]) );
  NANDN U8529 ( .A(n4366), .B(creg[40]), .Z(n6028) );
  NANDN U8530 ( .A(n6157), .B(m[40]), .Z(n6027) );
  NAND U8531 ( .A(n6028), .B(n6027), .Z(y[40]) );
  NANDN U8532 ( .A(n4366), .B(creg[41]), .Z(n6030) );
  NANDN U8533 ( .A(n6157), .B(m[41]), .Z(n6029) );
  NAND U8534 ( .A(n6030), .B(n6029), .Z(y[41]) );
  NANDN U8535 ( .A(n4366), .B(creg[42]), .Z(n6032) );
  NANDN U8536 ( .A(n6157), .B(m[42]), .Z(n6031) );
  NAND U8537 ( .A(n6032), .B(n6031), .Z(y[42]) );
  NANDN U8538 ( .A(n4366), .B(creg[43]), .Z(n6034) );
  NANDN U8539 ( .A(n6157), .B(m[43]), .Z(n6033) );
  NAND U8540 ( .A(n6034), .B(n6033), .Z(y[43]) );
  NANDN U8541 ( .A(n4366), .B(creg[44]), .Z(n6036) );
  NANDN U8542 ( .A(n6157), .B(m[44]), .Z(n6035) );
  NAND U8543 ( .A(n6036), .B(n6035), .Z(y[44]) );
  NANDN U8544 ( .A(n4366), .B(creg[45]), .Z(n6038) );
  NANDN U8545 ( .A(n6157), .B(m[45]), .Z(n6037) );
  NAND U8546 ( .A(n6038), .B(n6037), .Z(y[45]) );
  NANDN U8547 ( .A(n4366), .B(creg[46]), .Z(n6040) );
  NANDN U8548 ( .A(n6157), .B(m[46]), .Z(n6039) );
  NAND U8549 ( .A(n6040), .B(n6039), .Z(y[46]) );
  NANDN U8550 ( .A(n4366), .B(creg[47]), .Z(n6042) );
  NANDN U8551 ( .A(n6157), .B(m[47]), .Z(n6041) );
  NAND U8552 ( .A(n6042), .B(n6041), .Z(y[47]) );
  NANDN U8553 ( .A(n4366), .B(creg[48]), .Z(n6044) );
  NANDN U8554 ( .A(n6157), .B(m[48]), .Z(n6043) );
  NAND U8555 ( .A(n6044), .B(n6043), .Z(y[48]) );
  NANDN U8556 ( .A(n4366), .B(creg[49]), .Z(n6046) );
  NANDN U8557 ( .A(n6157), .B(m[49]), .Z(n6045) );
  NAND U8558 ( .A(n6046), .B(n6045), .Z(y[49]) );
  NANDN U8559 ( .A(n4366), .B(creg[4]), .Z(n6048) );
  NANDN U8560 ( .A(n6157), .B(m[4]), .Z(n6047) );
  NAND U8561 ( .A(n6048), .B(n6047), .Z(y[4]) );
  NANDN U8562 ( .A(n4366), .B(creg[50]), .Z(n6050) );
  NANDN U8563 ( .A(n6157), .B(m[50]), .Z(n6049) );
  NAND U8564 ( .A(n6050), .B(n6049), .Z(y[50]) );
  NANDN U8565 ( .A(n4366), .B(creg[51]), .Z(n6052) );
  NANDN U8566 ( .A(n6157), .B(m[51]), .Z(n6051) );
  NAND U8567 ( .A(n6052), .B(n6051), .Z(y[51]) );
  NANDN U8568 ( .A(n4366), .B(creg[52]), .Z(n6054) );
  NANDN U8569 ( .A(n6157), .B(m[52]), .Z(n6053) );
  NAND U8570 ( .A(n6054), .B(n6053), .Z(y[52]) );
  NANDN U8571 ( .A(n4366), .B(creg[53]), .Z(n6056) );
  NANDN U8572 ( .A(n6157), .B(m[53]), .Z(n6055) );
  NAND U8573 ( .A(n6056), .B(n6055), .Z(y[53]) );
  NANDN U8574 ( .A(n4366), .B(creg[54]), .Z(n6058) );
  NANDN U8575 ( .A(n6157), .B(m[54]), .Z(n6057) );
  NAND U8576 ( .A(n6058), .B(n6057), .Z(y[54]) );
  NANDN U8577 ( .A(n4366), .B(creg[55]), .Z(n6060) );
  NANDN U8578 ( .A(n6157), .B(m[55]), .Z(n6059) );
  NAND U8579 ( .A(n6060), .B(n6059), .Z(y[55]) );
  NANDN U8580 ( .A(n4366), .B(creg[56]), .Z(n6062) );
  NANDN U8581 ( .A(n6157), .B(m[56]), .Z(n6061) );
  NAND U8582 ( .A(n6062), .B(n6061), .Z(y[56]) );
  NANDN U8583 ( .A(n4366), .B(creg[57]), .Z(n6064) );
  NANDN U8584 ( .A(n6157), .B(m[57]), .Z(n6063) );
  NAND U8585 ( .A(n6064), .B(n6063), .Z(y[57]) );
  NANDN U8586 ( .A(n4366), .B(creg[58]), .Z(n6066) );
  NANDN U8587 ( .A(n6157), .B(m[58]), .Z(n6065) );
  NAND U8588 ( .A(n6066), .B(n6065), .Z(y[58]) );
  NANDN U8589 ( .A(n4366), .B(creg[59]), .Z(n6068) );
  NANDN U8590 ( .A(n6157), .B(m[59]), .Z(n6067) );
  NAND U8591 ( .A(n6068), .B(n6067), .Z(y[59]) );
  NANDN U8592 ( .A(n4366), .B(creg[5]), .Z(n6070) );
  NANDN U8593 ( .A(n6157), .B(m[5]), .Z(n6069) );
  NAND U8594 ( .A(n6070), .B(n6069), .Z(y[5]) );
  NANDN U8595 ( .A(n4366), .B(creg[60]), .Z(n6072) );
  NANDN U8596 ( .A(n6157), .B(m[60]), .Z(n6071) );
  NAND U8597 ( .A(n6072), .B(n6071), .Z(y[60]) );
  NANDN U8598 ( .A(n4366), .B(creg[61]), .Z(n6074) );
  NANDN U8599 ( .A(n6157), .B(m[61]), .Z(n6073) );
  NAND U8600 ( .A(n6074), .B(n6073), .Z(y[61]) );
  NANDN U8601 ( .A(n4366), .B(creg[62]), .Z(n6076) );
  NANDN U8602 ( .A(n6157), .B(m[62]), .Z(n6075) );
  NAND U8603 ( .A(n6076), .B(n6075), .Z(y[62]) );
  NANDN U8604 ( .A(n4366), .B(creg[63]), .Z(n6078) );
  NANDN U8605 ( .A(n6157), .B(m[63]), .Z(n6077) );
  NAND U8606 ( .A(n6078), .B(n6077), .Z(y[63]) );
  NANDN U8607 ( .A(n4366), .B(creg[64]), .Z(n6080) );
  NANDN U8608 ( .A(n6157), .B(m[64]), .Z(n6079) );
  NAND U8609 ( .A(n6080), .B(n6079), .Z(y[64]) );
  NANDN U8610 ( .A(n4366), .B(creg[65]), .Z(n6082) );
  NANDN U8611 ( .A(n6157), .B(m[65]), .Z(n6081) );
  NAND U8612 ( .A(n6082), .B(n6081), .Z(y[65]) );
  NANDN U8613 ( .A(n4366), .B(creg[66]), .Z(n6084) );
  NANDN U8614 ( .A(n6157), .B(m[66]), .Z(n6083) );
  NAND U8615 ( .A(n6084), .B(n6083), .Z(y[66]) );
  NANDN U8616 ( .A(n4366), .B(creg[67]), .Z(n6086) );
  NANDN U8617 ( .A(n6157), .B(m[67]), .Z(n6085) );
  NAND U8618 ( .A(n6086), .B(n6085), .Z(y[67]) );
  NANDN U8619 ( .A(n4366), .B(creg[68]), .Z(n6088) );
  NANDN U8620 ( .A(n6157), .B(m[68]), .Z(n6087) );
  NAND U8621 ( .A(n6088), .B(n6087), .Z(y[68]) );
  NANDN U8622 ( .A(n4366), .B(creg[69]), .Z(n6090) );
  NANDN U8623 ( .A(n6157), .B(m[69]), .Z(n6089) );
  NAND U8624 ( .A(n6090), .B(n6089), .Z(y[69]) );
  NANDN U8625 ( .A(n4366), .B(creg[6]), .Z(n6092) );
  NANDN U8626 ( .A(n6157), .B(m[6]), .Z(n6091) );
  NAND U8627 ( .A(n6092), .B(n6091), .Z(y[6]) );
  NANDN U8628 ( .A(n4366), .B(creg[70]), .Z(n6094) );
  NANDN U8629 ( .A(n6157), .B(m[70]), .Z(n6093) );
  NAND U8630 ( .A(n6094), .B(n6093), .Z(y[70]) );
  NANDN U8631 ( .A(n4366), .B(creg[71]), .Z(n6096) );
  NANDN U8632 ( .A(n6157), .B(m[71]), .Z(n6095) );
  NAND U8633 ( .A(n6096), .B(n6095), .Z(y[71]) );
  NANDN U8634 ( .A(n4366), .B(creg[72]), .Z(n6098) );
  NANDN U8635 ( .A(n6157), .B(m[72]), .Z(n6097) );
  NAND U8636 ( .A(n6098), .B(n6097), .Z(y[72]) );
  NANDN U8637 ( .A(n4366), .B(creg[73]), .Z(n6100) );
  NANDN U8638 ( .A(n6157), .B(m[73]), .Z(n6099) );
  NAND U8639 ( .A(n6100), .B(n6099), .Z(y[73]) );
  NANDN U8640 ( .A(n4366), .B(creg[74]), .Z(n6102) );
  NANDN U8641 ( .A(n6157), .B(m[74]), .Z(n6101) );
  NAND U8642 ( .A(n6102), .B(n6101), .Z(y[74]) );
  NANDN U8643 ( .A(n4366), .B(creg[75]), .Z(n6104) );
  NANDN U8644 ( .A(n6157), .B(m[75]), .Z(n6103) );
  NAND U8645 ( .A(n6104), .B(n6103), .Z(y[75]) );
  NANDN U8646 ( .A(n4366), .B(creg[76]), .Z(n6106) );
  NANDN U8647 ( .A(n6157), .B(m[76]), .Z(n6105) );
  NAND U8648 ( .A(n6106), .B(n6105), .Z(y[76]) );
  NANDN U8649 ( .A(n4366), .B(creg[77]), .Z(n6108) );
  NANDN U8650 ( .A(n6157), .B(m[77]), .Z(n6107) );
  NAND U8651 ( .A(n6108), .B(n6107), .Z(y[77]) );
  NANDN U8652 ( .A(n4366), .B(creg[78]), .Z(n6110) );
  NANDN U8653 ( .A(n6157), .B(m[78]), .Z(n6109) );
  NAND U8654 ( .A(n6110), .B(n6109), .Z(y[78]) );
  NANDN U8655 ( .A(n4366), .B(creg[79]), .Z(n6112) );
  NANDN U8656 ( .A(n6157), .B(m[79]), .Z(n6111) );
  NAND U8657 ( .A(n6112), .B(n6111), .Z(y[79]) );
  NANDN U8658 ( .A(n4366), .B(creg[7]), .Z(n6114) );
  NANDN U8659 ( .A(n6157), .B(m[7]), .Z(n6113) );
  NAND U8660 ( .A(n6114), .B(n6113), .Z(y[7]) );
  NANDN U8661 ( .A(n4366), .B(creg[80]), .Z(n6116) );
  NANDN U8662 ( .A(n6157), .B(m[80]), .Z(n6115) );
  NAND U8663 ( .A(n6116), .B(n6115), .Z(y[80]) );
  NANDN U8664 ( .A(n4366), .B(creg[81]), .Z(n6118) );
  NANDN U8665 ( .A(n6157), .B(m[81]), .Z(n6117) );
  NAND U8666 ( .A(n6118), .B(n6117), .Z(y[81]) );
  NANDN U8667 ( .A(n4366), .B(creg[82]), .Z(n6120) );
  NANDN U8668 ( .A(n6157), .B(m[82]), .Z(n6119) );
  NAND U8669 ( .A(n6120), .B(n6119), .Z(y[82]) );
  NANDN U8670 ( .A(n4366), .B(creg[83]), .Z(n6122) );
  NANDN U8671 ( .A(n6157), .B(m[83]), .Z(n6121) );
  NAND U8672 ( .A(n6122), .B(n6121), .Z(y[83]) );
  NANDN U8673 ( .A(n4366), .B(creg[84]), .Z(n6124) );
  NANDN U8674 ( .A(n6157), .B(m[84]), .Z(n6123) );
  NAND U8675 ( .A(n6124), .B(n6123), .Z(y[84]) );
  NANDN U8676 ( .A(n4366), .B(creg[85]), .Z(n6126) );
  NANDN U8677 ( .A(n6157), .B(m[85]), .Z(n6125) );
  NAND U8678 ( .A(n6126), .B(n6125), .Z(y[85]) );
  NANDN U8679 ( .A(n4366), .B(creg[86]), .Z(n6128) );
  NANDN U8680 ( .A(n6157), .B(m[86]), .Z(n6127) );
  NAND U8681 ( .A(n6128), .B(n6127), .Z(y[86]) );
  NANDN U8682 ( .A(n4366), .B(creg[87]), .Z(n6130) );
  NANDN U8683 ( .A(n6157), .B(m[87]), .Z(n6129) );
  NAND U8684 ( .A(n6130), .B(n6129), .Z(y[87]) );
  NANDN U8685 ( .A(n4366), .B(creg[88]), .Z(n6132) );
  NANDN U8686 ( .A(n6157), .B(m[88]), .Z(n6131) );
  NAND U8687 ( .A(n6132), .B(n6131), .Z(y[88]) );
  NANDN U8688 ( .A(n4366), .B(creg[89]), .Z(n6134) );
  NANDN U8689 ( .A(n6157), .B(m[89]), .Z(n6133) );
  NAND U8690 ( .A(n6134), .B(n6133), .Z(y[89]) );
  NANDN U8691 ( .A(n4366), .B(creg[8]), .Z(n6136) );
  NANDN U8692 ( .A(n6157), .B(m[8]), .Z(n6135) );
  NAND U8693 ( .A(n6136), .B(n6135), .Z(y[8]) );
  NANDN U8694 ( .A(n4366), .B(creg[90]), .Z(n6138) );
  NANDN U8695 ( .A(n6157), .B(m[90]), .Z(n6137) );
  NAND U8696 ( .A(n6138), .B(n6137), .Z(y[90]) );
  NANDN U8697 ( .A(n4366), .B(creg[91]), .Z(n6140) );
  NANDN U8698 ( .A(n6157), .B(m[91]), .Z(n6139) );
  NAND U8699 ( .A(n6140), .B(n6139), .Z(y[91]) );
  NANDN U8700 ( .A(n4366), .B(creg[92]), .Z(n6142) );
  NANDN U8701 ( .A(n6157), .B(m[92]), .Z(n6141) );
  NAND U8702 ( .A(n6142), .B(n6141), .Z(y[92]) );
  NANDN U8703 ( .A(n4366), .B(creg[93]), .Z(n6144) );
  NANDN U8704 ( .A(n6157), .B(m[93]), .Z(n6143) );
  NAND U8705 ( .A(n6144), .B(n6143), .Z(y[93]) );
  NANDN U8706 ( .A(n4366), .B(creg[94]), .Z(n6146) );
  NANDN U8707 ( .A(n6157), .B(m[94]), .Z(n6145) );
  NAND U8708 ( .A(n6146), .B(n6145), .Z(y[94]) );
  NANDN U8709 ( .A(n4366), .B(creg[95]), .Z(n6148) );
  NANDN U8710 ( .A(n6157), .B(m[95]), .Z(n6147) );
  NAND U8711 ( .A(n6148), .B(n6147), .Z(y[95]) );
  NANDN U8712 ( .A(n4366), .B(creg[96]), .Z(n6150) );
  NANDN U8713 ( .A(n6157), .B(m[96]), .Z(n6149) );
  NAND U8714 ( .A(n6150), .B(n6149), .Z(y[96]) );
  NANDN U8715 ( .A(n4366), .B(creg[97]), .Z(n6152) );
  NANDN U8716 ( .A(n6157), .B(m[97]), .Z(n6151) );
  NAND U8717 ( .A(n6152), .B(n6151), .Z(y[97]) );
  NANDN U8718 ( .A(n4366), .B(creg[98]), .Z(n6154) );
  NANDN U8719 ( .A(n6157), .B(m[98]), .Z(n6153) );
  NAND U8720 ( .A(n6154), .B(n6153), .Z(y[98]) );
  NANDN U8721 ( .A(n4366), .B(creg[99]), .Z(n6156) );
  NANDN U8722 ( .A(n6157), .B(m[99]), .Z(n6155) );
  NAND U8723 ( .A(n6156), .B(n6155), .Z(y[99]) );
  NANDN U8724 ( .A(n4366), .B(creg[9]), .Z(n6159) );
  NANDN U8725 ( .A(n6157), .B(m[9]), .Z(n6158) );
  NAND U8726 ( .A(n6159), .B(n6158), .Z(y[9]) );
  AND U8727 ( .A(start_reg[127]), .B(init), .Z(start_in[127]) );
  AND U8728 ( .A(first_one), .B(start_in[127]), .Z(n6161) );
  IV U8729 ( .A(mul_pow), .Z(n8214) );
  OR U8730 ( .A(ereg[255]), .B(n8214), .Z(n6160) );
  AND U8731 ( .A(n6161), .B(n6160), .Z(n7183) );
  NANDN U8732 ( .A(n7183), .B(init), .Z(n7182) );
  ANDN U8733 ( .B(creg[255]), .A(n7182), .Z(n6165) );
  NAND U8734 ( .A(o[255]), .B(n7183), .Z(n6163) );
  ANDN U8735 ( .B(n6163), .A(n6162), .Z(n6164) );
  NANDN U8736 ( .A(n6165), .B(n6164), .Z(n1801) );
  NANDN U8737 ( .A(n7182), .B(creg[254]), .Z(n6167) );
  NAND U8738 ( .A(n7183), .B(o[254]), .Z(n6166) );
  AND U8739 ( .A(n6167), .B(n6166), .Z(n6168) );
  NANDN U8740 ( .A(n6169), .B(n6168), .Z(n1802) );
  NANDN U8741 ( .A(n7182), .B(creg[253]), .Z(n6171) );
  NAND U8742 ( .A(n7183), .B(o[253]), .Z(n6170) );
  AND U8743 ( .A(n6171), .B(n6170), .Z(n6172) );
  NANDN U8744 ( .A(n6173), .B(n6172), .Z(n1803) );
  NANDN U8745 ( .A(n7182), .B(creg[252]), .Z(n6175) );
  NAND U8746 ( .A(n7183), .B(o[252]), .Z(n6174) );
  AND U8747 ( .A(n6175), .B(n6174), .Z(n6176) );
  NANDN U8748 ( .A(n6177), .B(n6176), .Z(n1804) );
  NANDN U8749 ( .A(n7182), .B(creg[251]), .Z(n6179) );
  NAND U8750 ( .A(n7183), .B(o[251]), .Z(n6178) );
  AND U8751 ( .A(n6179), .B(n6178), .Z(n6180) );
  NANDN U8752 ( .A(n6181), .B(n6180), .Z(n1805) );
  NANDN U8753 ( .A(n7182), .B(creg[250]), .Z(n6183) );
  NAND U8754 ( .A(n7183), .B(o[250]), .Z(n6182) );
  AND U8755 ( .A(n6183), .B(n6182), .Z(n6184) );
  NANDN U8756 ( .A(n6185), .B(n6184), .Z(n1806) );
  NANDN U8757 ( .A(n7182), .B(creg[249]), .Z(n6187) );
  NAND U8758 ( .A(n7183), .B(o[249]), .Z(n6186) );
  AND U8759 ( .A(n6187), .B(n6186), .Z(n6188) );
  NANDN U8760 ( .A(n6189), .B(n6188), .Z(n1807) );
  NANDN U8761 ( .A(n7182), .B(creg[248]), .Z(n6191) );
  NAND U8762 ( .A(n7183), .B(o[248]), .Z(n6190) );
  AND U8763 ( .A(n6191), .B(n6190), .Z(n6192) );
  NANDN U8764 ( .A(n6193), .B(n6192), .Z(n1808) );
  NANDN U8765 ( .A(n7182), .B(creg[247]), .Z(n6195) );
  NAND U8766 ( .A(n7183), .B(o[247]), .Z(n6194) );
  AND U8767 ( .A(n6195), .B(n6194), .Z(n6196) );
  NANDN U8768 ( .A(n6197), .B(n6196), .Z(n1809) );
  NANDN U8769 ( .A(n7182), .B(creg[246]), .Z(n6199) );
  NAND U8770 ( .A(n7183), .B(o[246]), .Z(n6198) );
  AND U8771 ( .A(n6199), .B(n6198), .Z(n6200) );
  NANDN U8772 ( .A(n6201), .B(n6200), .Z(n1810) );
  NANDN U8773 ( .A(n7182), .B(creg[245]), .Z(n6203) );
  NAND U8774 ( .A(n7183), .B(o[245]), .Z(n6202) );
  AND U8775 ( .A(n6203), .B(n6202), .Z(n6204) );
  NANDN U8776 ( .A(n6205), .B(n6204), .Z(n1811) );
  NANDN U8777 ( .A(n7182), .B(creg[244]), .Z(n6207) );
  NAND U8778 ( .A(n7183), .B(o[244]), .Z(n6206) );
  AND U8779 ( .A(n6207), .B(n6206), .Z(n6208) );
  NANDN U8780 ( .A(n6209), .B(n6208), .Z(n1812) );
  NANDN U8781 ( .A(n7182), .B(creg[243]), .Z(n6211) );
  NAND U8782 ( .A(n7183), .B(o[243]), .Z(n6210) );
  AND U8783 ( .A(n6211), .B(n6210), .Z(n6212) );
  NANDN U8784 ( .A(n6213), .B(n6212), .Z(n1813) );
  NANDN U8785 ( .A(n7182), .B(creg[242]), .Z(n6215) );
  NAND U8786 ( .A(n7183), .B(o[242]), .Z(n6214) );
  AND U8787 ( .A(n6215), .B(n6214), .Z(n6216) );
  NANDN U8788 ( .A(n6217), .B(n6216), .Z(n1814) );
  NANDN U8789 ( .A(n7182), .B(creg[241]), .Z(n6219) );
  NAND U8790 ( .A(n7183), .B(o[241]), .Z(n6218) );
  AND U8791 ( .A(n6219), .B(n6218), .Z(n6220) );
  NANDN U8792 ( .A(n6221), .B(n6220), .Z(n1815) );
  NANDN U8793 ( .A(n7182), .B(creg[240]), .Z(n6223) );
  NAND U8794 ( .A(n7183), .B(o[240]), .Z(n6222) );
  AND U8795 ( .A(n6223), .B(n6222), .Z(n6224) );
  NANDN U8796 ( .A(n6225), .B(n6224), .Z(n1816) );
  NANDN U8797 ( .A(n7182), .B(creg[239]), .Z(n6227) );
  NAND U8798 ( .A(n7183), .B(o[239]), .Z(n6226) );
  AND U8799 ( .A(n6227), .B(n6226), .Z(n6228) );
  NANDN U8800 ( .A(n6229), .B(n6228), .Z(n1817) );
  NANDN U8801 ( .A(n7182), .B(creg[238]), .Z(n6231) );
  NAND U8802 ( .A(n7183), .B(o[238]), .Z(n6230) );
  AND U8803 ( .A(n6231), .B(n6230), .Z(n6232) );
  NANDN U8804 ( .A(n6233), .B(n6232), .Z(n1818) );
  NANDN U8805 ( .A(n7182), .B(creg[237]), .Z(n6235) );
  NAND U8806 ( .A(n7183), .B(o[237]), .Z(n6234) );
  AND U8807 ( .A(n6235), .B(n6234), .Z(n6236) );
  NANDN U8808 ( .A(n6237), .B(n6236), .Z(n1819) );
  NANDN U8809 ( .A(n7182), .B(creg[236]), .Z(n6239) );
  NAND U8810 ( .A(n7183), .B(o[236]), .Z(n6238) );
  AND U8811 ( .A(n6239), .B(n6238), .Z(n6240) );
  NANDN U8812 ( .A(n6241), .B(n6240), .Z(n1820) );
  NANDN U8813 ( .A(n7182), .B(creg[235]), .Z(n6243) );
  NAND U8814 ( .A(n7183), .B(o[235]), .Z(n6242) );
  AND U8815 ( .A(n6243), .B(n6242), .Z(n6244) );
  NANDN U8816 ( .A(n6245), .B(n6244), .Z(n1821) );
  NANDN U8817 ( .A(n7182), .B(creg[234]), .Z(n6247) );
  NAND U8818 ( .A(n7183), .B(o[234]), .Z(n6246) );
  AND U8819 ( .A(n6247), .B(n6246), .Z(n6248) );
  NANDN U8820 ( .A(n6249), .B(n6248), .Z(n1822) );
  NANDN U8821 ( .A(n7182), .B(creg[233]), .Z(n6251) );
  NAND U8822 ( .A(n7183), .B(o[233]), .Z(n6250) );
  AND U8823 ( .A(n6251), .B(n6250), .Z(n6252) );
  NANDN U8824 ( .A(n6253), .B(n6252), .Z(n1823) );
  NANDN U8825 ( .A(n7182), .B(creg[232]), .Z(n6255) );
  NAND U8826 ( .A(n7183), .B(o[232]), .Z(n6254) );
  AND U8827 ( .A(n6255), .B(n6254), .Z(n6256) );
  NANDN U8828 ( .A(n6257), .B(n6256), .Z(n1824) );
  NANDN U8829 ( .A(n7182), .B(creg[231]), .Z(n6259) );
  NAND U8830 ( .A(n7183), .B(o[231]), .Z(n6258) );
  AND U8831 ( .A(n6259), .B(n6258), .Z(n6260) );
  NANDN U8832 ( .A(n6261), .B(n6260), .Z(n1825) );
  NANDN U8833 ( .A(n7182), .B(creg[230]), .Z(n6263) );
  NAND U8834 ( .A(n7183), .B(o[230]), .Z(n6262) );
  AND U8835 ( .A(n6263), .B(n6262), .Z(n6264) );
  NANDN U8836 ( .A(n6265), .B(n6264), .Z(n1826) );
  NANDN U8837 ( .A(n7182), .B(creg[229]), .Z(n6267) );
  NAND U8838 ( .A(n7183), .B(o[229]), .Z(n6266) );
  AND U8839 ( .A(n6267), .B(n6266), .Z(n6268) );
  NANDN U8840 ( .A(n6269), .B(n6268), .Z(n1827) );
  NANDN U8841 ( .A(n7182), .B(creg[228]), .Z(n6271) );
  NAND U8842 ( .A(n7183), .B(o[228]), .Z(n6270) );
  AND U8843 ( .A(n6271), .B(n6270), .Z(n6272) );
  NANDN U8844 ( .A(n6273), .B(n6272), .Z(n1828) );
  NANDN U8845 ( .A(n7182), .B(creg[227]), .Z(n6275) );
  NAND U8846 ( .A(n7183), .B(o[227]), .Z(n6274) );
  AND U8847 ( .A(n6275), .B(n6274), .Z(n6276) );
  NANDN U8848 ( .A(n6277), .B(n6276), .Z(n1829) );
  NANDN U8849 ( .A(n7182), .B(creg[226]), .Z(n6279) );
  NAND U8850 ( .A(n7183), .B(o[226]), .Z(n6278) );
  AND U8851 ( .A(n6279), .B(n6278), .Z(n6280) );
  NANDN U8852 ( .A(n6281), .B(n6280), .Z(n1830) );
  NANDN U8853 ( .A(n7182), .B(creg[225]), .Z(n6283) );
  NAND U8854 ( .A(n7183), .B(o[225]), .Z(n6282) );
  AND U8855 ( .A(n6283), .B(n6282), .Z(n6284) );
  NANDN U8856 ( .A(n6285), .B(n6284), .Z(n1831) );
  NANDN U8857 ( .A(n7182), .B(creg[224]), .Z(n6287) );
  NAND U8858 ( .A(n7183), .B(o[224]), .Z(n6286) );
  AND U8859 ( .A(n6287), .B(n6286), .Z(n6288) );
  NANDN U8860 ( .A(n6289), .B(n6288), .Z(n1832) );
  NANDN U8861 ( .A(n7182), .B(creg[223]), .Z(n6291) );
  NAND U8862 ( .A(n7183), .B(o[223]), .Z(n6290) );
  AND U8863 ( .A(n6291), .B(n6290), .Z(n6292) );
  NANDN U8864 ( .A(n6293), .B(n6292), .Z(n1833) );
  NANDN U8865 ( .A(n7182), .B(creg[222]), .Z(n6295) );
  NAND U8866 ( .A(n7183), .B(o[222]), .Z(n6294) );
  AND U8867 ( .A(n6295), .B(n6294), .Z(n6296) );
  NANDN U8868 ( .A(n6297), .B(n6296), .Z(n1834) );
  NANDN U8869 ( .A(n7182), .B(creg[221]), .Z(n6299) );
  NAND U8870 ( .A(n7183), .B(o[221]), .Z(n6298) );
  AND U8871 ( .A(n6299), .B(n6298), .Z(n6300) );
  NANDN U8872 ( .A(n6301), .B(n6300), .Z(n1835) );
  NANDN U8873 ( .A(n7182), .B(creg[220]), .Z(n6303) );
  NAND U8874 ( .A(n7183), .B(o[220]), .Z(n6302) );
  AND U8875 ( .A(n6303), .B(n6302), .Z(n6304) );
  NANDN U8876 ( .A(n6305), .B(n6304), .Z(n1836) );
  NANDN U8877 ( .A(n7182), .B(creg[219]), .Z(n6307) );
  NAND U8878 ( .A(n7183), .B(o[219]), .Z(n6306) );
  AND U8879 ( .A(n6307), .B(n6306), .Z(n6308) );
  NANDN U8880 ( .A(n6309), .B(n6308), .Z(n1837) );
  NANDN U8881 ( .A(n7182), .B(creg[218]), .Z(n6311) );
  NAND U8882 ( .A(n7183), .B(o[218]), .Z(n6310) );
  AND U8883 ( .A(n6311), .B(n6310), .Z(n6312) );
  NANDN U8884 ( .A(n6313), .B(n6312), .Z(n1838) );
  NANDN U8885 ( .A(n7182), .B(creg[217]), .Z(n6315) );
  NAND U8886 ( .A(n7183), .B(o[217]), .Z(n6314) );
  AND U8887 ( .A(n6315), .B(n6314), .Z(n6316) );
  NANDN U8888 ( .A(n6317), .B(n6316), .Z(n1839) );
  NANDN U8889 ( .A(n7182), .B(creg[216]), .Z(n6319) );
  NAND U8890 ( .A(n7183), .B(o[216]), .Z(n6318) );
  AND U8891 ( .A(n6319), .B(n6318), .Z(n6320) );
  NANDN U8892 ( .A(n6321), .B(n6320), .Z(n1840) );
  NANDN U8893 ( .A(n7182), .B(creg[215]), .Z(n6323) );
  NAND U8894 ( .A(n7183), .B(o[215]), .Z(n6322) );
  AND U8895 ( .A(n6323), .B(n6322), .Z(n6324) );
  NANDN U8896 ( .A(n6325), .B(n6324), .Z(n1841) );
  NANDN U8897 ( .A(n7182), .B(creg[214]), .Z(n6327) );
  NAND U8898 ( .A(n7183), .B(o[214]), .Z(n6326) );
  AND U8899 ( .A(n6327), .B(n6326), .Z(n6328) );
  NANDN U8900 ( .A(n6329), .B(n6328), .Z(n1842) );
  NANDN U8901 ( .A(n7182), .B(creg[213]), .Z(n6331) );
  NAND U8902 ( .A(n7183), .B(o[213]), .Z(n6330) );
  AND U8903 ( .A(n6331), .B(n6330), .Z(n6332) );
  NANDN U8904 ( .A(n6333), .B(n6332), .Z(n1843) );
  NANDN U8905 ( .A(n7182), .B(creg[212]), .Z(n6335) );
  NAND U8906 ( .A(n7183), .B(o[212]), .Z(n6334) );
  AND U8907 ( .A(n6335), .B(n6334), .Z(n6336) );
  NANDN U8908 ( .A(n6337), .B(n6336), .Z(n1844) );
  NANDN U8909 ( .A(n7182), .B(creg[211]), .Z(n6339) );
  NAND U8910 ( .A(n7183), .B(o[211]), .Z(n6338) );
  AND U8911 ( .A(n6339), .B(n6338), .Z(n6340) );
  NANDN U8912 ( .A(n6341), .B(n6340), .Z(n1845) );
  NANDN U8913 ( .A(n7182), .B(creg[210]), .Z(n6343) );
  NAND U8914 ( .A(n7183), .B(o[210]), .Z(n6342) );
  AND U8915 ( .A(n6343), .B(n6342), .Z(n6344) );
  NANDN U8916 ( .A(n6345), .B(n6344), .Z(n1846) );
  NANDN U8917 ( .A(n7182), .B(creg[209]), .Z(n6347) );
  NAND U8918 ( .A(n7183), .B(o[209]), .Z(n6346) );
  AND U8919 ( .A(n6347), .B(n6346), .Z(n6348) );
  NANDN U8920 ( .A(n6349), .B(n6348), .Z(n1847) );
  NANDN U8921 ( .A(n7182), .B(creg[208]), .Z(n6351) );
  NAND U8922 ( .A(n7183), .B(o[208]), .Z(n6350) );
  AND U8923 ( .A(n6351), .B(n6350), .Z(n6352) );
  NANDN U8924 ( .A(n6353), .B(n6352), .Z(n1848) );
  NANDN U8925 ( .A(n7182), .B(creg[207]), .Z(n6355) );
  NAND U8926 ( .A(n7183), .B(o[207]), .Z(n6354) );
  AND U8927 ( .A(n6355), .B(n6354), .Z(n6356) );
  NANDN U8928 ( .A(n6357), .B(n6356), .Z(n1849) );
  NANDN U8929 ( .A(n7182), .B(creg[206]), .Z(n6359) );
  NAND U8930 ( .A(n7183), .B(o[206]), .Z(n6358) );
  AND U8931 ( .A(n6359), .B(n6358), .Z(n6360) );
  NANDN U8932 ( .A(n6361), .B(n6360), .Z(n1850) );
  NANDN U8933 ( .A(n7182), .B(creg[205]), .Z(n6363) );
  NAND U8934 ( .A(n7183), .B(o[205]), .Z(n6362) );
  AND U8935 ( .A(n6363), .B(n6362), .Z(n6364) );
  NANDN U8936 ( .A(n6365), .B(n6364), .Z(n1851) );
  NANDN U8937 ( .A(n7182), .B(creg[204]), .Z(n6367) );
  NAND U8938 ( .A(n7183), .B(o[204]), .Z(n6366) );
  AND U8939 ( .A(n6367), .B(n6366), .Z(n6368) );
  NANDN U8940 ( .A(n6369), .B(n6368), .Z(n1852) );
  NANDN U8941 ( .A(n7182), .B(creg[203]), .Z(n6371) );
  NAND U8942 ( .A(n7183), .B(o[203]), .Z(n6370) );
  AND U8943 ( .A(n6371), .B(n6370), .Z(n6372) );
  NANDN U8944 ( .A(n6373), .B(n6372), .Z(n1853) );
  NANDN U8945 ( .A(n7182), .B(creg[202]), .Z(n6375) );
  NAND U8946 ( .A(n7183), .B(o[202]), .Z(n6374) );
  AND U8947 ( .A(n6375), .B(n6374), .Z(n6376) );
  NANDN U8948 ( .A(n6377), .B(n6376), .Z(n1854) );
  NANDN U8949 ( .A(n7182), .B(creg[201]), .Z(n6379) );
  NAND U8950 ( .A(n7183), .B(o[201]), .Z(n6378) );
  AND U8951 ( .A(n6379), .B(n6378), .Z(n6380) );
  NANDN U8952 ( .A(n6381), .B(n6380), .Z(n1855) );
  NANDN U8953 ( .A(n7182), .B(creg[200]), .Z(n6383) );
  NAND U8954 ( .A(n7183), .B(o[200]), .Z(n6382) );
  AND U8955 ( .A(n6383), .B(n6382), .Z(n6384) );
  NANDN U8956 ( .A(n6385), .B(n6384), .Z(n1856) );
  NANDN U8957 ( .A(n7182), .B(creg[199]), .Z(n6387) );
  NAND U8958 ( .A(n7183), .B(o[199]), .Z(n6386) );
  AND U8959 ( .A(n6387), .B(n6386), .Z(n6388) );
  NANDN U8960 ( .A(n6389), .B(n6388), .Z(n1857) );
  NANDN U8961 ( .A(n7182), .B(creg[198]), .Z(n6391) );
  NAND U8962 ( .A(n7183), .B(o[198]), .Z(n6390) );
  AND U8963 ( .A(n6391), .B(n6390), .Z(n6392) );
  NANDN U8964 ( .A(n6393), .B(n6392), .Z(n1858) );
  NANDN U8965 ( .A(n7182), .B(creg[197]), .Z(n6395) );
  NAND U8966 ( .A(n7183), .B(o[197]), .Z(n6394) );
  AND U8967 ( .A(n6395), .B(n6394), .Z(n6396) );
  NANDN U8968 ( .A(n6397), .B(n6396), .Z(n1859) );
  NANDN U8969 ( .A(n7182), .B(creg[196]), .Z(n6399) );
  NAND U8970 ( .A(n7183), .B(o[196]), .Z(n6398) );
  AND U8971 ( .A(n6399), .B(n6398), .Z(n6400) );
  NANDN U8972 ( .A(n6401), .B(n6400), .Z(n1860) );
  NANDN U8973 ( .A(n7182), .B(creg[195]), .Z(n6403) );
  NAND U8974 ( .A(n7183), .B(o[195]), .Z(n6402) );
  AND U8975 ( .A(n6403), .B(n6402), .Z(n6404) );
  NANDN U8976 ( .A(n6405), .B(n6404), .Z(n1861) );
  NANDN U8977 ( .A(n7182), .B(creg[194]), .Z(n6407) );
  NAND U8978 ( .A(n7183), .B(o[194]), .Z(n6406) );
  AND U8979 ( .A(n6407), .B(n6406), .Z(n6408) );
  NANDN U8980 ( .A(n6409), .B(n6408), .Z(n1862) );
  NANDN U8981 ( .A(n7182), .B(creg[193]), .Z(n6411) );
  NAND U8982 ( .A(n7183), .B(o[193]), .Z(n6410) );
  AND U8983 ( .A(n6411), .B(n6410), .Z(n6412) );
  NANDN U8984 ( .A(n6413), .B(n6412), .Z(n1863) );
  NANDN U8985 ( .A(n7182), .B(creg[192]), .Z(n6415) );
  NAND U8986 ( .A(n7183), .B(o[192]), .Z(n6414) );
  AND U8987 ( .A(n6415), .B(n6414), .Z(n6416) );
  NANDN U8988 ( .A(n6417), .B(n6416), .Z(n1864) );
  NANDN U8989 ( .A(n7182), .B(creg[191]), .Z(n6419) );
  NAND U8990 ( .A(n7183), .B(o[191]), .Z(n6418) );
  AND U8991 ( .A(n6419), .B(n6418), .Z(n6420) );
  NANDN U8992 ( .A(n6421), .B(n6420), .Z(n1865) );
  NANDN U8993 ( .A(n7182), .B(creg[190]), .Z(n6423) );
  NAND U8994 ( .A(n7183), .B(o[190]), .Z(n6422) );
  AND U8995 ( .A(n6423), .B(n6422), .Z(n6424) );
  NANDN U8996 ( .A(n6425), .B(n6424), .Z(n1866) );
  NANDN U8997 ( .A(n7182), .B(creg[189]), .Z(n6427) );
  NAND U8998 ( .A(n7183), .B(o[189]), .Z(n6426) );
  AND U8999 ( .A(n6427), .B(n6426), .Z(n6428) );
  NANDN U9000 ( .A(n6429), .B(n6428), .Z(n1867) );
  NANDN U9001 ( .A(n7182), .B(creg[188]), .Z(n6431) );
  NAND U9002 ( .A(n7183), .B(o[188]), .Z(n6430) );
  AND U9003 ( .A(n6431), .B(n6430), .Z(n6432) );
  NANDN U9004 ( .A(n6433), .B(n6432), .Z(n1868) );
  NANDN U9005 ( .A(n7182), .B(creg[187]), .Z(n6435) );
  NAND U9006 ( .A(n7183), .B(o[187]), .Z(n6434) );
  AND U9007 ( .A(n6435), .B(n6434), .Z(n6436) );
  NANDN U9008 ( .A(n6437), .B(n6436), .Z(n1869) );
  NANDN U9009 ( .A(n7182), .B(creg[186]), .Z(n6439) );
  NAND U9010 ( .A(n7183), .B(o[186]), .Z(n6438) );
  AND U9011 ( .A(n6439), .B(n6438), .Z(n6440) );
  NANDN U9012 ( .A(n6441), .B(n6440), .Z(n1870) );
  NANDN U9013 ( .A(n7182), .B(creg[185]), .Z(n6443) );
  NAND U9014 ( .A(n7183), .B(o[185]), .Z(n6442) );
  AND U9015 ( .A(n6443), .B(n6442), .Z(n6444) );
  NANDN U9016 ( .A(n6445), .B(n6444), .Z(n1871) );
  NANDN U9017 ( .A(n7182), .B(creg[184]), .Z(n6447) );
  NAND U9018 ( .A(n7183), .B(o[184]), .Z(n6446) );
  AND U9019 ( .A(n6447), .B(n6446), .Z(n6448) );
  NANDN U9020 ( .A(n6449), .B(n6448), .Z(n1872) );
  NANDN U9021 ( .A(n7182), .B(creg[183]), .Z(n6451) );
  NAND U9022 ( .A(n7183), .B(o[183]), .Z(n6450) );
  AND U9023 ( .A(n6451), .B(n6450), .Z(n6452) );
  NANDN U9024 ( .A(n6453), .B(n6452), .Z(n1873) );
  NANDN U9025 ( .A(n7182), .B(creg[182]), .Z(n6455) );
  NAND U9026 ( .A(n7183), .B(o[182]), .Z(n6454) );
  AND U9027 ( .A(n6455), .B(n6454), .Z(n6456) );
  NANDN U9028 ( .A(n6457), .B(n6456), .Z(n1874) );
  NANDN U9029 ( .A(n7182), .B(creg[181]), .Z(n6459) );
  NAND U9030 ( .A(n7183), .B(o[181]), .Z(n6458) );
  AND U9031 ( .A(n6459), .B(n6458), .Z(n6460) );
  NANDN U9032 ( .A(n6461), .B(n6460), .Z(n1875) );
  NANDN U9033 ( .A(n7182), .B(creg[180]), .Z(n6463) );
  NAND U9034 ( .A(n7183), .B(o[180]), .Z(n6462) );
  AND U9035 ( .A(n6463), .B(n6462), .Z(n6464) );
  NANDN U9036 ( .A(n6465), .B(n6464), .Z(n1876) );
  NANDN U9037 ( .A(n7182), .B(creg[179]), .Z(n6467) );
  NAND U9038 ( .A(n7183), .B(o[179]), .Z(n6466) );
  AND U9039 ( .A(n6467), .B(n6466), .Z(n6468) );
  NANDN U9040 ( .A(n6469), .B(n6468), .Z(n1877) );
  NANDN U9041 ( .A(n7182), .B(creg[178]), .Z(n6471) );
  NAND U9042 ( .A(n7183), .B(o[178]), .Z(n6470) );
  AND U9043 ( .A(n6471), .B(n6470), .Z(n6472) );
  NANDN U9044 ( .A(n6473), .B(n6472), .Z(n1878) );
  NANDN U9045 ( .A(n7182), .B(creg[177]), .Z(n6475) );
  NAND U9046 ( .A(n7183), .B(o[177]), .Z(n6474) );
  AND U9047 ( .A(n6475), .B(n6474), .Z(n6476) );
  NANDN U9048 ( .A(n6477), .B(n6476), .Z(n1879) );
  NANDN U9049 ( .A(n7182), .B(creg[176]), .Z(n6479) );
  NAND U9050 ( .A(n7183), .B(o[176]), .Z(n6478) );
  AND U9051 ( .A(n6479), .B(n6478), .Z(n6480) );
  NANDN U9052 ( .A(n6481), .B(n6480), .Z(n1880) );
  NANDN U9053 ( .A(n7182), .B(creg[175]), .Z(n6483) );
  NAND U9054 ( .A(n7183), .B(o[175]), .Z(n6482) );
  AND U9055 ( .A(n6483), .B(n6482), .Z(n6484) );
  NANDN U9056 ( .A(n6485), .B(n6484), .Z(n1881) );
  NANDN U9057 ( .A(n7182), .B(creg[174]), .Z(n6487) );
  NAND U9058 ( .A(n7183), .B(o[174]), .Z(n6486) );
  AND U9059 ( .A(n6487), .B(n6486), .Z(n6488) );
  NANDN U9060 ( .A(n6489), .B(n6488), .Z(n1882) );
  NANDN U9061 ( .A(n7182), .B(creg[173]), .Z(n6491) );
  NAND U9062 ( .A(n7183), .B(o[173]), .Z(n6490) );
  AND U9063 ( .A(n6491), .B(n6490), .Z(n6492) );
  NANDN U9064 ( .A(n6493), .B(n6492), .Z(n1883) );
  NANDN U9065 ( .A(n7182), .B(creg[172]), .Z(n6495) );
  NAND U9066 ( .A(n7183), .B(o[172]), .Z(n6494) );
  AND U9067 ( .A(n6495), .B(n6494), .Z(n6496) );
  NANDN U9068 ( .A(n6497), .B(n6496), .Z(n1884) );
  NANDN U9069 ( .A(n7182), .B(creg[171]), .Z(n6499) );
  NAND U9070 ( .A(n7183), .B(o[171]), .Z(n6498) );
  AND U9071 ( .A(n6499), .B(n6498), .Z(n6500) );
  NANDN U9072 ( .A(n6501), .B(n6500), .Z(n1885) );
  NANDN U9073 ( .A(n7182), .B(creg[170]), .Z(n6503) );
  NAND U9074 ( .A(n7183), .B(o[170]), .Z(n6502) );
  AND U9075 ( .A(n6503), .B(n6502), .Z(n6504) );
  NANDN U9076 ( .A(n6505), .B(n6504), .Z(n1886) );
  NANDN U9077 ( .A(n7182), .B(creg[169]), .Z(n6507) );
  NAND U9078 ( .A(n7183), .B(o[169]), .Z(n6506) );
  AND U9079 ( .A(n6507), .B(n6506), .Z(n6508) );
  NANDN U9080 ( .A(n6509), .B(n6508), .Z(n1887) );
  NANDN U9081 ( .A(n7182), .B(creg[168]), .Z(n6511) );
  NAND U9082 ( .A(n7183), .B(o[168]), .Z(n6510) );
  AND U9083 ( .A(n6511), .B(n6510), .Z(n6512) );
  NANDN U9084 ( .A(n6513), .B(n6512), .Z(n1888) );
  NANDN U9085 ( .A(n7182), .B(creg[167]), .Z(n6515) );
  NAND U9086 ( .A(n7183), .B(o[167]), .Z(n6514) );
  AND U9087 ( .A(n6515), .B(n6514), .Z(n6516) );
  NANDN U9088 ( .A(n6517), .B(n6516), .Z(n1889) );
  NANDN U9089 ( .A(n7182), .B(creg[166]), .Z(n6519) );
  NAND U9090 ( .A(n7183), .B(o[166]), .Z(n6518) );
  AND U9091 ( .A(n6519), .B(n6518), .Z(n6520) );
  NANDN U9092 ( .A(n6521), .B(n6520), .Z(n1890) );
  NANDN U9093 ( .A(n7182), .B(creg[165]), .Z(n6523) );
  NAND U9094 ( .A(n7183), .B(o[165]), .Z(n6522) );
  AND U9095 ( .A(n6523), .B(n6522), .Z(n6524) );
  NANDN U9096 ( .A(n6525), .B(n6524), .Z(n1891) );
  NANDN U9097 ( .A(n7182), .B(creg[164]), .Z(n6527) );
  NAND U9098 ( .A(n7183), .B(o[164]), .Z(n6526) );
  AND U9099 ( .A(n6527), .B(n6526), .Z(n6528) );
  NANDN U9100 ( .A(n6529), .B(n6528), .Z(n1892) );
  NANDN U9101 ( .A(n7182), .B(creg[163]), .Z(n6531) );
  NAND U9102 ( .A(n7183), .B(o[163]), .Z(n6530) );
  AND U9103 ( .A(n6531), .B(n6530), .Z(n6532) );
  NANDN U9104 ( .A(n6533), .B(n6532), .Z(n1893) );
  NANDN U9105 ( .A(n7182), .B(creg[162]), .Z(n6535) );
  NAND U9106 ( .A(n7183), .B(o[162]), .Z(n6534) );
  AND U9107 ( .A(n6535), .B(n6534), .Z(n6536) );
  NANDN U9108 ( .A(n6537), .B(n6536), .Z(n1894) );
  NANDN U9109 ( .A(n7182), .B(creg[161]), .Z(n6539) );
  NAND U9110 ( .A(n7183), .B(o[161]), .Z(n6538) );
  AND U9111 ( .A(n6539), .B(n6538), .Z(n6540) );
  NANDN U9112 ( .A(n6541), .B(n6540), .Z(n1895) );
  NANDN U9113 ( .A(n7182), .B(creg[160]), .Z(n6543) );
  NAND U9114 ( .A(n7183), .B(o[160]), .Z(n6542) );
  AND U9115 ( .A(n6543), .B(n6542), .Z(n6544) );
  NANDN U9116 ( .A(n6545), .B(n6544), .Z(n1896) );
  NANDN U9117 ( .A(n7182), .B(creg[159]), .Z(n6547) );
  NAND U9118 ( .A(n7183), .B(o[159]), .Z(n6546) );
  AND U9119 ( .A(n6547), .B(n6546), .Z(n6548) );
  NANDN U9120 ( .A(n6549), .B(n6548), .Z(n1897) );
  NANDN U9121 ( .A(n7182), .B(creg[158]), .Z(n6551) );
  NAND U9122 ( .A(n7183), .B(o[158]), .Z(n6550) );
  AND U9123 ( .A(n6551), .B(n6550), .Z(n6552) );
  NANDN U9124 ( .A(n6553), .B(n6552), .Z(n1898) );
  NANDN U9125 ( .A(n7182), .B(creg[157]), .Z(n6555) );
  NAND U9126 ( .A(n7183), .B(o[157]), .Z(n6554) );
  AND U9127 ( .A(n6555), .B(n6554), .Z(n6556) );
  NANDN U9128 ( .A(n6557), .B(n6556), .Z(n1899) );
  NANDN U9129 ( .A(n7182), .B(creg[156]), .Z(n6559) );
  NAND U9130 ( .A(n7183), .B(o[156]), .Z(n6558) );
  AND U9131 ( .A(n6559), .B(n6558), .Z(n6560) );
  NANDN U9132 ( .A(n6561), .B(n6560), .Z(n1900) );
  NANDN U9133 ( .A(n7182), .B(creg[155]), .Z(n6563) );
  NAND U9134 ( .A(n7183), .B(o[155]), .Z(n6562) );
  AND U9135 ( .A(n6563), .B(n6562), .Z(n6564) );
  NANDN U9136 ( .A(n6565), .B(n6564), .Z(n1901) );
  NANDN U9137 ( .A(n7182), .B(creg[154]), .Z(n6567) );
  NAND U9138 ( .A(n7183), .B(o[154]), .Z(n6566) );
  AND U9139 ( .A(n6567), .B(n6566), .Z(n6568) );
  NANDN U9140 ( .A(n6569), .B(n6568), .Z(n1902) );
  NANDN U9141 ( .A(n7182), .B(creg[153]), .Z(n6571) );
  NAND U9142 ( .A(n7183), .B(o[153]), .Z(n6570) );
  AND U9143 ( .A(n6571), .B(n6570), .Z(n6572) );
  NANDN U9144 ( .A(n6573), .B(n6572), .Z(n1903) );
  NANDN U9145 ( .A(n7182), .B(creg[152]), .Z(n6575) );
  NAND U9146 ( .A(n7183), .B(o[152]), .Z(n6574) );
  AND U9147 ( .A(n6575), .B(n6574), .Z(n6576) );
  NANDN U9148 ( .A(n6577), .B(n6576), .Z(n1904) );
  NANDN U9149 ( .A(n7182), .B(creg[151]), .Z(n6579) );
  NAND U9150 ( .A(n7183), .B(o[151]), .Z(n6578) );
  AND U9151 ( .A(n6579), .B(n6578), .Z(n6580) );
  NANDN U9152 ( .A(n6581), .B(n6580), .Z(n1905) );
  NANDN U9153 ( .A(n7182), .B(creg[150]), .Z(n6583) );
  NAND U9154 ( .A(n7183), .B(o[150]), .Z(n6582) );
  AND U9155 ( .A(n6583), .B(n6582), .Z(n6584) );
  NANDN U9156 ( .A(n6585), .B(n6584), .Z(n1906) );
  NANDN U9157 ( .A(n7182), .B(creg[149]), .Z(n6587) );
  NAND U9158 ( .A(n7183), .B(o[149]), .Z(n6586) );
  AND U9159 ( .A(n6587), .B(n6586), .Z(n6588) );
  NANDN U9160 ( .A(n6589), .B(n6588), .Z(n1907) );
  NANDN U9161 ( .A(n7182), .B(creg[148]), .Z(n6591) );
  NAND U9162 ( .A(n7183), .B(o[148]), .Z(n6590) );
  AND U9163 ( .A(n6591), .B(n6590), .Z(n6592) );
  NANDN U9164 ( .A(n6593), .B(n6592), .Z(n1908) );
  NANDN U9165 ( .A(n7182), .B(creg[147]), .Z(n6595) );
  NAND U9166 ( .A(n7183), .B(o[147]), .Z(n6594) );
  AND U9167 ( .A(n6595), .B(n6594), .Z(n6596) );
  NANDN U9168 ( .A(n6597), .B(n6596), .Z(n1909) );
  NANDN U9169 ( .A(n7182), .B(creg[146]), .Z(n6599) );
  NAND U9170 ( .A(n7183), .B(o[146]), .Z(n6598) );
  AND U9171 ( .A(n6599), .B(n6598), .Z(n6600) );
  NANDN U9172 ( .A(n6601), .B(n6600), .Z(n1910) );
  NANDN U9173 ( .A(n7182), .B(creg[145]), .Z(n6603) );
  NAND U9174 ( .A(n7183), .B(o[145]), .Z(n6602) );
  AND U9175 ( .A(n6603), .B(n6602), .Z(n6604) );
  NANDN U9176 ( .A(n6605), .B(n6604), .Z(n1911) );
  NANDN U9177 ( .A(n7182), .B(creg[144]), .Z(n6607) );
  NAND U9178 ( .A(n7183), .B(o[144]), .Z(n6606) );
  AND U9179 ( .A(n6607), .B(n6606), .Z(n6608) );
  NANDN U9180 ( .A(n6609), .B(n6608), .Z(n1912) );
  NANDN U9181 ( .A(n7182), .B(creg[143]), .Z(n6611) );
  NAND U9182 ( .A(n7183), .B(o[143]), .Z(n6610) );
  AND U9183 ( .A(n6611), .B(n6610), .Z(n6612) );
  NANDN U9184 ( .A(n6613), .B(n6612), .Z(n1913) );
  NANDN U9185 ( .A(n7182), .B(creg[142]), .Z(n6615) );
  NAND U9186 ( .A(n7183), .B(o[142]), .Z(n6614) );
  AND U9187 ( .A(n6615), .B(n6614), .Z(n6616) );
  NANDN U9188 ( .A(n6617), .B(n6616), .Z(n1914) );
  NANDN U9189 ( .A(n7182), .B(creg[141]), .Z(n6619) );
  NAND U9190 ( .A(n7183), .B(o[141]), .Z(n6618) );
  AND U9191 ( .A(n6619), .B(n6618), .Z(n6620) );
  NANDN U9192 ( .A(n6621), .B(n6620), .Z(n1915) );
  NANDN U9193 ( .A(n7182), .B(creg[140]), .Z(n6623) );
  NAND U9194 ( .A(n7183), .B(o[140]), .Z(n6622) );
  AND U9195 ( .A(n6623), .B(n6622), .Z(n6624) );
  NANDN U9196 ( .A(n6625), .B(n6624), .Z(n1916) );
  NANDN U9197 ( .A(n7182), .B(creg[139]), .Z(n6627) );
  NAND U9198 ( .A(n7183), .B(o[139]), .Z(n6626) );
  AND U9199 ( .A(n6627), .B(n6626), .Z(n6628) );
  NANDN U9200 ( .A(n6629), .B(n6628), .Z(n1917) );
  NANDN U9201 ( .A(n7182), .B(creg[138]), .Z(n6631) );
  NAND U9202 ( .A(n7183), .B(o[138]), .Z(n6630) );
  AND U9203 ( .A(n6631), .B(n6630), .Z(n6632) );
  NANDN U9204 ( .A(n6633), .B(n6632), .Z(n1918) );
  NANDN U9205 ( .A(n7182), .B(creg[137]), .Z(n6635) );
  NAND U9206 ( .A(n7183), .B(o[137]), .Z(n6634) );
  AND U9207 ( .A(n6635), .B(n6634), .Z(n6636) );
  NANDN U9208 ( .A(n6637), .B(n6636), .Z(n1919) );
  NANDN U9209 ( .A(n7182), .B(creg[136]), .Z(n6639) );
  NAND U9210 ( .A(n7183), .B(o[136]), .Z(n6638) );
  AND U9211 ( .A(n6639), .B(n6638), .Z(n6640) );
  NANDN U9212 ( .A(n6641), .B(n6640), .Z(n1920) );
  NANDN U9213 ( .A(n7182), .B(creg[135]), .Z(n6643) );
  NAND U9214 ( .A(n7183), .B(o[135]), .Z(n6642) );
  AND U9215 ( .A(n6643), .B(n6642), .Z(n6644) );
  NANDN U9216 ( .A(n6645), .B(n6644), .Z(n1921) );
  NANDN U9217 ( .A(n7182), .B(creg[134]), .Z(n6647) );
  NAND U9218 ( .A(n7183), .B(o[134]), .Z(n6646) );
  AND U9219 ( .A(n6647), .B(n6646), .Z(n6648) );
  NANDN U9220 ( .A(n6649), .B(n6648), .Z(n1922) );
  NANDN U9221 ( .A(n7182), .B(creg[133]), .Z(n6651) );
  NAND U9222 ( .A(n7183), .B(o[133]), .Z(n6650) );
  AND U9223 ( .A(n6651), .B(n6650), .Z(n6652) );
  NANDN U9224 ( .A(n6653), .B(n6652), .Z(n1923) );
  NANDN U9225 ( .A(n7182), .B(creg[132]), .Z(n6655) );
  NAND U9226 ( .A(n7183), .B(o[132]), .Z(n6654) );
  AND U9227 ( .A(n6655), .B(n6654), .Z(n6656) );
  NANDN U9228 ( .A(n6657), .B(n6656), .Z(n1924) );
  NANDN U9229 ( .A(n7182), .B(creg[131]), .Z(n6659) );
  NAND U9230 ( .A(n7183), .B(o[131]), .Z(n6658) );
  AND U9231 ( .A(n6659), .B(n6658), .Z(n6660) );
  NANDN U9232 ( .A(n6661), .B(n6660), .Z(n1925) );
  NANDN U9233 ( .A(n7182), .B(creg[130]), .Z(n6663) );
  NAND U9234 ( .A(n7183), .B(o[130]), .Z(n6662) );
  AND U9235 ( .A(n6663), .B(n6662), .Z(n6664) );
  NANDN U9236 ( .A(n6665), .B(n6664), .Z(n1926) );
  NANDN U9237 ( .A(n7182), .B(creg[129]), .Z(n6667) );
  NAND U9238 ( .A(n7183), .B(o[129]), .Z(n6666) );
  AND U9239 ( .A(n6667), .B(n6666), .Z(n6668) );
  NANDN U9240 ( .A(n6669), .B(n6668), .Z(n1927) );
  NANDN U9241 ( .A(n7182), .B(creg[128]), .Z(n6671) );
  NAND U9242 ( .A(n7183), .B(o[128]), .Z(n6670) );
  AND U9243 ( .A(n6671), .B(n6670), .Z(n6672) );
  NANDN U9244 ( .A(n6673), .B(n6672), .Z(n1928) );
  NANDN U9245 ( .A(n7182), .B(creg[127]), .Z(n6675) );
  NAND U9246 ( .A(n7183), .B(o[127]), .Z(n6674) );
  AND U9247 ( .A(n6675), .B(n6674), .Z(n6676) );
  NANDN U9248 ( .A(n6677), .B(n6676), .Z(n1929) );
  NANDN U9249 ( .A(n7182), .B(creg[126]), .Z(n6679) );
  NAND U9250 ( .A(n7183), .B(o[126]), .Z(n6678) );
  AND U9251 ( .A(n6679), .B(n6678), .Z(n6680) );
  NANDN U9252 ( .A(n6681), .B(n6680), .Z(n1930) );
  NANDN U9253 ( .A(n7182), .B(creg[125]), .Z(n6683) );
  NAND U9254 ( .A(n7183), .B(o[125]), .Z(n6682) );
  AND U9255 ( .A(n6683), .B(n6682), .Z(n6684) );
  NANDN U9256 ( .A(n6685), .B(n6684), .Z(n1931) );
  NANDN U9257 ( .A(n7182), .B(creg[124]), .Z(n6687) );
  NAND U9258 ( .A(n7183), .B(o[124]), .Z(n6686) );
  AND U9259 ( .A(n6687), .B(n6686), .Z(n6688) );
  NANDN U9260 ( .A(n6689), .B(n6688), .Z(n1932) );
  NANDN U9261 ( .A(n7182), .B(creg[123]), .Z(n6691) );
  NAND U9262 ( .A(n7183), .B(o[123]), .Z(n6690) );
  AND U9263 ( .A(n6691), .B(n6690), .Z(n6692) );
  NANDN U9264 ( .A(n6693), .B(n6692), .Z(n1933) );
  NANDN U9265 ( .A(n7182), .B(creg[122]), .Z(n6695) );
  NAND U9266 ( .A(n7183), .B(o[122]), .Z(n6694) );
  AND U9267 ( .A(n6695), .B(n6694), .Z(n6696) );
  NANDN U9268 ( .A(n6697), .B(n6696), .Z(n1934) );
  NANDN U9269 ( .A(n7182), .B(creg[121]), .Z(n6699) );
  NAND U9270 ( .A(n7183), .B(o[121]), .Z(n6698) );
  AND U9271 ( .A(n6699), .B(n6698), .Z(n6700) );
  NANDN U9272 ( .A(n6701), .B(n6700), .Z(n1935) );
  NANDN U9273 ( .A(n7182), .B(creg[120]), .Z(n6703) );
  NAND U9274 ( .A(n7183), .B(o[120]), .Z(n6702) );
  AND U9275 ( .A(n6703), .B(n6702), .Z(n6704) );
  NANDN U9276 ( .A(n6705), .B(n6704), .Z(n1936) );
  NANDN U9277 ( .A(n7182), .B(creg[119]), .Z(n6707) );
  NAND U9278 ( .A(n7183), .B(o[119]), .Z(n6706) );
  AND U9279 ( .A(n6707), .B(n6706), .Z(n6708) );
  NANDN U9280 ( .A(n6709), .B(n6708), .Z(n1937) );
  NANDN U9281 ( .A(n7182), .B(creg[118]), .Z(n6711) );
  NAND U9282 ( .A(n7183), .B(o[118]), .Z(n6710) );
  AND U9283 ( .A(n6711), .B(n6710), .Z(n6712) );
  NANDN U9284 ( .A(n6713), .B(n6712), .Z(n1938) );
  NANDN U9285 ( .A(n7182), .B(creg[117]), .Z(n6715) );
  NAND U9286 ( .A(n7183), .B(o[117]), .Z(n6714) );
  AND U9287 ( .A(n6715), .B(n6714), .Z(n6716) );
  NANDN U9288 ( .A(n6717), .B(n6716), .Z(n1939) );
  NANDN U9289 ( .A(n7182), .B(creg[116]), .Z(n6719) );
  NAND U9290 ( .A(n7183), .B(o[116]), .Z(n6718) );
  AND U9291 ( .A(n6719), .B(n6718), .Z(n6720) );
  NANDN U9292 ( .A(n6721), .B(n6720), .Z(n1940) );
  NANDN U9293 ( .A(n7182), .B(creg[115]), .Z(n6723) );
  NAND U9294 ( .A(n7183), .B(o[115]), .Z(n6722) );
  AND U9295 ( .A(n6723), .B(n6722), .Z(n6724) );
  NANDN U9296 ( .A(n6725), .B(n6724), .Z(n1941) );
  NANDN U9297 ( .A(n7182), .B(creg[114]), .Z(n6727) );
  NAND U9298 ( .A(n7183), .B(o[114]), .Z(n6726) );
  AND U9299 ( .A(n6727), .B(n6726), .Z(n6728) );
  NANDN U9300 ( .A(n6729), .B(n6728), .Z(n1942) );
  NANDN U9301 ( .A(n7182), .B(creg[113]), .Z(n6731) );
  NAND U9302 ( .A(n7183), .B(o[113]), .Z(n6730) );
  AND U9303 ( .A(n6731), .B(n6730), .Z(n6732) );
  NANDN U9304 ( .A(n6733), .B(n6732), .Z(n1943) );
  NANDN U9305 ( .A(n7182), .B(creg[112]), .Z(n6735) );
  NAND U9306 ( .A(n7183), .B(o[112]), .Z(n6734) );
  AND U9307 ( .A(n6735), .B(n6734), .Z(n6736) );
  NANDN U9308 ( .A(n6737), .B(n6736), .Z(n1944) );
  NANDN U9309 ( .A(n7182), .B(creg[111]), .Z(n6739) );
  NAND U9310 ( .A(n7183), .B(o[111]), .Z(n6738) );
  AND U9311 ( .A(n6739), .B(n6738), .Z(n6740) );
  NANDN U9312 ( .A(n6741), .B(n6740), .Z(n1945) );
  NANDN U9313 ( .A(n7182), .B(creg[110]), .Z(n6743) );
  NAND U9314 ( .A(n7183), .B(o[110]), .Z(n6742) );
  AND U9315 ( .A(n6743), .B(n6742), .Z(n6744) );
  NANDN U9316 ( .A(n6745), .B(n6744), .Z(n1946) );
  NANDN U9317 ( .A(n7182), .B(creg[109]), .Z(n6747) );
  NAND U9318 ( .A(n7183), .B(o[109]), .Z(n6746) );
  AND U9319 ( .A(n6747), .B(n6746), .Z(n6748) );
  NANDN U9320 ( .A(n6749), .B(n6748), .Z(n1947) );
  NANDN U9321 ( .A(n7182), .B(creg[108]), .Z(n6751) );
  NAND U9322 ( .A(n7183), .B(o[108]), .Z(n6750) );
  AND U9323 ( .A(n6751), .B(n6750), .Z(n6752) );
  NANDN U9324 ( .A(n6753), .B(n6752), .Z(n1948) );
  NANDN U9325 ( .A(n7182), .B(creg[107]), .Z(n6755) );
  NAND U9326 ( .A(n7183), .B(o[107]), .Z(n6754) );
  AND U9327 ( .A(n6755), .B(n6754), .Z(n6756) );
  NANDN U9328 ( .A(n6757), .B(n6756), .Z(n1949) );
  NANDN U9329 ( .A(n7182), .B(creg[106]), .Z(n6759) );
  NAND U9330 ( .A(n7183), .B(o[106]), .Z(n6758) );
  AND U9331 ( .A(n6759), .B(n6758), .Z(n6760) );
  NANDN U9332 ( .A(n6761), .B(n6760), .Z(n1950) );
  NANDN U9333 ( .A(n7182), .B(creg[105]), .Z(n6763) );
  NAND U9334 ( .A(n7183), .B(o[105]), .Z(n6762) );
  AND U9335 ( .A(n6763), .B(n6762), .Z(n6764) );
  NANDN U9336 ( .A(n6765), .B(n6764), .Z(n1951) );
  NANDN U9337 ( .A(n7182), .B(creg[104]), .Z(n6767) );
  NAND U9338 ( .A(n7183), .B(o[104]), .Z(n6766) );
  AND U9339 ( .A(n6767), .B(n6766), .Z(n6768) );
  NANDN U9340 ( .A(n6769), .B(n6768), .Z(n1952) );
  NANDN U9341 ( .A(n7182), .B(creg[103]), .Z(n6771) );
  NAND U9342 ( .A(n7183), .B(o[103]), .Z(n6770) );
  AND U9343 ( .A(n6771), .B(n6770), .Z(n6772) );
  NANDN U9344 ( .A(n6773), .B(n6772), .Z(n1953) );
  NANDN U9345 ( .A(n7182), .B(creg[102]), .Z(n6775) );
  NAND U9346 ( .A(n7183), .B(o[102]), .Z(n6774) );
  AND U9347 ( .A(n6775), .B(n6774), .Z(n6776) );
  NANDN U9348 ( .A(n6777), .B(n6776), .Z(n1954) );
  NANDN U9349 ( .A(n7182), .B(creg[101]), .Z(n6779) );
  NAND U9350 ( .A(n7183), .B(o[101]), .Z(n6778) );
  AND U9351 ( .A(n6779), .B(n6778), .Z(n6780) );
  NANDN U9352 ( .A(n6781), .B(n6780), .Z(n1955) );
  NANDN U9353 ( .A(n7182), .B(creg[100]), .Z(n6783) );
  NAND U9354 ( .A(n7183), .B(o[100]), .Z(n6782) );
  AND U9355 ( .A(n6783), .B(n6782), .Z(n6784) );
  NANDN U9356 ( .A(n6785), .B(n6784), .Z(n1956) );
  NANDN U9357 ( .A(n7182), .B(creg[99]), .Z(n6787) );
  NAND U9358 ( .A(n7183), .B(o[99]), .Z(n6786) );
  AND U9359 ( .A(n6787), .B(n6786), .Z(n6788) );
  NANDN U9360 ( .A(n6789), .B(n6788), .Z(n1957) );
  NANDN U9361 ( .A(n7182), .B(creg[98]), .Z(n6791) );
  NAND U9362 ( .A(n7183), .B(o[98]), .Z(n6790) );
  AND U9363 ( .A(n6791), .B(n6790), .Z(n6792) );
  NANDN U9364 ( .A(n6793), .B(n6792), .Z(n1958) );
  NANDN U9365 ( .A(n7182), .B(creg[97]), .Z(n6795) );
  NAND U9366 ( .A(n7183), .B(o[97]), .Z(n6794) );
  AND U9367 ( .A(n6795), .B(n6794), .Z(n6796) );
  NANDN U9368 ( .A(n6797), .B(n6796), .Z(n1959) );
  NANDN U9369 ( .A(n7182), .B(creg[96]), .Z(n6799) );
  NAND U9370 ( .A(n7183), .B(o[96]), .Z(n6798) );
  AND U9371 ( .A(n6799), .B(n6798), .Z(n6800) );
  NANDN U9372 ( .A(n6801), .B(n6800), .Z(n1960) );
  NANDN U9373 ( .A(n7182), .B(creg[95]), .Z(n6803) );
  NAND U9374 ( .A(n7183), .B(o[95]), .Z(n6802) );
  AND U9375 ( .A(n6803), .B(n6802), .Z(n6804) );
  NANDN U9376 ( .A(n6805), .B(n6804), .Z(n1961) );
  NANDN U9377 ( .A(n7182), .B(creg[94]), .Z(n6807) );
  NAND U9378 ( .A(n7183), .B(o[94]), .Z(n6806) );
  AND U9379 ( .A(n6807), .B(n6806), .Z(n6808) );
  NANDN U9380 ( .A(n6809), .B(n6808), .Z(n1962) );
  NANDN U9381 ( .A(n7182), .B(creg[93]), .Z(n6811) );
  NAND U9382 ( .A(n7183), .B(o[93]), .Z(n6810) );
  AND U9383 ( .A(n6811), .B(n6810), .Z(n6812) );
  NANDN U9384 ( .A(n6813), .B(n6812), .Z(n1963) );
  NANDN U9385 ( .A(n7182), .B(creg[92]), .Z(n6815) );
  NAND U9386 ( .A(n7183), .B(o[92]), .Z(n6814) );
  AND U9387 ( .A(n6815), .B(n6814), .Z(n6816) );
  NANDN U9388 ( .A(n6817), .B(n6816), .Z(n1964) );
  NANDN U9389 ( .A(n7182), .B(creg[91]), .Z(n6819) );
  NAND U9390 ( .A(n7183), .B(o[91]), .Z(n6818) );
  AND U9391 ( .A(n6819), .B(n6818), .Z(n6820) );
  NANDN U9392 ( .A(n6821), .B(n6820), .Z(n1965) );
  NANDN U9393 ( .A(n7182), .B(creg[90]), .Z(n6823) );
  NAND U9394 ( .A(n7183), .B(o[90]), .Z(n6822) );
  AND U9395 ( .A(n6823), .B(n6822), .Z(n6824) );
  NANDN U9396 ( .A(n6825), .B(n6824), .Z(n1966) );
  NANDN U9397 ( .A(n7182), .B(creg[89]), .Z(n6827) );
  NAND U9398 ( .A(n7183), .B(o[89]), .Z(n6826) );
  AND U9399 ( .A(n6827), .B(n6826), .Z(n6828) );
  NANDN U9400 ( .A(n6829), .B(n6828), .Z(n1967) );
  NANDN U9401 ( .A(n7182), .B(creg[88]), .Z(n6831) );
  NAND U9402 ( .A(n7183), .B(o[88]), .Z(n6830) );
  AND U9403 ( .A(n6831), .B(n6830), .Z(n6832) );
  NANDN U9404 ( .A(n6833), .B(n6832), .Z(n1968) );
  NANDN U9405 ( .A(n7182), .B(creg[87]), .Z(n6835) );
  NAND U9406 ( .A(n7183), .B(o[87]), .Z(n6834) );
  AND U9407 ( .A(n6835), .B(n6834), .Z(n6836) );
  NANDN U9408 ( .A(n6837), .B(n6836), .Z(n1969) );
  NANDN U9409 ( .A(n7182), .B(creg[86]), .Z(n6839) );
  NAND U9410 ( .A(n7183), .B(o[86]), .Z(n6838) );
  AND U9411 ( .A(n6839), .B(n6838), .Z(n6840) );
  NANDN U9412 ( .A(n6841), .B(n6840), .Z(n1970) );
  NANDN U9413 ( .A(n7182), .B(creg[85]), .Z(n6843) );
  NAND U9414 ( .A(n7183), .B(o[85]), .Z(n6842) );
  AND U9415 ( .A(n6843), .B(n6842), .Z(n6844) );
  NANDN U9416 ( .A(n6845), .B(n6844), .Z(n1971) );
  NANDN U9417 ( .A(n7182), .B(creg[84]), .Z(n6847) );
  NAND U9418 ( .A(n7183), .B(o[84]), .Z(n6846) );
  AND U9419 ( .A(n6847), .B(n6846), .Z(n6848) );
  NANDN U9420 ( .A(n6849), .B(n6848), .Z(n1972) );
  NANDN U9421 ( .A(n7182), .B(creg[83]), .Z(n6851) );
  NAND U9422 ( .A(n7183), .B(o[83]), .Z(n6850) );
  AND U9423 ( .A(n6851), .B(n6850), .Z(n6852) );
  NANDN U9424 ( .A(n6853), .B(n6852), .Z(n1973) );
  NANDN U9425 ( .A(n7182), .B(creg[82]), .Z(n6855) );
  NAND U9426 ( .A(n7183), .B(o[82]), .Z(n6854) );
  AND U9427 ( .A(n6855), .B(n6854), .Z(n6856) );
  NANDN U9428 ( .A(n6857), .B(n6856), .Z(n1974) );
  NANDN U9429 ( .A(n7182), .B(creg[81]), .Z(n6859) );
  NAND U9430 ( .A(n7183), .B(o[81]), .Z(n6858) );
  AND U9431 ( .A(n6859), .B(n6858), .Z(n6860) );
  NANDN U9432 ( .A(n6861), .B(n6860), .Z(n1975) );
  NANDN U9433 ( .A(n7182), .B(creg[80]), .Z(n6863) );
  NAND U9434 ( .A(n7183), .B(o[80]), .Z(n6862) );
  AND U9435 ( .A(n6863), .B(n6862), .Z(n6864) );
  NANDN U9436 ( .A(n6865), .B(n6864), .Z(n1976) );
  NANDN U9437 ( .A(n7182), .B(creg[79]), .Z(n6867) );
  NAND U9438 ( .A(n7183), .B(o[79]), .Z(n6866) );
  AND U9439 ( .A(n6867), .B(n6866), .Z(n6868) );
  NANDN U9440 ( .A(n6869), .B(n6868), .Z(n1977) );
  NANDN U9441 ( .A(n7182), .B(creg[78]), .Z(n6871) );
  NAND U9442 ( .A(n7183), .B(o[78]), .Z(n6870) );
  AND U9443 ( .A(n6871), .B(n6870), .Z(n6872) );
  NANDN U9444 ( .A(n6873), .B(n6872), .Z(n1978) );
  NANDN U9445 ( .A(n7182), .B(creg[77]), .Z(n6875) );
  NAND U9446 ( .A(n7183), .B(o[77]), .Z(n6874) );
  AND U9447 ( .A(n6875), .B(n6874), .Z(n6876) );
  NANDN U9448 ( .A(n6877), .B(n6876), .Z(n1979) );
  NANDN U9449 ( .A(n7182), .B(creg[76]), .Z(n6879) );
  NAND U9450 ( .A(n7183), .B(o[76]), .Z(n6878) );
  AND U9451 ( .A(n6879), .B(n6878), .Z(n6880) );
  NANDN U9452 ( .A(n6881), .B(n6880), .Z(n1980) );
  NANDN U9453 ( .A(n7182), .B(creg[75]), .Z(n6883) );
  NAND U9454 ( .A(n7183), .B(o[75]), .Z(n6882) );
  AND U9455 ( .A(n6883), .B(n6882), .Z(n6884) );
  NANDN U9456 ( .A(n6885), .B(n6884), .Z(n1981) );
  NANDN U9457 ( .A(n7182), .B(creg[74]), .Z(n6887) );
  NAND U9458 ( .A(n7183), .B(o[74]), .Z(n6886) );
  AND U9459 ( .A(n6887), .B(n6886), .Z(n6888) );
  NANDN U9460 ( .A(n6889), .B(n6888), .Z(n1982) );
  NANDN U9461 ( .A(n7182), .B(creg[73]), .Z(n6891) );
  NAND U9462 ( .A(n7183), .B(o[73]), .Z(n6890) );
  AND U9463 ( .A(n6891), .B(n6890), .Z(n6892) );
  NANDN U9464 ( .A(n6893), .B(n6892), .Z(n1983) );
  NANDN U9465 ( .A(n7182), .B(creg[72]), .Z(n6895) );
  NAND U9466 ( .A(n7183), .B(o[72]), .Z(n6894) );
  AND U9467 ( .A(n6895), .B(n6894), .Z(n6896) );
  NANDN U9468 ( .A(n6897), .B(n6896), .Z(n1984) );
  NANDN U9469 ( .A(n7182), .B(creg[71]), .Z(n6899) );
  NAND U9470 ( .A(n7183), .B(o[71]), .Z(n6898) );
  AND U9471 ( .A(n6899), .B(n6898), .Z(n6900) );
  NANDN U9472 ( .A(n6901), .B(n6900), .Z(n1985) );
  NANDN U9473 ( .A(n7182), .B(creg[70]), .Z(n6903) );
  NAND U9474 ( .A(n7183), .B(o[70]), .Z(n6902) );
  AND U9475 ( .A(n6903), .B(n6902), .Z(n6904) );
  NANDN U9476 ( .A(n6905), .B(n6904), .Z(n1986) );
  NANDN U9477 ( .A(n7182), .B(creg[69]), .Z(n6907) );
  NAND U9478 ( .A(n7183), .B(o[69]), .Z(n6906) );
  AND U9479 ( .A(n6907), .B(n6906), .Z(n6908) );
  NANDN U9480 ( .A(n6909), .B(n6908), .Z(n1987) );
  NANDN U9481 ( .A(n7182), .B(creg[68]), .Z(n6911) );
  NAND U9482 ( .A(n7183), .B(o[68]), .Z(n6910) );
  AND U9483 ( .A(n6911), .B(n6910), .Z(n6912) );
  NANDN U9484 ( .A(n6913), .B(n6912), .Z(n1988) );
  NANDN U9485 ( .A(n7182), .B(creg[67]), .Z(n6915) );
  NAND U9486 ( .A(n7183), .B(o[67]), .Z(n6914) );
  AND U9487 ( .A(n6915), .B(n6914), .Z(n6916) );
  NANDN U9488 ( .A(n6917), .B(n6916), .Z(n1989) );
  NANDN U9489 ( .A(n7182), .B(creg[66]), .Z(n6919) );
  NAND U9490 ( .A(n7183), .B(o[66]), .Z(n6918) );
  AND U9491 ( .A(n6919), .B(n6918), .Z(n6920) );
  NANDN U9492 ( .A(n6921), .B(n6920), .Z(n1990) );
  NANDN U9493 ( .A(n7182), .B(creg[65]), .Z(n6923) );
  NAND U9494 ( .A(n7183), .B(o[65]), .Z(n6922) );
  AND U9495 ( .A(n6923), .B(n6922), .Z(n6924) );
  NANDN U9496 ( .A(n6925), .B(n6924), .Z(n1991) );
  NANDN U9497 ( .A(n7182), .B(creg[64]), .Z(n6927) );
  NAND U9498 ( .A(n7183), .B(o[64]), .Z(n6926) );
  AND U9499 ( .A(n6927), .B(n6926), .Z(n6928) );
  NANDN U9500 ( .A(n6929), .B(n6928), .Z(n1992) );
  NANDN U9501 ( .A(n7182), .B(creg[63]), .Z(n6931) );
  NAND U9502 ( .A(n7183), .B(o[63]), .Z(n6930) );
  AND U9503 ( .A(n6931), .B(n6930), .Z(n6932) );
  NANDN U9504 ( .A(n6933), .B(n6932), .Z(n1993) );
  NANDN U9505 ( .A(n7182), .B(creg[62]), .Z(n6935) );
  NAND U9506 ( .A(n7183), .B(o[62]), .Z(n6934) );
  AND U9507 ( .A(n6935), .B(n6934), .Z(n6936) );
  NANDN U9508 ( .A(n6937), .B(n6936), .Z(n1994) );
  NANDN U9509 ( .A(n7182), .B(creg[61]), .Z(n6939) );
  NAND U9510 ( .A(n7183), .B(o[61]), .Z(n6938) );
  AND U9511 ( .A(n6939), .B(n6938), .Z(n6940) );
  NANDN U9512 ( .A(n6941), .B(n6940), .Z(n1995) );
  NANDN U9513 ( .A(n7182), .B(creg[60]), .Z(n6943) );
  NAND U9514 ( .A(n7183), .B(o[60]), .Z(n6942) );
  AND U9515 ( .A(n6943), .B(n6942), .Z(n6944) );
  NANDN U9516 ( .A(n6945), .B(n6944), .Z(n1996) );
  NANDN U9517 ( .A(n7182), .B(creg[59]), .Z(n6947) );
  NAND U9518 ( .A(n7183), .B(o[59]), .Z(n6946) );
  AND U9519 ( .A(n6947), .B(n6946), .Z(n6948) );
  NANDN U9520 ( .A(n6949), .B(n6948), .Z(n1997) );
  NANDN U9521 ( .A(n7182), .B(creg[58]), .Z(n6951) );
  NAND U9522 ( .A(n7183), .B(o[58]), .Z(n6950) );
  AND U9523 ( .A(n6951), .B(n6950), .Z(n6952) );
  NANDN U9524 ( .A(n6953), .B(n6952), .Z(n1998) );
  NANDN U9525 ( .A(n7182), .B(creg[57]), .Z(n6955) );
  NAND U9526 ( .A(n7183), .B(o[57]), .Z(n6954) );
  AND U9527 ( .A(n6955), .B(n6954), .Z(n6956) );
  NANDN U9528 ( .A(n6957), .B(n6956), .Z(n1999) );
  NANDN U9529 ( .A(n7182), .B(creg[56]), .Z(n6959) );
  NAND U9530 ( .A(n7183), .B(o[56]), .Z(n6958) );
  AND U9531 ( .A(n6959), .B(n6958), .Z(n6960) );
  NANDN U9532 ( .A(n6961), .B(n6960), .Z(n2000) );
  NANDN U9533 ( .A(n7182), .B(creg[55]), .Z(n6963) );
  NAND U9534 ( .A(n7183), .B(o[55]), .Z(n6962) );
  AND U9535 ( .A(n6963), .B(n6962), .Z(n6964) );
  NANDN U9536 ( .A(n6965), .B(n6964), .Z(n2001) );
  NANDN U9537 ( .A(n7182), .B(creg[54]), .Z(n6967) );
  NAND U9538 ( .A(n7183), .B(o[54]), .Z(n6966) );
  AND U9539 ( .A(n6967), .B(n6966), .Z(n6968) );
  NANDN U9540 ( .A(n6969), .B(n6968), .Z(n2002) );
  NANDN U9541 ( .A(n7182), .B(creg[53]), .Z(n6971) );
  NAND U9542 ( .A(n7183), .B(o[53]), .Z(n6970) );
  AND U9543 ( .A(n6971), .B(n6970), .Z(n6972) );
  NANDN U9544 ( .A(n6973), .B(n6972), .Z(n2003) );
  NANDN U9545 ( .A(n7182), .B(creg[52]), .Z(n6975) );
  NAND U9546 ( .A(n7183), .B(o[52]), .Z(n6974) );
  AND U9547 ( .A(n6975), .B(n6974), .Z(n6976) );
  NANDN U9548 ( .A(n6977), .B(n6976), .Z(n2004) );
  NANDN U9549 ( .A(n7182), .B(creg[51]), .Z(n6979) );
  NAND U9550 ( .A(n7183), .B(o[51]), .Z(n6978) );
  AND U9551 ( .A(n6979), .B(n6978), .Z(n6980) );
  NANDN U9552 ( .A(n6981), .B(n6980), .Z(n2005) );
  NANDN U9553 ( .A(n7182), .B(creg[50]), .Z(n6983) );
  NAND U9554 ( .A(n7183), .B(o[50]), .Z(n6982) );
  AND U9555 ( .A(n6983), .B(n6982), .Z(n6984) );
  NANDN U9556 ( .A(n6985), .B(n6984), .Z(n2006) );
  NANDN U9557 ( .A(n7182), .B(creg[49]), .Z(n6987) );
  NAND U9558 ( .A(n7183), .B(o[49]), .Z(n6986) );
  AND U9559 ( .A(n6987), .B(n6986), .Z(n6988) );
  NANDN U9560 ( .A(n6989), .B(n6988), .Z(n2007) );
  NANDN U9561 ( .A(n7182), .B(creg[48]), .Z(n6991) );
  NAND U9562 ( .A(n7183), .B(o[48]), .Z(n6990) );
  AND U9563 ( .A(n6991), .B(n6990), .Z(n6992) );
  NANDN U9564 ( .A(n6993), .B(n6992), .Z(n2008) );
  NANDN U9565 ( .A(n7182), .B(creg[47]), .Z(n6995) );
  NAND U9566 ( .A(n7183), .B(o[47]), .Z(n6994) );
  AND U9567 ( .A(n6995), .B(n6994), .Z(n6996) );
  NANDN U9568 ( .A(n6997), .B(n6996), .Z(n2009) );
  NANDN U9569 ( .A(n7182), .B(creg[46]), .Z(n6999) );
  NAND U9570 ( .A(n7183), .B(o[46]), .Z(n6998) );
  AND U9571 ( .A(n6999), .B(n6998), .Z(n7000) );
  NANDN U9572 ( .A(n7001), .B(n7000), .Z(n2010) );
  NANDN U9573 ( .A(n7182), .B(creg[45]), .Z(n7003) );
  NAND U9574 ( .A(n7183), .B(o[45]), .Z(n7002) );
  AND U9575 ( .A(n7003), .B(n7002), .Z(n7004) );
  NANDN U9576 ( .A(n7005), .B(n7004), .Z(n2011) );
  NANDN U9577 ( .A(n7182), .B(creg[44]), .Z(n7007) );
  NAND U9578 ( .A(n7183), .B(o[44]), .Z(n7006) );
  AND U9579 ( .A(n7007), .B(n7006), .Z(n7008) );
  NANDN U9580 ( .A(n7009), .B(n7008), .Z(n2012) );
  NANDN U9581 ( .A(n7182), .B(creg[43]), .Z(n7011) );
  NAND U9582 ( .A(n7183), .B(o[43]), .Z(n7010) );
  AND U9583 ( .A(n7011), .B(n7010), .Z(n7012) );
  NANDN U9584 ( .A(n7013), .B(n7012), .Z(n2013) );
  NANDN U9585 ( .A(n7182), .B(creg[42]), .Z(n7015) );
  NAND U9586 ( .A(n7183), .B(o[42]), .Z(n7014) );
  AND U9587 ( .A(n7015), .B(n7014), .Z(n7016) );
  NANDN U9588 ( .A(n7017), .B(n7016), .Z(n2014) );
  NANDN U9589 ( .A(n7182), .B(creg[41]), .Z(n7019) );
  NAND U9590 ( .A(n7183), .B(o[41]), .Z(n7018) );
  AND U9591 ( .A(n7019), .B(n7018), .Z(n7020) );
  NANDN U9592 ( .A(n7021), .B(n7020), .Z(n2015) );
  NANDN U9593 ( .A(n7182), .B(creg[40]), .Z(n7023) );
  NAND U9594 ( .A(n7183), .B(o[40]), .Z(n7022) );
  AND U9595 ( .A(n7023), .B(n7022), .Z(n7024) );
  NANDN U9596 ( .A(n7025), .B(n7024), .Z(n2016) );
  NANDN U9597 ( .A(n7182), .B(creg[39]), .Z(n7027) );
  NAND U9598 ( .A(n7183), .B(o[39]), .Z(n7026) );
  AND U9599 ( .A(n7027), .B(n7026), .Z(n7028) );
  NANDN U9600 ( .A(n7029), .B(n7028), .Z(n2017) );
  NANDN U9601 ( .A(n7182), .B(creg[38]), .Z(n7031) );
  NAND U9602 ( .A(n7183), .B(o[38]), .Z(n7030) );
  AND U9603 ( .A(n7031), .B(n7030), .Z(n7032) );
  NANDN U9604 ( .A(n7033), .B(n7032), .Z(n2018) );
  NANDN U9605 ( .A(n7182), .B(creg[37]), .Z(n7035) );
  NAND U9606 ( .A(n7183), .B(o[37]), .Z(n7034) );
  AND U9607 ( .A(n7035), .B(n7034), .Z(n7036) );
  NANDN U9608 ( .A(n7037), .B(n7036), .Z(n2019) );
  NANDN U9609 ( .A(n7182), .B(creg[36]), .Z(n7039) );
  NAND U9610 ( .A(n7183), .B(o[36]), .Z(n7038) );
  AND U9611 ( .A(n7039), .B(n7038), .Z(n7040) );
  NANDN U9612 ( .A(n7041), .B(n7040), .Z(n2020) );
  NANDN U9613 ( .A(n7182), .B(creg[35]), .Z(n7043) );
  NAND U9614 ( .A(n7183), .B(o[35]), .Z(n7042) );
  AND U9615 ( .A(n7043), .B(n7042), .Z(n7044) );
  NANDN U9616 ( .A(n7045), .B(n7044), .Z(n2021) );
  NANDN U9617 ( .A(n7182), .B(creg[34]), .Z(n7047) );
  NAND U9618 ( .A(n7183), .B(o[34]), .Z(n7046) );
  AND U9619 ( .A(n7047), .B(n7046), .Z(n7048) );
  NANDN U9620 ( .A(n7049), .B(n7048), .Z(n2022) );
  NANDN U9621 ( .A(n7182), .B(creg[33]), .Z(n7051) );
  NAND U9622 ( .A(n7183), .B(o[33]), .Z(n7050) );
  AND U9623 ( .A(n7051), .B(n7050), .Z(n7052) );
  NANDN U9624 ( .A(n7053), .B(n7052), .Z(n2023) );
  NANDN U9625 ( .A(n7182), .B(creg[32]), .Z(n7055) );
  NAND U9626 ( .A(n7183), .B(o[32]), .Z(n7054) );
  AND U9627 ( .A(n7055), .B(n7054), .Z(n7056) );
  NANDN U9628 ( .A(n7057), .B(n7056), .Z(n2024) );
  NANDN U9629 ( .A(n7182), .B(creg[31]), .Z(n7059) );
  NAND U9630 ( .A(n7183), .B(o[31]), .Z(n7058) );
  AND U9631 ( .A(n7059), .B(n7058), .Z(n7060) );
  NANDN U9632 ( .A(n7061), .B(n7060), .Z(n2025) );
  NANDN U9633 ( .A(n7182), .B(creg[30]), .Z(n7063) );
  NAND U9634 ( .A(n7183), .B(o[30]), .Z(n7062) );
  AND U9635 ( .A(n7063), .B(n7062), .Z(n7064) );
  NANDN U9636 ( .A(n7065), .B(n7064), .Z(n2026) );
  NANDN U9637 ( .A(n7182), .B(creg[29]), .Z(n7067) );
  NAND U9638 ( .A(n7183), .B(o[29]), .Z(n7066) );
  AND U9639 ( .A(n7067), .B(n7066), .Z(n7068) );
  NANDN U9640 ( .A(n7069), .B(n7068), .Z(n2027) );
  NANDN U9641 ( .A(n7182), .B(creg[28]), .Z(n7071) );
  NAND U9642 ( .A(n7183), .B(o[28]), .Z(n7070) );
  AND U9643 ( .A(n7071), .B(n7070), .Z(n7072) );
  NANDN U9644 ( .A(n7073), .B(n7072), .Z(n2028) );
  NANDN U9645 ( .A(n7182), .B(creg[27]), .Z(n7075) );
  NAND U9646 ( .A(n7183), .B(o[27]), .Z(n7074) );
  AND U9647 ( .A(n7075), .B(n7074), .Z(n7076) );
  NANDN U9648 ( .A(n7077), .B(n7076), .Z(n2029) );
  NANDN U9649 ( .A(n7182), .B(creg[26]), .Z(n7079) );
  NAND U9650 ( .A(n7183), .B(o[26]), .Z(n7078) );
  AND U9651 ( .A(n7079), .B(n7078), .Z(n7080) );
  NANDN U9652 ( .A(n7081), .B(n7080), .Z(n2030) );
  NANDN U9653 ( .A(n7182), .B(creg[25]), .Z(n7083) );
  NAND U9654 ( .A(n7183), .B(o[25]), .Z(n7082) );
  AND U9655 ( .A(n7083), .B(n7082), .Z(n7084) );
  NANDN U9656 ( .A(n7085), .B(n7084), .Z(n2031) );
  NANDN U9657 ( .A(n7182), .B(creg[24]), .Z(n7087) );
  NAND U9658 ( .A(n7183), .B(o[24]), .Z(n7086) );
  AND U9659 ( .A(n7087), .B(n7086), .Z(n7088) );
  NANDN U9660 ( .A(n7089), .B(n7088), .Z(n2032) );
  NANDN U9661 ( .A(n7182), .B(creg[23]), .Z(n7091) );
  NAND U9662 ( .A(n7183), .B(o[23]), .Z(n7090) );
  AND U9663 ( .A(n7091), .B(n7090), .Z(n7092) );
  NANDN U9664 ( .A(n7093), .B(n7092), .Z(n2033) );
  NANDN U9665 ( .A(n7182), .B(creg[22]), .Z(n7095) );
  NAND U9666 ( .A(n7183), .B(o[22]), .Z(n7094) );
  AND U9667 ( .A(n7095), .B(n7094), .Z(n7096) );
  NANDN U9668 ( .A(n7097), .B(n7096), .Z(n2034) );
  NANDN U9669 ( .A(n7182), .B(creg[21]), .Z(n7099) );
  NAND U9670 ( .A(n7183), .B(o[21]), .Z(n7098) );
  AND U9671 ( .A(n7099), .B(n7098), .Z(n7100) );
  NANDN U9672 ( .A(n7101), .B(n7100), .Z(n2035) );
  NANDN U9673 ( .A(n7182), .B(creg[20]), .Z(n7103) );
  NAND U9674 ( .A(n7183), .B(o[20]), .Z(n7102) );
  AND U9675 ( .A(n7103), .B(n7102), .Z(n7104) );
  NANDN U9676 ( .A(n7105), .B(n7104), .Z(n2036) );
  NANDN U9677 ( .A(n7182), .B(creg[19]), .Z(n7107) );
  NAND U9678 ( .A(n7183), .B(o[19]), .Z(n7106) );
  AND U9679 ( .A(n7107), .B(n7106), .Z(n7108) );
  NANDN U9680 ( .A(n7109), .B(n7108), .Z(n2037) );
  NANDN U9681 ( .A(n7182), .B(creg[18]), .Z(n7111) );
  NAND U9682 ( .A(n7183), .B(o[18]), .Z(n7110) );
  AND U9683 ( .A(n7111), .B(n7110), .Z(n7112) );
  NANDN U9684 ( .A(n7113), .B(n7112), .Z(n2038) );
  NANDN U9685 ( .A(n7182), .B(creg[17]), .Z(n7115) );
  NAND U9686 ( .A(n7183), .B(o[17]), .Z(n7114) );
  AND U9687 ( .A(n7115), .B(n7114), .Z(n7116) );
  NANDN U9688 ( .A(n7117), .B(n7116), .Z(n2039) );
  NANDN U9689 ( .A(n7182), .B(creg[16]), .Z(n7119) );
  NAND U9690 ( .A(n7183), .B(o[16]), .Z(n7118) );
  AND U9691 ( .A(n7119), .B(n7118), .Z(n7120) );
  NANDN U9692 ( .A(n7121), .B(n7120), .Z(n2040) );
  NANDN U9693 ( .A(n7182), .B(creg[15]), .Z(n7123) );
  NAND U9694 ( .A(n7183), .B(o[15]), .Z(n7122) );
  AND U9695 ( .A(n7123), .B(n7122), .Z(n7124) );
  NANDN U9696 ( .A(n7125), .B(n7124), .Z(n2041) );
  NANDN U9697 ( .A(n7182), .B(creg[14]), .Z(n7127) );
  NAND U9698 ( .A(n7183), .B(o[14]), .Z(n7126) );
  AND U9699 ( .A(n7127), .B(n7126), .Z(n7128) );
  NANDN U9700 ( .A(n7129), .B(n7128), .Z(n2042) );
  NANDN U9701 ( .A(n7182), .B(creg[13]), .Z(n7131) );
  NAND U9702 ( .A(n7183), .B(o[13]), .Z(n7130) );
  AND U9703 ( .A(n7131), .B(n7130), .Z(n7132) );
  NANDN U9704 ( .A(n7133), .B(n7132), .Z(n2043) );
  NANDN U9705 ( .A(n7182), .B(creg[12]), .Z(n7135) );
  NAND U9706 ( .A(n7183), .B(o[12]), .Z(n7134) );
  AND U9707 ( .A(n7135), .B(n7134), .Z(n7136) );
  NANDN U9708 ( .A(n7137), .B(n7136), .Z(n2044) );
  NANDN U9709 ( .A(n7182), .B(creg[11]), .Z(n7139) );
  NAND U9710 ( .A(n7183), .B(o[11]), .Z(n7138) );
  AND U9711 ( .A(n7139), .B(n7138), .Z(n7140) );
  NANDN U9712 ( .A(n7141), .B(n7140), .Z(n2045) );
  NANDN U9713 ( .A(n7182), .B(creg[10]), .Z(n7143) );
  NAND U9714 ( .A(n7183), .B(o[10]), .Z(n7142) );
  AND U9715 ( .A(n7143), .B(n7142), .Z(n7144) );
  NANDN U9716 ( .A(n7145), .B(n7144), .Z(n2046) );
  NANDN U9717 ( .A(n7182), .B(creg[9]), .Z(n7147) );
  NAND U9718 ( .A(n7183), .B(o[9]), .Z(n7146) );
  AND U9719 ( .A(n7147), .B(n7146), .Z(n7148) );
  NANDN U9720 ( .A(n7149), .B(n7148), .Z(n2047) );
  NANDN U9721 ( .A(n7182), .B(creg[8]), .Z(n7151) );
  NAND U9722 ( .A(n7183), .B(o[8]), .Z(n7150) );
  AND U9723 ( .A(n7151), .B(n7150), .Z(n7152) );
  NANDN U9724 ( .A(n7153), .B(n7152), .Z(n2048) );
  NANDN U9725 ( .A(n7182), .B(creg[7]), .Z(n7155) );
  NAND U9726 ( .A(n7183), .B(o[7]), .Z(n7154) );
  AND U9727 ( .A(n7155), .B(n7154), .Z(n7156) );
  NANDN U9728 ( .A(n7157), .B(n7156), .Z(n2049) );
  NANDN U9729 ( .A(n7182), .B(creg[6]), .Z(n7159) );
  NAND U9730 ( .A(n7183), .B(o[6]), .Z(n7158) );
  AND U9731 ( .A(n7159), .B(n7158), .Z(n7160) );
  NANDN U9732 ( .A(n7161), .B(n7160), .Z(n2050) );
  NANDN U9733 ( .A(n7182), .B(creg[5]), .Z(n7163) );
  NAND U9734 ( .A(n7183), .B(o[5]), .Z(n7162) );
  AND U9735 ( .A(n7163), .B(n7162), .Z(n7164) );
  NANDN U9736 ( .A(n7165), .B(n7164), .Z(n2051) );
  NANDN U9737 ( .A(n7182), .B(creg[4]), .Z(n7167) );
  NAND U9738 ( .A(n7183), .B(o[4]), .Z(n7166) );
  AND U9739 ( .A(n7167), .B(n7166), .Z(n7168) );
  NANDN U9740 ( .A(n7169), .B(n7168), .Z(n2052) );
  NANDN U9741 ( .A(n7182), .B(creg[3]), .Z(n7171) );
  NAND U9742 ( .A(n7183), .B(o[3]), .Z(n7170) );
  AND U9743 ( .A(n7171), .B(n7170), .Z(n7172) );
  NANDN U9744 ( .A(n7173), .B(n7172), .Z(n2053) );
  NANDN U9745 ( .A(n7182), .B(creg[2]), .Z(n7175) );
  NAND U9746 ( .A(n7183), .B(o[2]), .Z(n7174) );
  AND U9747 ( .A(n7175), .B(n7174), .Z(n7176) );
  NANDN U9748 ( .A(n7177), .B(n7176), .Z(n2054) );
  NANDN U9749 ( .A(n7182), .B(creg[1]), .Z(n7179) );
  NAND U9750 ( .A(n7183), .B(o[1]), .Z(n7178) );
  AND U9751 ( .A(n7179), .B(n7178), .Z(n7180) );
  NANDN U9752 ( .A(n7181), .B(n7180), .Z(n2055) );
  NANDN U9753 ( .A(n7182), .B(creg[0]), .Z(n7185) );
  NAND U9754 ( .A(n7183), .B(o[0]), .Z(n7184) );
  AND U9755 ( .A(n7185), .B(n7184), .Z(n7186) );
  NANDN U9756 ( .A(n7187), .B(n7186), .Z(n2056) );
  AND U9757 ( .A(start_in[127]), .B(mul_pow), .Z(n8206) );
  NANDN U9758 ( .A(n7188), .B(n8206), .Z(n7189) );
  NANDN U9759 ( .A(first_one), .B(n7189), .Z(n2057) );
  NAND U9760 ( .A(n8206), .B(ereg[254]), .Z(n7191) );
  NANDN U9761 ( .A(n8206), .B(init), .Z(n8211) );
  NANDN U9762 ( .A(n8211), .B(ereg[255]), .Z(n7190) );
  AND U9763 ( .A(n7191), .B(n7190), .Z(n7192) );
  NANDN U9764 ( .A(n7193), .B(n7192), .Z(n2058) );
  NAND U9765 ( .A(n8206), .B(ereg[253]), .Z(n7195) );
  NANDN U9766 ( .A(init), .B(e[254]), .Z(n7194) );
  AND U9767 ( .A(n7195), .B(n7194), .Z(n7197) );
  NANDN U9768 ( .A(n8211), .B(ereg[254]), .Z(n7196) );
  NAND U9769 ( .A(n7197), .B(n7196), .Z(n2059) );
  NAND U9770 ( .A(n8206), .B(ereg[252]), .Z(n7199) );
  NANDN U9771 ( .A(init), .B(e[253]), .Z(n7198) );
  AND U9772 ( .A(n7199), .B(n7198), .Z(n7201) );
  NANDN U9773 ( .A(n8211), .B(ereg[253]), .Z(n7200) );
  NAND U9774 ( .A(n7201), .B(n7200), .Z(n2060) );
  NAND U9775 ( .A(n8206), .B(ereg[251]), .Z(n7203) );
  NANDN U9776 ( .A(init), .B(e[252]), .Z(n7202) );
  AND U9777 ( .A(n7203), .B(n7202), .Z(n7205) );
  NANDN U9778 ( .A(n8211), .B(ereg[252]), .Z(n7204) );
  NAND U9779 ( .A(n7205), .B(n7204), .Z(n2061) );
  NAND U9780 ( .A(n8206), .B(ereg[250]), .Z(n7207) );
  NANDN U9781 ( .A(init), .B(e[251]), .Z(n7206) );
  AND U9782 ( .A(n7207), .B(n7206), .Z(n7209) );
  NANDN U9783 ( .A(n8211), .B(ereg[251]), .Z(n7208) );
  NAND U9784 ( .A(n7209), .B(n7208), .Z(n2062) );
  NAND U9785 ( .A(n8206), .B(ereg[249]), .Z(n7211) );
  NANDN U9786 ( .A(init), .B(e[250]), .Z(n7210) );
  AND U9787 ( .A(n7211), .B(n7210), .Z(n7213) );
  NANDN U9788 ( .A(n8211), .B(ereg[250]), .Z(n7212) );
  NAND U9789 ( .A(n7213), .B(n7212), .Z(n2063) );
  NAND U9790 ( .A(n8206), .B(ereg[248]), .Z(n7215) );
  NANDN U9791 ( .A(init), .B(e[249]), .Z(n7214) );
  AND U9792 ( .A(n7215), .B(n7214), .Z(n7217) );
  NANDN U9793 ( .A(n8211), .B(ereg[249]), .Z(n7216) );
  NAND U9794 ( .A(n7217), .B(n7216), .Z(n2064) );
  NAND U9795 ( .A(n8206), .B(ereg[247]), .Z(n7219) );
  NANDN U9796 ( .A(init), .B(e[248]), .Z(n7218) );
  AND U9797 ( .A(n7219), .B(n7218), .Z(n7221) );
  NANDN U9798 ( .A(n8211), .B(ereg[248]), .Z(n7220) );
  NAND U9799 ( .A(n7221), .B(n7220), .Z(n2065) );
  NAND U9800 ( .A(n8206), .B(ereg[246]), .Z(n7223) );
  NANDN U9801 ( .A(init), .B(e[247]), .Z(n7222) );
  AND U9802 ( .A(n7223), .B(n7222), .Z(n7225) );
  NANDN U9803 ( .A(n8211), .B(ereg[247]), .Z(n7224) );
  NAND U9804 ( .A(n7225), .B(n7224), .Z(n2066) );
  NAND U9805 ( .A(n8206), .B(ereg[245]), .Z(n7227) );
  NANDN U9806 ( .A(init), .B(e[246]), .Z(n7226) );
  AND U9807 ( .A(n7227), .B(n7226), .Z(n7229) );
  NANDN U9808 ( .A(n8211), .B(ereg[246]), .Z(n7228) );
  NAND U9809 ( .A(n7229), .B(n7228), .Z(n2067) );
  NAND U9810 ( .A(n8206), .B(ereg[244]), .Z(n7231) );
  NANDN U9811 ( .A(init), .B(e[245]), .Z(n7230) );
  AND U9812 ( .A(n7231), .B(n7230), .Z(n7233) );
  NANDN U9813 ( .A(n8211), .B(ereg[245]), .Z(n7232) );
  NAND U9814 ( .A(n7233), .B(n7232), .Z(n2068) );
  NAND U9815 ( .A(n8206), .B(ereg[243]), .Z(n7235) );
  NANDN U9816 ( .A(init), .B(e[244]), .Z(n7234) );
  AND U9817 ( .A(n7235), .B(n7234), .Z(n7237) );
  NANDN U9818 ( .A(n8211), .B(ereg[244]), .Z(n7236) );
  NAND U9819 ( .A(n7237), .B(n7236), .Z(n2069) );
  NAND U9820 ( .A(n8206), .B(ereg[242]), .Z(n7239) );
  NANDN U9821 ( .A(init), .B(e[243]), .Z(n7238) );
  AND U9822 ( .A(n7239), .B(n7238), .Z(n7241) );
  NANDN U9823 ( .A(n8211), .B(ereg[243]), .Z(n7240) );
  NAND U9824 ( .A(n7241), .B(n7240), .Z(n2070) );
  NAND U9825 ( .A(n8206), .B(ereg[241]), .Z(n7243) );
  NANDN U9826 ( .A(init), .B(e[242]), .Z(n7242) );
  AND U9827 ( .A(n7243), .B(n7242), .Z(n7245) );
  NANDN U9828 ( .A(n8211), .B(ereg[242]), .Z(n7244) );
  NAND U9829 ( .A(n7245), .B(n7244), .Z(n2071) );
  NAND U9830 ( .A(n8206), .B(ereg[240]), .Z(n7247) );
  NANDN U9831 ( .A(init), .B(e[241]), .Z(n7246) );
  AND U9832 ( .A(n7247), .B(n7246), .Z(n7249) );
  NANDN U9833 ( .A(n8211), .B(ereg[241]), .Z(n7248) );
  NAND U9834 ( .A(n7249), .B(n7248), .Z(n2072) );
  NAND U9835 ( .A(n8206), .B(ereg[239]), .Z(n7251) );
  NANDN U9836 ( .A(init), .B(e[240]), .Z(n7250) );
  AND U9837 ( .A(n7251), .B(n7250), .Z(n7253) );
  NANDN U9838 ( .A(n8211), .B(ereg[240]), .Z(n7252) );
  NAND U9839 ( .A(n7253), .B(n7252), .Z(n2073) );
  NAND U9840 ( .A(n8206), .B(ereg[238]), .Z(n7255) );
  NANDN U9841 ( .A(init), .B(e[239]), .Z(n7254) );
  AND U9842 ( .A(n7255), .B(n7254), .Z(n7257) );
  NANDN U9843 ( .A(n8211), .B(ereg[239]), .Z(n7256) );
  NAND U9844 ( .A(n7257), .B(n7256), .Z(n2074) );
  NAND U9845 ( .A(n8206), .B(ereg[237]), .Z(n7259) );
  NANDN U9846 ( .A(init), .B(e[238]), .Z(n7258) );
  AND U9847 ( .A(n7259), .B(n7258), .Z(n7261) );
  NANDN U9848 ( .A(n8211), .B(ereg[238]), .Z(n7260) );
  NAND U9849 ( .A(n7261), .B(n7260), .Z(n2075) );
  NAND U9850 ( .A(n8206), .B(ereg[236]), .Z(n7263) );
  NANDN U9851 ( .A(init), .B(e[237]), .Z(n7262) );
  AND U9852 ( .A(n7263), .B(n7262), .Z(n7265) );
  NANDN U9853 ( .A(n8211), .B(ereg[237]), .Z(n7264) );
  NAND U9854 ( .A(n7265), .B(n7264), .Z(n2076) );
  NAND U9855 ( .A(n8206), .B(ereg[235]), .Z(n7267) );
  NANDN U9856 ( .A(init), .B(e[236]), .Z(n7266) );
  AND U9857 ( .A(n7267), .B(n7266), .Z(n7269) );
  NANDN U9858 ( .A(n8211), .B(ereg[236]), .Z(n7268) );
  NAND U9859 ( .A(n7269), .B(n7268), .Z(n2077) );
  NAND U9860 ( .A(n8206), .B(ereg[234]), .Z(n7271) );
  NANDN U9861 ( .A(init), .B(e[235]), .Z(n7270) );
  AND U9862 ( .A(n7271), .B(n7270), .Z(n7273) );
  NANDN U9863 ( .A(n8211), .B(ereg[235]), .Z(n7272) );
  NAND U9864 ( .A(n7273), .B(n7272), .Z(n2078) );
  NAND U9865 ( .A(n8206), .B(ereg[233]), .Z(n7275) );
  NANDN U9866 ( .A(init), .B(e[234]), .Z(n7274) );
  AND U9867 ( .A(n7275), .B(n7274), .Z(n7277) );
  NANDN U9868 ( .A(n8211), .B(ereg[234]), .Z(n7276) );
  NAND U9869 ( .A(n7277), .B(n7276), .Z(n2079) );
  NAND U9870 ( .A(n8206), .B(ereg[232]), .Z(n7279) );
  NANDN U9871 ( .A(init), .B(e[233]), .Z(n7278) );
  AND U9872 ( .A(n7279), .B(n7278), .Z(n7281) );
  NANDN U9873 ( .A(n8211), .B(ereg[233]), .Z(n7280) );
  NAND U9874 ( .A(n7281), .B(n7280), .Z(n2080) );
  NAND U9875 ( .A(n8206), .B(ereg[231]), .Z(n7283) );
  NANDN U9876 ( .A(init), .B(e[232]), .Z(n7282) );
  AND U9877 ( .A(n7283), .B(n7282), .Z(n7285) );
  NANDN U9878 ( .A(n8211), .B(ereg[232]), .Z(n7284) );
  NAND U9879 ( .A(n7285), .B(n7284), .Z(n2081) );
  NAND U9880 ( .A(n8206), .B(ereg[230]), .Z(n7287) );
  NANDN U9881 ( .A(init), .B(e[231]), .Z(n7286) );
  AND U9882 ( .A(n7287), .B(n7286), .Z(n7289) );
  NANDN U9883 ( .A(n8211), .B(ereg[231]), .Z(n7288) );
  NAND U9884 ( .A(n7289), .B(n7288), .Z(n2082) );
  NAND U9885 ( .A(n8206), .B(ereg[229]), .Z(n7291) );
  NANDN U9886 ( .A(init), .B(e[230]), .Z(n7290) );
  AND U9887 ( .A(n7291), .B(n7290), .Z(n7293) );
  NANDN U9888 ( .A(n8211), .B(ereg[230]), .Z(n7292) );
  NAND U9889 ( .A(n7293), .B(n7292), .Z(n2083) );
  NAND U9890 ( .A(n8206), .B(ereg[228]), .Z(n7295) );
  NANDN U9891 ( .A(init), .B(e[229]), .Z(n7294) );
  AND U9892 ( .A(n7295), .B(n7294), .Z(n7297) );
  NANDN U9893 ( .A(n8211), .B(ereg[229]), .Z(n7296) );
  NAND U9894 ( .A(n7297), .B(n7296), .Z(n2084) );
  NAND U9895 ( .A(n8206), .B(ereg[227]), .Z(n7299) );
  NANDN U9896 ( .A(init), .B(e[228]), .Z(n7298) );
  AND U9897 ( .A(n7299), .B(n7298), .Z(n7301) );
  NANDN U9898 ( .A(n8211), .B(ereg[228]), .Z(n7300) );
  NAND U9899 ( .A(n7301), .B(n7300), .Z(n2085) );
  NAND U9900 ( .A(n8206), .B(ereg[226]), .Z(n7303) );
  NANDN U9901 ( .A(init), .B(e[227]), .Z(n7302) );
  AND U9902 ( .A(n7303), .B(n7302), .Z(n7305) );
  NANDN U9903 ( .A(n8211), .B(ereg[227]), .Z(n7304) );
  NAND U9904 ( .A(n7305), .B(n7304), .Z(n2086) );
  NAND U9905 ( .A(n8206), .B(ereg[225]), .Z(n7307) );
  NANDN U9906 ( .A(init), .B(e[226]), .Z(n7306) );
  AND U9907 ( .A(n7307), .B(n7306), .Z(n7309) );
  NANDN U9908 ( .A(n8211), .B(ereg[226]), .Z(n7308) );
  NAND U9909 ( .A(n7309), .B(n7308), .Z(n2087) );
  NAND U9910 ( .A(n8206), .B(ereg[224]), .Z(n7311) );
  NANDN U9911 ( .A(init), .B(e[225]), .Z(n7310) );
  AND U9912 ( .A(n7311), .B(n7310), .Z(n7313) );
  NANDN U9913 ( .A(n8211), .B(ereg[225]), .Z(n7312) );
  NAND U9914 ( .A(n7313), .B(n7312), .Z(n2088) );
  NAND U9915 ( .A(n8206), .B(ereg[223]), .Z(n7315) );
  NANDN U9916 ( .A(init), .B(e[224]), .Z(n7314) );
  AND U9917 ( .A(n7315), .B(n7314), .Z(n7317) );
  NANDN U9918 ( .A(n8211), .B(ereg[224]), .Z(n7316) );
  NAND U9919 ( .A(n7317), .B(n7316), .Z(n2089) );
  NAND U9920 ( .A(n8206), .B(ereg[222]), .Z(n7319) );
  NANDN U9921 ( .A(init), .B(e[223]), .Z(n7318) );
  AND U9922 ( .A(n7319), .B(n7318), .Z(n7321) );
  NANDN U9923 ( .A(n8211), .B(ereg[223]), .Z(n7320) );
  NAND U9924 ( .A(n7321), .B(n7320), .Z(n2090) );
  NAND U9925 ( .A(n8206), .B(ereg[221]), .Z(n7323) );
  NANDN U9926 ( .A(init), .B(e[222]), .Z(n7322) );
  AND U9927 ( .A(n7323), .B(n7322), .Z(n7325) );
  NANDN U9928 ( .A(n8211), .B(ereg[222]), .Z(n7324) );
  NAND U9929 ( .A(n7325), .B(n7324), .Z(n2091) );
  NAND U9930 ( .A(n8206), .B(ereg[220]), .Z(n7327) );
  NANDN U9931 ( .A(init), .B(e[221]), .Z(n7326) );
  AND U9932 ( .A(n7327), .B(n7326), .Z(n7329) );
  NANDN U9933 ( .A(n8211), .B(ereg[221]), .Z(n7328) );
  NAND U9934 ( .A(n7329), .B(n7328), .Z(n2092) );
  NAND U9935 ( .A(n8206), .B(ereg[219]), .Z(n7331) );
  NANDN U9936 ( .A(init), .B(e[220]), .Z(n7330) );
  AND U9937 ( .A(n7331), .B(n7330), .Z(n7333) );
  NANDN U9938 ( .A(n8211), .B(ereg[220]), .Z(n7332) );
  NAND U9939 ( .A(n7333), .B(n7332), .Z(n2093) );
  NAND U9940 ( .A(n8206), .B(ereg[218]), .Z(n7335) );
  NANDN U9941 ( .A(init), .B(e[219]), .Z(n7334) );
  AND U9942 ( .A(n7335), .B(n7334), .Z(n7337) );
  NANDN U9943 ( .A(n8211), .B(ereg[219]), .Z(n7336) );
  NAND U9944 ( .A(n7337), .B(n7336), .Z(n2094) );
  NAND U9945 ( .A(n8206), .B(ereg[217]), .Z(n7339) );
  NANDN U9946 ( .A(init), .B(e[218]), .Z(n7338) );
  AND U9947 ( .A(n7339), .B(n7338), .Z(n7341) );
  NANDN U9948 ( .A(n8211), .B(ereg[218]), .Z(n7340) );
  NAND U9949 ( .A(n7341), .B(n7340), .Z(n2095) );
  NAND U9950 ( .A(n8206), .B(ereg[216]), .Z(n7343) );
  NANDN U9951 ( .A(init), .B(e[217]), .Z(n7342) );
  AND U9952 ( .A(n7343), .B(n7342), .Z(n7345) );
  NANDN U9953 ( .A(n8211), .B(ereg[217]), .Z(n7344) );
  NAND U9954 ( .A(n7345), .B(n7344), .Z(n2096) );
  NAND U9955 ( .A(n8206), .B(ereg[215]), .Z(n7347) );
  NANDN U9956 ( .A(init), .B(e[216]), .Z(n7346) );
  AND U9957 ( .A(n7347), .B(n7346), .Z(n7349) );
  NANDN U9958 ( .A(n8211), .B(ereg[216]), .Z(n7348) );
  NAND U9959 ( .A(n7349), .B(n7348), .Z(n2097) );
  NAND U9960 ( .A(n8206), .B(ereg[214]), .Z(n7351) );
  NANDN U9961 ( .A(init), .B(e[215]), .Z(n7350) );
  AND U9962 ( .A(n7351), .B(n7350), .Z(n7353) );
  NANDN U9963 ( .A(n8211), .B(ereg[215]), .Z(n7352) );
  NAND U9964 ( .A(n7353), .B(n7352), .Z(n2098) );
  NAND U9965 ( .A(n8206), .B(ereg[213]), .Z(n7355) );
  NANDN U9966 ( .A(init), .B(e[214]), .Z(n7354) );
  AND U9967 ( .A(n7355), .B(n7354), .Z(n7357) );
  NANDN U9968 ( .A(n8211), .B(ereg[214]), .Z(n7356) );
  NAND U9969 ( .A(n7357), .B(n7356), .Z(n2099) );
  NAND U9970 ( .A(n8206), .B(ereg[212]), .Z(n7359) );
  NANDN U9971 ( .A(init), .B(e[213]), .Z(n7358) );
  AND U9972 ( .A(n7359), .B(n7358), .Z(n7361) );
  NANDN U9973 ( .A(n8211), .B(ereg[213]), .Z(n7360) );
  NAND U9974 ( .A(n7361), .B(n7360), .Z(n2100) );
  NAND U9975 ( .A(n8206), .B(ereg[211]), .Z(n7363) );
  NANDN U9976 ( .A(init), .B(e[212]), .Z(n7362) );
  AND U9977 ( .A(n7363), .B(n7362), .Z(n7365) );
  NANDN U9978 ( .A(n8211), .B(ereg[212]), .Z(n7364) );
  NAND U9979 ( .A(n7365), .B(n7364), .Z(n2101) );
  NAND U9980 ( .A(n8206), .B(ereg[210]), .Z(n7367) );
  NANDN U9981 ( .A(init), .B(e[211]), .Z(n7366) );
  AND U9982 ( .A(n7367), .B(n7366), .Z(n7369) );
  NANDN U9983 ( .A(n8211), .B(ereg[211]), .Z(n7368) );
  NAND U9984 ( .A(n7369), .B(n7368), .Z(n2102) );
  NAND U9985 ( .A(n8206), .B(ereg[209]), .Z(n7371) );
  NANDN U9986 ( .A(init), .B(e[210]), .Z(n7370) );
  AND U9987 ( .A(n7371), .B(n7370), .Z(n7373) );
  NANDN U9988 ( .A(n8211), .B(ereg[210]), .Z(n7372) );
  NAND U9989 ( .A(n7373), .B(n7372), .Z(n2103) );
  NAND U9990 ( .A(n8206), .B(ereg[208]), .Z(n7375) );
  NANDN U9991 ( .A(init), .B(e[209]), .Z(n7374) );
  AND U9992 ( .A(n7375), .B(n7374), .Z(n7377) );
  NANDN U9993 ( .A(n8211), .B(ereg[209]), .Z(n7376) );
  NAND U9994 ( .A(n7377), .B(n7376), .Z(n2104) );
  NAND U9995 ( .A(n8206), .B(ereg[207]), .Z(n7379) );
  NANDN U9996 ( .A(init), .B(e[208]), .Z(n7378) );
  AND U9997 ( .A(n7379), .B(n7378), .Z(n7381) );
  NANDN U9998 ( .A(n8211), .B(ereg[208]), .Z(n7380) );
  NAND U9999 ( .A(n7381), .B(n7380), .Z(n2105) );
  NAND U10000 ( .A(n8206), .B(ereg[206]), .Z(n7383) );
  NANDN U10001 ( .A(init), .B(e[207]), .Z(n7382) );
  AND U10002 ( .A(n7383), .B(n7382), .Z(n7385) );
  NANDN U10003 ( .A(n8211), .B(ereg[207]), .Z(n7384) );
  NAND U10004 ( .A(n7385), .B(n7384), .Z(n2106) );
  NAND U10005 ( .A(n8206), .B(ereg[205]), .Z(n7387) );
  NANDN U10006 ( .A(init), .B(e[206]), .Z(n7386) );
  AND U10007 ( .A(n7387), .B(n7386), .Z(n7389) );
  NANDN U10008 ( .A(n8211), .B(ereg[206]), .Z(n7388) );
  NAND U10009 ( .A(n7389), .B(n7388), .Z(n2107) );
  NAND U10010 ( .A(n8206), .B(ereg[204]), .Z(n7391) );
  NANDN U10011 ( .A(init), .B(e[205]), .Z(n7390) );
  AND U10012 ( .A(n7391), .B(n7390), .Z(n7393) );
  NANDN U10013 ( .A(n8211), .B(ereg[205]), .Z(n7392) );
  NAND U10014 ( .A(n7393), .B(n7392), .Z(n2108) );
  NAND U10015 ( .A(n8206), .B(ereg[203]), .Z(n7395) );
  NANDN U10016 ( .A(init), .B(e[204]), .Z(n7394) );
  AND U10017 ( .A(n7395), .B(n7394), .Z(n7397) );
  NANDN U10018 ( .A(n8211), .B(ereg[204]), .Z(n7396) );
  NAND U10019 ( .A(n7397), .B(n7396), .Z(n2109) );
  NAND U10020 ( .A(n8206), .B(ereg[202]), .Z(n7399) );
  NANDN U10021 ( .A(init), .B(e[203]), .Z(n7398) );
  AND U10022 ( .A(n7399), .B(n7398), .Z(n7401) );
  NANDN U10023 ( .A(n8211), .B(ereg[203]), .Z(n7400) );
  NAND U10024 ( .A(n7401), .B(n7400), .Z(n2110) );
  NAND U10025 ( .A(n8206), .B(ereg[201]), .Z(n7403) );
  NANDN U10026 ( .A(init), .B(e[202]), .Z(n7402) );
  AND U10027 ( .A(n7403), .B(n7402), .Z(n7405) );
  NANDN U10028 ( .A(n8211), .B(ereg[202]), .Z(n7404) );
  NAND U10029 ( .A(n7405), .B(n7404), .Z(n2111) );
  NAND U10030 ( .A(n8206), .B(ereg[200]), .Z(n7407) );
  NANDN U10031 ( .A(init), .B(e[201]), .Z(n7406) );
  AND U10032 ( .A(n7407), .B(n7406), .Z(n7409) );
  NANDN U10033 ( .A(n8211), .B(ereg[201]), .Z(n7408) );
  NAND U10034 ( .A(n7409), .B(n7408), .Z(n2112) );
  NAND U10035 ( .A(n8206), .B(ereg[199]), .Z(n7411) );
  NANDN U10036 ( .A(init), .B(e[200]), .Z(n7410) );
  AND U10037 ( .A(n7411), .B(n7410), .Z(n7413) );
  NANDN U10038 ( .A(n8211), .B(ereg[200]), .Z(n7412) );
  NAND U10039 ( .A(n7413), .B(n7412), .Z(n2113) );
  NAND U10040 ( .A(n8206), .B(ereg[198]), .Z(n7415) );
  NANDN U10041 ( .A(init), .B(e[199]), .Z(n7414) );
  AND U10042 ( .A(n7415), .B(n7414), .Z(n7417) );
  NANDN U10043 ( .A(n8211), .B(ereg[199]), .Z(n7416) );
  NAND U10044 ( .A(n7417), .B(n7416), .Z(n2114) );
  NAND U10045 ( .A(n8206), .B(ereg[197]), .Z(n7419) );
  NANDN U10046 ( .A(init), .B(e[198]), .Z(n7418) );
  AND U10047 ( .A(n7419), .B(n7418), .Z(n7421) );
  NANDN U10048 ( .A(n8211), .B(ereg[198]), .Z(n7420) );
  NAND U10049 ( .A(n7421), .B(n7420), .Z(n2115) );
  NAND U10050 ( .A(n8206), .B(ereg[196]), .Z(n7423) );
  NANDN U10051 ( .A(init), .B(e[197]), .Z(n7422) );
  AND U10052 ( .A(n7423), .B(n7422), .Z(n7425) );
  NANDN U10053 ( .A(n8211), .B(ereg[197]), .Z(n7424) );
  NAND U10054 ( .A(n7425), .B(n7424), .Z(n2116) );
  NAND U10055 ( .A(n8206), .B(ereg[195]), .Z(n7427) );
  NANDN U10056 ( .A(init), .B(e[196]), .Z(n7426) );
  AND U10057 ( .A(n7427), .B(n7426), .Z(n7429) );
  NANDN U10058 ( .A(n8211), .B(ereg[196]), .Z(n7428) );
  NAND U10059 ( .A(n7429), .B(n7428), .Z(n2117) );
  NAND U10060 ( .A(n8206), .B(ereg[194]), .Z(n7431) );
  NANDN U10061 ( .A(init), .B(e[195]), .Z(n7430) );
  AND U10062 ( .A(n7431), .B(n7430), .Z(n7433) );
  NANDN U10063 ( .A(n8211), .B(ereg[195]), .Z(n7432) );
  NAND U10064 ( .A(n7433), .B(n7432), .Z(n2118) );
  NAND U10065 ( .A(n8206), .B(ereg[193]), .Z(n7435) );
  NANDN U10066 ( .A(init), .B(e[194]), .Z(n7434) );
  AND U10067 ( .A(n7435), .B(n7434), .Z(n7437) );
  NANDN U10068 ( .A(n8211), .B(ereg[194]), .Z(n7436) );
  NAND U10069 ( .A(n7437), .B(n7436), .Z(n2119) );
  NAND U10070 ( .A(n8206), .B(ereg[192]), .Z(n7439) );
  NANDN U10071 ( .A(init), .B(e[193]), .Z(n7438) );
  AND U10072 ( .A(n7439), .B(n7438), .Z(n7441) );
  NANDN U10073 ( .A(n8211), .B(ereg[193]), .Z(n7440) );
  NAND U10074 ( .A(n7441), .B(n7440), .Z(n2120) );
  NAND U10075 ( .A(n8206), .B(ereg[191]), .Z(n7443) );
  NANDN U10076 ( .A(init), .B(e[192]), .Z(n7442) );
  AND U10077 ( .A(n7443), .B(n7442), .Z(n7445) );
  NANDN U10078 ( .A(n8211), .B(ereg[192]), .Z(n7444) );
  NAND U10079 ( .A(n7445), .B(n7444), .Z(n2121) );
  NAND U10080 ( .A(n8206), .B(ereg[190]), .Z(n7447) );
  NANDN U10081 ( .A(init), .B(e[191]), .Z(n7446) );
  AND U10082 ( .A(n7447), .B(n7446), .Z(n7449) );
  NANDN U10083 ( .A(n8211), .B(ereg[191]), .Z(n7448) );
  NAND U10084 ( .A(n7449), .B(n7448), .Z(n2122) );
  NAND U10085 ( .A(n8206), .B(ereg[189]), .Z(n7451) );
  NANDN U10086 ( .A(init), .B(e[190]), .Z(n7450) );
  AND U10087 ( .A(n7451), .B(n7450), .Z(n7453) );
  NANDN U10088 ( .A(n8211), .B(ereg[190]), .Z(n7452) );
  NAND U10089 ( .A(n7453), .B(n7452), .Z(n2123) );
  NAND U10090 ( .A(n8206), .B(ereg[188]), .Z(n7455) );
  NANDN U10091 ( .A(init), .B(e[189]), .Z(n7454) );
  AND U10092 ( .A(n7455), .B(n7454), .Z(n7457) );
  NANDN U10093 ( .A(n8211), .B(ereg[189]), .Z(n7456) );
  NAND U10094 ( .A(n7457), .B(n7456), .Z(n2124) );
  NAND U10095 ( .A(n8206), .B(ereg[187]), .Z(n7459) );
  NANDN U10096 ( .A(init), .B(e[188]), .Z(n7458) );
  AND U10097 ( .A(n7459), .B(n7458), .Z(n7461) );
  NANDN U10098 ( .A(n8211), .B(ereg[188]), .Z(n7460) );
  NAND U10099 ( .A(n7461), .B(n7460), .Z(n2125) );
  NAND U10100 ( .A(n8206), .B(ereg[186]), .Z(n7463) );
  NANDN U10101 ( .A(init), .B(e[187]), .Z(n7462) );
  AND U10102 ( .A(n7463), .B(n7462), .Z(n7465) );
  NANDN U10103 ( .A(n8211), .B(ereg[187]), .Z(n7464) );
  NAND U10104 ( .A(n7465), .B(n7464), .Z(n2126) );
  NAND U10105 ( .A(n8206), .B(ereg[185]), .Z(n7467) );
  NANDN U10106 ( .A(init), .B(e[186]), .Z(n7466) );
  AND U10107 ( .A(n7467), .B(n7466), .Z(n7469) );
  NANDN U10108 ( .A(n8211), .B(ereg[186]), .Z(n7468) );
  NAND U10109 ( .A(n7469), .B(n7468), .Z(n2127) );
  NAND U10110 ( .A(n8206), .B(ereg[184]), .Z(n7471) );
  NANDN U10111 ( .A(init), .B(e[185]), .Z(n7470) );
  AND U10112 ( .A(n7471), .B(n7470), .Z(n7473) );
  NANDN U10113 ( .A(n8211), .B(ereg[185]), .Z(n7472) );
  NAND U10114 ( .A(n7473), .B(n7472), .Z(n2128) );
  NAND U10115 ( .A(n8206), .B(ereg[183]), .Z(n7475) );
  NANDN U10116 ( .A(init), .B(e[184]), .Z(n7474) );
  AND U10117 ( .A(n7475), .B(n7474), .Z(n7477) );
  NANDN U10118 ( .A(n8211), .B(ereg[184]), .Z(n7476) );
  NAND U10119 ( .A(n7477), .B(n7476), .Z(n2129) );
  NAND U10120 ( .A(n8206), .B(ereg[182]), .Z(n7479) );
  NANDN U10121 ( .A(init), .B(e[183]), .Z(n7478) );
  AND U10122 ( .A(n7479), .B(n7478), .Z(n7481) );
  NANDN U10123 ( .A(n8211), .B(ereg[183]), .Z(n7480) );
  NAND U10124 ( .A(n7481), .B(n7480), .Z(n2130) );
  NAND U10125 ( .A(n8206), .B(ereg[181]), .Z(n7483) );
  NANDN U10126 ( .A(init), .B(e[182]), .Z(n7482) );
  AND U10127 ( .A(n7483), .B(n7482), .Z(n7485) );
  NANDN U10128 ( .A(n8211), .B(ereg[182]), .Z(n7484) );
  NAND U10129 ( .A(n7485), .B(n7484), .Z(n2131) );
  NAND U10130 ( .A(n8206), .B(ereg[180]), .Z(n7487) );
  NANDN U10131 ( .A(init), .B(e[181]), .Z(n7486) );
  AND U10132 ( .A(n7487), .B(n7486), .Z(n7489) );
  NANDN U10133 ( .A(n8211), .B(ereg[181]), .Z(n7488) );
  NAND U10134 ( .A(n7489), .B(n7488), .Z(n2132) );
  NAND U10135 ( .A(n8206), .B(ereg[179]), .Z(n7491) );
  NANDN U10136 ( .A(init), .B(e[180]), .Z(n7490) );
  AND U10137 ( .A(n7491), .B(n7490), .Z(n7493) );
  NANDN U10138 ( .A(n8211), .B(ereg[180]), .Z(n7492) );
  NAND U10139 ( .A(n7493), .B(n7492), .Z(n2133) );
  NAND U10140 ( .A(n8206), .B(ereg[178]), .Z(n7495) );
  NANDN U10141 ( .A(init), .B(e[179]), .Z(n7494) );
  AND U10142 ( .A(n7495), .B(n7494), .Z(n7497) );
  NANDN U10143 ( .A(n8211), .B(ereg[179]), .Z(n7496) );
  NAND U10144 ( .A(n7497), .B(n7496), .Z(n2134) );
  NAND U10145 ( .A(n8206), .B(ereg[177]), .Z(n7499) );
  NANDN U10146 ( .A(init), .B(e[178]), .Z(n7498) );
  AND U10147 ( .A(n7499), .B(n7498), .Z(n7501) );
  NANDN U10148 ( .A(n8211), .B(ereg[178]), .Z(n7500) );
  NAND U10149 ( .A(n7501), .B(n7500), .Z(n2135) );
  NAND U10150 ( .A(n8206), .B(ereg[176]), .Z(n7503) );
  NANDN U10151 ( .A(init), .B(e[177]), .Z(n7502) );
  AND U10152 ( .A(n7503), .B(n7502), .Z(n7505) );
  NANDN U10153 ( .A(n8211), .B(ereg[177]), .Z(n7504) );
  NAND U10154 ( .A(n7505), .B(n7504), .Z(n2136) );
  NAND U10155 ( .A(n8206), .B(ereg[175]), .Z(n7507) );
  NANDN U10156 ( .A(init), .B(e[176]), .Z(n7506) );
  AND U10157 ( .A(n7507), .B(n7506), .Z(n7509) );
  NANDN U10158 ( .A(n8211), .B(ereg[176]), .Z(n7508) );
  NAND U10159 ( .A(n7509), .B(n7508), .Z(n2137) );
  NAND U10160 ( .A(n8206), .B(ereg[174]), .Z(n7511) );
  NANDN U10161 ( .A(init), .B(e[175]), .Z(n7510) );
  AND U10162 ( .A(n7511), .B(n7510), .Z(n7513) );
  NANDN U10163 ( .A(n8211), .B(ereg[175]), .Z(n7512) );
  NAND U10164 ( .A(n7513), .B(n7512), .Z(n2138) );
  NAND U10165 ( .A(n8206), .B(ereg[173]), .Z(n7515) );
  NANDN U10166 ( .A(init), .B(e[174]), .Z(n7514) );
  AND U10167 ( .A(n7515), .B(n7514), .Z(n7517) );
  NANDN U10168 ( .A(n8211), .B(ereg[174]), .Z(n7516) );
  NAND U10169 ( .A(n7517), .B(n7516), .Z(n2139) );
  NAND U10170 ( .A(n8206), .B(ereg[172]), .Z(n7519) );
  NANDN U10171 ( .A(init), .B(e[173]), .Z(n7518) );
  AND U10172 ( .A(n7519), .B(n7518), .Z(n7521) );
  NANDN U10173 ( .A(n8211), .B(ereg[173]), .Z(n7520) );
  NAND U10174 ( .A(n7521), .B(n7520), .Z(n2140) );
  NAND U10175 ( .A(n8206), .B(ereg[171]), .Z(n7523) );
  NANDN U10176 ( .A(init), .B(e[172]), .Z(n7522) );
  AND U10177 ( .A(n7523), .B(n7522), .Z(n7525) );
  NANDN U10178 ( .A(n8211), .B(ereg[172]), .Z(n7524) );
  NAND U10179 ( .A(n7525), .B(n7524), .Z(n2141) );
  NAND U10180 ( .A(n8206), .B(ereg[170]), .Z(n7527) );
  NANDN U10181 ( .A(init), .B(e[171]), .Z(n7526) );
  AND U10182 ( .A(n7527), .B(n7526), .Z(n7529) );
  NANDN U10183 ( .A(n8211), .B(ereg[171]), .Z(n7528) );
  NAND U10184 ( .A(n7529), .B(n7528), .Z(n2142) );
  NAND U10185 ( .A(n8206), .B(ereg[169]), .Z(n7531) );
  NANDN U10186 ( .A(init), .B(e[170]), .Z(n7530) );
  AND U10187 ( .A(n7531), .B(n7530), .Z(n7533) );
  NANDN U10188 ( .A(n8211), .B(ereg[170]), .Z(n7532) );
  NAND U10189 ( .A(n7533), .B(n7532), .Z(n2143) );
  NAND U10190 ( .A(n8206), .B(ereg[168]), .Z(n7535) );
  NANDN U10191 ( .A(init), .B(e[169]), .Z(n7534) );
  AND U10192 ( .A(n7535), .B(n7534), .Z(n7537) );
  NANDN U10193 ( .A(n8211), .B(ereg[169]), .Z(n7536) );
  NAND U10194 ( .A(n7537), .B(n7536), .Z(n2144) );
  NAND U10195 ( .A(n8206), .B(ereg[167]), .Z(n7539) );
  NANDN U10196 ( .A(init), .B(e[168]), .Z(n7538) );
  AND U10197 ( .A(n7539), .B(n7538), .Z(n7541) );
  NANDN U10198 ( .A(n8211), .B(ereg[168]), .Z(n7540) );
  NAND U10199 ( .A(n7541), .B(n7540), .Z(n2145) );
  NAND U10200 ( .A(n8206), .B(ereg[166]), .Z(n7543) );
  NANDN U10201 ( .A(init), .B(e[167]), .Z(n7542) );
  AND U10202 ( .A(n7543), .B(n7542), .Z(n7545) );
  NANDN U10203 ( .A(n8211), .B(ereg[167]), .Z(n7544) );
  NAND U10204 ( .A(n7545), .B(n7544), .Z(n2146) );
  NAND U10205 ( .A(n8206), .B(ereg[165]), .Z(n7547) );
  NANDN U10206 ( .A(init), .B(e[166]), .Z(n7546) );
  AND U10207 ( .A(n7547), .B(n7546), .Z(n7549) );
  NANDN U10208 ( .A(n8211), .B(ereg[166]), .Z(n7548) );
  NAND U10209 ( .A(n7549), .B(n7548), .Z(n2147) );
  NAND U10210 ( .A(n8206), .B(ereg[164]), .Z(n7551) );
  NANDN U10211 ( .A(init), .B(e[165]), .Z(n7550) );
  AND U10212 ( .A(n7551), .B(n7550), .Z(n7553) );
  NANDN U10213 ( .A(n8211), .B(ereg[165]), .Z(n7552) );
  NAND U10214 ( .A(n7553), .B(n7552), .Z(n2148) );
  NAND U10215 ( .A(n8206), .B(ereg[163]), .Z(n7555) );
  NANDN U10216 ( .A(init), .B(e[164]), .Z(n7554) );
  AND U10217 ( .A(n7555), .B(n7554), .Z(n7557) );
  NANDN U10218 ( .A(n8211), .B(ereg[164]), .Z(n7556) );
  NAND U10219 ( .A(n7557), .B(n7556), .Z(n2149) );
  NAND U10220 ( .A(n8206), .B(ereg[162]), .Z(n7559) );
  NANDN U10221 ( .A(init), .B(e[163]), .Z(n7558) );
  AND U10222 ( .A(n7559), .B(n7558), .Z(n7561) );
  NANDN U10223 ( .A(n8211), .B(ereg[163]), .Z(n7560) );
  NAND U10224 ( .A(n7561), .B(n7560), .Z(n2150) );
  NAND U10225 ( .A(n8206), .B(ereg[161]), .Z(n7563) );
  NANDN U10226 ( .A(init), .B(e[162]), .Z(n7562) );
  AND U10227 ( .A(n7563), .B(n7562), .Z(n7565) );
  NANDN U10228 ( .A(n8211), .B(ereg[162]), .Z(n7564) );
  NAND U10229 ( .A(n7565), .B(n7564), .Z(n2151) );
  NAND U10230 ( .A(n8206), .B(ereg[160]), .Z(n7567) );
  NANDN U10231 ( .A(init), .B(e[161]), .Z(n7566) );
  AND U10232 ( .A(n7567), .B(n7566), .Z(n7569) );
  NANDN U10233 ( .A(n8211), .B(ereg[161]), .Z(n7568) );
  NAND U10234 ( .A(n7569), .B(n7568), .Z(n2152) );
  NAND U10235 ( .A(n8206), .B(ereg[159]), .Z(n7571) );
  NANDN U10236 ( .A(init), .B(e[160]), .Z(n7570) );
  AND U10237 ( .A(n7571), .B(n7570), .Z(n7573) );
  NANDN U10238 ( .A(n8211), .B(ereg[160]), .Z(n7572) );
  NAND U10239 ( .A(n7573), .B(n7572), .Z(n2153) );
  NAND U10240 ( .A(n8206), .B(ereg[158]), .Z(n7575) );
  NANDN U10241 ( .A(init), .B(e[159]), .Z(n7574) );
  AND U10242 ( .A(n7575), .B(n7574), .Z(n7577) );
  NANDN U10243 ( .A(n8211), .B(ereg[159]), .Z(n7576) );
  NAND U10244 ( .A(n7577), .B(n7576), .Z(n2154) );
  NAND U10245 ( .A(n8206), .B(ereg[157]), .Z(n7579) );
  NANDN U10246 ( .A(init), .B(e[158]), .Z(n7578) );
  AND U10247 ( .A(n7579), .B(n7578), .Z(n7581) );
  NANDN U10248 ( .A(n8211), .B(ereg[158]), .Z(n7580) );
  NAND U10249 ( .A(n7581), .B(n7580), .Z(n2155) );
  NAND U10250 ( .A(n8206), .B(ereg[156]), .Z(n7583) );
  NANDN U10251 ( .A(init), .B(e[157]), .Z(n7582) );
  AND U10252 ( .A(n7583), .B(n7582), .Z(n7585) );
  NANDN U10253 ( .A(n8211), .B(ereg[157]), .Z(n7584) );
  NAND U10254 ( .A(n7585), .B(n7584), .Z(n2156) );
  NAND U10255 ( .A(n8206), .B(ereg[155]), .Z(n7587) );
  NANDN U10256 ( .A(init), .B(e[156]), .Z(n7586) );
  AND U10257 ( .A(n7587), .B(n7586), .Z(n7589) );
  NANDN U10258 ( .A(n8211), .B(ereg[156]), .Z(n7588) );
  NAND U10259 ( .A(n7589), .B(n7588), .Z(n2157) );
  NAND U10260 ( .A(n8206), .B(ereg[154]), .Z(n7591) );
  NANDN U10261 ( .A(init), .B(e[155]), .Z(n7590) );
  AND U10262 ( .A(n7591), .B(n7590), .Z(n7593) );
  NANDN U10263 ( .A(n8211), .B(ereg[155]), .Z(n7592) );
  NAND U10264 ( .A(n7593), .B(n7592), .Z(n2158) );
  NAND U10265 ( .A(n8206), .B(ereg[153]), .Z(n7595) );
  NANDN U10266 ( .A(init), .B(e[154]), .Z(n7594) );
  AND U10267 ( .A(n7595), .B(n7594), .Z(n7597) );
  NANDN U10268 ( .A(n8211), .B(ereg[154]), .Z(n7596) );
  NAND U10269 ( .A(n7597), .B(n7596), .Z(n2159) );
  NAND U10270 ( .A(n8206), .B(ereg[152]), .Z(n7599) );
  NANDN U10271 ( .A(init), .B(e[153]), .Z(n7598) );
  AND U10272 ( .A(n7599), .B(n7598), .Z(n7601) );
  NANDN U10273 ( .A(n8211), .B(ereg[153]), .Z(n7600) );
  NAND U10274 ( .A(n7601), .B(n7600), .Z(n2160) );
  NAND U10275 ( .A(n8206), .B(ereg[151]), .Z(n7603) );
  NANDN U10276 ( .A(init), .B(e[152]), .Z(n7602) );
  AND U10277 ( .A(n7603), .B(n7602), .Z(n7605) );
  NANDN U10278 ( .A(n8211), .B(ereg[152]), .Z(n7604) );
  NAND U10279 ( .A(n7605), .B(n7604), .Z(n2161) );
  NAND U10280 ( .A(n8206), .B(ereg[150]), .Z(n7607) );
  NANDN U10281 ( .A(init), .B(e[151]), .Z(n7606) );
  AND U10282 ( .A(n7607), .B(n7606), .Z(n7609) );
  NANDN U10283 ( .A(n8211), .B(ereg[151]), .Z(n7608) );
  NAND U10284 ( .A(n7609), .B(n7608), .Z(n2162) );
  NAND U10285 ( .A(n8206), .B(ereg[149]), .Z(n7611) );
  NANDN U10286 ( .A(init), .B(e[150]), .Z(n7610) );
  AND U10287 ( .A(n7611), .B(n7610), .Z(n7613) );
  NANDN U10288 ( .A(n8211), .B(ereg[150]), .Z(n7612) );
  NAND U10289 ( .A(n7613), .B(n7612), .Z(n2163) );
  NAND U10290 ( .A(n8206), .B(ereg[148]), .Z(n7615) );
  NANDN U10291 ( .A(init), .B(e[149]), .Z(n7614) );
  AND U10292 ( .A(n7615), .B(n7614), .Z(n7617) );
  NANDN U10293 ( .A(n8211), .B(ereg[149]), .Z(n7616) );
  NAND U10294 ( .A(n7617), .B(n7616), .Z(n2164) );
  NAND U10295 ( .A(n8206), .B(ereg[147]), .Z(n7619) );
  NANDN U10296 ( .A(init), .B(e[148]), .Z(n7618) );
  AND U10297 ( .A(n7619), .B(n7618), .Z(n7621) );
  NANDN U10298 ( .A(n8211), .B(ereg[148]), .Z(n7620) );
  NAND U10299 ( .A(n7621), .B(n7620), .Z(n2165) );
  NAND U10300 ( .A(n8206), .B(ereg[146]), .Z(n7623) );
  NANDN U10301 ( .A(init), .B(e[147]), .Z(n7622) );
  AND U10302 ( .A(n7623), .B(n7622), .Z(n7625) );
  NANDN U10303 ( .A(n8211), .B(ereg[147]), .Z(n7624) );
  NAND U10304 ( .A(n7625), .B(n7624), .Z(n2166) );
  NAND U10305 ( .A(n8206), .B(ereg[145]), .Z(n7627) );
  NANDN U10306 ( .A(init), .B(e[146]), .Z(n7626) );
  AND U10307 ( .A(n7627), .B(n7626), .Z(n7629) );
  NANDN U10308 ( .A(n8211), .B(ereg[146]), .Z(n7628) );
  NAND U10309 ( .A(n7629), .B(n7628), .Z(n2167) );
  NAND U10310 ( .A(n8206), .B(ereg[144]), .Z(n7631) );
  NANDN U10311 ( .A(init), .B(e[145]), .Z(n7630) );
  AND U10312 ( .A(n7631), .B(n7630), .Z(n7633) );
  NANDN U10313 ( .A(n8211), .B(ereg[145]), .Z(n7632) );
  NAND U10314 ( .A(n7633), .B(n7632), .Z(n2168) );
  NAND U10315 ( .A(n8206), .B(ereg[143]), .Z(n7635) );
  NANDN U10316 ( .A(init), .B(e[144]), .Z(n7634) );
  AND U10317 ( .A(n7635), .B(n7634), .Z(n7637) );
  NANDN U10318 ( .A(n8211), .B(ereg[144]), .Z(n7636) );
  NAND U10319 ( .A(n7637), .B(n7636), .Z(n2169) );
  NAND U10320 ( .A(n8206), .B(ereg[142]), .Z(n7639) );
  NANDN U10321 ( .A(init), .B(e[143]), .Z(n7638) );
  AND U10322 ( .A(n7639), .B(n7638), .Z(n7641) );
  NANDN U10323 ( .A(n8211), .B(ereg[143]), .Z(n7640) );
  NAND U10324 ( .A(n7641), .B(n7640), .Z(n2170) );
  NAND U10325 ( .A(n8206), .B(ereg[141]), .Z(n7643) );
  NANDN U10326 ( .A(init), .B(e[142]), .Z(n7642) );
  AND U10327 ( .A(n7643), .B(n7642), .Z(n7645) );
  NANDN U10328 ( .A(n8211), .B(ereg[142]), .Z(n7644) );
  NAND U10329 ( .A(n7645), .B(n7644), .Z(n2171) );
  NAND U10330 ( .A(n8206), .B(ereg[140]), .Z(n7647) );
  NANDN U10331 ( .A(init), .B(e[141]), .Z(n7646) );
  AND U10332 ( .A(n7647), .B(n7646), .Z(n7649) );
  NANDN U10333 ( .A(n8211), .B(ereg[141]), .Z(n7648) );
  NAND U10334 ( .A(n7649), .B(n7648), .Z(n2172) );
  NAND U10335 ( .A(n8206), .B(ereg[139]), .Z(n7651) );
  NANDN U10336 ( .A(init), .B(e[140]), .Z(n7650) );
  AND U10337 ( .A(n7651), .B(n7650), .Z(n7653) );
  NANDN U10338 ( .A(n8211), .B(ereg[140]), .Z(n7652) );
  NAND U10339 ( .A(n7653), .B(n7652), .Z(n2173) );
  NAND U10340 ( .A(n8206), .B(ereg[138]), .Z(n7655) );
  NANDN U10341 ( .A(init), .B(e[139]), .Z(n7654) );
  AND U10342 ( .A(n7655), .B(n7654), .Z(n7657) );
  NANDN U10343 ( .A(n8211), .B(ereg[139]), .Z(n7656) );
  NAND U10344 ( .A(n7657), .B(n7656), .Z(n2174) );
  NAND U10345 ( .A(n8206), .B(ereg[137]), .Z(n7659) );
  NANDN U10346 ( .A(init), .B(e[138]), .Z(n7658) );
  AND U10347 ( .A(n7659), .B(n7658), .Z(n7661) );
  NANDN U10348 ( .A(n8211), .B(ereg[138]), .Z(n7660) );
  NAND U10349 ( .A(n7661), .B(n7660), .Z(n2175) );
  NAND U10350 ( .A(n8206), .B(ereg[136]), .Z(n7663) );
  NANDN U10351 ( .A(init), .B(e[137]), .Z(n7662) );
  AND U10352 ( .A(n7663), .B(n7662), .Z(n7665) );
  NANDN U10353 ( .A(n8211), .B(ereg[137]), .Z(n7664) );
  NAND U10354 ( .A(n7665), .B(n7664), .Z(n2176) );
  NAND U10355 ( .A(n8206), .B(ereg[135]), .Z(n7667) );
  NANDN U10356 ( .A(init), .B(e[136]), .Z(n7666) );
  AND U10357 ( .A(n7667), .B(n7666), .Z(n7669) );
  NANDN U10358 ( .A(n8211), .B(ereg[136]), .Z(n7668) );
  NAND U10359 ( .A(n7669), .B(n7668), .Z(n2177) );
  NAND U10360 ( .A(n8206), .B(ereg[134]), .Z(n7671) );
  NANDN U10361 ( .A(init), .B(e[135]), .Z(n7670) );
  AND U10362 ( .A(n7671), .B(n7670), .Z(n7673) );
  NANDN U10363 ( .A(n8211), .B(ereg[135]), .Z(n7672) );
  NAND U10364 ( .A(n7673), .B(n7672), .Z(n2178) );
  NAND U10365 ( .A(n8206), .B(ereg[133]), .Z(n7675) );
  NANDN U10366 ( .A(init), .B(e[134]), .Z(n7674) );
  AND U10367 ( .A(n7675), .B(n7674), .Z(n7677) );
  NANDN U10368 ( .A(n8211), .B(ereg[134]), .Z(n7676) );
  NAND U10369 ( .A(n7677), .B(n7676), .Z(n2179) );
  NAND U10370 ( .A(n8206), .B(ereg[132]), .Z(n7679) );
  NANDN U10371 ( .A(init), .B(e[133]), .Z(n7678) );
  AND U10372 ( .A(n7679), .B(n7678), .Z(n7681) );
  NANDN U10373 ( .A(n8211), .B(ereg[133]), .Z(n7680) );
  NAND U10374 ( .A(n7681), .B(n7680), .Z(n2180) );
  NAND U10375 ( .A(n8206), .B(ereg[131]), .Z(n7683) );
  NANDN U10376 ( .A(init), .B(e[132]), .Z(n7682) );
  AND U10377 ( .A(n7683), .B(n7682), .Z(n7685) );
  NANDN U10378 ( .A(n8211), .B(ereg[132]), .Z(n7684) );
  NAND U10379 ( .A(n7685), .B(n7684), .Z(n2181) );
  NAND U10380 ( .A(n8206), .B(ereg[130]), .Z(n7687) );
  NANDN U10381 ( .A(init), .B(e[131]), .Z(n7686) );
  AND U10382 ( .A(n7687), .B(n7686), .Z(n7689) );
  NANDN U10383 ( .A(n8211), .B(ereg[131]), .Z(n7688) );
  NAND U10384 ( .A(n7689), .B(n7688), .Z(n2182) );
  NAND U10385 ( .A(n8206), .B(ereg[129]), .Z(n7691) );
  NANDN U10386 ( .A(init), .B(e[130]), .Z(n7690) );
  AND U10387 ( .A(n7691), .B(n7690), .Z(n7693) );
  NANDN U10388 ( .A(n8211), .B(ereg[130]), .Z(n7692) );
  NAND U10389 ( .A(n7693), .B(n7692), .Z(n2183) );
  NAND U10390 ( .A(n8206), .B(ereg[128]), .Z(n7695) );
  NANDN U10391 ( .A(init), .B(e[129]), .Z(n7694) );
  AND U10392 ( .A(n7695), .B(n7694), .Z(n7697) );
  NANDN U10393 ( .A(n8211), .B(ereg[129]), .Z(n7696) );
  NAND U10394 ( .A(n7697), .B(n7696), .Z(n2184) );
  NAND U10395 ( .A(n8206), .B(ereg[127]), .Z(n7699) );
  NANDN U10396 ( .A(init), .B(e[128]), .Z(n7698) );
  AND U10397 ( .A(n7699), .B(n7698), .Z(n7701) );
  NANDN U10398 ( .A(n8211), .B(ereg[128]), .Z(n7700) );
  NAND U10399 ( .A(n7701), .B(n7700), .Z(n2185) );
  NAND U10400 ( .A(n8206), .B(ereg[126]), .Z(n7703) );
  NANDN U10401 ( .A(init), .B(e[127]), .Z(n7702) );
  AND U10402 ( .A(n7703), .B(n7702), .Z(n7705) );
  NANDN U10403 ( .A(n8211), .B(ereg[127]), .Z(n7704) );
  NAND U10404 ( .A(n7705), .B(n7704), .Z(n2186) );
  NAND U10405 ( .A(n8206), .B(ereg[125]), .Z(n7707) );
  NANDN U10406 ( .A(init), .B(e[126]), .Z(n7706) );
  AND U10407 ( .A(n7707), .B(n7706), .Z(n7709) );
  NANDN U10408 ( .A(n8211), .B(ereg[126]), .Z(n7708) );
  NAND U10409 ( .A(n7709), .B(n7708), .Z(n2187) );
  NAND U10410 ( .A(n8206), .B(ereg[124]), .Z(n7711) );
  NANDN U10411 ( .A(init), .B(e[125]), .Z(n7710) );
  AND U10412 ( .A(n7711), .B(n7710), .Z(n7713) );
  NANDN U10413 ( .A(n8211), .B(ereg[125]), .Z(n7712) );
  NAND U10414 ( .A(n7713), .B(n7712), .Z(n2188) );
  NAND U10415 ( .A(n8206), .B(ereg[123]), .Z(n7715) );
  NANDN U10416 ( .A(init), .B(e[124]), .Z(n7714) );
  AND U10417 ( .A(n7715), .B(n7714), .Z(n7717) );
  NANDN U10418 ( .A(n8211), .B(ereg[124]), .Z(n7716) );
  NAND U10419 ( .A(n7717), .B(n7716), .Z(n2189) );
  NAND U10420 ( .A(n8206), .B(ereg[122]), .Z(n7719) );
  NANDN U10421 ( .A(init), .B(e[123]), .Z(n7718) );
  AND U10422 ( .A(n7719), .B(n7718), .Z(n7721) );
  NANDN U10423 ( .A(n8211), .B(ereg[123]), .Z(n7720) );
  NAND U10424 ( .A(n7721), .B(n7720), .Z(n2190) );
  NAND U10425 ( .A(n8206), .B(ereg[121]), .Z(n7723) );
  NANDN U10426 ( .A(init), .B(e[122]), .Z(n7722) );
  AND U10427 ( .A(n7723), .B(n7722), .Z(n7725) );
  NANDN U10428 ( .A(n8211), .B(ereg[122]), .Z(n7724) );
  NAND U10429 ( .A(n7725), .B(n7724), .Z(n2191) );
  NAND U10430 ( .A(n8206), .B(ereg[120]), .Z(n7727) );
  NANDN U10431 ( .A(init), .B(e[121]), .Z(n7726) );
  AND U10432 ( .A(n7727), .B(n7726), .Z(n7729) );
  NANDN U10433 ( .A(n8211), .B(ereg[121]), .Z(n7728) );
  NAND U10434 ( .A(n7729), .B(n7728), .Z(n2192) );
  NAND U10435 ( .A(n8206), .B(ereg[119]), .Z(n7731) );
  NANDN U10436 ( .A(init), .B(e[120]), .Z(n7730) );
  AND U10437 ( .A(n7731), .B(n7730), .Z(n7733) );
  NANDN U10438 ( .A(n8211), .B(ereg[120]), .Z(n7732) );
  NAND U10439 ( .A(n7733), .B(n7732), .Z(n2193) );
  NAND U10440 ( .A(n8206), .B(ereg[118]), .Z(n7735) );
  NANDN U10441 ( .A(init), .B(e[119]), .Z(n7734) );
  AND U10442 ( .A(n7735), .B(n7734), .Z(n7737) );
  NANDN U10443 ( .A(n8211), .B(ereg[119]), .Z(n7736) );
  NAND U10444 ( .A(n7737), .B(n7736), .Z(n2194) );
  NAND U10445 ( .A(n8206), .B(ereg[117]), .Z(n7739) );
  NANDN U10446 ( .A(init), .B(e[118]), .Z(n7738) );
  AND U10447 ( .A(n7739), .B(n7738), .Z(n7741) );
  NANDN U10448 ( .A(n8211), .B(ereg[118]), .Z(n7740) );
  NAND U10449 ( .A(n7741), .B(n7740), .Z(n2195) );
  NAND U10450 ( .A(n8206), .B(ereg[116]), .Z(n7743) );
  NANDN U10451 ( .A(init), .B(e[117]), .Z(n7742) );
  AND U10452 ( .A(n7743), .B(n7742), .Z(n7745) );
  NANDN U10453 ( .A(n8211), .B(ereg[117]), .Z(n7744) );
  NAND U10454 ( .A(n7745), .B(n7744), .Z(n2196) );
  NAND U10455 ( .A(n8206), .B(ereg[115]), .Z(n7747) );
  NANDN U10456 ( .A(init), .B(e[116]), .Z(n7746) );
  AND U10457 ( .A(n7747), .B(n7746), .Z(n7749) );
  NANDN U10458 ( .A(n8211), .B(ereg[116]), .Z(n7748) );
  NAND U10459 ( .A(n7749), .B(n7748), .Z(n2197) );
  NAND U10460 ( .A(n8206), .B(ereg[114]), .Z(n7751) );
  NANDN U10461 ( .A(init), .B(e[115]), .Z(n7750) );
  AND U10462 ( .A(n7751), .B(n7750), .Z(n7753) );
  NANDN U10463 ( .A(n8211), .B(ereg[115]), .Z(n7752) );
  NAND U10464 ( .A(n7753), .B(n7752), .Z(n2198) );
  NAND U10465 ( .A(n8206), .B(ereg[113]), .Z(n7755) );
  NANDN U10466 ( .A(init), .B(e[114]), .Z(n7754) );
  AND U10467 ( .A(n7755), .B(n7754), .Z(n7757) );
  NANDN U10468 ( .A(n8211), .B(ereg[114]), .Z(n7756) );
  NAND U10469 ( .A(n7757), .B(n7756), .Z(n2199) );
  NAND U10470 ( .A(n8206), .B(ereg[112]), .Z(n7759) );
  NANDN U10471 ( .A(init), .B(e[113]), .Z(n7758) );
  AND U10472 ( .A(n7759), .B(n7758), .Z(n7761) );
  NANDN U10473 ( .A(n8211), .B(ereg[113]), .Z(n7760) );
  NAND U10474 ( .A(n7761), .B(n7760), .Z(n2200) );
  NAND U10475 ( .A(n8206), .B(ereg[111]), .Z(n7763) );
  NANDN U10476 ( .A(init), .B(e[112]), .Z(n7762) );
  AND U10477 ( .A(n7763), .B(n7762), .Z(n7765) );
  NANDN U10478 ( .A(n8211), .B(ereg[112]), .Z(n7764) );
  NAND U10479 ( .A(n7765), .B(n7764), .Z(n2201) );
  NAND U10480 ( .A(n8206), .B(ereg[110]), .Z(n7767) );
  NANDN U10481 ( .A(init), .B(e[111]), .Z(n7766) );
  AND U10482 ( .A(n7767), .B(n7766), .Z(n7769) );
  NANDN U10483 ( .A(n8211), .B(ereg[111]), .Z(n7768) );
  NAND U10484 ( .A(n7769), .B(n7768), .Z(n2202) );
  NAND U10485 ( .A(n8206), .B(ereg[109]), .Z(n7771) );
  NANDN U10486 ( .A(init), .B(e[110]), .Z(n7770) );
  AND U10487 ( .A(n7771), .B(n7770), .Z(n7773) );
  NANDN U10488 ( .A(n8211), .B(ereg[110]), .Z(n7772) );
  NAND U10489 ( .A(n7773), .B(n7772), .Z(n2203) );
  NAND U10490 ( .A(n8206), .B(ereg[108]), .Z(n7775) );
  NANDN U10491 ( .A(init), .B(e[109]), .Z(n7774) );
  AND U10492 ( .A(n7775), .B(n7774), .Z(n7777) );
  NANDN U10493 ( .A(n8211), .B(ereg[109]), .Z(n7776) );
  NAND U10494 ( .A(n7777), .B(n7776), .Z(n2204) );
  NAND U10495 ( .A(n8206), .B(ereg[107]), .Z(n7779) );
  NANDN U10496 ( .A(init), .B(e[108]), .Z(n7778) );
  AND U10497 ( .A(n7779), .B(n7778), .Z(n7781) );
  NANDN U10498 ( .A(n8211), .B(ereg[108]), .Z(n7780) );
  NAND U10499 ( .A(n7781), .B(n7780), .Z(n2205) );
  NAND U10500 ( .A(n8206), .B(ereg[106]), .Z(n7783) );
  NANDN U10501 ( .A(init), .B(e[107]), .Z(n7782) );
  AND U10502 ( .A(n7783), .B(n7782), .Z(n7785) );
  NANDN U10503 ( .A(n8211), .B(ereg[107]), .Z(n7784) );
  NAND U10504 ( .A(n7785), .B(n7784), .Z(n2206) );
  NAND U10505 ( .A(n8206), .B(ereg[105]), .Z(n7787) );
  NANDN U10506 ( .A(init), .B(e[106]), .Z(n7786) );
  AND U10507 ( .A(n7787), .B(n7786), .Z(n7789) );
  NANDN U10508 ( .A(n8211), .B(ereg[106]), .Z(n7788) );
  NAND U10509 ( .A(n7789), .B(n7788), .Z(n2207) );
  NAND U10510 ( .A(n8206), .B(ereg[104]), .Z(n7791) );
  NANDN U10511 ( .A(init), .B(e[105]), .Z(n7790) );
  AND U10512 ( .A(n7791), .B(n7790), .Z(n7793) );
  NANDN U10513 ( .A(n8211), .B(ereg[105]), .Z(n7792) );
  NAND U10514 ( .A(n7793), .B(n7792), .Z(n2208) );
  NAND U10515 ( .A(n8206), .B(ereg[103]), .Z(n7795) );
  NANDN U10516 ( .A(init), .B(e[104]), .Z(n7794) );
  AND U10517 ( .A(n7795), .B(n7794), .Z(n7797) );
  NANDN U10518 ( .A(n8211), .B(ereg[104]), .Z(n7796) );
  NAND U10519 ( .A(n7797), .B(n7796), .Z(n2209) );
  NAND U10520 ( .A(n8206), .B(ereg[102]), .Z(n7799) );
  NANDN U10521 ( .A(init), .B(e[103]), .Z(n7798) );
  AND U10522 ( .A(n7799), .B(n7798), .Z(n7801) );
  NANDN U10523 ( .A(n8211), .B(ereg[103]), .Z(n7800) );
  NAND U10524 ( .A(n7801), .B(n7800), .Z(n2210) );
  NAND U10525 ( .A(n8206), .B(ereg[101]), .Z(n7803) );
  NANDN U10526 ( .A(init), .B(e[102]), .Z(n7802) );
  AND U10527 ( .A(n7803), .B(n7802), .Z(n7805) );
  NANDN U10528 ( .A(n8211), .B(ereg[102]), .Z(n7804) );
  NAND U10529 ( .A(n7805), .B(n7804), .Z(n2211) );
  NAND U10530 ( .A(n8206), .B(ereg[100]), .Z(n7807) );
  NANDN U10531 ( .A(init), .B(e[101]), .Z(n7806) );
  AND U10532 ( .A(n7807), .B(n7806), .Z(n7809) );
  NANDN U10533 ( .A(n8211), .B(ereg[101]), .Z(n7808) );
  NAND U10534 ( .A(n7809), .B(n7808), .Z(n2212) );
  NAND U10535 ( .A(n8206), .B(ereg[99]), .Z(n7811) );
  NANDN U10536 ( .A(init), .B(e[100]), .Z(n7810) );
  AND U10537 ( .A(n7811), .B(n7810), .Z(n7813) );
  NANDN U10538 ( .A(n8211), .B(ereg[100]), .Z(n7812) );
  NAND U10539 ( .A(n7813), .B(n7812), .Z(n2213) );
  NAND U10540 ( .A(n8206), .B(ereg[98]), .Z(n7815) );
  NANDN U10541 ( .A(init), .B(e[99]), .Z(n7814) );
  AND U10542 ( .A(n7815), .B(n7814), .Z(n7817) );
  NANDN U10543 ( .A(n8211), .B(ereg[99]), .Z(n7816) );
  NAND U10544 ( .A(n7817), .B(n7816), .Z(n2214) );
  NAND U10545 ( .A(n8206), .B(ereg[97]), .Z(n7819) );
  NANDN U10546 ( .A(init), .B(e[98]), .Z(n7818) );
  AND U10547 ( .A(n7819), .B(n7818), .Z(n7821) );
  NANDN U10548 ( .A(n8211), .B(ereg[98]), .Z(n7820) );
  NAND U10549 ( .A(n7821), .B(n7820), .Z(n2215) );
  NAND U10550 ( .A(n8206), .B(ereg[96]), .Z(n7823) );
  NANDN U10551 ( .A(init), .B(e[97]), .Z(n7822) );
  AND U10552 ( .A(n7823), .B(n7822), .Z(n7825) );
  NANDN U10553 ( .A(n8211), .B(ereg[97]), .Z(n7824) );
  NAND U10554 ( .A(n7825), .B(n7824), .Z(n2216) );
  NAND U10555 ( .A(n8206), .B(ereg[95]), .Z(n7827) );
  NANDN U10556 ( .A(init), .B(e[96]), .Z(n7826) );
  AND U10557 ( .A(n7827), .B(n7826), .Z(n7829) );
  NANDN U10558 ( .A(n8211), .B(ereg[96]), .Z(n7828) );
  NAND U10559 ( .A(n7829), .B(n7828), .Z(n2217) );
  NAND U10560 ( .A(n8206), .B(ereg[94]), .Z(n7831) );
  NANDN U10561 ( .A(init), .B(e[95]), .Z(n7830) );
  AND U10562 ( .A(n7831), .B(n7830), .Z(n7833) );
  NANDN U10563 ( .A(n8211), .B(ereg[95]), .Z(n7832) );
  NAND U10564 ( .A(n7833), .B(n7832), .Z(n2218) );
  NAND U10565 ( .A(n8206), .B(ereg[93]), .Z(n7835) );
  NANDN U10566 ( .A(init), .B(e[94]), .Z(n7834) );
  AND U10567 ( .A(n7835), .B(n7834), .Z(n7837) );
  NANDN U10568 ( .A(n8211), .B(ereg[94]), .Z(n7836) );
  NAND U10569 ( .A(n7837), .B(n7836), .Z(n2219) );
  NAND U10570 ( .A(n8206), .B(ereg[92]), .Z(n7839) );
  NANDN U10571 ( .A(init), .B(e[93]), .Z(n7838) );
  AND U10572 ( .A(n7839), .B(n7838), .Z(n7841) );
  NANDN U10573 ( .A(n8211), .B(ereg[93]), .Z(n7840) );
  NAND U10574 ( .A(n7841), .B(n7840), .Z(n2220) );
  NAND U10575 ( .A(n8206), .B(ereg[91]), .Z(n7843) );
  NANDN U10576 ( .A(init), .B(e[92]), .Z(n7842) );
  AND U10577 ( .A(n7843), .B(n7842), .Z(n7845) );
  NANDN U10578 ( .A(n8211), .B(ereg[92]), .Z(n7844) );
  NAND U10579 ( .A(n7845), .B(n7844), .Z(n2221) );
  NAND U10580 ( .A(n8206), .B(ereg[90]), .Z(n7847) );
  NANDN U10581 ( .A(init), .B(e[91]), .Z(n7846) );
  AND U10582 ( .A(n7847), .B(n7846), .Z(n7849) );
  NANDN U10583 ( .A(n8211), .B(ereg[91]), .Z(n7848) );
  NAND U10584 ( .A(n7849), .B(n7848), .Z(n2222) );
  NAND U10585 ( .A(n8206), .B(ereg[89]), .Z(n7851) );
  NANDN U10586 ( .A(init), .B(e[90]), .Z(n7850) );
  AND U10587 ( .A(n7851), .B(n7850), .Z(n7853) );
  NANDN U10588 ( .A(n8211), .B(ereg[90]), .Z(n7852) );
  NAND U10589 ( .A(n7853), .B(n7852), .Z(n2223) );
  NAND U10590 ( .A(n8206), .B(ereg[88]), .Z(n7855) );
  NANDN U10591 ( .A(init), .B(e[89]), .Z(n7854) );
  AND U10592 ( .A(n7855), .B(n7854), .Z(n7857) );
  NANDN U10593 ( .A(n8211), .B(ereg[89]), .Z(n7856) );
  NAND U10594 ( .A(n7857), .B(n7856), .Z(n2224) );
  NAND U10595 ( .A(n8206), .B(ereg[87]), .Z(n7859) );
  NANDN U10596 ( .A(init), .B(e[88]), .Z(n7858) );
  AND U10597 ( .A(n7859), .B(n7858), .Z(n7861) );
  NANDN U10598 ( .A(n8211), .B(ereg[88]), .Z(n7860) );
  NAND U10599 ( .A(n7861), .B(n7860), .Z(n2225) );
  NAND U10600 ( .A(n8206), .B(ereg[86]), .Z(n7863) );
  NANDN U10601 ( .A(init), .B(e[87]), .Z(n7862) );
  AND U10602 ( .A(n7863), .B(n7862), .Z(n7865) );
  NANDN U10603 ( .A(n8211), .B(ereg[87]), .Z(n7864) );
  NAND U10604 ( .A(n7865), .B(n7864), .Z(n2226) );
  NAND U10605 ( .A(n8206), .B(ereg[85]), .Z(n7867) );
  NANDN U10606 ( .A(init), .B(e[86]), .Z(n7866) );
  AND U10607 ( .A(n7867), .B(n7866), .Z(n7869) );
  NANDN U10608 ( .A(n8211), .B(ereg[86]), .Z(n7868) );
  NAND U10609 ( .A(n7869), .B(n7868), .Z(n2227) );
  NAND U10610 ( .A(n8206), .B(ereg[84]), .Z(n7871) );
  NANDN U10611 ( .A(init), .B(e[85]), .Z(n7870) );
  AND U10612 ( .A(n7871), .B(n7870), .Z(n7873) );
  NANDN U10613 ( .A(n8211), .B(ereg[85]), .Z(n7872) );
  NAND U10614 ( .A(n7873), .B(n7872), .Z(n2228) );
  NAND U10615 ( .A(n8206), .B(ereg[83]), .Z(n7875) );
  NANDN U10616 ( .A(init), .B(e[84]), .Z(n7874) );
  AND U10617 ( .A(n7875), .B(n7874), .Z(n7877) );
  NANDN U10618 ( .A(n8211), .B(ereg[84]), .Z(n7876) );
  NAND U10619 ( .A(n7877), .B(n7876), .Z(n2229) );
  NAND U10620 ( .A(n8206), .B(ereg[82]), .Z(n7879) );
  NANDN U10621 ( .A(init), .B(e[83]), .Z(n7878) );
  AND U10622 ( .A(n7879), .B(n7878), .Z(n7881) );
  NANDN U10623 ( .A(n8211), .B(ereg[83]), .Z(n7880) );
  NAND U10624 ( .A(n7881), .B(n7880), .Z(n2230) );
  NAND U10625 ( .A(n8206), .B(ereg[81]), .Z(n7883) );
  NANDN U10626 ( .A(init), .B(e[82]), .Z(n7882) );
  AND U10627 ( .A(n7883), .B(n7882), .Z(n7885) );
  NANDN U10628 ( .A(n8211), .B(ereg[82]), .Z(n7884) );
  NAND U10629 ( .A(n7885), .B(n7884), .Z(n2231) );
  NAND U10630 ( .A(n8206), .B(ereg[80]), .Z(n7887) );
  NANDN U10631 ( .A(init), .B(e[81]), .Z(n7886) );
  AND U10632 ( .A(n7887), .B(n7886), .Z(n7889) );
  NANDN U10633 ( .A(n8211), .B(ereg[81]), .Z(n7888) );
  NAND U10634 ( .A(n7889), .B(n7888), .Z(n2232) );
  NAND U10635 ( .A(n8206), .B(ereg[79]), .Z(n7891) );
  NANDN U10636 ( .A(init), .B(e[80]), .Z(n7890) );
  AND U10637 ( .A(n7891), .B(n7890), .Z(n7893) );
  NANDN U10638 ( .A(n8211), .B(ereg[80]), .Z(n7892) );
  NAND U10639 ( .A(n7893), .B(n7892), .Z(n2233) );
  NAND U10640 ( .A(n8206), .B(ereg[78]), .Z(n7895) );
  NANDN U10641 ( .A(init), .B(e[79]), .Z(n7894) );
  AND U10642 ( .A(n7895), .B(n7894), .Z(n7897) );
  NANDN U10643 ( .A(n8211), .B(ereg[79]), .Z(n7896) );
  NAND U10644 ( .A(n7897), .B(n7896), .Z(n2234) );
  NAND U10645 ( .A(n8206), .B(ereg[77]), .Z(n7899) );
  NANDN U10646 ( .A(init), .B(e[78]), .Z(n7898) );
  AND U10647 ( .A(n7899), .B(n7898), .Z(n7901) );
  NANDN U10648 ( .A(n8211), .B(ereg[78]), .Z(n7900) );
  NAND U10649 ( .A(n7901), .B(n7900), .Z(n2235) );
  NAND U10650 ( .A(n8206), .B(ereg[76]), .Z(n7903) );
  NANDN U10651 ( .A(init), .B(e[77]), .Z(n7902) );
  AND U10652 ( .A(n7903), .B(n7902), .Z(n7905) );
  NANDN U10653 ( .A(n8211), .B(ereg[77]), .Z(n7904) );
  NAND U10654 ( .A(n7905), .B(n7904), .Z(n2236) );
  NAND U10655 ( .A(n8206), .B(ereg[75]), .Z(n7907) );
  NANDN U10656 ( .A(init), .B(e[76]), .Z(n7906) );
  AND U10657 ( .A(n7907), .B(n7906), .Z(n7909) );
  NANDN U10658 ( .A(n8211), .B(ereg[76]), .Z(n7908) );
  NAND U10659 ( .A(n7909), .B(n7908), .Z(n2237) );
  NAND U10660 ( .A(n8206), .B(ereg[74]), .Z(n7911) );
  NANDN U10661 ( .A(init), .B(e[75]), .Z(n7910) );
  AND U10662 ( .A(n7911), .B(n7910), .Z(n7913) );
  NANDN U10663 ( .A(n8211), .B(ereg[75]), .Z(n7912) );
  NAND U10664 ( .A(n7913), .B(n7912), .Z(n2238) );
  NAND U10665 ( .A(n8206), .B(ereg[73]), .Z(n7915) );
  NANDN U10666 ( .A(init), .B(e[74]), .Z(n7914) );
  AND U10667 ( .A(n7915), .B(n7914), .Z(n7917) );
  NANDN U10668 ( .A(n8211), .B(ereg[74]), .Z(n7916) );
  NAND U10669 ( .A(n7917), .B(n7916), .Z(n2239) );
  NAND U10670 ( .A(n8206), .B(ereg[72]), .Z(n7919) );
  NANDN U10671 ( .A(init), .B(e[73]), .Z(n7918) );
  AND U10672 ( .A(n7919), .B(n7918), .Z(n7921) );
  NANDN U10673 ( .A(n8211), .B(ereg[73]), .Z(n7920) );
  NAND U10674 ( .A(n7921), .B(n7920), .Z(n2240) );
  NAND U10675 ( .A(n8206), .B(ereg[71]), .Z(n7923) );
  NANDN U10676 ( .A(init), .B(e[72]), .Z(n7922) );
  AND U10677 ( .A(n7923), .B(n7922), .Z(n7925) );
  NANDN U10678 ( .A(n8211), .B(ereg[72]), .Z(n7924) );
  NAND U10679 ( .A(n7925), .B(n7924), .Z(n2241) );
  NAND U10680 ( .A(n8206), .B(ereg[70]), .Z(n7927) );
  NANDN U10681 ( .A(init), .B(e[71]), .Z(n7926) );
  AND U10682 ( .A(n7927), .B(n7926), .Z(n7929) );
  NANDN U10683 ( .A(n8211), .B(ereg[71]), .Z(n7928) );
  NAND U10684 ( .A(n7929), .B(n7928), .Z(n2242) );
  NAND U10685 ( .A(n8206), .B(ereg[69]), .Z(n7931) );
  NANDN U10686 ( .A(init), .B(e[70]), .Z(n7930) );
  AND U10687 ( .A(n7931), .B(n7930), .Z(n7933) );
  NANDN U10688 ( .A(n8211), .B(ereg[70]), .Z(n7932) );
  NAND U10689 ( .A(n7933), .B(n7932), .Z(n2243) );
  NAND U10690 ( .A(n8206), .B(ereg[68]), .Z(n7935) );
  NANDN U10691 ( .A(init), .B(e[69]), .Z(n7934) );
  AND U10692 ( .A(n7935), .B(n7934), .Z(n7937) );
  NANDN U10693 ( .A(n8211), .B(ereg[69]), .Z(n7936) );
  NAND U10694 ( .A(n7937), .B(n7936), .Z(n2244) );
  NAND U10695 ( .A(n8206), .B(ereg[67]), .Z(n7939) );
  NANDN U10696 ( .A(init), .B(e[68]), .Z(n7938) );
  AND U10697 ( .A(n7939), .B(n7938), .Z(n7941) );
  NANDN U10698 ( .A(n8211), .B(ereg[68]), .Z(n7940) );
  NAND U10699 ( .A(n7941), .B(n7940), .Z(n2245) );
  NAND U10700 ( .A(n8206), .B(ereg[66]), .Z(n7943) );
  NANDN U10701 ( .A(init), .B(e[67]), .Z(n7942) );
  AND U10702 ( .A(n7943), .B(n7942), .Z(n7945) );
  NANDN U10703 ( .A(n8211), .B(ereg[67]), .Z(n7944) );
  NAND U10704 ( .A(n7945), .B(n7944), .Z(n2246) );
  NAND U10705 ( .A(n8206), .B(ereg[65]), .Z(n7947) );
  NANDN U10706 ( .A(init), .B(e[66]), .Z(n7946) );
  AND U10707 ( .A(n7947), .B(n7946), .Z(n7949) );
  NANDN U10708 ( .A(n8211), .B(ereg[66]), .Z(n7948) );
  NAND U10709 ( .A(n7949), .B(n7948), .Z(n2247) );
  NAND U10710 ( .A(n8206), .B(ereg[64]), .Z(n7951) );
  NANDN U10711 ( .A(init), .B(e[65]), .Z(n7950) );
  AND U10712 ( .A(n7951), .B(n7950), .Z(n7953) );
  NANDN U10713 ( .A(n8211), .B(ereg[65]), .Z(n7952) );
  NAND U10714 ( .A(n7953), .B(n7952), .Z(n2248) );
  NAND U10715 ( .A(n8206), .B(ereg[63]), .Z(n7955) );
  NANDN U10716 ( .A(init), .B(e[64]), .Z(n7954) );
  AND U10717 ( .A(n7955), .B(n7954), .Z(n7957) );
  NANDN U10718 ( .A(n8211), .B(ereg[64]), .Z(n7956) );
  NAND U10719 ( .A(n7957), .B(n7956), .Z(n2249) );
  NAND U10720 ( .A(n8206), .B(ereg[62]), .Z(n7959) );
  NANDN U10721 ( .A(init), .B(e[63]), .Z(n7958) );
  AND U10722 ( .A(n7959), .B(n7958), .Z(n7961) );
  NANDN U10723 ( .A(n8211), .B(ereg[63]), .Z(n7960) );
  NAND U10724 ( .A(n7961), .B(n7960), .Z(n2250) );
  NAND U10725 ( .A(n8206), .B(ereg[61]), .Z(n7963) );
  NANDN U10726 ( .A(init), .B(e[62]), .Z(n7962) );
  AND U10727 ( .A(n7963), .B(n7962), .Z(n7965) );
  NANDN U10728 ( .A(n8211), .B(ereg[62]), .Z(n7964) );
  NAND U10729 ( .A(n7965), .B(n7964), .Z(n2251) );
  NAND U10730 ( .A(n8206), .B(ereg[60]), .Z(n7967) );
  NANDN U10731 ( .A(init), .B(e[61]), .Z(n7966) );
  AND U10732 ( .A(n7967), .B(n7966), .Z(n7969) );
  NANDN U10733 ( .A(n8211), .B(ereg[61]), .Z(n7968) );
  NAND U10734 ( .A(n7969), .B(n7968), .Z(n2252) );
  NAND U10735 ( .A(n8206), .B(ereg[59]), .Z(n7971) );
  NANDN U10736 ( .A(init), .B(e[60]), .Z(n7970) );
  AND U10737 ( .A(n7971), .B(n7970), .Z(n7973) );
  NANDN U10738 ( .A(n8211), .B(ereg[60]), .Z(n7972) );
  NAND U10739 ( .A(n7973), .B(n7972), .Z(n2253) );
  NAND U10740 ( .A(n8206), .B(ereg[58]), .Z(n7975) );
  NANDN U10741 ( .A(init), .B(e[59]), .Z(n7974) );
  AND U10742 ( .A(n7975), .B(n7974), .Z(n7977) );
  NANDN U10743 ( .A(n8211), .B(ereg[59]), .Z(n7976) );
  NAND U10744 ( .A(n7977), .B(n7976), .Z(n2254) );
  NAND U10745 ( .A(n8206), .B(ereg[57]), .Z(n7979) );
  NANDN U10746 ( .A(init), .B(e[58]), .Z(n7978) );
  AND U10747 ( .A(n7979), .B(n7978), .Z(n7981) );
  NANDN U10748 ( .A(n8211), .B(ereg[58]), .Z(n7980) );
  NAND U10749 ( .A(n7981), .B(n7980), .Z(n2255) );
  NAND U10750 ( .A(n8206), .B(ereg[56]), .Z(n7983) );
  NANDN U10751 ( .A(init), .B(e[57]), .Z(n7982) );
  AND U10752 ( .A(n7983), .B(n7982), .Z(n7985) );
  NANDN U10753 ( .A(n8211), .B(ereg[57]), .Z(n7984) );
  NAND U10754 ( .A(n7985), .B(n7984), .Z(n2256) );
  NAND U10755 ( .A(n8206), .B(ereg[55]), .Z(n7987) );
  NANDN U10756 ( .A(init), .B(e[56]), .Z(n7986) );
  AND U10757 ( .A(n7987), .B(n7986), .Z(n7989) );
  NANDN U10758 ( .A(n8211), .B(ereg[56]), .Z(n7988) );
  NAND U10759 ( .A(n7989), .B(n7988), .Z(n2257) );
  NAND U10760 ( .A(n8206), .B(ereg[54]), .Z(n7991) );
  NANDN U10761 ( .A(init), .B(e[55]), .Z(n7990) );
  AND U10762 ( .A(n7991), .B(n7990), .Z(n7993) );
  NANDN U10763 ( .A(n8211), .B(ereg[55]), .Z(n7992) );
  NAND U10764 ( .A(n7993), .B(n7992), .Z(n2258) );
  NAND U10765 ( .A(n8206), .B(ereg[53]), .Z(n7995) );
  NANDN U10766 ( .A(init), .B(e[54]), .Z(n7994) );
  AND U10767 ( .A(n7995), .B(n7994), .Z(n7997) );
  NANDN U10768 ( .A(n8211), .B(ereg[54]), .Z(n7996) );
  NAND U10769 ( .A(n7997), .B(n7996), .Z(n2259) );
  NAND U10770 ( .A(n8206), .B(ereg[52]), .Z(n7999) );
  NANDN U10771 ( .A(init), .B(e[53]), .Z(n7998) );
  AND U10772 ( .A(n7999), .B(n7998), .Z(n8001) );
  NANDN U10773 ( .A(n8211), .B(ereg[53]), .Z(n8000) );
  NAND U10774 ( .A(n8001), .B(n8000), .Z(n2260) );
  NAND U10775 ( .A(n8206), .B(ereg[51]), .Z(n8003) );
  NANDN U10776 ( .A(init), .B(e[52]), .Z(n8002) );
  AND U10777 ( .A(n8003), .B(n8002), .Z(n8005) );
  NANDN U10778 ( .A(n8211), .B(ereg[52]), .Z(n8004) );
  NAND U10779 ( .A(n8005), .B(n8004), .Z(n2261) );
  NAND U10780 ( .A(n8206), .B(ereg[50]), .Z(n8007) );
  NANDN U10781 ( .A(init), .B(e[51]), .Z(n8006) );
  AND U10782 ( .A(n8007), .B(n8006), .Z(n8009) );
  NANDN U10783 ( .A(n8211), .B(ereg[51]), .Z(n8008) );
  NAND U10784 ( .A(n8009), .B(n8008), .Z(n2262) );
  NAND U10785 ( .A(n8206), .B(ereg[49]), .Z(n8011) );
  NANDN U10786 ( .A(init), .B(e[50]), .Z(n8010) );
  AND U10787 ( .A(n8011), .B(n8010), .Z(n8013) );
  NANDN U10788 ( .A(n8211), .B(ereg[50]), .Z(n8012) );
  NAND U10789 ( .A(n8013), .B(n8012), .Z(n2263) );
  NAND U10790 ( .A(n8206), .B(ereg[48]), .Z(n8015) );
  NANDN U10791 ( .A(init), .B(e[49]), .Z(n8014) );
  AND U10792 ( .A(n8015), .B(n8014), .Z(n8017) );
  NANDN U10793 ( .A(n8211), .B(ereg[49]), .Z(n8016) );
  NAND U10794 ( .A(n8017), .B(n8016), .Z(n2264) );
  NAND U10795 ( .A(n8206), .B(ereg[47]), .Z(n8019) );
  NANDN U10796 ( .A(init), .B(e[48]), .Z(n8018) );
  AND U10797 ( .A(n8019), .B(n8018), .Z(n8021) );
  NANDN U10798 ( .A(n8211), .B(ereg[48]), .Z(n8020) );
  NAND U10799 ( .A(n8021), .B(n8020), .Z(n2265) );
  NAND U10800 ( .A(n8206), .B(ereg[46]), .Z(n8023) );
  NANDN U10801 ( .A(init), .B(e[47]), .Z(n8022) );
  AND U10802 ( .A(n8023), .B(n8022), .Z(n8025) );
  NANDN U10803 ( .A(n8211), .B(ereg[47]), .Z(n8024) );
  NAND U10804 ( .A(n8025), .B(n8024), .Z(n2266) );
  NAND U10805 ( .A(n8206), .B(ereg[45]), .Z(n8027) );
  NANDN U10806 ( .A(init), .B(e[46]), .Z(n8026) );
  AND U10807 ( .A(n8027), .B(n8026), .Z(n8029) );
  NANDN U10808 ( .A(n8211), .B(ereg[46]), .Z(n8028) );
  NAND U10809 ( .A(n8029), .B(n8028), .Z(n2267) );
  NAND U10810 ( .A(n8206), .B(ereg[44]), .Z(n8031) );
  NANDN U10811 ( .A(init), .B(e[45]), .Z(n8030) );
  AND U10812 ( .A(n8031), .B(n8030), .Z(n8033) );
  NANDN U10813 ( .A(n8211), .B(ereg[45]), .Z(n8032) );
  NAND U10814 ( .A(n8033), .B(n8032), .Z(n2268) );
  NAND U10815 ( .A(n8206), .B(ereg[43]), .Z(n8035) );
  NANDN U10816 ( .A(init), .B(e[44]), .Z(n8034) );
  AND U10817 ( .A(n8035), .B(n8034), .Z(n8037) );
  NANDN U10818 ( .A(n8211), .B(ereg[44]), .Z(n8036) );
  NAND U10819 ( .A(n8037), .B(n8036), .Z(n2269) );
  NAND U10820 ( .A(n8206), .B(ereg[42]), .Z(n8039) );
  NANDN U10821 ( .A(init), .B(e[43]), .Z(n8038) );
  AND U10822 ( .A(n8039), .B(n8038), .Z(n8041) );
  NANDN U10823 ( .A(n8211), .B(ereg[43]), .Z(n8040) );
  NAND U10824 ( .A(n8041), .B(n8040), .Z(n2270) );
  NAND U10825 ( .A(n8206), .B(ereg[41]), .Z(n8043) );
  NANDN U10826 ( .A(init), .B(e[42]), .Z(n8042) );
  AND U10827 ( .A(n8043), .B(n8042), .Z(n8045) );
  NANDN U10828 ( .A(n8211), .B(ereg[42]), .Z(n8044) );
  NAND U10829 ( .A(n8045), .B(n8044), .Z(n2271) );
  NAND U10830 ( .A(n8206), .B(ereg[40]), .Z(n8047) );
  NANDN U10831 ( .A(init), .B(e[41]), .Z(n8046) );
  AND U10832 ( .A(n8047), .B(n8046), .Z(n8049) );
  NANDN U10833 ( .A(n8211), .B(ereg[41]), .Z(n8048) );
  NAND U10834 ( .A(n8049), .B(n8048), .Z(n2272) );
  NAND U10835 ( .A(n8206), .B(ereg[39]), .Z(n8051) );
  NANDN U10836 ( .A(init), .B(e[40]), .Z(n8050) );
  AND U10837 ( .A(n8051), .B(n8050), .Z(n8053) );
  NANDN U10838 ( .A(n8211), .B(ereg[40]), .Z(n8052) );
  NAND U10839 ( .A(n8053), .B(n8052), .Z(n2273) );
  NAND U10840 ( .A(n8206), .B(ereg[38]), .Z(n8055) );
  NANDN U10841 ( .A(init), .B(e[39]), .Z(n8054) );
  AND U10842 ( .A(n8055), .B(n8054), .Z(n8057) );
  NANDN U10843 ( .A(n8211), .B(ereg[39]), .Z(n8056) );
  NAND U10844 ( .A(n8057), .B(n8056), .Z(n2274) );
  NAND U10845 ( .A(n8206), .B(ereg[37]), .Z(n8059) );
  NANDN U10846 ( .A(init), .B(e[38]), .Z(n8058) );
  AND U10847 ( .A(n8059), .B(n8058), .Z(n8061) );
  NANDN U10848 ( .A(n8211), .B(ereg[38]), .Z(n8060) );
  NAND U10849 ( .A(n8061), .B(n8060), .Z(n2275) );
  NAND U10850 ( .A(n8206), .B(ereg[36]), .Z(n8063) );
  NANDN U10851 ( .A(init), .B(e[37]), .Z(n8062) );
  AND U10852 ( .A(n8063), .B(n8062), .Z(n8065) );
  NANDN U10853 ( .A(n8211), .B(ereg[37]), .Z(n8064) );
  NAND U10854 ( .A(n8065), .B(n8064), .Z(n2276) );
  NAND U10855 ( .A(n8206), .B(ereg[35]), .Z(n8067) );
  NANDN U10856 ( .A(init), .B(e[36]), .Z(n8066) );
  AND U10857 ( .A(n8067), .B(n8066), .Z(n8069) );
  NANDN U10858 ( .A(n8211), .B(ereg[36]), .Z(n8068) );
  NAND U10859 ( .A(n8069), .B(n8068), .Z(n2277) );
  NAND U10860 ( .A(n8206), .B(ereg[34]), .Z(n8071) );
  NANDN U10861 ( .A(init), .B(e[35]), .Z(n8070) );
  AND U10862 ( .A(n8071), .B(n8070), .Z(n8073) );
  NANDN U10863 ( .A(n8211), .B(ereg[35]), .Z(n8072) );
  NAND U10864 ( .A(n8073), .B(n8072), .Z(n2278) );
  NAND U10865 ( .A(n8206), .B(ereg[33]), .Z(n8075) );
  NANDN U10866 ( .A(init), .B(e[34]), .Z(n8074) );
  AND U10867 ( .A(n8075), .B(n8074), .Z(n8077) );
  NANDN U10868 ( .A(n8211), .B(ereg[34]), .Z(n8076) );
  NAND U10869 ( .A(n8077), .B(n8076), .Z(n2279) );
  NAND U10870 ( .A(n8206), .B(ereg[32]), .Z(n8079) );
  NANDN U10871 ( .A(init), .B(e[33]), .Z(n8078) );
  AND U10872 ( .A(n8079), .B(n8078), .Z(n8081) );
  NANDN U10873 ( .A(n8211), .B(ereg[33]), .Z(n8080) );
  NAND U10874 ( .A(n8081), .B(n8080), .Z(n2280) );
  NAND U10875 ( .A(n8206), .B(ereg[31]), .Z(n8083) );
  NANDN U10876 ( .A(init), .B(e[32]), .Z(n8082) );
  AND U10877 ( .A(n8083), .B(n8082), .Z(n8085) );
  NANDN U10878 ( .A(n8211), .B(ereg[32]), .Z(n8084) );
  NAND U10879 ( .A(n8085), .B(n8084), .Z(n2281) );
  NAND U10880 ( .A(n8206), .B(ereg[30]), .Z(n8087) );
  NANDN U10881 ( .A(init), .B(e[31]), .Z(n8086) );
  AND U10882 ( .A(n8087), .B(n8086), .Z(n8089) );
  NANDN U10883 ( .A(n8211), .B(ereg[31]), .Z(n8088) );
  NAND U10884 ( .A(n8089), .B(n8088), .Z(n2282) );
  NAND U10885 ( .A(n8206), .B(ereg[29]), .Z(n8091) );
  NANDN U10886 ( .A(init), .B(e[30]), .Z(n8090) );
  AND U10887 ( .A(n8091), .B(n8090), .Z(n8093) );
  NANDN U10888 ( .A(n8211), .B(ereg[30]), .Z(n8092) );
  NAND U10889 ( .A(n8093), .B(n8092), .Z(n2283) );
  NAND U10890 ( .A(n8206), .B(ereg[28]), .Z(n8095) );
  NANDN U10891 ( .A(init), .B(e[29]), .Z(n8094) );
  AND U10892 ( .A(n8095), .B(n8094), .Z(n8097) );
  NANDN U10893 ( .A(n8211), .B(ereg[29]), .Z(n8096) );
  NAND U10894 ( .A(n8097), .B(n8096), .Z(n2284) );
  NAND U10895 ( .A(n8206), .B(ereg[27]), .Z(n8099) );
  NANDN U10896 ( .A(init), .B(e[28]), .Z(n8098) );
  AND U10897 ( .A(n8099), .B(n8098), .Z(n8101) );
  NANDN U10898 ( .A(n8211), .B(ereg[28]), .Z(n8100) );
  NAND U10899 ( .A(n8101), .B(n8100), .Z(n2285) );
  NAND U10900 ( .A(n8206), .B(ereg[26]), .Z(n8103) );
  NANDN U10901 ( .A(init), .B(e[27]), .Z(n8102) );
  AND U10902 ( .A(n8103), .B(n8102), .Z(n8105) );
  NANDN U10903 ( .A(n8211), .B(ereg[27]), .Z(n8104) );
  NAND U10904 ( .A(n8105), .B(n8104), .Z(n2286) );
  NAND U10905 ( .A(n8206), .B(ereg[25]), .Z(n8107) );
  NANDN U10906 ( .A(init), .B(e[26]), .Z(n8106) );
  AND U10907 ( .A(n8107), .B(n8106), .Z(n8109) );
  NANDN U10908 ( .A(n8211), .B(ereg[26]), .Z(n8108) );
  NAND U10909 ( .A(n8109), .B(n8108), .Z(n2287) );
  NAND U10910 ( .A(n8206), .B(ereg[24]), .Z(n8111) );
  NANDN U10911 ( .A(init), .B(e[25]), .Z(n8110) );
  AND U10912 ( .A(n8111), .B(n8110), .Z(n8113) );
  NANDN U10913 ( .A(n8211), .B(ereg[25]), .Z(n8112) );
  NAND U10914 ( .A(n8113), .B(n8112), .Z(n2288) );
  NAND U10915 ( .A(n8206), .B(ereg[23]), .Z(n8115) );
  NANDN U10916 ( .A(init), .B(e[24]), .Z(n8114) );
  AND U10917 ( .A(n8115), .B(n8114), .Z(n8117) );
  NANDN U10918 ( .A(n8211), .B(ereg[24]), .Z(n8116) );
  NAND U10919 ( .A(n8117), .B(n8116), .Z(n2289) );
  NAND U10920 ( .A(n8206), .B(ereg[22]), .Z(n8119) );
  NANDN U10921 ( .A(init), .B(e[23]), .Z(n8118) );
  AND U10922 ( .A(n8119), .B(n8118), .Z(n8121) );
  NANDN U10923 ( .A(n8211), .B(ereg[23]), .Z(n8120) );
  NAND U10924 ( .A(n8121), .B(n8120), .Z(n2290) );
  NAND U10925 ( .A(n8206), .B(ereg[21]), .Z(n8123) );
  NANDN U10926 ( .A(init), .B(e[22]), .Z(n8122) );
  AND U10927 ( .A(n8123), .B(n8122), .Z(n8125) );
  NANDN U10928 ( .A(n8211), .B(ereg[22]), .Z(n8124) );
  NAND U10929 ( .A(n8125), .B(n8124), .Z(n2291) );
  NAND U10930 ( .A(n8206), .B(ereg[20]), .Z(n8127) );
  NANDN U10931 ( .A(init), .B(e[21]), .Z(n8126) );
  AND U10932 ( .A(n8127), .B(n8126), .Z(n8129) );
  NANDN U10933 ( .A(n8211), .B(ereg[21]), .Z(n8128) );
  NAND U10934 ( .A(n8129), .B(n8128), .Z(n2292) );
  NAND U10935 ( .A(n8206), .B(ereg[19]), .Z(n8131) );
  NANDN U10936 ( .A(init), .B(e[20]), .Z(n8130) );
  AND U10937 ( .A(n8131), .B(n8130), .Z(n8133) );
  NANDN U10938 ( .A(n8211), .B(ereg[20]), .Z(n8132) );
  NAND U10939 ( .A(n8133), .B(n8132), .Z(n2293) );
  NAND U10940 ( .A(n8206), .B(ereg[18]), .Z(n8135) );
  NANDN U10941 ( .A(init), .B(e[19]), .Z(n8134) );
  AND U10942 ( .A(n8135), .B(n8134), .Z(n8137) );
  NANDN U10943 ( .A(n8211), .B(ereg[19]), .Z(n8136) );
  NAND U10944 ( .A(n8137), .B(n8136), .Z(n2294) );
  NAND U10945 ( .A(n8206), .B(ereg[17]), .Z(n8139) );
  NANDN U10946 ( .A(init), .B(e[18]), .Z(n8138) );
  AND U10947 ( .A(n8139), .B(n8138), .Z(n8141) );
  NANDN U10948 ( .A(n8211), .B(ereg[18]), .Z(n8140) );
  NAND U10949 ( .A(n8141), .B(n8140), .Z(n2295) );
  NAND U10950 ( .A(n8206), .B(ereg[16]), .Z(n8143) );
  NANDN U10951 ( .A(init), .B(e[17]), .Z(n8142) );
  AND U10952 ( .A(n8143), .B(n8142), .Z(n8145) );
  NANDN U10953 ( .A(n8211), .B(ereg[17]), .Z(n8144) );
  NAND U10954 ( .A(n8145), .B(n8144), .Z(n2296) );
  NAND U10955 ( .A(n8206), .B(ereg[15]), .Z(n8147) );
  NANDN U10956 ( .A(init), .B(e[16]), .Z(n8146) );
  AND U10957 ( .A(n8147), .B(n8146), .Z(n8149) );
  NANDN U10958 ( .A(n8211), .B(ereg[16]), .Z(n8148) );
  NAND U10959 ( .A(n8149), .B(n8148), .Z(n2297) );
  NAND U10960 ( .A(n8206), .B(ereg[14]), .Z(n8151) );
  NANDN U10961 ( .A(init), .B(e[15]), .Z(n8150) );
  AND U10962 ( .A(n8151), .B(n8150), .Z(n8153) );
  NANDN U10963 ( .A(n8211), .B(ereg[15]), .Z(n8152) );
  NAND U10964 ( .A(n8153), .B(n8152), .Z(n2298) );
  NAND U10965 ( .A(n8206), .B(ereg[13]), .Z(n8155) );
  NANDN U10966 ( .A(init), .B(e[14]), .Z(n8154) );
  AND U10967 ( .A(n8155), .B(n8154), .Z(n8157) );
  NANDN U10968 ( .A(n8211), .B(ereg[14]), .Z(n8156) );
  NAND U10969 ( .A(n8157), .B(n8156), .Z(n2299) );
  NAND U10970 ( .A(n8206), .B(ereg[12]), .Z(n8159) );
  NANDN U10971 ( .A(init), .B(e[13]), .Z(n8158) );
  AND U10972 ( .A(n8159), .B(n8158), .Z(n8161) );
  NANDN U10973 ( .A(n8211), .B(ereg[13]), .Z(n8160) );
  NAND U10974 ( .A(n8161), .B(n8160), .Z(n2300) );
  NAND U10975 ( .A(n8206), .B(ereg[11]), .Z(n8163) );
  NANDN U10976 ( .A(init), .B(e[12]), .Z(n8162) );
  AND U10977 ( .A(n8163), .B(n8162), .Z(n8165) );
  NANDN U10978 ( .A(n8211), .B(ereg[12]), .Z(n8164) );
  NAND U10979 ( .A(n8165), .B(n8164), .Z(n2301) );
  NAND U10980 ( .A(n8206), .B(ereg[10]), .Z(n8167) );
  NANDN U10981 ( .A(init), .B(e[11]), .Z(n8166) );
  AND U10982 ( .A(n8167), .B(n8166), .Z(n8169) );
  NANDN U10983 ( .A(n8211), .B(ereg[11]), .Z(n8168) );
  NAND U10984 ( .A(n8169), .B(n8168), .Z(n2302) );
  NAND U10985 ( .A(n8206), .B(ereg[9]), .Z(n8171) );
  NANDN U10986 ( .A(init), .B(e[10]), .Z(n8170) );
  AND U10987 ( .A(n8171), .B(n8170), .Z(n8173) );
  NANDN U10988 ( .A(n8211), .B(ereg[10]), .Z(n8172) );
  NAND U10989 ( .A(n8173), .B(n8172), .Z(n2303) );
  NAND U10990 ( .A(n8206), .B(ereg[8]), .Z(n8175) );
  NANDN U10991 ( .A(init), .B(e[9]), .Z(n8174) );
  AND U10992 ( .A(n8175), .B(n8174), .Z(n8177) );
  NANDN U10993 ( .A(n8211), .B(ereg[9]), .Z(n8176) );
  NAND U10994 ( .A(n8177), .B(n8176), .Z(n2304) );
  NAND U10995 ( .A(n8206), .B(ereg[7]), .Z(n8179) );
  NANDN U10996 ( .A(init), .B(e[8]), .Z(n8178) );
  AND U10997 ( .A(n8179), .B(n8178), .Z(n8181) );
  NANDN U10998 ( .A(n8211), .B(ereg[8]), .Z(n8180) );
  NAND U10999 ( .A(n8181), .B(n8180), .Z(n2305) );
  NAND U11000 ( .A(n8206), .B(ereg[6]), .Z(n8183) );
  NANDN U11001 ( .A(init), .B(e[7]), .Z(n8182) );
  AND U11002 ( .A(n8183), .B(n8182), .Z(n8185) );
  NANDN U11003 ( .A(n8211), .B(ereg[7]), .Z(n8184) );
  NAND U11004 ( .A(n8185), .B(n8184), .Z(n2306) );
  NAND U11005 ( .A(n8206), .B(ereg[5]), .Z(n8187) );
  NANDN U11006 ( .A(init), .B(e[6]), .Z(n8186) );
  AND U11007 ( .A(n8187), .B(n8186), .Z(n8189) );
  NANDN U11008 ( .A(n8211), .B(ereg[6]), .Z(n8188) );
  NAND U11009 ( .A(n8189), .B(n8188), .Z(n2307) );
  NAND U11010 ( .A(n8206), .B(ereg[4]), .Z(n8191) );
  NANDN U11011 ( .A(init), .B(e[5]), .Z(n8190) );
  AND U11012 ( .A(n8191), .B(n8190), .Z(n8193) );
  NANDN U11013 ( .A(n8211), .B(ereg[5]), .Z(n8192) );
  NAND U11014 ( .A(n8193), .B(n8192), .Z(n2308) );
  NAND U11015 ( .A(n8206), .B(ereg[3]), .Z(n8195) );
  NANDN U11016 ( .A(init), .B(e[4]), .Z(n8194) );
  AND U11017 ( .A(n8195), .B(n8194), .Z(n8197) );
  NANDN U11018 ( .A(n8211), .B(ereg[4]), .Z(n8196) );
  NAND U11019 ( .A(n8197), .B(n8196), .Z(n2309) );
  NAND U11020 ( .A(n8206), .B(ereg[2]), .Z(n8199) );
  NANDN U11021 ( .A(init), .B(e[3]), .Z(n8198) );
  AND U11022 ( .A(n8199), .B(n8198), .Z(n8201) );
  NANDN U11023 ( .A(n8211), .B(ereg[3]), .Z(n8200) );
  NAND U11024 ( .A(n8201), .B(n8200), .Z(n2310) );
  NAND U11025 ( .A(n8206), .B(ereg[1]), .Z(n8203) );
  NANDN U11026 ( .A(init), .B(e[2]), .Z(n8202) );
  AND U11027 ( .A(n8203), .B(n8202), .Z(n8205) );
  NANDN U11028 ( .A(n8211), .B(ereg[2]), .Z(n8204) );
  NAND U11029 ( .A(n8205), .B(n8204), .Z(n2311) );
  NAND U11030 ( .A(n8206), .B(ereg[0]), .Z(n8208) );
  NANDN U11031 ( .A(init), .B(e[1]), .Z(n8207) );
  AND U11032 ( .A(n8208), .B(n8207), .Z(n8210) );
  NANDN U11033 ( .A(n8211), .B(ereg[1]), .Z(n8209) );
  NAND U11034 ( .A(n8210), .B(n8209), .Z(n2312) );
  NANDN U11035 ( .A(init), .B(e[0]), .Z(n8213) );
  NANDN U11036 ( .A(n8211), .B(ereg[0]), .Z(n8212) );
  NAND U11037 ( .A(n8213), .B(n8212), .Z(n2313) );
  XNOR U11038 ( .A(start_in[127]), .B(n8214), .Z(n2314) );
endmodule

