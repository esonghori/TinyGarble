
module matrixMult_N_M_1_N5_M32 ( clk, rst, x, y, o );
  input [159:0] x;
  input [799:0] y;
  output [159:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903;

  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  DFF \oi_reg[3][31]  ( .D(N256), .CLK(clk), .RST(rst), .Q(o[127]) );
  DFF \oi_reg[3][30]  ( .D(N255), .CLK(clk), .RST(rst), .Q(o[126]) );
  DFF \oi_reg[3][29]  ( .D(N254), .CLK(clk), .RST(rst), .Q(o[125]) );
  DFF \oi_reg[3][28]  ( .D(N253), .CLK(clk), .RST(rst), .Q(o[124]) );
  DFF \oi_reg[3][27]  ( .D(N252), .CLK(clk), .RST(rst), .Q(o[123]) );
  DFF \oi_reg[3][26]  ( .D(N251), .CLK(clk), .RST(rst), .Q(o[122]) );
  DFF \oi_reg[3][25]  ( .D(N250), .CLK(clk), .RST(rst), .Q(o[121]) );
  DFF \oi_reg[3][24]  ( .D(N249), .CLK(clk), .RST(rst), .Q(o[120]) );
  DFF \oi_reg[3][23]  ( .D(N248), .CLK(clk), .RST(rst), .Q(o[119]) );
  DFF \oi_reg[3][22]  ( .D(N247), .CLK(clk), .RST(rst), .Q(o[118]) );
  DFF \oi_reg[3][21]  ( .D(N246), .CLK(clk), .RST(rst), .Q(o[117]) );
  DFF \oi_reg[3][20]  ( .D(N245), .CLK(clk), .RST(rst), .Q(o[116]) );
  DFF \oi_reg[3][19]  ( .D(N244), .CLK(clk), .RST(rst), .Q(o[115]) );
  DFF \oi_reg[3][18]  ( .D(N243), .CLK(clk), .RST(rst), .Q(o[114]) );
  DFF \oi_reg[3][17]  ( .D(N242), .CLK(clk), .RST(rst), .Q(o[113]) );
  DFF \oi_reg[3][16]  ( .D(N241), .CLK(clk), .RST(rst), .Q(o[112]) );
  DFF \oi_reg[3][15]  ( .D(N240), .CLK(clk), .RST(rst), .Q(o[111]) );
  DFF \oi_reg[3][14]  ( .D(N239), .CLK(clk), .RST(rst), .Q(o[110]) );
  DFF \oi_reg[3][13]  ( .D(N238), .CLK(clk), .RST(rst), .Q(o[109]) );
  DFF \oi_reg[3][12]  ( .D(N237), .CLK(clk), .RST(rst), .Q(o[108]) );
  DFF \oi_reg[3][11]  ( .D(N236), .CLK(clk), .RST(rst), .Q(o[107]) );
  DFF \oi_reg[3][10]  ( .D(N235), .CLK(clk), .RST(rst), .Q(o[106]) );
  DFF \oi_reg[3][9]  ( .D(N234), .CLK(clk), .RST(rst), .Q(o[105]) );
  DFF \oi_reg[3][8]  ( .D(N233), .CLK(clk), .RST(rst), .Q(o[104]) );
  DFF \oi_reg[3][7]  ( .D(N232), .CLK(clk), .RST(rst), .Q(o[103]) );
  DFF \oi_reg[3][6]  ( .D(N231), .CLK(clk), .RST(rst), .Q(o[102]) );
  DFF \oi_reg[3][5]  ( .D(N230), .CLK(clk), .RST(rst), .Q(o[101]) );
  DFF \oi_reg[3][4]  ( .D(N229), .CLK(clk), .RST(rst), .Q(o[100]) );
  DFF \oi_reg[3][3]  ( .D(N228), .CLK(clk), .RST(rst), .Q(o[99]) );
  DFF \oi_reg[3][2]  ( .D(N227), .CLK(clk), .RST(rst), .Q(o[98]) );
  DFF \oi_reg[3][1]  ( .D(N226), .CLK(clk), .RST(rst), .Q(o[97]) );
  DFF \oi_reg[3][0]  ( .D(N225), .CLK(clk), .RST(rst), .Q(o[96]) );
  DFF \oi_reg[4][31]  ( .D(N320), .CLK(clk), .RST(rst), .Q(o[159]) );
  DFF \oi_reg[4][30]  ( .D(N319), .CLK(clk), .RST(rst), .Q(o[158]) );
  DFF \oi_reg[4][29]  ( .D(N318), .CLK(clk), .RST(rst), .Q(o[157]) );
  DFF \oi_reg[4][28]  ( .D(N317), .CLK(clk), .RST(rst), .Q(o[156]) );
  DFF \oi_reg[4][27]  ( .D(N316), .CLK(clk), .RST(rst), .Q(o[155]) );
  DFF \oi_reg[4][26]  ( .D(N315), .CLK(clk), .RST(rst), .Q(o[154]) );
  DFF \oi_reg[4][25]  ( .D(N314), .CLK(clk), .RST(rst), .Q(o[153]) );
  DFF \oi_reg[4][24]  ( .D(N313), .CLK(clk), .RST(rst), .Q(o[152]) );
  DFF \oi_reg[4][23]  ( .D(N312), .CLK(clk), .RST(rst), .Q(o[151]) );
  DFF \oi_reg[4][22]  ( .D(N311), .CLK(clk), .RST(rst), .Q(o[150]) );
  DFF \oi_reg[4][21]  ( .D(N310), .CLK(clk), .RST(rst), .Q(o[149]) );
  DFF \oi_reg[4][20]  ( .D(N309), .CLK(clk), .RST(rst), .Q(o[148]) );
  DFF \oi_reg[4][19]  ( .D(N308), .CLK(clk), .RST(rst), .Q(o[147]) );
  DFF \oi_reg[4][18]  ( .D(N307), .CLK(clk), .RST(rst), .Q(o[146]) );
  DFF \oi_reg[4][17]  ( .D(N306), .CLK(clk), .RST(rst), .Q(o[145]) );
  DFF \oi_reg[4][16]  ( .D(N305), .CLK(clk), .RST(rst), .Q(o[144]) );
  DFF \oi_reg[4][15]  ( .D(N304), .CLK(clk), .RST(rst), .Q(o[143]) );
  DFF \oi_reg[4][14]  ( .D(N303), .CLK(clk), .RST(rst), .Q(o[142]) );
  DFF \oi_reg[4][13]  ( .D(N302), .CLK(clk), .RST(rst), .Q(o[141]) );
  DFF \oi_reg[4][12]  ( .D(N301), .CLK(clk), .RST(rst), .Q(o[140]) );
  DFF \oi_reg[4][11]  ( .D(N300), .CLK(clk), .RST(rst), .Q(o[139]) );
  DFF \oi_reg[4][10]  ( .D(N299), .CLK(clk), .RST(rst), .Q(o[138]) );
  DFF \oi_reg[4][9]  ( .D(N298), .CLK(clk), .RST(rst), .Q(o[137]) );
  DFF \oi_reg[4][8]  ( .D(N297), .CLK(clk), .RST(rst), .Q(o[136]) );
  DFF \oi_reg[4][7]  ( .D(N296), .CLK(clk), .RST(rst), .Q(o[135]) );
  DFF \oi_reg[4][6]  ( .D(N295), .CLK(clk), .RST(rst), .Q(o[134]) );
  DFF \oi_reg[4][5]  ( .D(N294), .CLK(clk), .RST(rst), .Q(o[133]) );
  DFF \oi_reg[4][4]  ( .D(N293), .CLK(clk), .RST(rst), .Q(o[132]) );
  DFF \oi_reg[4][3]  ( .D(N292), .CLK(clk), .RST(rst), .Q(o[131]) );
  DFF \oi_reg[4][2]  ( .D(N291), .CLK(clk), .RST(rst), .Q(o[130]) );
  DFF \oi_reg[4][1]  ( .D(N290), .CLK(clk), .RST(rst), .Q(o[129]) );
  DFF \oi_reg[4][0]  ( .D(N289), .CLK(clk), .RST(rst), .Q(o[128]) );
  ANDN U3 ( .B(y[714]), .A(n169), .Z(n8423) );
  XOR U4 ( .A(n10845), .B(n10846), .Z(n10848) );
  OR U5 ( .A(n1563), .B(n1564), .Z(n1) );
  OR U6 ( .A(n1852), .B(n1562), .Z(n2) );
  NAND U7 ( .A(n1), .B(n2), .Z(n1666) );
  XOR U8 ( .A(n13661), .B(n13662), .Z(n13655) );
  OR U9 ( .A(n13909), .B(n13910), .Z(n3) );
  NANDN U10 ( .A(n13908), .B(n13907), .Z(n4) );
  NAND U11 ( .A(n3), .B(n4), .Z(n14086) );
  XNOR U12 ( .A(n6473), .B(n6474), .Z(n6446) );
  OR U13 ( .A(n8008), .B(n8009), .Z(n5) );
  NANDN U14 ( .A(n8010), .B(n8011), .Z(n6) );
  AND U15 ( .A(n5), .B(n6), .Z(n8151) );
  XNOR U16 ( .A(n3513), .B(n3514), .Z(n3502) );
  XNOR U17 ( .A(n3830), .B(n3831), .Z(n3833) );
  XNOR U18 ( .A(n3961), .B(n3962), .Z(n3964) );
  XOR U19 ( .A(n4837), .B(n4838), .Z(n4831) );
  OR U20 ( .A(n5181), .B(n5182), .Z(n7) );
  OR U21 ( .A(n5179), .B(n5180), .Z(n8) );
  AND U22 ( .A(n7), .B(n8), .Z(n5373) );
  XNOR U23 ( .A(n10381), .B(n10382), .Z(n10383) );
  XOR U24 ( .A(n7832), .B(n7833), .Z(n7871) );
  XNOR U25 ( .A(n10851), .B(n10852), .Z(n10853) );
  XOR U26 ( .A(n10903), .B(n10904), .Z(n10905) );
  XNOR U27 ( .A(n10969), .B(n10970), .Z(n10971) );
  XNOR U28 ( .A(n6691), .B(n6692), .Z(n6693) );
  XNOR U29 ( .A(n7332), .B(n7333), .Z(n7292) );
  OR U30 ( .A(n7464), .B(n7465), .Z(n9) );
  OR U31 ( .A(n7743), .B(n7463), .Z(n10) );
  NAND U32 ( .A(n9), .B(n10), .Z(n7585) );
  XOR U33 ( .A(n7704), .B(n7705), .Z(n7706) );
  XOR U34 ( .A(n7815), .B(n7814), .Z(n7882) );
  XOR U35 ( .A(n8020), .B(n8021), .Z(n8025) );
  XNOR U36 ( .A(n4041), .B(n4042), .Z(n4065) );
  XNOR U37 ( .A(n4396), .B(n4397), .Z(n4388) );
  ANDN U38 ( .B(y[777]), .A(n152), .Z(n13212) );
  XNOR U39 ( .A(n12478), .B(n12479), .Z(n12467) );
  XOR U40 ( .A(n13607), .B(n13608), .Z(n13539) );
  XNOR U41 ( .A(n13659), .B(n13660), .Z(n13661) );
  XOR U42 ( .A(n14037), .B(n14038), .Z(n14026) );
  OR U43 ( .A(n13911), .B(n13912), .Z(n11) );
  NANDN U44 ( .A(n13913), .B(n13914), .Z(n12) );
  NAND U45 ( .A(n11), .B(n12), .Z(n14089) );
  ANDN U46 ( .B(y[742]), .A(n153), .Z(n9726) );
  XNOR U47 ( .A(n9540), .B(n9541), .Z(n9529) );
  XNOR U48 ( .A(n9652), .B(n9653), .Z(n9654) );
  XNOR U49 ( .A(n10201), .B(n10202), .Z(n10204) );
  XNOR U50 ( .A(n10241), .B(n10242), .Z(n10244) );
  XOR U51 ( .A(n10671), .B(n10670), .Z(n10682) );
  XOR U52 ( .A(n10847), .B(n10848), .Z(n10795) );
  NAND U53 ( .A(y[754]), .B(x[136]), .Z(n11155) );
  XNOR U54 ( .A(n11108), .B(n11109), .Z(n11079) );
  XOR U55 ( .A(n6446), .B(n6445), .Z(n6447) );
  XNOR U56 ( .A(n6604), .B(n6605), .Z(n6593) );
  XNOR U57 ( .A(n7319), .B(n7320), .Z(n7322) );
  XNOR U58 ( .A(n7279), .B(n7280), .Z(n7282) );
  OR U59 ( .A(n7998), .B(n7999), .Z(n13) );
  NANDN U60 ( .A(n8000), .B(n8001), .Z(n14) );
  NAND U61 ( .A(n13), .B(n14), .Z(n8104) );
  XNOR U62 ( .A(n8162), .B(n8163), .Z(n8090) );
  XNOR U63 ( .A(n3654), .B(n3655), .Z(n3643) );
  XOR U64 ( .A(n3502), .B(n3501), .Z(n3503) );
  XOR U65 ( .A(n3569), .B(n3570), .Z(n3554) );
  XNOR U66 ( .A(n3767), .B(n3768), .Z(n3769) );
  XOR U67 ( .A(n3833), .B(n3832), .Z(n3839) );
  XOR U68 ( .A(n3955), .B(n3956), .Z(n3957) );
  XNOR U69 ( .A(n3897), .B(n3898), .Z(n3899) );
  XOR U70 ( .A(n4790), .B(n4789), .Z(n4712) );
  XNOR U71 ( .A(n4835), .B(n4836), .Z(n4837) );
  XOR U72 ( .A(n5093), .B(n5094), .Z(n5013) );
  XNOR U73 ( .A(n689), .B(n690), .Z(n678) );
  XNOR U74 ( .A(n755), .B(n756), .Z(n771) );
  XOR U75 ( .A(n1409), .B(n1408), .Z(n1367) );
  XNOR U76 ( .A(n1431), .B(n1432), .Z(n1442) );
  XOR U77 ( .A(n2207), .B(n2208), .Z(n2210) );
  XNOR U78 ( .A(n12337), .B(n12338), .Z(n12321) );
  OR U79 ( .A(n14082), .B(n14083), .Z(n15) );
  NANDN U80 ( .A(n14084), .B(n14085), .Z(n16) );
  AND U81 ( .A(n15), .B(n16), .Z(n14242) );
  XNOR U82 ( .A(n9399), .B(n9400), .Z(n9383) );
  XNOR U83 ( .A(n11179), .B(n11180), .Z(n11182) );
  XNOR U84 ( .A(n8239), .B(n8240), .Z(n8242) );
  XNOR U85 ( .A(n4100), .B(n4101), .Z(n4173) );
  XNOR U86 ( .A(n4970), .B(n4971), .Z(n4973) );
  ANDN U87 ( .B(y[682]), .A(n169), .Z(n5530) );
  XNOR U88 ( .A(n5381), .B(n5382), .Z(n5425) );
  XOR U89 ( .A(n1769), .B(n1770), .Z(n1746) );
  XOR U90 ( .A(n14313), .B(n14314), .Z(n14278) );
  OR U91 ( .A(n14126), .B(n14127), .Z(n17) );
  NANDN U92 ( .A(n14125), .B(n14124), .Z(n18) );
  NAND U93 ( .A(n17), .B(n18), .Z(n14416) );
  OR U94 ( .A(n14370), .B(n14371), .Z(n19) );
  OR U95 ( .A(n14368), .B(n14369), .Z(n20) );
  NAND U96 ( .A(n19), .B(n20), .Z(n14483) );
  XNOR U97 ( .A(n11559), .B(n11560), .Z(n11551) );
  XNOR U98 ( .A(n11344), .B(n11345), .Z(n11475) );
  OR U99 ( .A(n11304), .B(n11305), .Z(n21) );
  OR U100 ( .A(n11302), .B(n11303), .Z(n22) );
  AND U101 ( .A(n21), .B(n22), .Z(n11472) );
  OR U102 ( .A(n8946), .B(n8682), .Z(n23) );
  OR U103 ( .A(n8680), .B(n8681), .Z(n24) );
  AND U104 ( .A(n23), .B(n24), .Z(n8768) );
  XNOR U105 ( .A(n8521), .B(n8522), .Z(n8535) );
  OR U106 ( .A(n8365), .B(n8366), .Z(n25) );
  NANDN U107 ( .A(n8364), .B(n8363), .Z(n26) );
  NAND U108 ( .A(n25), .B(n26), .Z(n8532) );
  XOR U109 ( .A(n5708), .B(n5709), .Z(n5726) );
  OR U110 ( .A(n5423), .B(n5424), .Z(n27) );
  NANDN U111 ( .A(n5422), .B(n5421), .Z(n28) );
  AND U112 ( .A(n27), .B(n28), .Z(n5601) );
  XNOR U113 ( .A(n5499), .B(n5500), .Z(n5595) );
  XOR U114 ( .A(n14447), .B(n14446), .Z(n14458) );
  XNOR U115 ( .A(n13371), .B(n13372), .Z(n13373) );
  XOR U116 ( .A(n13689), .B(n13690), .Z(n13691) );
  XOR U117 ( .A(n13763), .B(n13764), .Z(n13766) );
  XOR U118 ( .A(n10785), .B(n10786), .Z(n10826) );
  XOR U119 ( .A(n13217), .B(n13218), .Z(n13220) );
  XOR U120 ( .A(n13223), .B(n13224), .Z(n13226) );
  XOR U121 ( .A(n13418), .B(n13417), .Z(n13450) );
  XOR U122 ( .A(n13720), .B(n13721), .Z(n13723) );
  XNOR U123 ( .A(n13925), .B(n13926), .Z(n13928) );
  XNOR U124 ( .A(n13862), .B(n13861), .Z(n13867) );
  XOR U125 ( .A(n9793), .B(n9792), .Z(n9794) );
  XNOR U126 ( .A(n10009), .B(n10010), .Z(n9996) );
  XNOR U127 ( .A(n10152), .B(n10249), .Z(n10104) );
  XOR U128 ( .A(n10965), .B(n10966), .Z(n10972) );
  XOR U129 ( .A(n10893), .B(n10894), .Z(n10896) );
  XOR U130 ( .A(n6399), .B(n6400), .Z(n6401) );
  NAND U131 ( .A(y[717]), .B(x[129]), .Z(n6711) );
  XNOR U132 ( .A(n6815), .B(n6816), .Z(n6817) );
  XOR U133 ( .A(n7355), .B(n7354), .Z(n7356) );
  XNOR U134 ( .A(n7339), .B(n7340), .Z(n7293) );
  XNOR U135 ( .A(n7420), .B(n7421), .Z(n7422) );
  XOR U136 ( .A(n7744), .B(n7745), .Z(n7693) );
  XOR U137 ( .A(n7892), .B(n7893), .Z(n7895) );
  XOR U138 ( .A(n8024), .B(n8025), .Z(n8026) );
  XOR U139 ( .A(n3449), .B(n3450), .Z(n3451) );
  XNOR U140 ( .A(n4244), .B(n4245), .Z(n4246) );
  XOR U141 ( .A(n4382), .B(n4383), .Z(n4385) );
  XNOR U142 ( .A(n4366), .B(n4367), .Z(n4389) );
  XNOR U143 ( .A(n4471), .B(n4472), .Z(n4473) );
  XNOR U144 ( .A(n4787), .B(n4788), .Z(n4790) );
  XOR U145 ( .A(n4896), .B(n4897), .Z(n4899) );
  XOR U146 ( .A(n4952), .B(n4953), .Z(n4954) );
  NAND U147 ( .A(y[681]), .B(x[144]), .Z(n5063) );
  XNOR U148 ( .A(n5030), .B(n5031), .Z(n5032) );
  XNOR U149 ( .A(n1426), .B(n1427), .Z(n1379) );
  XNOR U150 ( .A(n1585), .B(n1586), .Z(n1588) );
  XOR U151 ( .A(n1853), .B(n1854), .Z(n1804) );
  XOR U152 ( .A(n2057), .B(n2058), .Z(n2059) );
  XOR U153 ( .A(n12273), .B(n12274), .Z(n12275) );
  XNOR U154 ( .A(n12571), .B(n12572), .Z(n12573) );
  XNOR U155 ( .A(n12461), .B(n12462), .Z(n12463) );
  XNOR U156 ( .A(n12561), .B(n12562), .Z(n12597) );
  XOR U157 ( .A(n12733), .B(n12734), .Z(n12716) );
  XOR U158 ( .A(n13656), .B(n13655), .Z(n13560) );
  XOR U159 ( .A(n13648), .B(n13647), .Z(n13649) );
  XOR U160 ( .A(n13983), .B(n13984), .Z(n13985) );
  XOR U161 ( .A(n14025), .B(n14026), .Z(n13975) );
  XOR U162 ( .A(n9335), .B(n9336), .Z(n9337) );
  XOR U163 ( .A(n9523), .B(n9524), .Z(n9526) );
  XOR U164 ( .A(n9479), .B(n9480), .Z(n9474) );
  NAND U165 ( .A(y[749]), .B(x[129]), .Z(n9614) );
  XNOR U166 ( .A(n9605), .B(n9606), .Z(n9620) );
  XNOR U167 ( .A(n10167), .B(n10168), .Z(n10133) );
  XOR U168 ( .A(n10209), .B(n10210), .Z(n10235) );
  XOR U169 ( .A(n10244), .B(n10243), .Z(n10203) );
  XNOR U170 ( .A(n10474), .B(n10475), .Z(n10467) );
  XOR U171 ( .A(n10686), .B(n10687), .Z(n10689) );
  XOR U172 ( .A(n10622), .B(n10623), .Z(n10605) );
  XNOR U173 ( .A(n10668), .B(n10669), .Z(n10671) );
  XOR U174 ( .A(n10792), .B(n10791), .Z(n10798) );
  NAND U175 ( .A(y[753]), .B(x[137]), .Z(n11156) );
  OR U176 ( .A(n10948), .B(n10949), .Z(n29) );
  NANDN U177 ( .A(n10950), .B(n10951), .Z(n30) );
  NAND U178 ( .A(n29), .B(n30), .Z(n11034) );
  OR U179 ( .A(n10944), .B(n10945), .Z(n31) );
  NANDN U180 ( .A(n10946), .B(n10947), .Z(n32) );
  AND U181 ( .A(n31), .B(n32), .Z(n11030) );
  OR U182 ( .A(n10934), .B(n10935), .Z(n33) );
  NANDN U183 ( .A(n10936), .B(n10937), .Z(n34) );
  NAND U184 ( .A(n33), .B(n34), .Z(n11090) );
  NAND U185 ( .A(y[712]), .B(x[130]), .Z(n6379) );
  XNOR U186 ( .A(n6675), .B(n6676), .Z(n6717) );
  XOR U187 ( .A(n7700), .B(n7701), .Z(n7671) );
  XOR U188 ( .A(n7888), .B(n7889), .Z(n7842) );
  NAND U189 ( .A(y[722]), .B(x[136]), .Z(n8216) );
  XNOR U190 ( .A(n8122), .B(n8123), .Z(n8093) );
  XOR U191 ( .A(n3637), .B(n3638), .Z(n3639) );
  XOR U192 ( .A(n3679), .B(n3678), .Z(n3680) );
  XNOR U193 ( .A(n3751), .B(n3752), .Z(n3734) );
  XNOR U194 ( .A(n3815), .B(n3816), .Z(n3817) );
  XNOR U195 ( .A(n3836), .B(n3837), .Z(n3838) );
  XOR U196 ( .A(n4120), .B(n4119), .Z(n4121) );
  XNOR U197 ( .A(n4167), .B(n4168), .Z(n4169) );
  XOR U198 ( .A(n4783), .B(n4784), .Z(n4715) );
  XNOR U199 ( .A(n4829), .B(n4830), .Z(n4832) );
  XOR U200 ( .A(n4754), .B(n4753), .Z(n4838) );
  XOR U201 ( .A(n5215), .B(n5216), .Z(n5221) );
  XNOR U202 ( .A(n543), .B(n544), .Z(n545) );
  XOR U203 ( .A(n624), .B(n625), .Z(n603) );
  XOR U204 ( .A(n672), .B(n673), .Z(n675) );
  XOR U205 ( .A(n634), .B(n635), .Z(n629) );
  NAND U206 ( .A(y[653]), .B(x[129]), .Z(n764) );
  XNOR U207 ( .A(n799), .B(n800), .Z(n770) );
  XOR U208 ( .A(n972), .B(n971), .Z(n964) );
  XNOR U209 ( .A(n1319), .B(n1320), .Z(n1285) );
  XOR U210 ( .A(n1373), .B(n1374), .Z(n1400) );
  XNOR U211 ( .A(n1365), .B(n1366), .Z(n1368) );
  XOR U212 ( .A(n1442), .B(n1441), .Z(n1443) );
  XOR U213 ( .A(n2051), .B(n2052), .Z(n2054) );
  XOR U214 ( .A(n2447), .B(n2448), .Z(n2466) );
  XOR U215 ( .A(n2231), .B(n2232), .Z(n2234) );
  OR U216 ( .A(n12665), .B(n12152), .Z(n35) );
  OR U217 ( .A(n12150), .B(n12151), .Z(n36) );
  NAND U218 ( .A(n35), .B(n36), .Z(n12213) );
  OR U219 ( .A(n13155), .B(n12255), .Z(n37) );
  NANDN U220 ( .A(n13212), .B(n12256), .Z(n38) );
  NAND U221 ( .A(n37), .B(n38), .Z(n12331) );
  XOR U222 ( .A(n12321), .B(n12320), .Z(n12322) );
  XOR U223 ( .A(n12468), .B(n12467), .Z(n12469) );
  XNOR U224 ( .A(n13490), .B(n13491), .Z(n13401) );
  XOR U225 ( .A(n13538), .B(n13539), .Z(n13549) );
  XNOR U226 ( .A(n13744), .B(n13745), .Z(n13746) );
  XNOR U227 ( .A(n14090), .B(n14091), .Z(n14092) );
  OR U228 ( .A(n13979), .B(n13980), .Z(n39) );
  NANDN U229 ( .A(n13981), .B(n13982), .Z(n40) );
  NAND U230 ( .A(n39), .B(n40), .Z(n14129) );
  OR U231 ( .A(n14233), .B(n14234), .Z(n41) );
  OR U232 ( .A(n14231), .B(n14232), .Z(n42) );
  NAND U233 ( .A(n41), .B(n42), .Z(n14375) );
  OR U234 ( .A(n9726), .B(n9200), .Z(n43) );
  OR U235 ( .A(n9198), .B(n9199), .Z(n44) );
  NAND U236 ( .A(n43), .B(n44), .Z(n9273) );
  XOR U237 ( .A(n9383), .B(n9382), .Z(n9384) );
  XOR U238 ( .A(n9594), .B(n9595), .Z(n9597) );
  XOR U239 ( .A(n10082), .B(n10083), .Z(n10086) );
  XNOR U240 ( .A(n10303), .B(n10304), .Z(n10295) );
  XNOR U241 ( .A(n10426), .B(n10427), .Z(n10337) );
  XNOR U242 ( .A(n10574), .B(n10575), .Z(n10460) );
  XNOR U243 ( .A(n10921), .B(n10922), .Z(n10924) );
  XNOR U244 ( .A(n11242), .B(n11243), .Z(n11244) );
  XNOR U245 ( .A(n11250), .B(n11251), .Z(n11256) );
  OR U246 ( .A(n11540), .B(n11541), .Z(n45) );
  OR U247 ( .A(n11766), .B(n11539), .Z(n46) );
  AND U248 ( .A(n45), .B(n46), .Z(n11795) );
  XNOR U249 ( .A(n11320), .B(n11321), .Z(n11315) );
  OR U250 ( .A(n6789), .B(n6292), .Z(n47) );
  OR U251 ( .A(n6290), .B(n6291), .Z(n48) );
  AND U252 ( .A(n47), .B(n48), .Z(n6337) );
  XNOR U253 ( .A(n6533), .B(n6534), .Z(n6557) );
  XNOR U254 ( .A(n6563), .B(n6564), .Z(n6565) );
  XOR U255 ( .A(n6664), .B(n6665), .Z(n6667) );
  XOR U256 ( .A(n6822), .B(n6821), .Z(n6823) );
  XOR U257 ( .A(n7118), .B(n7119), .Z(n7044) );
  XOR U258 ( .A(n7282), .B(n7281), .Z(n7369) );
  XNOR U259 ( .A(n7402), .B(n7403), .Z(n7404) );
  XOR U260 ( .A(n7664), .B(n7665), .Z(n7768) );
  XOR U261 ( .A(n7773), .B(n7774), .Z(n7656) );
  XNOR U262 ( .A(n7982), .B(n7983), .Z(n8051) );
  XOR U263 ( .A(n8311), .B(n8312), .Z(n8318) );
  XNOR U264 ( .A(n3613), .B(n3614), .Z(n3615) );
  XOR U265 ( .A(n3555), .B(n3556), .Z(n3607) );
  XOR U266 ( .A(n3708), .B(n3709), .Z(n3711) );
  XNOR U267 ( .A(n3919), .B(n3920), .Z(n3921) );
  XOR U268 ( .A(n3964), .B(n3963), .Z(n3891) );
  XOR U269 ( .A(n4033), .B(n4032), .Z(n3991) );
  XOR U270 ( .A(n4314), .B(n4315), .Z(n4307) );
  XOR U271 ( .A(n4720), .B(n4721), .Z(n4730) );
  XNOR U272 ( .A(n5018), .B(n5019), .Z(n5020) );
  XNOR U273 ( .A(n5280), .B(n5281), .Z(n5282) );
  OR U274 ( .A(n859), .B(n351), .Z(n49) );
  OR U275 ( .A(n349), .B(n350), .Z(n50) );
  NAND U276 ( .A(n49), .B(n50), .Z(n425) );
  XOR U277 ( .A(n782), .B(n783), .Z(n785) );
  XOR U278 ( .A(n1198), .B(n1199), .Z(n1222) );
  XNOR U279 ( .A(n1226), .B(n1227), .Z(n1228) );
  XOR U280 ( .A(n1234), .B(n1235), .Z(n1238) );
  XNOR U281 ( .A(n1461), .B(n1462), .Z(n1465) );
  XOR U282 ( .A(n1745), .B(n1746), .Z(n1755) );
  XOR U283 ( .A(n1879), .B(n1880), .Z(n1884) );
  XNOR U284 ( .A(n12029), .B(n12030), .Z(n12015) );
  XOR U285 ( .A(n14277), .B(n14278), .Z(n14399) );
  XOR U286 ( .A(n14271), .B(n14272), .Z(n14411) );
  OR U287 ( .A(n14243), .B(n14244), .Z(n51) );
  OR U288 ( .A(n14241), .B(n14242), .Z(n52) );
  AND U289 ( .A(n51), .B(n52), .Z(n14423) );
  OR U290 ( .A(n14121), .B(n14120), .Z(n53) );
  NANDN U291 ( .A(n14123), .B(n14122), .Z(n54) );
  NAND U292 ( .A(n53), .B(n54), .Z(n14417) );
  XOR U293 ( .A(n14501), .B(n14502), .Z(n14506) );
  XOR U294 ( .A(n14650), .B(n14651), .Z(n14649) );
  XNOR U295 ( .A(n10068), .B(n10069), .Z(n10070) );
  XNOR U296 ( .A(n10331), .B(n10332), .Z(n10334) );
  OR U297 ( .A(n11238), .B(n11239), .Z(n55) );
  NANDN U298 ( .A(n11240), .B(n11241), .Z(n56) );
  NAND U299 ( .A(n55), .B(n56), .Z(n11342) );
  XOR U300 ( .A(n11386), .B(n11387), .Z(n11351) );
  XOR U301 ( .A(n11639), .B(n11640), .Z(n11644) );
  XNOR U302 ( .A(n6155), .B(n6156), .Z(n6141) );
  OR U303 ( .A(n8299), .B(n8300), .Z(n57) );
  NANDN U304 ( .A(n8301), .B(n8302), .Z(n58) );
  NAND U305 ( .A(n57), .B(n58), .Z(n8519) );
  XOR U306 ( .A(n8454), .B(n8455), .Z(n8515) );
  OR U307 ( .A(n8425), .B(n8426), .Z(n59) );
  OR U308 ( .A(n8423), .B(n8424), .Z(n60) );
  NAND U309 ( .A(n59), .B(n60), .Z(n8583) );
  XNOR U310 ( .A(n3203), .B(n3204), .Z(n3189) );
  XNOR U311 ( .A(n5133), .B(n5134), .Z(n5135) );
  OR U312 ( .A(n5363), .B(n5364), .Z(n61) );
  NANDN U313 ( .A(n5365), .B(n5366), .Z(n62) );
  NAND U314 ( .A(n61), .B(n62), .Z(n5497) );
  OR U315 ( .A(n5871), .B(n5697), .Z(n63) );
  OR U316 ( .A(n5695), .B(n5696), .Z(n64) );
  AND U317 ( .A(n63), .B(n64), .Z(n5832) );
  XOR U318 ( .A(n5763), .B(n5764), .Z(n5768) );
  XOR U319 ( .A(n2508), .B(n2509), .Z(n2637) );
  OR U320 ( .A(n2956), .B(n2808), .Z(n65) );
  OR U321 ( .A(n2806), .B(n2807), .Z(n66) );
  AND U322 ( .A(n65), .B(n66), .Z(n2882) );
  XOR U323 ( .A(n2728), .B(n2729), .Z(n2733) );
  OR U324 ( .A(n14486), .B(n14696), .Z(n67) );
  NANDN U325 ( .A(n14488), .B(n14487), .Z(n68) );
  NAND U326 ( .A(n67), .B(n68), .Z(n14639) );
  XNOR U327 ( .A(n11673), .B(n11674), .Z(n11943) );
  OR U328 ( .A(n11471), .B(n11472), .Z(n69) );
  NANDN U329 ( .A(n11474), .B(n11473), .Z(n70) );
  AND U330 ( .A(n69), .B(n70), .Z(n11505) );
  OR U331 ( .A(n8588), .B(n8589), .Z(n71) );
  OR U332 ( .A(n8813), .B(n8587), .Z(n72) );
  NAND U333 ( .A(n71), .B(n72), .Z(n8756) );
  OR U334 ( .A(n8531), .B(n8532), .Z(n73) );
  NANDN U335 ( .A(n8534), .B(n8533), .Z(n74) );
  AND U336 ( .A(n73), .B(n74), .Z(n8565) );
  XNOR U337 ( .A(n5635), .B(n5636), .Z(n5709) );
  OR U338 ( .A(n5602), .B(n5601), .Z(n75) );
  NANDN U339 ( .A(n5604), .B(n5603), .Z(n76) );
  NAND U340 ( .A(n75), .B(n76), .Z(n5629) );
  XNOR U341 ( .A(n14610), .B(n14611), .Z(n14898) );
  XOR U342 ( .A(n11959), .B(n11960), .Z(n11956) );
  XOR U343 ( .A(n8735), .B(n8736), .Z(n8734) );
  ANDN U344 ( .B(y[771]), .A(n162), .Z(n12680) );
  XOR U345 ( .A(n7868), .B(n7869), .Z(n7870) );
  XOR U346 ( .A(n4911), .B(n4910), .Z(n4940) );
  XOR U347 ( .A(n1945), .B(n1946), .Z(n1913) );
  XOR U348 ( .A(n12565), .B(n12566), .Z(n12568) );
  XNOR U349 ( .A(n12691), .B(n12692), .Z(n12693) );
  XOR U350 ( .A(n12786), .B(n12785), .Z(n12761) );
  XNOR U351 ( .A(n12865), .B(n12866), .Z(n12867) );
  XNOR U352 ( .A(n12820), .B(n12821), .Z(n12822) );
  XOR U353 ( .A(n13068), .B(n13069), .Z(n13071) );
  XOR U354 ( .A(n13062), .B(n13063), .Z(n13065) );
  XOR U355 ( .A(n13715), .B(n13329), .Z(n13302) );
  XNOR U356 ( .A(n13407), .B(n13408), .Z(n13409) );
  XNOR U357 ( .A(n13464), .B(n13465), .Z(n13508) );
  XOR U358 ( .A(n13468), .B(n13469), .Z(n13470) );
  XNOR U359 ( .A(n13611), .B(n13612), .Z(n13613) );
  XOR U360 ( .A(n13775), .B(n13776), .Z(n13777) );
  XNOR U361 ( .A(n9776), .B(n9777), .Z(n9778) );
  XNOR U362 ( .A(n9876), .B(n9877), .Z(n9878) );
  XNOR U363 ( .A(n10139), .B(n10140), .Z(n10141) );
  XOR U364 ( .A(n10213), .B(n10214), .Z(n10216) );
  XOR U365 ( .A(n10509), .B(n10510), .Z(n10512) );
  XOR U366 ( .A(n10552), .B(n10553), .Z(n10554) );
  XNOR U367 ( .A(n10626), .B(n10627), .Z(n10628) );
  XOR U368 ( .A(n10887), .B(n10888), .Z(n10890) );
  XOR U369 ( .A(n10987), .B(n10988), .Z(n10990) );
  XOR U370 ( .A(n6688), .B(n6687), .Z(n6694) );
  XNOR U371 ( .A(n6950), .B(n6951), .Z(n6952) );
  XNOR U372 ( .A(n7212), .B(n7331), .Z(n7166) );
  XNOR U373 ( .A(n7344), .B(n7345), .Z(n7355) );
  XNOR U374 ( .A(n7348), .B(n7349), .Z(n7350) );
  XNOR U375 ( .A(n7408), .B(n7409), .Z(n7410) );
  XOR U376 ( .A(n7432), .B(n7433), .Z(n7435) );
  ANDN U377 ( .B(y[718]), .A(n158), .Z(n7743) );
  XOR U378 ( .A(n7740), .B(n7739), .Z(n7694) );
  XOR U379 ( .A(n7880), .B(n7881), .Z(n7883) );
  XNOR U380 ( .A(n7856), .B(n7857), .Z(n7874) );
  XOR U381 ( .A(n7986), .B(n7987), .Z(n7988) );
  XOR U382 ( .A(n7962), .B(n7963), .Z(n7964) );
  XNOR U383 ( .A(n3430), .B(n4365), .Z(n3438) );
  XOR U384 ( .A(n4145), .B(n4223), .Z(n4125) );
  XNOR U385 ( .A(n4132), .B(n4133), .Z(n4120) );
  XOR U386 ( .A(n4483), .B(n4484), .Z(n4485) );
  XNOR U387 ( .A(n4589), .B(n4590), .Z(n4591) );
  XNOR U388 ( .A(n4646), .B(n4647), .Z(n4690) );
  XOR U389 ( .A(n4664), .B(n4665), .Z(n4666) );
  XOR U390 ( .A(n4946), .B(n4947), .Z(n4949) );
  NAND U391 ( .A(y[672]), .B(x[153]), .Z(n5103) );
  XNOR U392 ( .A(n5109), .B(n5110), .Z(n5112) );
  XOR U393 ( .A(n5115), .B(n5116), .Z(n5118) );
  XNOR U394 ( .A(n952), .B(n953), .Z(n933) );
  XNOR U395 ( .A(n1027), .B(n1028), .Z(n1075) );
  XOR U396 ( .A(n1069), .B(n1070), .Z(n1072) );
  XOR U397 ( .A(n1161), .B(n1162), .Z(n1149) );
  XNOR U398 ( .A(n1298), .B(n1418), .Z(n1275) );
  XOR U399 ( .A(n1377), .B(n1378), .Z(n1380) );
  XOR U400 ( .A(n1588), .B(n1587), .Z(n1509) );
  XOR U401 ( .A(n1815), .B(n1816), .Z(n1817) );
  XNOR U402 ( .A(n1665), .B(n1666), .Z(n1678) );
  XOR U403 ( .A(n1859), .B(n1860), .Z(n1805) );
  XOR U404 ( .A(n1919), .B(n1920), .Z(n1921) );
  XOR U405 ( .A(n1980), .B(n1981), .Z(n1928) );
  XOR U406 ( .A(n12245), .B(n12246), .Z(n12248) );
  XOR U407 ( .A(n12502), .B(n12503), .Z(n12505) );
  XOR U408 ( .A(n12598), .B(n12597), .Z(n12599) );
  XNOR U409 ( .A(n12670), .B(n12671), .Z(n12672) );
  XOR U410 ( .A(n12985), .B(n12986), .Z(n12988) );
  XOR U411 ( .A(n13196), .B(n13195), .Z(n13197) );
  XNOR U412 ( .A(n13297), .B(n13298), .Z(n13309) );
  XOR U413 ( .A(n13183), .B(n13184), .Z(n13186) );
  XOR U414 ( .A(n13283), .B(n13284), .Z(n13286) );
  XNOR U415 ( .A(n13653), .B(n13654), .Z(n13656) );
  XOR U416 ( .A(n13578), .B(n13577), .Z(n13662) );
  XOR U417 ( .A(n13835), .B(n13836), .Z(n13838) );
  XOR U418 ( .A(n13847), .B(n13848), .Z(n13850) );
  OR U419 ( .A(n13917), .B(n13918), .Z(n77) );
  NANDN U420 ( .A(n13916), .B(n13915), .Z(n78) );
  AND U421 ( .A(n77), .B(n78), .Z(n14082) );
  XOR U422 ( .A(n9469), .B(n9470), .Z(n9447) );
  XOR U423 ( .A(n9565), .B(n9564), .Z(n9566) );
  XOR U424 ( .A(n9649), .B(n9648), .Z(n9655) );
  XOR U425 ( .A(n9620), .B(n9619), .Z(n9621) );
  XNOR U426 ( .A(n9996), .B(n9997), .Z(n9998) );
  XOR U427 ( .A(n10134), .B(n10133), .Z(n10135) );
  XOR U428 ( .A(n10278), .B(n10277), .Z(n10279) );
  XNOR U429 ( .A(n10271), .B(n10272), .Z(n10273) );
  XOR U430 ( .A(n10467), .B(n10466), .Z(n10468) );
  XOR U431 ( .A(n10662), .B(n10663), .Z(n10665) );
  XOR U432 ( .A(n10740), .B(n10741), .Z(n10743) );
  XNOR U433 ( .A(n10909), .B(n10910), .Z(n10911) );
  XNOR U434 ( .A(n11139), .B(n11138), .Z(n11035) );
  OR U435 ( .A(n10899), .B(n10900), .Z(n79) );
  NANDN U436 ( .A(n10901), .B(n10902), .Z(n80) );
  NAND U437 ( .A(n79), .B(n80), .Z(n11083) );
  XNOR U438 ( .A(n11066), .B(n11067), .Z(n11076) );
  XNOR U439 ( .A(n6434), .B(n6435), .Z(n6436) );
  XOR U440 ( .A(n6587), .B(n6588), .Z(n6590) );
  XNOR U441 ( .A(n6537), .B(n6538), .Z(n6531) );
  XOR U442 ( .A(n6612), .B(n6611), .Z(n6613) );
  XOR U443 ( .A(n6718), .B(n6717), .Z(n6719) );
  XNOR U444 ( .A(n6794), .B(n6795), .Z(n6796) );
  OR U445 ( .A(n6902), .B(n6765), .Z(n81) );
  NANDN U446 ( .A(n6767), .B(n6766), .Z(n82) );
  AND U447 ( .A(n81), .B(n82), .Z(n6872) );
  XNOR U448 ( .A(n7193), .B(n7194), .Z(n7195) );
  XOR U449 ( .A(n7287), .B(n7288), .Z(n7313) );
  XOR U450 ( .A(n7322), .B(n7321), .Z(n7281) );
  XNOR U451 ( .A(n7426), .B(n7427), .Z(n7428) );
  XNOR U452 ( .A(n7614), .B(n7615), .Z(n7616) );
  XNOR U453 ( .A(n8199), .B(n8198), .Z(n8146) );
  OR U454 ( .A(n7960), .B(n7961), .Z(n83) );
  OR U455 ( .A(n7958), .B(n7959), .Z(n84) );
  NAND U456 ( .A(n83), .B(n84), .Z(n8097) );
  XNOR U457 ( .A(n3490), .B(n3491), .Z(n3492) );
  XOR U458 ( .A(n3597), .B(n3598), .Z(n3581) );
  XOR U459 ( .A(n3764), .B(n3763), .Z(n3770) );
  XOR U460 ( .A(n3735), .B(n3734), .Z(n3736) );
  XNOR U461 ( .A(n3843), .B(n3844), .Z(n3832) );
  XNOR U462 ( .A(n4058), .B(n4059), .Z(n4060) );
  XOR U463 ( .A(n4065), .B(n4064), .Z(n4066) );
  XNOR U464 ( .A(n4030), .B(n4031), .Z(n4033) );
  XOR U465 ( .A(n4251), .B(n4250), .Z(n4252) );
  XNOR U466 ( .A(n4330), .B(n4331), .Z(n4332) );
  XOR U467 ( .A(n4561), .B(n4562), .Z(n4554) );
  XOR U468 ( .A(n4832), .B(n4831), .Z(n4736) );
  XOR U469 ( .A(n4824), .B(n4823), .Z(n4825) );
  XOR U470 ( .A(n5012), .B(n5013), .Z(n5015) );
  XNOR U471 ( .A(n5258), .B(n5259), .Z(n5163) );
  XNOR U472 ( .A(n5185), .B(n5186), .Z(n5225) );
  XOR U473 ( .A(n565), .B(n566), .Z(n532) );
  XOR U474 ( .A(n714), .B(n713), .Z(n715) );
  XOR U475 ( .A(n771), .B(n770), .Z(n772) );
  XNOR U476 ( .A(n969), .B(n970), .Z(n972) );
  XOR U477 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U478 ( .A(n1435), .B(n1436), .Z(n1437) );
  XNOR U479 ( .A(n1406), .B(n1407), .Z(n1409) );
  XNOR U480 ( .A(n1695), .B(n1696), .Z(n1697) );
  XNOR U481 ( .A(n1811), .B(n1812), .Z(n1793) );
  XNOR U482 ( .A(n1823), .B(n1824), .Z(n1785) );
  ANDN U483 ( .B(y[656]), .A(n162), .Z(n2447) );
  XNOR U484 ( .A(n2283), .B(n2284), .Z(n2197) );
  XNOR U485 ( .A(n2253), .B(n2254), .Z(n2192) );
  XNOR U486 ( .A(n2221), .B(n2222), .Z(n2257) );
  XOR U487 ( .A(n12265), .B(n12264), .Z(n12285) );
  XNOR U488 ( .A(n12331), .B(n12332), .Z(n12333) );
  XNOR U489 ( .A(n12314), .B(n12315), .Z(n12316) );
  XNOR U490 ( .A(n12546), .B(n12547), .Z(n12533) );
  XOR U491 ( .A(n13003), .B(n13004), .Z(n13006) );
  XNOR U492 ( .A(n13279), .B(n13280), .Z(n13271) );
  XNOR U493 ( .A(n13677), .B(n13678), .Z(n13679) );
  XNOR U494 ( .A(n13841), .B(n13842), .Z(n13843) );
  XNOR U495 ( .A(n13793), .B(n13794), .Z(n13795) );
  OR U496 ( .A(n14067), .B(n14068), .Z(n85) );
  OR U497 ( .A(n14065), .B(n14066), .Z(n86) );
  NAND U498 ( .A(n85), .B(n86), .Z(n14172) );
  XNOR U499 ( .A(n14203), .B(n14204), .Z(n14128) );
  OR U500 ( .A(n14087), .B(n14086), .Z(n87) );
  NANDN U501 ( .A(n14089), .B(n14088), .Z(n88) );
  NAND U502 ( .A(n87), .B(n88), .Z(n14243) );
  OR U503 ( .A(n14013), .B(n14014), .Z(n89) );
  NANDN U504 ( .A(n14016), .B(n14015), .Z(n90) );
  AND U505 ( .A(n89), .B(n90), .Z(n14120) );
  XNOR U506 ( .A(n9393), .B(n9394), .Z(n9395) );
  XNOR U507 ( .A(n9376), .B(n9377), .Z(n9378) );
  XOR U508 ( .A(n9475), .B(n9476), .Z(n9499) );
  XOR U509 ( .A(n9530), .B(n9529), .Z(n9531) );
  XOR U510 ( .A(n9800), .B(n9801), .Z(n9807) );
  XNOR U511 ( .A(n9733), .B(n9734), .Z(n9694) );
  XOR U512 ( .A(n9690), .B(n9691), .Z(n9683) );
  OR U513 ( .A(n9910), .B(n9911), .Z(n91) );
  OR U514 ( .A(n9983), .B(n9909), .Z(n92) );
  NAND U515 ( .A(n91), .B(n92), .Z(n10064) );
  XOR U516 ( .A(n9978), .B(n9977), .Z(n10050) );
  XOR U517 ( .A(n10204), .B(n10203), .Z(n10292) );
  XNOR U518 ( .A(n10610), .B(n10611), .Z(n10614) );
  XNOR U519 ( .A(n10734), .B(n10735), .Z(n10736) );
  XNOR U520 ( .A(n11234), .B(n11235), .Z(n11263) );
  XNOR U521 ( .A(n11392), .B(n11393), .Z(n11356) );
  AND U522 ( .A(x[146]), .B(y[746]), .Z(n11442) );
  XOR U523 ( .A(n11454), .B(n11455), .Z(n11461) );
  OR U524 ( .A(n11029), .B(n11030), .Z(n93) );
  NANDN U525 ( .A(n11032), .B(n11031), .Z(n94) );
  AND U526 ( .A(n93), .B(n94), .Z(n11304) );
  XOR U527 ( .A(n11182), .B(n11181), .Z(n11307) );
  XNOR U528 ( .A(n6485), .B(n6486), .Z(n6487) );
  XOR U529 ( .A(n6594), .B(n6593), .Z(n6595) );
  XOR U530 ( .A(n6755), .B(n6756), .Z(n6748) );
  XOR U531 ( .A(n6862), .B(n6863), .Z(n6869) );
  XOR U532 ( .A(n7050), .B(n7049), .Z(n7122) );
  XOR U533 ( .A(n7380), .B(n7381), .Z(n7373) );
  XNOR U534 ( .A(n7900), .B(n7901), .Z(n7910) );
  XOR U535 ( .A(n8092), .B(n8093), .Z(n8167) );
  XNOR U536 ( .A(n8460), .B(n8461), .Z(n8497) );
  XOR U537 ( .A(n8441), .B(n8442), .Z(n8429) );
  OR U538 ( .A(n8151), .B(n8150), .Z(n95) );
  NANDN U539 ( .A(n8153), .B(n8152), .Z(n96) );
  NAND U540 ( .A(n95), .B(n96), .Z(n8365) );
  XOR U541 ( .A(n8242), .B(n8241), .Z(n8368) );
  OR U542 ( .A(n3868), .B(n3340), .Z(n97) );
  OR U543 ( .A(n3338), .B(n3339), .Z(n98) );
  AND U544 ( .A(n97), .B(n98), .Z(n3387) );
  XNOR U545 ( .A(n3507), .B(n3508), .Z(n3509) );
  XOR U546 ( .A(n3644), .B(n3643), .Z(n3645) );
  XNOR U547 ( .A(n4076), .B(n4077), .Z(n4078) );
  XNOR U548 ( .A(n4187), .B(n4188), .Z(n4094) );
  XOR U549 ( .A(n4306), .B(n4307), .Z(n4309) );
  XOR U550 ( .A(n4431), .B(n4432), .Z(n4424) );
  XNOR U551 ( .A(n4672), .B(n4673), .Z(n4577) );
  XOR U552 ( .A(n4853), .B(n4854), .Z(n4856) );
  XNOR U553 ( .A(n4920), .B(n4921), .Z(n4922) );
  XNOR U554 ( .A(n4861), .B(n4862), .Z(n4972) );
  XNOR U555 ( .A(n5560), .B(n5561), .Z(n5481) );
  OR U556 ( .A(n5158), .B(n5157), .Z(n99) );
  NANDN U557 ( .A(n5160), .B(n5159), .Z(n100) );
  NAND U558 ( .A(n99), .B(n100), .Z(n5427) );
  XOR U559 ( .A(n5310), .B(n5311), .Z(n5313) );
  XOR U560 ( .A(n679), .B(n678), .Z(n680) );
  XOR U561 ( .A(n841), .B(n842), .Z(n834) );
  XOR U562 ( .A(n1131), .B(n1130), .Z(n1202) );
  XNOR U563 ( .A(n2150), .B(n2149), .Z(n2143) );
  XOR U564 ( .A(n2119), .B(n2120), .Z(n2130) );
  XNOR U565 ( .A(n2271), .B(n2272), .Z(n2178) );
  XNOR U566 ( .A(n2314), .B(n2315), .Z(n2263) );
  XOR U567 ( .A(n2586), .B(n2587), .Z(n2593) );
  XOR U568 ( .A(n2958), .B(n2957), .Z(n2926) );
  XNOR U569 ( .A(n2544), .B(n2545), .Z(n2520) );
  XNOR U570 ( .A(n2435), .B(n2436), .Z(n2360) );
  XOR U571 ( .A(n2342), .B(n2343), .Z(n2345) );
  XNOR U572 ( .A(n12437), .B(n12438), .Z(n12439) );
  XNOR U573 ( .A(n12377), .B(n12378), .Z(n12379) );
  XOR U574 ( .A(n12893), .B(n12894), .Z(n12896) );
  XOR U575 ( .A(n14251), .B(n14252), .Z(n14254) );
  XOR U576 ( .A(n14400), .B(n14401), .Z(n14412) );
  XOR U577 ( .A(n14476), .B(n14477), .Z(n14599) );
  ANDN U578 ( .B(y[788]), .A(n160), .Z(n14696) );
  OR U579 ( .A(n14703), .B(n14575), .Z(n101) );
  OR U580 ( .A(n14573), .B(n14574), .Z(n102) );
  AND U581 ( .A(n101), .B(n102), .Z(n14651) );
  XOR U582 ( .A(n14684), .B(n14685), .Z(n14682) );
  XNOR U583 ( .A(n9348), .B(n9349), .Z(n9299) );
  XNOR U584 ( .A(n9439), .B(n9440), .Z(n9441) );
  XOR U585 ( .A(n9665), .B(n9664), .Z(n9666) );
  XNOR U586 ( .A(n10339), .B(n10340), .Z(n10333) );
  XOR U587 ( .A(n10924), .B(n10923), .Z(n10881) );
  XOR U588 ( .A(n11374), .B(n11375), .Z(n11380) );
  OR U589 ( .A(n11229), .B(n11228), .Z(n103) );
  NANDN U590 ( .A(n11231), .B(n11230), .Z(n104) );
  NAND U591 ( .A(n103), .B(n104), .Z(n11345) );
  XOR U592 ( .A(n11614), .B(n11615), .Z(n11597) );
  XNOR U593 ( .A(n11758), .B(n11759), .Z(n11739) );
  XOR U594 ( .A(n11721), .B(n11722), .Z(n11719) );
  XOR U595 ( .A(n11713), .B(n11714), .Z(n11712) );
  OR U596 ( .A(n11450), .B(n11451), .Z(n105) );
  NANDN U597 ( .A(n11449), .B(n11448), .Z(n106) );
  AND U598 ( .A(n105), .B(n106), .Z(n11557) );
  OR U599 ( .A(n6328), .B(n6329), .Z(n107) );
  OR U600 ( .A(n6670), .B(n6995), .Z(n108) );
  NAND U601 ( .A(n107), .B(n108), .Z(n6416) );
  XNOR U602 ( .A(n7396), .B(n7397), .Z(n7398) );
  XOR U603 ( .A(n8050), .B(n8051), .Z(n8066) );
  XNOR U604 ( .A(n8223), .B(n8224), .Z(n8078) );
  XOR U605 ( .A(n8509), .B(n8510), .Z(n8527) );
  OR U606 ( .A(n8290), .B(n8289), .Z(n109) );
  NAND U607 ( .A(n8292), .B(n8291), .Z(n110) );
  NAND U608 ( .A(n109), .B(n110), .Z(n8522) );
  XOR U609 ( .A(n8602), .B(n8603), .Z(n8607) );
  XOR U610 ( .A(n8571), .B(n8572), .Z(n8706) );
  XNOR U611 ( .A(n8620), .B(n8621), .Z(n8693) );
  XOR U612 ( .A(n8781), .B(n8782), .Z(n8779) );
  XOR U613 ( .A(n8767), .B(n8768), .Z(n8766) );
  XOR U614 ( .A(n3633), .B(n3634), .Z(n3627) );
  XOR U615 ( .A(n3780), .B(n3779), .Z(n3781) );
  XOR U616 ( .A(n3893), .B(n3894), .Z(n3885) );
  XNOR U617 ( .A(n3985), .B(n3986), .Z(n3987) );
  XOR U618 ( .A(n5021), .B(n5020), .Z(n5000) );
  XOR U619 ( .A(n5443), .B(n5444), .Z(n5446) );
  OR U620 ( .A(n5354), .B(n5353), .Z(n111) );
  NANDN U621 ( .A(n5356), .B(n5355), .Z(n112) );
  NAND U622 ( .A(n111), .B(n112), .Z(n5500) );
  XOR U623 ( .A(n5585), .B(n5586), .Z(n5470) );
  XOR U624 ( .A(n5493), .B(n5494), .Z(n5591) );
  XOR U625 ( .A(n5511), .B(n5512), .Z(n5518) );
  XOR U626 ( .A(n5732), .B(n5733), .Z(n5720) );
  XNOR U627 ( .A(n5700), .B(n5699), .Z(n5737) );
  OR U628 ( .A(n5532), .B(n5533), .Z(n113) );
  OR U629 ( .A(n5530), .B(n5531), .Z(n114) );
  NAND U630 ( .A(n113), .B(n114), .Z(n5745) );
  XOR U631 ( .A(n5865), .B(n5866), .Z(n5863) );
  XOR U632 ( .A(n5831), .B(n5832), .Z(n5830) );
  XNOR U633 ( .A(n5451), .B(n5452), .Z(n5611) );
  XOR U634 ( .A(n744), .B(n743), .Z(n745) );
  XOR U635 ( .A(n1010), .B(n1011), .Z(n1112) );
  XOR U636 ( .A(n1593), .B(n1594), .Z(n1485) );
  XOR U637 ( .A(n2568), .B(n2569), .Z(n2532) );
  XNOR U638 ( .A(n2811), .B(n2810), .Z(n2702) );
  XOR U639 ( .A(n2895), .B(n2896), .Z(n2893) );
  XOR U640 ( .A(n2881), .B(n2882), .Z(n2880) );
  XOR U641 ( .A(n2697), .B(n2698), .Z(n2832) );
  XNOR U642 ( .A(n2538), .B(n2539), .Z(n2647) );
  XNOR U643 ( .A(n2661), .B(n2662), .Z(n2494) );
  NAND U644 ( .A(n12028), .B(n11998), .Z(n115) );
  XOR U645 ( .A(n11998), .B(n12028), .Z(n116) );
  NANDN U646 ( .A(n11999), .B(n116), .Z(n117) );
  NAND U647 ( .A(n115), .B(n117), .Z(n12010) );
  XOR U648 ( .A(n12016), .B(n12015), .Z(n12017) );
  XOR U649 ( .A(n12214), .B(n12215), .Z(n12192) );
  XOR U650 ( .A(n13801), .B(n13802), .Z(n13674) );
  XNOR U651 ( .A(n13961), .B(n13962), .Z(n13963) );
  XNOR U652 ( .A(n14108), .B(n14109), .Z(n14110) );
  XOR U653 ( .A(n14880), .B(n14881), .Z(n14879) );
  XOR U654 ( .A(n14657), .B(n14656), .Z(n14858) );
  XNOR U655 ( .A(n14622), .B(n14623), .Z(n14619) );
  NAND U656 ( .A(n9088), .B(n9058), .Z(n118) );
  XOR U657 ( .A(n9058), .B(n9088), .Z(n119) );
  NANDN U658 ( .A(n9059), .B(n119), .Z(n120) );
  NAND U659 ( .A(n118), .B(n120), .Z(n9070) );
  XNOR U660 ( .A(n9075), .B(n9076), .Z(n9078) );
  XOR U661 ( .A(n9274), .B(n9275), .Z(n9252) );
  XNOR U662 ( .A(n9676), .B(n9677), .Z(n9678) );
  XNOR U663 ( .A(n10195), .B(n10196), .Z(n10197) );
  XOR U664 ( .A(n10313), .B(n10314), .Z(n10316) );
  XNOR U665 ( .A(n10454), .B(n10455), .Z(n10456) );
  XOR U666 ( .A(n10859), .B(n10860), .Z(n10731) );
  XOR U667 ( .A(n11663), .B(n11664), .Z(n11650) );
  XOR U668 ( .A(n11937), .B(n11938), .Z(n11936) );
  OR U669 ( .A(n11625), .B(n11626), .Z(n121) );
  OR U670 ( .A(n11747), .B(n11624), .Z(n122) );
  NAND U671 ( .A(n121), .B(n122), .Z(n11702) );
  XOR U672 ( .A(n11705), .B(n11706), .Z(n11688) );
  XNOR U673 ( .A(n6126), .B(n6127), .Z(n6122) );
  XOR U674 ( .A(n6142), .B(n6141), .Z(n6143) );
  XNOR U675 ( .A(n6640), .B(n6641), .Z(n6642) );
  XNOR U676 ( .A(n6741), .B(n6742), .Z(n6743) );
  XNOR U677 ( .A(n7516), .B(n7517), .Z(n7518) );
  XOR U678 ( .A(n7659), .B(n7658), .Z(n7652) );
  XNOR U679 ( .A(n7785), .B(n7786), .Z(n7924) );
  XNOR U680 ( .A(n8711), .B(n8712), .Z(n8715) );
  XOR U681 ( .A(n8774), .B(n8773), .Z(n8982) );
  NAND U682 ( .A(n3202), .B(n3172), .Z(n123) );
  XOR U683 ( .A(n3172), .B(n3202), .Z(n124) );
  NANDN U684 ( .A(n3173), .B(n124), .Z(n125) );
  NAND U685 ( .A(n123), .B(n125), .Z(n3184) );
  XOR U686 ( .A(n3190), .B(n3189), .Z(n3191) );
  XNOR U687 ( .A(n3690), .B(n3691), .Z(n3692) );
  XNOR U688 ( .A(n3791), .B(n3792), .Z(n3793) );
  XOR U689 ( .A(n4733), .B(n4732), .Z(n4708) );
  XOR U690 ( .A(n4978), .B(n4979), .Z(n4850) );
  XNOR U691 ( .A(n5145), .B(n5146), .Z(n5147) );
  XNOR U692 ( .A(n5298), .B(n5299), .Z(n5300) );
  XNOR U693 ( .A(n6061), .B(n6062), .Z(n6059) );
  OR U694 ( .A(n5749), .B(n5750), .Z(n126) );
  OR U695 ( .A(n5921), .B(n5748), .Z(n127) );
  NAND U696 ( .A(n126), .B(n127), .Z(n5826) );
  XOR U697 ( .A(n5838), .B(n5837), .Z(n5812) );
  XNOR U698 ( .A(n211), .B(n212), .Z(n207) );
  XNOR U699 ( .A(n226), .B(n227), .Z(n228) );
  XOR U700 ( .A(n426), .B(n427), .Z(n404) );
  XNOR U701 ( .A(n583), .B(n584), .Z(n585) );
  XOR U702 ( .A(n662), .B(n663), .Z(n728) );
  XNOR U703 ( .A(n1347), .B(n1348), .Z(n1349) );
  XOR U704 ( .A(n1359), .B(n1360), .Z(n1362) );
  XOR U705 ( .A(n1873), .B(n1874), .Z(n2012) );
  XOR U706 ( .A(n3117), .B(n3118), .Z(n3116) );
  OR U707 ( .A(n2714), .B(n2715), .Z(n128) );
  OR U708 ( .A(n2927), .B(n2713), .Z(n129) );
  NAND U709 ( .A(n128), .B(n129), .Z(n2870) );
  XOR U710 ( .A(n2888), .B(n2887), .Z(n2862) );
  XNOR U711 ( .A(n2691), .B(n2692), .Z(n2838) );
  XOR U712 ( .A(n12072), .B(n12073), .Z(n12067) );
  XOR U713 ( .A(n13532), .B(n13533), .Z(n13527) );
  OR U714 ( .A(n14436), .B(n14437), .Z(n130) );
  NANDN U715 ( .A(n14434), .B(n14435), .Z(n131) );
  AND U716 ( .A(n130), .B(n131), .Z(n14602) );
  XOR U717 ( .A(n9132), .B(n9133), .Z(n9127) );
  XOR U718 ( .A(n10592), .B(n10593), .Z(n10587) );
  XOR U719 ( .A(n11175), .B(n11176), .Z(n11170) );
  OR U720 ( .A(n11507), .B(n11508), .Z(n132) );
  NANDN U721 ( .A(n11505), .B(n11506), .Z(n133) );
  AND U722 ( .A(n132), .B(n133), .Z(n11953) );
  XOR U723 ( .A(n6198), .B(n6199), .Z(n6193) );
  XOR U724 ( .A(n7263), .B(n7264), .Z(n7258) );
  XOR U725 ( .A(n8235), .B(n8236), .Z(n8230) );
  OR U726 ( .A(n8567), .B(n8568), .Z(n134) );
  NANDN U727 ( .A(n8565), .B(n8566), .Z(n135) );
  AND U728 ( .A(n134), .B(n135), .Z(n9013) );
  XOR U729 ( .A(n3246), .B(n3247), .Z(n3241) );
  NANDN U730 ( .A(n5632), .B(n5631), .Z(n136) );
  NANDN U731 ( .A(n5629), .B(n5630), .Z(n137) );
  AND U732 ( .A(n136), .B(n137), .Z(n6080) );
  XOR U733 ( .A(n283), .B(n284), .Z(n278) );
  XOR U734 ( .A(n1739), .B(n1740), .Z(n1734) );
  IV U735 ( .A(y[640]), .Z(n138) );
  IV U736 ( .A(y[641]), .Z(n139) );
  IV U737 ( .A(y[642]), .Z(n140) );
  IV U738 ( .A(y[643]), .Z(n141) );
  IV U739 ( .A(y[645]), .Z(n142) );
  IV U740 ( .A(y[647]), .Z(n143) );
  IV U741 ( .A(y[648]), .Z(n144) );
  IV U742 ( .A(y[675]), .Z(n145) );
  IV U743 ( .A(y[678]), .Z(n146) );
  IV U744 ( .A(y[707]), .Z(n147) );
  IV U745 ( .A(y[710]), .Z(n148) );
  IV U746 ( .A(y[739]), .Z(n149) );
  IV U747 ( .A(y[774]), .Z(n150) );
  IV U748 ( .A(x[128]), .Z(n151) );
  IV U749 ( .A(x[129]), .Z(n152) );
  IV U750 ( .A(x[130]), .Z(n153) );
  IV U751 ( .A(x[131]), .Z(n154) );
  IV U752 ( .A(x[132]), .Z(n155) );
  IV U753 ( .A(x[133]), .Z(n156) );
  IV U754 ( .A(x[134]), .Z(n157) );
  IV U755 ( .A(x[135]), .Z(n158) );
  IV U756 ( .A(x[136]), .Z(n159) );
  IV U757 ( .A(x[137]), .Z(n160) );
  IV U758 ( .A(x[138]), .Z(n161) );
  IV U759 ( .A(x[139]), .Z(n162) );
  IV U760 ( .A(x[140]), .Z(n163) );
  IV U761 ( .A(x[141]), .Z(n164) );
  IV U762 ( .A(x[142]), .Z(n165) );
  IV U763 ( .A(x[143]), .Z(n166) );
  IV U764 ( .A(x[144]), .Z(n167) );
  IV U765 ( .A(x[145]), .Z(n168) );
  IV U766 ( .A(x[146]), .Z(n169) );
  IV U767 ( .A(x[147]), .Z(n170) );
  IV U768 ( .A(x[148]), .Z(n171) );
  IV U769 ( .A(x[149]), .Z(n172) );
  IV U770 ( .A(x[150]), .Z(n173) );
  IV U771 ( .A(x[151]), .Z(n174) );
  IV U772 ( .A(x[152]), .Z(n175) );
  IV U773 ( .A(x[154]), .Z(n176) );
  IV U774 ( .A(x[155]), .Z(n177) );
  AND U775 ( .A(y[640]), .B(x[128]), .Z(n877) );
  XOR U776 ( .A(n877), .B(o[0]), .Z(N33) );
  AND U777 ( .A(x[129]), .B(y[640]), .Z(n178) );
  NAND U778 ( .A(y[641]), .B(x[128]), .Z(n184) );
  XNOR U779 ( .A(n184), .B(o[1]), .Z(n179) );
  XOR U780 ( .A(n178), .B(n179), .Z(n180) );
  AND U781 ( .A(o[0]), .B(n877), .Z(n181) );
  XOR U782 ( .A(n180), .B(n181), .Z(N34) );
  OR U783 ( .A(n179), .B(n178), .Z(n183) );
  NANDN U784 ( .A(n181), .B(n180), .Z(n182) );
  NAND U785 ( .A(n183), .B(n182), .Z(n186) );
  NAND U786 ( .A(x[128]), .B(y[642]), .Z(n197) );
  XOR U787 ( .A(n197), .B(o[2]), .Z(n185) );
  XNOR U788 ( .A(n186), .B(n185), .Z(n188) );
  ANDN U789 ( .B(o[1]), .A(n184), .Z(n191) );
  ANDN U790 ( .B(y[640]), .A(n153), .Z(n192) );
  XNOR U791 ( .A(n191), .B(n192), .Z(n194) );
  ANDN U792 ( .B(y[641]), .A(n152), .Z(n193) );
  XNOR U793 ( .A(n194), .B(n193), .Z(n187) );
  XNOR U794 ( .A(n188), .B(n187), .Z(N35) );
  NAND U795 ( .A(n186), .B(n185), .Z(n190) );
  OR U796 ( .A(n188), .B(n187), .Z(n189) );
  NAND U797 ( .A(n190), .B(n189), .Z(n200) );
  OR U798 ( .A(n192), .B(n191), .Z(n196) );
  OR U799 ( .A(n194), .B(n193), .Z(n195) );
  AND U800 ( .A(n196), .B(n195), .Z(n201) );
  XNOR U801 ( .A(n200), .B(n201), .Z(n202) );
  AND U802 ( .A(y[642]), .B(x[129]), .Z(n239) );
  NAND U803 ( .A(y[641]), .B(x[130]), .Z(n217) );
  XOR U804 ( .A(o[3]), .B(n217), .Z(n206) );
  XOR U805 ( .A(n239), .B(n206), .Z(n208) );
  NANDN U806 ( .A(n197), .B(o[2]), .Z(n212) );
  AND U807 ( .A(y[640]), .B(x[131]), .Z(n199) );
  NAND U808 ( .A(y[643]), .B(x[128]), .Z(n198) );
  XNOR U809 ( .A(n199), .B(n198), .Z(n211) );
  XNOR U810 ( .A(n208), .B(n207), .Z(n203) );
  XOR U811 ( .A(n202), .B(n203), .Z(N36) );
  NANDN U812 ( .A(n201), .B(n200), .Z(n205) );
  NANDN U813 ( .A(n203), .B(n202), .Z(n204) );
  NAND U814 ( .A(n205), .B(n204), .Z(n220) );
  NANDN U815 ( .A(n206), .B(n239), .Z(n210) );
  NANDN U816 ( .A(n208), .B(n207), .Z(n209) );
  NAND U817 ( .A(n210), .B(n209), .Z(n221) );
  XNOR U818 ( .A(n220), .B(n221), .Z(n222) );
  ANDN U819 ( .B(x[131]), .A(n141), .Z(n287) );
  NAND U820 ( .A(n877), .B(n287), .Z(n214) );
  NANDN U821 ( .A(n212), .B(n211), .Z(n213) );
  NAND U822 ( .A(n214), .B(n213), .Z(n226) );
  AND U823 ( .A(y[643]), .B(x[129]), .Z(n216) );
  NAND U824 ( .A(x[130]), .B(y[642]), .Z(n215) );
  XOR U825 ( .A(n216), .B(n215), .Z(n241) );
  NAND U826 ( .A(y[641]), .B(x[131]), .Z(n232) );
  XNOR U827 ( .A(n232), .B(o[4]), .Z(n240) );
  XOR U828 ( .A(n241), .B(n240), .Z(n227) );
  NANDN U829 ( .A(n217), .B(o[3]), .Z(n236) );
  AND U830 ( .A(y[640]), .B(x[132]), .Z(n219) );
  AND U831 ( .A(y[644]), .B(x[128]), .Z(n218) );
  XNOR U832 ( .A(n219), .B(n218), .Z(n235) );
  XOR U833 ( .A(n236), .B(n235), .Z(n229) );
  XOR U834 ( .A(n228), .B(n229), .Z(n223) );
  XOR U835 ( .A(n222), .B(n223), .Z(N37) );
  NANDN U836 ( .A(n221), .B(n220), .Z(n225) );
  NANDN U837 ( .A(n223), .B(n222), .Z(n224) );
  NAND U838 ( .A(n225), .B(n224), .Z(n244) );
  NANDN U839 ( .A(n227), .B(n226), .Z(n231) );
  NAND U840 ( .A(n229), .B(n228), .Z(n230) );
  NAND U841 ( .A(n231), .B(n230), .Z(n245) );
  XNOR U842 ( .A(n244), .B(n245), .Z(n246) );
  NANDN U843 ( .A(n232), .B(o[4]), .Z(n263) );
  AND U844 ( .A(x[128]), .B(y[645]), .Z(n234) );
  AND U845 ( .A(y[640]), .B(x[133]), .Z(n233) );
  XNOR U846 ( .A(n234), .B(n233), .Z(n262) );
  XOR U847 ( .A(n263), .B(n262), .Z(n258) );
  ANDN U848 ( .B(y[643]), .A(n153), .Z(n256) );
  IV U849 ( .A(y[644]), .Z(n2634) );
  ANDN U850 ( .B(x[129]), .A(n2634), .Z(n271) );
  ANDN U851 ( .B(x[132]), .A(n139), .Z(n266) );
  XOR U852 ( .A(o[5]), .B(n266), .Z(n269) );
  ANDN U853 ( .B(x[131]), .A(n140), .Z(n270) );
  XNOR U854 ( .A(n269), .B(n270), .Z(n272) );
  XNOR U855 ( .A(n271), .B(n272), .Z(n257) );
  XNOR U856 ( .A(n256), .B(n257), .Z(n259) );
  XNOR U857 ( .A(n258), .B(n259), .Z(n253) );
  ANDN U858 ( .B(x[132]), .A(n2634), .Z(n349) );
  NAND U859 ( .A(n877), .B(n349), .Z(n238) );
  OR U860 ( .A(n236), .B(n235), .Z(n237) );
  NAND U861 ( .A(n238), .B(n237), .Z(n251) );
  NAND U862 ( .A(n239), .B(n256), .Z(n243) );
  NANDN U863 ( .A(n241), .B(n240), .Z(n242) );
  NAND U864 ( .A(n243), .B(n242), .Z(n250) );
  XNOR U865 ( .A(n251), .B(n250), .Z(n252) );
  XNOR U866 ( .A(n253), .B(n252), .Z(n247) );
  XOR U867 ( .A(n246), .B(n247), .Z(N38) );
  NANDN U868 ( .A(n245), .B(n244), .Z(n249) );
  NANDN U869 ( .A(n247), .B(n246), .Z(n248) );
  NAND U870 ( .A(n249), .B(n248), .Z(n275) );
  OR U871 ( .A(n251), .B(n250), .Z(n255) );
  OR U872 ( .A(n253), .B(n252), .Z(n254) );
  AND U873 ( .A(n255), .B(n254), .Z(n276) );
  XNOR U874 ( .A(n275), .B(n276), .Z(n277) );
  OR U875 ( .A(n257), .B(n256), .Z(n261) );
  OR U876 ( .A(n259), .B(n258), .Z(n260) );
  AND U877 ( .A(n261), .B(n260), .Z(n281) );
  NAND U878 ( .A(x[133]), .B(y[645]), .Z(n617) );
  NANDN U879 ( .A(n617), .B(n877), .Z(n265) );
  OR U880 ( .A(n263), .B(n262), .Z(n264) );
  NAND U881 ( .A(n265), .B(n264), .Z(n303) );
  NAND U882 ( .A(n266), .B(o[5]), .Z(n293) );
  AND U883 ( .A(y[646]), .B(x[128]), .Z(n268) );
  AND U884 ( .A(y[640]), .B(x[134]), .Z(n267) );
  XNOR U885 ( .A(n268), .B(n267), .Z(n292) );
  XOR U886 ( .A(n293), .B(n292), .Z(n302) );
  XNOR U887 ( .A(n303), .B(n302), .Z(n305) );
  AND U888 ( .A(y[645]), .B(x[129]), .Z(n560) );
  NAND U889 ( .A(y[641]), .B(x[133]), .Z(n296) );
  XNOR U890 ( .A(n296), .B(o[6]), .Z(n297) );
  XNOR U891 ( .A(n560), .B(n297), .Z(n299) );
  AND U892 ( .A(x[132]), .B(y[642]), .Z(n298) );
  XOR U893 ( .A(n299), .B(n298), .Z(n288) );
  AND U894 ( .A(x[130]), .B(y[644]), .Z(n607) );
  XNOR U895 ( .A(n287), .B(n607), .Z(n289) );
  XOR U896 ( .A(n288), .B(n289), .Z(n304) );
  XNOR U897 ( .A(n305), .B(n304), .Z(n282) );
  XOR U898 ( .A(n281), .B(n282), .Z(n283) );
  OR U899 ( .A(n270), .B(n269), .Z(n274) );
  OR U900 ( .A(n272), .B(n271), .Z(n273) );
  AND U901 ( .A(n274), .B(n273), .Z(n284) );
  XOR U902 ( .A(n277), .B(n278), .Z(N39) );
  NANDN U903 ( .A(n276), .B(n275), .Z(n280) );
  NANDN U904 ( .A(n278), .B(n277), .Z(n279) );
  NAND U905 ( .A(n280), .B(n279), .Z(n337) );
  OR U906 ( .A(n282), .B(n281), .Z(n286) );
  NANDN U907 ( .A(n284), .B(n283), .Z(n285) );
  AND U908 ( .A(n286), .B(n285), .Z(n338) );
  XNOR U909 ( .A(n337), .B(n338), .Z(n339) );
  OR U910 ( .A(n287), .B(n607), .Z(n291) );
  NANDN U911 ( .A(n289), .B(n288), .Z(n290) );
  NAND U912 ( .A(n291), .B(n290), .Z(n334) );
  AND U913 ( .A(x[134]), .B(y[646]), .Z(n576) );
  NAND U914 ( .A(n877), .B(n576), .Z(n295) );
  OR U915 ( .A(n293), .B(n292), .Z(n294) );
  AND U916 ( .A(n295), .B(n294), .Z(n332) );
  ANDN U917 ( .B(y[642]), .A(n156), .Z(n464) );
  AND U918 ( .A(y[646]), .B(x[129]), .Z(n687) );
  NAND U919 ( .A(y[641]), .B(x[134]), .Z(n320) );
  XNOR U920 ( .A(o[7]), .B(n320), .Z(n321) );
  XNOR U921 ( .A(n687), .B(n321), .Z(n322) );
  XNOR U922 ( .A(n464), .B(n322), .Z(n331) );
  XOR U923 ( .A(n332), .B(n331), .Z(n333) );
  XNOR U924 ( .A(n334), .B(n333), .Z(n343) );
  ANDN U925 ( .B(y[645]), .A(n153), .Z(n749) );
  ANDN U926 ( .B(x[132]), .A(n141), .Z(n475) );
  ANDN U927 ( .B(x[131]), .A(n2634), .Z(n316) );
  XNOR U928 ( .A(n475), .B(n316), .Z(n317) );
  XOR U929 ( .A(n749), .B(n317), .Z(n325) );
  NAND U930 ( .A(x[128]), .B(y[647]), .Z(n312) );
  ANDN U931 ( .B(o[6]), .A(n296), .Z(n311) );
  NAND U932 ( .A(y[640]), .B(x[135]), .Z(n310) );
  XOR U933 ( .A(n311), .B(n310), .Z(n313) );
  XNOR U934 ( .A(n312), .B(n313), .Z(n326) );
  XNOR U935 ( .A(n325), .B(n326), .Z(n328) );
  NAND U936 ( .A(n560), .B(n297), .Z(n301) );
  NANDN U937 ( .A(n299), .B(n298), .Z(n300) );
  AND U938 ( .A(n301), .B(n300), .Z(n327) );
  XOR U939 ( .A(n328), .B(n327), .Z(n344) );
  XOR U940 ( .A(n343), .B(n344), .Z(n346) );
  OR U941 ( .A(n303), .B(n302), .Z(n307) );
  OR U942 ( .A(n305), .B(n304), .Z(n306) );
  AND U943 ( .A(n307), .B(n306), .Z(n345) );
  XOR U944 ( .A(n346), .B(n345), .Z(n340) );
  XNOR U945 ( .A(n339), .B(n340), .Z(N40) );
  AND U946 ( .A(x[128]), .B(y[648]), .Z(n309) );
  NAND U947 ( .A(y[640]), .B(x[136]), .Z(n308) );
  XOR U948 ( .A(n309), .B(n308), .Z(n358) );
  NAND U949 ( .A(x[135]), .B(y[641]), .Z(n361) );
  XOR U950 ( .A(n361), .B(o[8]), .Z(n357) );
  XNOR U951 ( .A(n358), .B(n357), .Z(n379) );
  NANDN U952 ( .A(n311), .B(n310), .Z(n315) );
  NANDN U953 ( .A(n313), .B(n312), .Z(n314) );
  NAND U954 ( .A(n315), .B(n314), .Z(n378) );
  XOR U955 ( .A(n379), .B(n378), .Z(n380) );
  OR U956 ( .A(n316), .B(n475), .Z(n319) );
  OR U957 ( .A(n317), .B(n749), .Z(n318) );
  NAND U958 ( .A(n319), .B(n318), .Z(n381) );
  XNOR U959 ( .A(n380), .B(n381), .Z(n392) );
  ANDN U960 ( .B(x[134]), .A(n140), .Z(n350) );
  XNOR U961 ( .A(n349), .B(n350), .Z(n351) );
  IV U962 ( .A(y[646]), .Z(n2618) );
  NOR U963 ( .A(n153), .B(n2618), .Z(n859) );
  XNOR U964 ( .A(n351), .B(n859), .Z(n352) );
  ANDN U965 ( .B(x[131]), .A(n142), .Z(n1173) );
  XNOR U966 ( .A(n352), .B(n1173), .Z(n354) );
  NANDN U967 ( .A(n320), .B(o[7]), .Z(n369) );
  AND U968 ( .A(y[643]), .B(x[133]), .Z(n959) );
  AND U969 ( .A(y[647]), .B(x[129]), .Z(n872) );
  XNOR U970 ( .A(n959), .B(n872), .Z(n368) );
  XOR U971 ( .A(n369), .B(n368), .Z(n353) );
  XNOR U972 ( .A(n354), .B(n353), .Z(n372) );
  NAND U973 ( .A(n687), .B(n321), .Z(n324) );
  NANDN U974 ( .A(n322), .B(n464), .Z(n323) );
  AND U975 ( .A(n324), .B(n323), .Z(n373) );
  XOR U976 ( .A(n372), .B(n373), .Z(n375) );
  OR U977 ( .A(n326), .B(n325), .Z(n330) );
  OR U978 ( .A(n328), .B(n327), .Z(n329) );
  AND U979 ( .A(n330), .B(n329), .Z(n374) );
  XOR U980 ( .A(n375), .B(n374), .Z(n390) );
  NANDN U981 ( .A(n332), .B(n331), .Z(n336) );
  OR U982 ( .A(n334), .B(n333), .Z(n335) );
  NAND U983 ( .A(n336), .B(n335), .Z(n391) );
  XNOR U984 ( .A(n390), .B(n391), .Z(n393) );
  XNOR U985 ( .A(n392), .B(n393), .Z(n387) );
  NANDN U986 ( .A(n338), .B(n337), .Z(n342) );
  NAND U987 ( .A(n340), .B(n339), .Z(n341) );
  NAND U988 ( .A(n342), .B(n341), .Z(n384) );
  NANDN U989 ( .A(n344), .B(n343), .Z(n348) );
  OR U990 ( .A(n346), .B(n345), .Z(n347) );
  AND U991 ( .A(n348), .B(n347), .Z(n385) );
  XNOR U992 ( .A(n384), .B(n385), .Z(n386) );
  XOR U993 ( .A(n387), .B(n386), .Z(N41) );
  OR U994 ( .A(n352), .B(n1173), .Z(n356) );
  OR U995 ( .A(n354), .B(n353), .Z(n355) );
  NAND U996 ( .A(n356), .B(n355), .Z(n424) );
  XOR U997 ( .A(n425), .B(n424), .Z(n426) );
  AND U998 ( .A(y[648]), .B(x[136]), .Z(n866) );
  NAND U999 ( .A(n877), .B(n866), .Z(n360) );
  OR U1000 ( .A(n358), .B(n357), .Z(n359) );
  NAND U1001 ( .A(n360), .B(n359), .Z(n411) );
  NANDN U1002 ( .A(n361), .B(o[8]), .Z(n440) );
  AND U1003 ( .A(x[135]), .B(y[642]), .Z(n754) );
  NAND U1004 ( .A(y[644]), .B(x[133]), .Z(n362) );
  XNOR U1005 ( .A(n754), .B(n362), .Z(n439) );
  XNOR U1006 ( .A(n440), .B(n439), .Z(n409) );
  AND U1007 ( .A(x[128]), .B(y[649]), .Z(n364) );
  NAND U1008 ( .A(y[640]), .B(x[137]), .Z(n363) );
  XOR U1009 ( .A(n364), .B(n363), .Z(n436) );
  NAND U1010 ( .A(y[641]), .B(x[136]), .Z(n430) );
  XOR U1011 ( .A(n430), .B(o[9]), .Z(n435) );
  XNOR U1012 ( .A(n436), .B(n435), .Z(n408) );
  XOR U1013 ( .A(n409), .B(n408), .Z(n410) );
  XNOR U1014 ( .A(n411), .B(n410), .Z(n420) );
  AND U1015 ( .A(y[645]), .B(x[132]), .Z(n884) );
  AND U1016 ( .A(x[129]), .B(y[648]), .Z(n366) );
  NAND U1017 ( .A(y[643]), .B(x[134]), .Z(n365) );
  XNOR U1018 ( .A(n366), .B(n365), .Z(n432) );
  XOR U1019 ( .A(n884), .B(n432), .Z(n414) );
  ANDN U1020 ( .B(y[647]), .A(n153), .Z(n1052) );
  NAND U1021 ( .A(x[131]), .B(y[646]), .Z(n794) );
  XOR U1022 ( .A(n1052), .B(n794), .Z(n415) );
  XNOR U1023 ( .A(n414), .B(n415), .Z(n418) );
  NAND U1024 ( .A(y[643]), .B(x[129]), .Z(n431) );
  AND U1025 ( .A(x[133]), .B(y[647]), .Z(n367) );
  NANDN U1026 ( .A(n431), .B(n367), .Z(n371) );
  OR U1027 ( .A(n369), .B(n368), .Z(n370) );
  AND U1028 ( .A(n371), .B(n370), .Z(n419) );
  XOR U1029 ( .A(n418), .B(n419), .Z(n421) );
  XOR U1030 ( .A(n420), .B(n421), .Z(n427) );
  NANDN U1031 ( .A(n373), .B(n372), .Z(n377) );
  OR U1032 ( .A(n375), .B(n374), .Z(n376) );
  NAND U1033 ( .A(n377), .B(n376), .Z(n403) );
  OR U1034 ( .A(n379), .B(n378), .Z(n383) );
  NANDN U1035 ( .A(n381), .B(n380), .Z(n382) );
  NAND U1036 ( .A(n383), .B(n382), .Z(n402) );
  XOR U1037 ( .A(n403), .B(n402), .Z(n405) );
  XNOR U1038 ( .A(n404), .B(n405), .Z(n399) );
  NANDN U1039 ( .A(n385), .B(n384), .Z(n389) );
  NANDN U1040 ( .A(n387), .B(n386), .Z(n388) );
  NAND U1041 ( .A(n389), .B(n388), .Z(n396) );
  OR U1042 ( .A(n391), .B(n390), .Z(n395) );
  OR U1043 ( .A(n393), .B(n392), .Z(n394) );
  AND U1044 ( .A(n395), .B(n394), .Z(n397) );
  XNOR U1045 ( .A(n396), .B(n397), .Z(n398) );
  XOR U1046 ( .A(n399), .B(n398), .Z(N42) );
  NANDN U1047 ( .A(n397), .B(n396), .Z(n401) );
  NANDN U1048 ( .A(n399), .B(n398), .Z(n400) );
  NAND U1049 ( .A(n401), .B(n400), .Z(n445) );
  OR U1050 ( .A(n403), .B(n402), .Z(n407) );
  NAND U1051 ( .A(n405), .B(n404), .Z(n406) );
  AND U1052 ( .A(n407), .B(n406), .Z(n446) );
  XNOR U1053 ( .A(n445), .B(n446), .Z(n447) );
  NANDN U1054 ( .A(n409), .B(n408), .Z(n413) );
  OR U1055 ( .A(n411), .B(n410), .Z(n412) );
  NAND U1056 ( .A(n413), .B(n412), .Z(n503) );
  NANDN U1057 ( .A(n1052), .B(n794), .Z(n417) );
  OR U1058 ( .A(n415), .B(n414), .Z(n416) );
  NAND U1059 ( .A(n417), .B(n416), .Z(n502) );
  XOR U1060 ( .A(n503), .B(n502), .Z(n504) );
  NANDN U1061 ( .A(n419), .B(n418), .Z(n423) );
  NANDN U1062 ( .A(n421), .B(n420), .Z(n422) );
  AND U1063 ( .A(n423), .B(n422), .Z(n505) );
  XNOR U1064 ( .A(n504), .B(n505), .Z(n453) );
  OR U1065 ( .A(n425), .B(n424), .Z(n429) );
  NANDN U1066 ( .A(n427), .B(n426), .Z(n428) );
  NAND U1067 ( .A(n429), .B(n428), .Z(n452) );
  NAND U1068 ( .A(y[650]), .B(x[128]), .Z(n481) );
  NANDN U1069 ( .A(n430), .B(o[9]), .Z(n479) );
  NAND U1070 ( .A(x[138]), .B(y[640]), .Z(n480) );
  XNOR U1071 ( .A(n479), .B(n480), .Z(n482) );
  XNOR U1072 ( .A(n481), .B(n482), .Z(n472) );
  ANDN U1073 ( .B(y[649]), .A(n152), .Z(n1395) );
  ANDN U1074 ( .B(x[131]), .A(n143), .Z(n1425) );
  NANDN U1075 ( .A(n144), .B(x[130]), .Z(n460) );
  XNOR U1076 ( .A(n1425), .B(n460), .Z(n461) );
  XNOR U1077 ( .A(n1395), .B(n461), .Z(n470) );
  ANDN U1078 ( .B(x[134]), .A(n144), .Z(n767) );
  NANDN U1079 ( .A(n431), .B(n767), .Z(n434) );
  NAND U1080 ( .A(n432), .B(n884), .Z(n433) );
  AND U1081 ( .A(n434), .B(n433), .Z(n469) );
  XOR U1082 ( .A(n470), .B(n469), .Z(n471) );
  XNOR U1083 ( .A(n472), .B(n471), .Z(n496) );
  AND U1084 ( .A(x[137]), .B(y[649]), .Z(n1021) );
  NAND U1085 ( .A(n877), .B(n1021), .Z(n438) );
  OR U1086 ( .A(n436), .B(n435), .Z(n437) );
  NAND U1087 ( .A(n438), .B(n437), .Z(n497) );
  XNOR U1088 ( .A(n496), .B(n497), .Z(n499) );
  ANDN U1089 ( .B(x[135]), .A(n2634), .Z(n570) );
  NAND U1090 ( .A(n570), .B(n464), .Z(n442) );
  NANDN U1091 ( .A(n440), .B(n439), .Z(n441) );
  NAND U1092 ( .A(n442), .B(n441), .Z(n493) );
  ANDN U1093 ( .B(x[134]), .A(n2634), .Z(n704) );
  AND U1094 ( .A(x[132]), .B(y[646]), .Z(n444) );
  NAND U1095 ( .A(y[643]), .B(x[135]), .Z(n443) );
  XOR U1096 ( .A(n444), .B(n443), .Z(n476) );
  XOR U1097 ( .A(n704), .B(n476), .Z(n490) );
  AND U1098 ( .A(x[136]), .B(y[642]), .Z(n569) );
  XOR U1099 ( .A(n569), .B(n617), .Z(n466) );
  NAND U1100 ( .A(x[137]), .B(y[641]), .Z(n487) );
  XOR U1101 ( .A(o[10]), .B(n487), .Z(n465) );
  XOR U1102 ( .A(n466), .B(n465), .Z(n491) );
  XNOR U1103 ( .A(n490), .B(n491), .Z(n492) );
  XOR U1104 ( .A(n493), .B(n492), .Z(n498) );
  XOR U1105 ( .A(n499), .B(n498), .Z(n451) );
  XOR U1106 ( .A(n452), .B(n451), .Z(n454) );
  XNOR U1107 ( .A(n453), .B(n454), .Z(n448) );
  XOR U1108 ( .A(n447), .B(n448), .Z(N43) );
  NANDN U1109 ( .A(n446), .B(n445), .Z(n450) );
  NANDN U1110 ( .A(n448), .B(n447), .Z(n449) );
  NAND U1111 ( .A(n450), .B(n449), .Z(n508) );
  NANDN U1112 ( .A(n452), .B(n451), .Z(n456) );
  OR U1113 ( .A(n454), .B(n453), .Z(n455) );
  AND U1114 ( .A(n456), .B(n455), .Z(n509) );
  XNOR U1115 ( .A(n508), .B(n509), .Z(n510) );
  AND U1116 ( .A(x[131]), .B(y[648]), .Z(n1557) );
  NAND U1117 ( .A(y[647]), .B(x[132]), .Z(n557) );
  AND U1118 ( .A(x[133]), .B(y[646]), .Z(n458) );
  NAND U1119 ( .A(x[130]), .B(y[649]), .Z(n457) );
  XOR U1120 ( .A(n458), .B(n457), .Z(n556) );
  XNOR U1121 ( .A(n557), .B(n556), .Z(n526) );
  XOR U1122 ( .A(n1557), .B(n526), .Z(n528) );
  AND U1123 ( .A(x[137]), .B(y[642]), .Z(n645) );
  NAND U1124 ( .A(y[643]), .B(x[136]), .Z(n459) );
  XNOR U1125 ( .A(n645), .B(n459), .Z(n571) );
  XNOR U1126 ( .A(n570), .B(n571), .Z(n527) );
  XNOR U1127 ( .A(n528), .B(n527), .Z(n546) );
  NANDN U1128 ( .A(n1425), .B(n460), .Z(n463) );
  NANDN U1129 ( .A(n1395), .B(n461), .Z(n462) );
  NAND U1130 ( .A(n463), .B(n462), .Z(n543) );
  ANDN U1131 ( .B(y[645]), .A(n159), .Z(n1313) );
  NAND U1132 ( .A(n1313), .B(n464), .Z(n468) );
  OR U1133 ( .A(n466), .B(n465), .Z(n467) );
  NAND U1134 ( .A(n468), .B(n467), .Z(n544) );
  XOR U1135 ( .A(n546), .B(n545), .Z(n539) );
  OR U1136 ( .A(n470), .B(n469), .Z(n474) );
  NANDN U1137 ( .A(n472), .B(n471), .Z(n473) );
  NAND U1138 ( .A(n474), .B(n473), .Z(n523) );
  AND U1139 ( .A(y[646]), .B(x[135]), .Z(n615) );
  NAND U1140 ( .A(n615), .B(n475), .Z(n478) );
  NANDN U1141 ( .A(n476), .B(n704), .Z(n477) );
  NAND U1142 ( .A(n478), .B(n477), .Z(n521) );
  NAND U1143 ( .A(n480), .B(n479), .Z(n484) );
  NANDN U1144 ( .A(n482), .B(n481), .Z(n483) );
  NAND U1145 ( .A(n484), .B(n483), .Z(n534) );
  AND U1146 ( .A(x[134]), .B(y[645]), .Z(n486) );
  NAND U1147 ( .A(x[129]), .B(y[650]), .Z(n485) );
  XOR U1148 ( .A(n486), .B(n485), .Z(n562) );
  NAND U1149 ( .A(x[138]), .B(y[641]), .Z(n574) );
  XOR U1150 ( .A(o[11]), .B(n574), .Z(n561) );
  XOR U1151 ( .A(n562), .B(n561), .Z(n531) );
  NANDN U1152 ( .A(n487), .B(o[10]), .Z(n566) );
  AND U1153 ( .A(x[128]), .B(y[651]), .Z(n489) );
  NAND U1154 ( .A(y[640]), .B(x[139]), .Z(n488) );
  XNOR U1155 ( .A(n489), .B(n488), .Z(n565) );
  XOR U1156 ( .A(n531), .B(n532), .Z(n533) );
  XOR U1157 ( .A(n534), .B(n533), .Z(n520) );
  XNOR U1158 ( .A(n521), .B(n520), .Z(n522) );
  XNOR U1159 ( .A(n523), .B(n522), .Z(n537) );
  NANDN U1160 ( .A(n491), .B(n490), .Z(n495) );
  NANDN U1161 ( .A(n493), .B(n492), .Z(n494) );
  NAND U1162 ( .A(n495), .B(n494), .Z(n538) );
  XOR U1163 ( .A(n537), .B(n538), .Z(n540) );
  XOR U1164 ( .A(n539), .B(n540), .Z(n514) );
  OR U1165 ( .A(n497), .B(n496), .Z(n501) );
  OR U1166 ( .A(n499), .B(n498), .Z(n500) );
  AND U1167 ( .A(n501), .B(n500), .Z(n515) );
  XNOR U1168 ( .A(n514), .B(n515), .Z(n517) );
  OR U1169 ( .A(n503), .B(n502), .Z(n507) );
  NANDN U1170 ( .A(n505), .B(n504), .Z(n506) );
  NAND U1171 ( .A(n507), .B(n506), .Z(n516) );
  XOR U1172 ( .A(n517), .B(n516), .Z(n511) );
  XNOR U1173 ( .A(n510), .B(n511), .Z(N44) );
  NANDN U1174 ( .A(n509), .B(n508), .Z(n513) );
  NAND U1175 ( .A(n511), .B(n510), .Z(n512) );
  NAND U1176 ( .A(n513), .B(n512), .Z(n577) );
  OR U1177 ( .A(n515), .B(n514), .Z(n519) );
  OR U1178 ( .A(n517), .B(n516), .Z(n518) );
  AND U1179 ( .A(n519), .B(n518), .Z(n578) );
  XNOR U1180 ( .A(n577), .B(n578), .Z(n579) );
  OR U1181 ( .A(n521), .B(n520), .Z(n525) );
  OR U1182 ( .A(n523), .B(n522), .Z(n524) );
  AND U1183 ( .A(n525), .B(n524), .Z(n592) );
  NANDN U1184 ( .A(n526), .B(n1557), .Z(n530) );
  OR U1185 ( .A(n528), .B(n527), .Z(n529) );
  NAND U1186 ( .A(n530), .B(n529), .Z(n590) );
  NANDN U1187 ( .A(n532), .B(n531), .Z(n536) );
  OR U1188 ( .A(n534), .B(n533), .Z(n535) );
  NAND U1189 ( .A(n536), .B(n535), .Z(n589) );
  XOR U1190 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U1191 ( .A(n592), .B(n591), .Z(n586) );
  NANDN U1192 ( .A(n538), .B(n537), .Z(n542) );
  OR U1193 ( .A(n540), .B(n539), .Z(n541) );
  NAND U1194 ( .A(n542), .B(n541), .Z(n583) );
  NANDN U1195 ( .A(n544), .B(n543), .Z(n548) );
  NAND U1196 ( .A(n546), .B(n545), .Z(n547) );
  NAND U1197 ( .A(n548), .B(n547), .Z(n598) );
  AND U1198 ( .A(x[135]), .B(y[645]), .Z(n550) );
  NAND U1199 ( .A(y[647]), .B(x[133]), .Z(n549) );
  XOR U1200 ( .A(n550), .B(n549), .Z(n619) );
  AND U1201 ( .A(x[138]), .B(y[642]), .Z(n551) );
  NAND U1202 ( .A(y[643]), .B(x[137]), .Z(n1250) );
  XOR U1203 ( .A(n551), .B(n1250), .Z(n647) );
  NAND U1204 ( .A(x[132]), .B(y[648]), .Z(n646) );
  XNOR U1205 ( .A(n647), .B(n646), .Z(n618) );
  XOR U1206 ( .A(n619), .B(n618), .Z(n624) );
  AND U1207 ( .A(y[640]), .B(x[140]), .Z(n553) );
  NAND U1208 ( .A(y[652]), .B(x[128]), .Z(n552) );
  XOR U1209 ( .A(n553), .B(n552), .Z(n639) );
  NAND U1210 ( .A(x[139]), .B(y[641]), .Z(n613) );
  XOR U1211 ( .A(o[12]), .B(n613), .Z(n638) );
  XOR U1212 ( .A(n639), .B(n638), .Z(n622) );
  AND U1213 ( .A(y[644]), .B(x[136]), .Z(n555) );
  NAND U1214 ( .A(x[130]), .B(y[650]), .Z(n554) );
  XOR U1215 ( .A(n555), .B(n554), .Z(n609) );
  NAND U1216 ( .A(x[131]), .B(y[649]), .Z(n608) );
  XNOR U1217 ( .A(n609), .B(n608), .Z(n623) );
  XOR U1218 ( .A(n622), .B(n623), .Z(n625) );
  ANDN U1219 ( .B(y[649]), .A(n156), .Z(n795) );
  NAND U1220 ( .A(n859), .B(n795), .Z(n559) );
  OR U1221 ( .A(n557), .B(n556), .Z(n558) );
  NAND U1222 ( .A(n559), .B(n558), .Z(n602) );
  AND U1223 ( .A(x[134]), .B(y[650]), .Z(n883) );
  NAND U1224 ( .A(n883), .B(n560), .Z(n564) );
  OR U1225 ( .A(n562), .B(n561), .Z(n563) );
  NAND U1226 ( .A(n564), .B(n563), .Z(n601) );
  XOR U1227 ( .A(n602), .B(n601), .Z(n604) );
  XNOR U1228 ( .A(n603), .B(n604), .Z(n595) );
  AND U1229 ( .A(y[651]), .B(x[139]), .Z(n1682) );
  NAND U1230 ( .A(n877), .B(n1682), .Z(n568) );
  NANDN U1231 ( .A(n566), .B(n565), .Z(n567) );
  NAND U1232 ( .A(n568), .B(n567), .Z(n630) );
  NANDN U1233 ( .A(n1250), .B(n569), .Z(n573) );
  NAND U1234 ( .A(n571), .B(n570), .Z(n572) );
  NAND U1235 ( .A(n573), .B(n572), .Z(n628) );
  NANDN U1236 ( .A(n574), .B(o[11]), .Z(n635) );
  NAND U1237 ( .A(x[129]), .B(y[651]), .Z(n575) );
  XNOR U1238 ( .A(n576), .B(n575), .Z(n634) );
  XOR U1239 ( .A(n628), .B(n629), .Z(n631) );
  XOR U1240 ( .A(n630), .B(n631), .Z(n596) );
  XNOR U1241 ( .A(n595), .B(n596), .Z(n597) );
  XOR U1242 ( .A(n598), .B(n597), .Z(n584) );
  XNOR U1243 ( .A(n586), .B(n585), .Z(n580) );
  XOR U1244 ( .A(n579), .B(n580), .Z(N45) );
  NANDN U1245 ( .A(n578), .B(n577), .Z(n582) );
  NANDN U1246 ( .A(n580), .B(n579), .Z(n581) );
  NAND U1247 ( .A(n582), .B(n581), .Z(n719) );
  NANDN U1248 ( .A(n584), .B(n583), .Z(n588) );
  NANDN U1249 ( .A(n586), .B(n585), .Z(n587) );
  NAND U1250 ( .A(n588), .B(n587), .Z(n720) );
  XNOR U1251 ( .A(n719), .B(n720), .Z(n721) );
  OR U1252 ( .A(n590), .B(n589), .Z(n594) );
  NANDN U1253 ( .A(n592), .B(n591), .Z(n593) );
  AND U1254 ( .A(n594), .B(n593), .Z(n725) );
  NANDN U1255 ( .A(n596), .B(n595), .Z(n600) );
  NANDN U1256 ( .A(n598), .B(n597), .Z(n599) );
  NAND U1257 ( .A(n600), .B(n599), .Z(n726) );
  XOR U1258 ( .A(n725), .B(n726), .Z(n727) );
  OR U1259 ( .A(n602), .B(n601), .Z(n606) );
  NAND U1260 ( .A(n604), .B(n603), .Z(n605) );
  AND U1261 ( .A(n606), .B(n605), .Z(n660) );
  AND U1262 ( .A(x[136]), .B(y[650]), .Z(n1032) );
  NAND U1263 ( .A(n1032), .B(n607), .Z(n611) );
  OR U1264 ( .A(n609), .B(n608), .Z(n610) );
  NAND U1265 ( .A(n611), .B(n610), .Z(n681) );
  NAND U1266 ( .A(x[130]), .B(y[651]), .Z(n706) );
  AND U1267 ( .A(y[647]), .B(x[134]), .Z(n612) );
  AND U1268 ( .A(y[644]), .B(x[137]), .Z(n1136) );
  XNOR U1269 ( .A(n612), .B(n1136), .Z(n705) );
  XOR U1270 ( .A(n706), .B(n705), .Z(n679) );
  NANDN U1271 ( .A(n613), .B(o[12]), .Z(n690) );
  NAND U1272 ( .A(y[652]), .B(x[129]), .Z(n614) );
  XNOR U1273 ( .A(n615), .B(n614), .Z(n689) );
  XNOR U1274 ( .A(n681), .B(n680), .Z(n655) );
  AND U1275 ( .A(x[135]), .B(y[647]), .Z(n616) );
  NANDN U1276 ( .A(n617), .B(n616), .Z(n621) );
  OR U1277 ( .A(n619), .B(n618), .Z(n620) );
  AND U1278 ( .A(n621), .B(n620), .Z(n654) );
  XOR U1279 ( .A(n655), .B(n654), .Z(n656) );
  NANDN U1280 ( .A(n623), .B(n622), .Z(n627) );
  NANDN U1281 ( .A(n625), .B(n624), .Z(n626) );
  AND U1282 ( .A(n627), .B(n626), .Z(n657) );
  XNOR U1283 ( .A(n656), .B(n657), .Z(n661) );
  XOR U1284 ( .A(n660), .B(n661), .Z(n662) );
  NANDN U1285 ( .A(n629), .B(n628), .Z(n633) );
  NANDN U1286 ( .A(n631), .B(n630), .Z(n632) );
  NAND U1287 ( .A(n633), .B(n632), .Z(n669) );
  ANDN U1288 ( .B(y[651]), .A(n157), .Z(n1059) );
  NAND U1289 ( .A(n687), .B(n1059), .Z(n637) );
  NANDN U1290 ( .A(n635), .B(n634), .Z(n636) );
  NAND U1291 ( .A(n637), .B(n636), .Z(n674) );
  ANDN U1292 ( .B(y[652]), .A(n163), .Z(n1980) );
  NAND U1293 ( .A(n1980), .B(n877), .Z(n641) );
  OR U1294 ( .A(n639), .B(n638), .Z(n640) );
  NAND U1295 ( .A(n641), .B(n640), .Z(n672) );
  AND U1296 ( .A(y[642]), .B(x[139]), .Z(n643) );
  NAND U1297 ( .A(y[643]), .B(x[138]), .Z(n642) );
  XNOR U1298 ( .A(n643), .B(n642), .Z(n693) );
  XNOR U1299 ( .A(n1313), .B(n693), .Z(n673) );
  XOR U1300 ( .A(n674), .B(n675), .Z(n666) );
  AND U1301 ( .A(x[138]), .B(y[643]), .Z(n644) );
  NAND U1302 ( .A(n645), .B(n644), .Z(n649) );
  OR U1303 ( .A(n647), .B(n646), .Z(n648) );
  NAND U1304 ( .A(n649), .B(n648), .Z(n716) );
  AND U1305 ( .A(x[128]), .B(y[653]), .Z(n651) );
  NAND U1306 ( .A(y[640]), .B(x[141]), .Z(n650) );
  XOR U1307 ( .A(n651), .B(n650), .Z(n701) );
  NAND U1308 ( .A(x[140]), .B(y[641]), .Z(n710) );
  XOR U1309 ( .A(o[13]), .B(n710), .Z(n700) );
  XOR U1310 ( .A(n701), .B(n700), .Z(n714) );
  AND U1311 ( .A(x[133]), .B(y[648]), .Z(n653) );
  NAND U1312 ( .A(y[650]), .B(x[131]), .Z(n652) );
  XOR U1313 ( .A(n653), .B(n652), .Z(n697) );
  NAND U1314 ( .A(y[649]), .B(x[132]), .Z(n696) );
  XOR U1315 ( .A(n697), .B(n696), .Z(n713) );
  XOR U1316 ( .A(n716), .B(n715), .Z(n667) );
  XNOR U1317 ( .A(n666), .B(n667), .Z(n668) );
  XOR U1318 ( .A(n669), .B(n668), .Z(n663) );
  XOR U1319 ( .A(n727), .B(n728), .Z(n722) );
  XOR U1320 ( .A(n721), .B(n722), .Z(N46) );
  OR U1321 ( .A(n655), .B(n654), .Z(n659) );
  NANDN U1322 ( .A(n657), .B(n656), .Z(n658) );
  NAND U1323 ( .A(n659), .B(n658), .Z(n740) );
  OR U1324 ( .A(n661), .B(n660), .Z(n665) );
  NANDN U1325 ( .A(n663), .B(n662), .Z(n664) );
  AND U1326 ( .A(n665), .B(n664), .Z(n737) );
  NANDN U1327 ( .A(n667), .B(n666), .Z(n671) );
  NANDN U1328 ( .A(n669), .B(n668), .Z(n670) );
  AND U1329 ( .A(n671), .B(n670), .Z(n746) );
  NANDN U1330 ( .A(n673), .B(n672), .Z(n677) );
  NANDN U1331 ( .A(n675), .B(n674), .Z(n676) );
  NAND U1332 ( .A(n677), .B(n676), .Z(n784) );
  NAND U1333 ( .A(n679), .B(n678), .Z(n683) );
  NAND U1334 ( .A(n681), .B(n680), .Z(n682) );
  NAND U1335 ( .A(n683), .B(n682), .Z(n782) );
  AND U1336 ( .A(x[131]), .B(y[651]), .Z(n685) );
  AND U1337 ( .A(y[646]), .B(x[136]), .Z(n684) );
  XNOR U1338 ( .A(n685), .B(n684), .Z(n796) );
  XNOR U1339 ( .A(n795), .B(n796), .Z(n805) );
  IV U1340 ( .A(y[650]), .Z(n2627) );
  ANDN U1341 ( .B(x[132]), .A(n2627), .Z(n803) );
  AND U1342 ( .A(x[138]), .B(y[644]), .Z(n1430) );
  AND U1343 ( .A(x[137]), .B(y[645]), .Z(n1389) );
  NAND U1344 ( .A(y[652]), .B(x[130]), .Z(n686) );
  XOR U1345 ( .A(n1389), .B(n686), .Z(n750) );
  XNOR U1346 ( .A(n1430), .B(n750), .Z(n804) );
  XNOR U1347 ( .A(n803), .B(n804), .Z(n806) );
  XNOR U1348 ( .A(n805), .B(n806), .Z(n811) );
  AND U1349 ( .A(x[135]), .B(y[652]), .Z(n688) );
  NAND U1350 ( .A(n688), .B(n687), .Z(n692) );
  NANDN U1351 ( .A(n690), .B(n689), .Z(n691) );
  AND U1352 ( .A(n692), .B(n691), .Z(n809) );
  NAND U1353 ( .A(x[138]), .B(y[642]), .Z(n1318) );
  NOR U1354 ( .A(n141), .B(n162), .Z(n894) );
  NANDN U1355 ( .A(n1318), .B(n894), .Z(n695) );
  NAND U1356 ( .A(n693), .B(n1313), .Z(n694) );
  AND U1357 ( .A(n695), .B(n694), .Z(n810) );
  XOR U1358 ( .A(n809), .B(n810), .Z(n812) );
  XNOR U1359 ( .A(n811), .B(n812), .Z(n783) );
  XOR U1360 ( .A(n784), .B(n785), .Z(n743) );
  ANDN U1361 ( .B(x[133]), .A(n2627), .Z(n867) );
  NAND U1362 ( .A(n1557), .B(n867), .Z(n699) );
  OR U1363 ( .A(n697), .B(n696), .Z(n698) );
  NAND U1364 ( .A(n699), .B(n698), .Z(n778) );
  IV U1365 ( .A(n894), .Z(n765) );
  XNOR U1366 ( .A(n765), .B(n764), .Z(n766) );
  XOR U1367 ( .A(n767), .B(n766), .Z(n777) );
  ANDN U1368 ( .B(y[653]), .A(n164), .Z(n2293) );
  NAND U1369 ( .A(n877), .B(n2293), .Z(n703) );
  OR U1370 ( .A(n701), .B(n700), .Z(n702) );
  AND U1371 ( .A(n703), .B(n702), .Z(n776) );
  XNOR U1372 ( .A(n777), .B(n776), .Z(n779) );
  XOR U1373 ( .A(n778), .B(n779), .Z(n817) );
  AND U1374 ( .A(x[137]), .B(y[647]), .Z(n900) );
  NAND U1375 ( .A(n900), .B(n704), .Z(n708) );
  OR U1376 ( .A(n706), .B(n705), .Z(n707) );
  AND U1377 ( .A(n708), .B(n707), .Z(n773) );
  NAND U1378 ( .A(x[141]), .B(y[641]), .Z(n761) );
  XOR U1379 ( .A(o[14]), .B(n761), .Z(n756) );
  AND U1380 ( .A(y[642]), .B(x[140]), .Z(n1383) );
  NAND U1381 ( .A(y[647]), .B(x[135]), .Z(n709) );
  XNOR U1382 ( .A(n1383), .B(n709), .Z(n755) );
  NANDN U1383 ( .A(n710), .B(o[13]), .Z(n800) );
  AND U1384 ( .A(y[654]), .B(x[128]), .Z(n712) );
  NAND U1385 ( .A(x[142]), .B(y[640]), .Z(n711) );
  XNOR U1386 ( .A(n712), .B(n711), .Z(n799) );
  XOR U1387 ( .A(n773), .B(n772), .Z(n815) );
  NAND U1388 ( .A(n714), .B(n713), .Z(n718) );
  NAND U1389 ( .A(n716), .B(n715), .Z(n717) );
  NAND U1390 ( .A(n718), .B(n717), .Z(n816) );
  XOR U1391 ( .A(n815), .B(n816), .Z(n818) );
  XNOR U1392 ( .A(n817), .B(n818), .Z(n744) );
  XOR U1393 ( .A(n746), .B(n745), .Z(n738) );
  XNOR U1394 ( .A(n737), .B(n738), .Z(n739) );
  XNOR U1395 ( .A(n740), .B(n739), .Z(n734) );
  NANDN U1396 ( .A(n720), .B(n719), .Z(n724) );
  NANDN U1397 ( .A(n722), .B(n721), .Z(n723) );
  NAND U1398 ( .A(n724), .B(n723), .Z(n731) );
  OR U1399 ( .A(n726), .B(n725), .Z(n730) );
  NANDN U1400 ( .A(n728), .B(n727), .Z(n729) );
  AND U1401 ( .A(n730), .B(n729), .Z(n732) );
  XNOR U1402 ( .A(n731), .B(n732), .Z(n733) );
  XOR U1403 ( .A(n734), .B(n733), .Z(N47) );
  NANDN U1404 ( .A(n732), .B(n731), .Z(n736) );
  NANDN U1405 ( .A(n734), .B(n733), .Z(n735) );
  NAND U1406 ( .A(n736), .B(n735), .Z(n821) );
  OR U1407 ( .A(n738), .B(n737), .Z(n742) );
  OR U1408 ( .A(n740), .B(n739), .Z(n741) );
  AND U1409 ( .A(n742), .B(n741), .Z(n822) );
  XNOR U1410 ( .A(n821), .B(n822), .Z(n823) );
  NAND U1411 ( .A(n744), .B(n743), .Z(n748) );
  NANDN U1412 ( .A(n746), .B(n745), .Z(n747) );
  NAND U1413 ( .A(n748), .B(n747), .Z(n830) );
  IV U1414 ( .A(y[652]), .Z(n2617) );
  ANDN U1415 ( .B(x[137]), .A(n2617), .Z(n1531) );
  NAND U1416 ( .A(n749), .B(n1531), .Z(n752) );
  NANDN U1417 ( .A(n750), .B(n1430), .Z(n751) );
  AND U1418 ( .A(n752), .B(n751), .Z(n839) );
  AND U1419 ( .A(x[140]), .B(y[647]), .Z(n753) );
  NAND U1420 ( .A(n754), .B(n753), .Z(n758) );
  NANDN U1421 ( .A(n756), .B(n755), .Z(n757) );
  NAND U1422 ( .A(n758), .B(n757), .Z(n891) );
  AND U1423 ( .A(y[643]), .B(x[140]), .Z(n760) );
  NAND U1424 ( .A(y[644]), .B(x[139]), .Z(n759) );
  XOR U1425 ( .A(n760), .B(n759), .Z(n896) );
  NAND U1426 ( .A(x[141]), .B(y[642]), .Z(n895) );
  XOR U1427 ( .A(n896), .B(n895), .Z(n888) );
  NANDN U1428 ( .A(n761), .B(o[14]), .Z(n879) );
  AND U1429 ( .A(x[128]), .B(y[655]), .Z(n763) );
  NAND U1430 ( .A(y[640]), .B(x[143]), .Z(n762) );
  XOR U1431 ( .A(n763), .B(n762), .Z(n878) );
  XOR U1432 ( .A(n879), .B(n878), .Z(n889) );
  XNOR U1433 ( .A(n888), .B(n889), .Z(n890) );
  XOR U1434 ( .A(n891), .B(n890), .Z(n840) );
  XOR U1435 ( .A(n839), .B(n840), .Z(n841) );
  NAND U1436 ( .A(n765), .B(n764), .Z(n769) );
  OR U1437 ( .A(n767), .B(n766), .Z(n768) );
  NAND U1438 ( .A(n769), .B(n768), .Z(n842) );
  NAND U1439 ( .A(n771), .B(n770), .Z(n775) );
  NANDN U1440 ( .A(n773), .B(n772), .Z(n774) );
  AND U1441 ( .A(n775), .B(n774), .Z(n833) );
  XNOR U1442 ( .A(n834), .B(n833), .Z(n836) );
  OR U1443 ( .A(n777), .B(n776), .Z(n781) );
  NANDN U1444 ( .A(n779), .B(n778), .Z(n780) );
  AND U1445 ( .A(n781), .B(n780), .Z(n835) );
  XOR U1446 ( .A(n836), .B(n835), .Z(n911) );
  NANDN U1447 ( .A(n783), .B(n782), .Z(n787) );
  NANDN U1448 ( .A(n785), .B(n784), .Z(n786) );
  NAND U1449 ( .A(n787), .B(n786), .Z(n910) );
  NAND U1450 ( .A(y[641]), .B(x[142]), .Z(n864) );
  XOR U1451 ( .A(o[15]), .B(n864), .Z(n874) );
  AND U1452 ( .A(y[654]), .B(x[129]), .Z(n789) );
  NAND U1453 ( .A(y[647]), .B(x[136]), .Z(n788) );
  XNOR U1454 ( .A(n789), .B(n788), .Z(n873) );
  XNOR U1455 ( .A(n874), .B(n873), .Z(n903) );
  NAND U1456 ( .A(y[652]), .B(x[131]), .Z(n861) );
  AND U1457 ( .A(y[646]), .B(x[137]), .Z(n791) );
  NAND U1458 ( .A(x[130]), .B(y[653]), .Z(n790) );
  XOR U1459 ( .A(n791), .B(n790), .Z(n860) );
  XOR U1460 ( .A(n861), .B(n860), .Z(n904) );
  XNOR U1461 ( .A(n903), .B(n904), .Z(n906) );
  NAND U1462 ( .A(x[135]), .B(y[648]), .Z(n1265) );
  AND U1463 ( .A(x[138]), .B(y[645]), .Z(n793) );
  NAND U1464 ( .A(x[132]), .B(y[651]), .Z(n792) );
  XOR U1465 ( .A(n793), .B(n792), .Z(n885) );
  XNOR U1466 ( .A(n1265), .B(n885), .Z(n868) );
  AND U1467 ( .A(y[649]), .B(x[134]), .Z(n951) );
  XNOR U1468 ( .A(n867), .B(n951), .Z(n869) );
  XNOR U1469 ( .A(n868), .B(n869), .Z(n905) );
  XOR U1470 ( .A(n906), .B(n905), .Z(n854) );
  NAND U1471 ( .A(x[136]), .B(y[651]), .Z(n1182) );
  OR U1472 ( .A(n1182), .B(n794), .Z(n798) );
  NANDN U1473 ( .A(n796), .B(n795), .Z(n797) );
  NAND U1474 ( .A(n798), .B(n797), .Z(n852) );
  ANDN U1475 ( .B(y[654]), .A(n165), .Z(n2599) );
  NAND U1476 ( .A(n877), .B(n2599), .Z(n802) );
  NANDN U1477 ( .A(n800), .B(n799), .Z(n801) );
  NAND U1478 ( .A(n802), .B(n801), .Z(n851) );
  XNOR U1479 ( .A(n852), .B(n851), .Z(n853) );
  XNOR U1480 ( .A(n854), .B(n853), .Z(n846) );
  OR U1481 ( .A(n804), .B(n803), .Z(n808) );
  OR U1482 ( .A(n806), .B(n805), .Z(n807) );
  AND U1483 ( .A(n808), .B(n807), .Z(n845) );
  XNOR U1484 ( .A(n846), .B(n845), .Z(n847) );
  OR U1485 ( .A(n810), .B(n809), .Z(n814) );
  NAND U1486 ( .A(n812), .B(n811), .Z(n813) );
  NAND U1487 ( .A(n814), .B(n813), .Z(n848) );
  XOR U1488 ( .A(n847), .B(n848), .Z(n909) );
  XOR U1489 ( .A(n910), .B(n909), .Z(n912) );
  XOR U1490 ( .A(n911), .B(n912), .Z(n827) );
  NANDN U1491 ( .A(n816), .B(n815), .Z(n820) );
  NANDN U1492 ( .A(n818), .B(n817), .Z(n819) );
  NAND U1493 ( .A(n820), .B(n819), .Z(n828) );
  XOR U1494 ( .A(n827), .B(n828), .Z(n829) );
  XNOR U1495 ( .A(n830), .B(n829), .Z(n824) );
  XOR U1496 ( .A(n823), .B(n824), .Z(N48) );
  NANDN U1497 ( .A(n822), .B(n821), .Z(n826) );
  NANDN U1498 ( .A(n824), .B(n823), .Z(n825) );
  NAND U1499 ( .A(n826), .B(n825), .Z(n915) );
  OR U1500 ( .A(n828), .B(n827), .Z(n832) );
  NANDN U1501 ( .A(n830), .B(n829), .Z(n831) );
  NAND U1502 ( .A(n832), .B(n831), .Z(n916) );
  XNOR U1503 ( .A(n915), .B(n916), .Z(n917) );
  OR U1504 ( .A(n834), .B(n833), .Z(n838) );
  OR U1505 ( .A(n836), .B(n835), .Z(n837) );
  NAND U1506 ( .A(n838), .B(n837), .Z(n1005) );
  OR U1507 ( .A(n840), .B(n839), .Z(n844) );
  NANDN U1508 ( .A(n842), .B(n841), .Z(n843) );
  NAND U1509 ( .A(n844), .B(n843), .Z(n1003) );
  OR U1510 ( .A(n846), .B(n845), .Z(n850) );
  OR U1511 ( .A(n848), .B(n847), .Z(n849) );
  AND U1512 ( .A(n850), .B(n849), .Z(n1002) );
  XOR U1513 ( .A(n1003), .B(n1002), .Z(n1004) );
  XNOR U1514 ( .A(n1005), .B(n1004), .Z(n924) );
  OR U1515 ( .A(n852), .B(n851), .Z(n856) );
  OR U1516 ( .A(n854), .B(n853), .Z(n855) );
  AND U1517 ( .A(n856), .B(n855), .Z(n996) );
  AND U1518 ( .A(y[645]), .B(x[139]), .Z(n858) );
  NAND U1519 ( .A(x[142]), .B(y[642]), .Z(n857) );
  XOR U1520 ( .A(n858), .B(n857), .Z(n977) );
  NAND U1521 ( .A(x[132]), .B(y[652]), .Z(n976) );
  XOR U1522 ( .A(n977), .B(n976), .Z(n927) );
  AND U1523 ( .A(y[653]), .B(x[137]), .Z(n1629) );
  NAND U1524 ( .A(n859), .B(n1629), .Z(n863) );
  OR U1525 ( .A(n861), .B(n860), .Z(n862) );
  NAND U1526 ( .A(n863), .B(n862), .Z(n928) );
  XNOR U1527 ( .A(n927), .B(n928), .Z(n930) );
  NANDN U1528 ( .A(n864), .B(o[15]), .Z(n948) );
  NAND U1529 ( .A(x[129]), .B(y[655]), .Z(n865) );
  XNOR U1530 ( .A(n866), .B(n865), .Z(n947) );
  XNOR U1531 ( .A(n948), .B(n947), .Z(n929) );
  XNOR U1532 ( .A(n930), .B(n929), .Z(n966) );
  OR U1533 ( .A(n867), .B(n951), .Z(n871) );
  NANDN U1534 ( .A(n869), .B(n868), .Z(n870) );
  AND U1535 ( .A(n871), .B(n870), .Z(n963) );
  AND U1536 ( .A(x[136]), .B(y[654]), .Z(n1566) );
  NAND U1537 ( .A(n872), .B(n1566), .Z(n876) );
  NANDN U1538 ( .A(n874), .B(n873), .Z(n875) );
  NAND U1539 ( .A(n876), .B(n875), .Z(n969) );
  AND U1540 ( .A(x[143]), .B(y[655]), .Z(n3051) );
  NAND U1541 ( .A(n877), .B(n3051), .Z(n881) );
  OR U1542 ( .A(n879), .B(n878), .Z(n880) );
  AND U1543 ( .A(n881), .B(n880), .Z(n970) );
  NAND U1544 ( .A(x[128]), .B(y[656]), .Z(n942) );
  NAND U1545 ( .A(y[640]), .B(x[144]), .Z(n941) );
  XOR U1546 ( .A(n942), .B(n941), .Z(n943) );
  NAND U1547 ( .A(x[143]), .B(y[641]), .Z(n956) );
  XOR U1548 ( .A(o[16]), .B(n956), .Z(n944) );
  XOR U1549 ( .A(n943), .B(n944), .Z(n934) );
  NAND U1550 ( .A(y[646]), .B(x[138]), .Z(n953) );
  NAND U1551 ( .A(x[135]), .B(y[649]), .Z(n882) );
  XNOR U1552 ( .A(n883), .B(n882), .Z(n952) );
  XOR U1553 ( .A(n934), .B(n933), .Z(n935) );
  ANDN U1554 ( .B(y[651]), .A(n161), .Z(n1575) );
  NAND U1555 ( .A(n884), .B(n1575), .Z(n887) );
  OR U1556 ( .A(n1265), .B(n885), .Z(n886) );
  AND U1557 ( .A(n887), .B(n886), .Z(n936) );
  XOR U1558 ( .A(n935), .B(n936), .Z(n971) );
  XNOR U1559 ( .A(n963), .B(n964), .Z(n965) );
  XNOR U1560 ( .A(n966), .B(n965), .Z(n997) );
  XOR U1561 ( .A(n996), .B(n997), .Z(n999) );
  OR U1562 ( .A(n889), .B(n888), .Z(n893) );
  OR U1563 ( .A(n891), .B(n890), .Z(n892) );
  AND U1564 ( .A(n893), .B(n892), .Z(n992) );
  ANDN U1565 ( .B(x[140]), .A(n2634), .Z(n1633) );
  NAND U1566 ( .A(n894), .B(n1633), .Z(n898) );
  OR U1567 ( .A(n896), .B(n895), .Z(n897) );
  NAND U1568 ( .A(n898), .B(n897), .Z(n986) );
  NAND U1569 ( .A(x[130]), .B(y[654]), .Z(n899) );
  XOR U1570 ( .A(n900), .B(n899), .Z(n981) );
  NAND U1571 ( .A(y[653]), .B(x[131]), .Z(n980) );
  XOR U1572 ( .A(n981), .B(n980), .Z(n984) );
  AND U1573 ( .A(x[133]), .B(y[651]), .Z(n902) );
  NAND U1574 ( .A(y[643]), .B(x[141]), .Z(n901) );
  XNOR U1575 ( .A(n902), .B(n901), .Z(n960) );
  XNOR U1576 ( .A(n1633), .B(n960), .Z(n985) );
  XOR U1577 ( .A(n984), .B(n985), .Z(n987) );
  XNOR U1578 ( .A(n986), .B(n987), .Z(n990) );
  OR U1579 ( .A(n904), .B(n903), .Z(n908) );
  NANDN U1580 ( .A(n906), .B(n905), .Z(n907) );
  AND U1581 ( .A(n908), .B(n907), .Z(n991) );
  XNOR U1582 ( .A(n990), .B(n991), .Z(n993) );
  XOR U1583 ( .A(n992), .B(n993), .Z(n998) );
  XOR U1584 ( .A(n999), .B(n998), .Z(n921) );
  NANDN U1585 ( .A(n910), .B(n909), .Z(n914) );
  OR U1586 ( .A(n912), .B(n911), .Z(n913) );
  NAND U1587 ( .A(n914), .B(n913), .Z(n922) );
  XOR U1588 ( .A(n921), .B(n922), .Z(n923) );
  XNOR U1589 ( .A(n924), .B(n923), .Z(n918) );
  XOR U1590 ( .A(n917), .B(n918), .Z(N49) );
  NANDN U1591 ( .A(n916), .B(n915), .Z(n920) );
  NANDN U1592 ( .A(n918), .B(n917), .Z(n919) );
  NAND U1593 ( .A(n920), .B(n919), .Z(n1105) );
  OR U1594 ( .A(n922), .B(n921), .Z(n926) );
  NANDN U1595 ( .A(n924), .B(n923), .Z(n925) );
  NAND U1596 ( .A(n926), .B(n925), .Z(n1106) );
  XNOR U1597 ( .A(n1105), .B(n1106), .Z(n1107) );
  OR U1598 ( .A(n928), .B(n927), .Z(n932) );
  OR U1599 ( .A(n930), .B(n929), .Z(n931) );
  AND U1600 ( .A(n932), .B(n931), .Z(n1008) );
  NANDN U1601 ( .A(n934), .B(n933), .Z(n938) );
  OR U1602 ( .A(n936), .B(n935), .Z(n937) );
  NAND U1603 ( .A(n938), .B(n937), .Z(n1090) );
  NAND U1604 ( .A(y[654]), .B(x[131]), .Z(n1054) );
  AND U1605 ( .A(x[138]), .B(y[647]), .Z(n940) );
  AND U1606 ( .A(x[130]), .B(y[655]), .Z(n939) );
  XNOR U1607 ( .A(n940), .B(n939), .Z(n1053) );
  XOR U1608 ( .A(n1054), .B(n1053), .Z(n1076) );
  NAND U1609 ( .A(x[128]), .B(y[657]), .Z(n1028) );
  NAND U1610 ( .A(y[641]), .B(x[144]), .Z(n1022) );
  XOR U1611 ( .A(o[17]), .B(n1022), .Z(n1026) );
  AND U1612 ( .A(y[640]), .B(x[145]), .Z(n1025) );
  XNOR U1613 ( .A(n1026), .B(n1025), .Z(n1027) );
  XNOR U1614 ( .A(n1076), .B(n1075), .Z(n1078) );
  OR U1615 ( .A(n942), .B(n941), .Z(n946) );
  NANDN U1616 ( .A(n944), .B(n943), .Z(n945) );
  AND U1617 ( .A(n946), .B(n945), .Z(n1077) );
  XOR U1618 ( .A(n1078), .B(n1077), .Z(n1084) );
  IV U1619 ( .A(y[655]), .Z(n2237) );
  ANDN U1620 ( .B(x[136]), .A(n2237), .Z(n1853) );
  ANDN U1621 ( .B(y[648]), .A(n152), .Z(n1160) );
  NAND U1622 ( .A(n1853), .B(n1160), .Z(n950) );
  NANDN U1623 ( .A(n948), .B(n947), .Z(n949) );
  NAND U1624 ( .A(n950), .B(n949), .Z(n1082) );
  ANDN U1625 ( .B(y[650]), .A(n158), .Z(n1181) );
  NAND U1626 ( .A(n1181), .B(n951), .Z(n955) );
  NANDN U1627 ( .A(n953), .B(n952), .Z(n954) );
  NAND U1628 ( .A(n955), .B(n954), .Z(n1081) );
  XNOR U1629 ( .A(n1082), .B(n1081), .Z(n1083) );
  XOR U1630 ( .A(n1084), .B(n1083), .Z(n1087) );
  ANDN U1631 ( .B(x[140]), .A(n142), .Z(n1037) );
  ANDN U1632 ( .B(x[142]), .A(n141), .Z(n1035) );
  ANDN U1633 ( .B(x[143]), .A(n140), .Z(n1036) );
  XNOR U1634 ( .A(n1035), .B(n1036), .Z(n1038) );
  XOR U1635 ( .A(n1037), .B(n1038), .Z(n1071) );
  NANDN U1636 ( .A(n956), .B(o[16]), .Z(n1066) );
  AND U1637 ( .A(y[648]), .B(x[137]), .Z(n958) );
  AND U1638 ( .A(x[129]), .B(y[656]), .Z(n957) );
  XNOR U1639 ( .A(n958), .B(n957), .Z(n1065) );
  XOR U1640 ( .A(n1066), .B(n1065), .Z(n1069) );
  ANDN U1641 ( .B(y[651]), .A(n164), .Z(n1973) );
  NAND U1642 ( .A(n959), .B(n1973), .Z(n962) );
  NAND U1643 ( .A(n960), .B(n1633), .Z(n961) );
  AND U1644 ( .A(n962), .B(n961), .Z(n1070) );
  XNOR U1645 ( .A(n1071), .B(n1072), .Z(n1088) );
  XOR U1646 ( .A(n1087), .B(n1088), .Z(n1089) );
  XOR U1647 ( .A(n1090), .B(n1089), .Z(n1009) );
  XOR U1648 ( .A(n1008), .B(n1009), .Z(n1010) );
  OR U1649 ( .A(n964), .B(n963), .Z(n968) );
  OR U1650 ( .A(n966), .B(n965), .Z(n967) );
  AND U1651 ( .A(n968), .B(n967), .Z(n1011) );
  NANDN U1652 ( .A(n970), .B(n969), .Z(n974) );
  NAND U1653 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1654 ( .A(n974), .B(n973), .Z(n1096) );
  IV U1655 ( .A(y[649]), .Z(n2457) );
  ANDN U1656 ( .B(x[136]), .A(n2457), .Z(n1060) );
  XNOR U1657 ( .A(n1059), .B(n1060), .Z(n1062) );
  ANDN U1658 ( .B(x[133]), .A(n2617), .Z(n1061) );
  XOR U1659 ( .A(n1062), .B(n1061), .Z(n1048) );
  ANDN U1660 ( .B(y[653]), .A(n155), .Z(n1016) );
  ANDN U1661 ( .B(x[139]), .A(n2618), .Z(n1014) );
  ANDN U1662 ( .B(x[141]), .A(n2634), .Z(n1015) );
  XNOR U1663 ( .A(n1014), .B(n1015), .Z(n1017) );
  XNOR U1664 ( .A(n1016), .B(n1017), .Z(n1047) );
  XOR U1665 ( .A(n1048), .B(n1047), .Z(n1049) );
  XNOR U1666 ( .A(n1181), .B(n1049), .Z(n1044) );
  NAND U1667 ( .A(y[642]), .B(x[139]), .Z(n1143) );
  AND U1668 ( .A(y[645]), .B(x[142]), .Z(n975) );
  NANDN U1669 ( .A(n1143), .B(n975), .Z(n979) );
  OR U1670 ( .A(n977), .B(n976), .Z(n978) );
  NAND U1671 ( .A(n979), .B(n978), .Z(n1042) );
  AND U1672 ( .A(x[137]), .B(y[654]), .Z(n1694) );
  NAND U1673 ( .A(n1694), .B(n1052), .Z(n983) );
  OR U1674 ( .A(n981), .B(n980), .Z(n982) );
  NAND U1675 ( .A(n983), .B(n982), .Z(n1041) );
  XNOR U1676 ( .A(n1042), .B(n1041), .Z(n1043) );
  XOR U1677 ( .A(n1044), .B(n1043), .Z(n1094) );
  NANDN U1678 ( .A(n985), .B(n984), .Z(n989) );
  NANDN U1679 ( .A(n987), .B(n986), .Z(n988) );
  AND U1680 ( .A(n989), .B(n988), .Z(n1093) );
  XOR U1681 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1682 ( .A(n1096), .B(n1095), .Z(n1100) );
  OR U1683 ( .A(n991), .B(n990), .Z(n995) );
  OR U1684 ( .A(n993), .B(n992), .Z(n994) );
  NAND U1685 ( .A(n995), .B(n994), .Z(n1099) );
  XOR U1686 ( .A(n1100), .B(n1099), .Z(n1101) );
  OR U1687 ( .A(n997), .B(n996), .Z(n1001) );
  NAND U1688 ( .A(n999), .B(n998), .Z(n1000) );
  NAND U1689 ( .A(n1001), .B(n1000), .Z(n1102) );
  XNOR U1690 ( .A(n1101), .B(n1102), .Z(n1111) );
  XNOR U1691 ( .A(n1112), .B(n1111), .Z(n1114) );
  OR U1692 ( .A(n1003), .B(n1002), .Z(n1007) );
  NANDN U1693 ( .A(n1005), .B(n1004), .Z(n1006) );
  AND U1694 ( .A(n1007), .B(n1006), .Z(n1113) );
  XOR U1695 ( .A(n1114), .B(n1113), .Z(n1108) );
  XNOR U1696 ( .A(n1107), .B(n1108), .Z(N50) );
  OR U1697 ( .A(n1009), .B(n1008), .Z(n1013) );
  NANDN U1698 ( .A(n1011), .B(n1010), .Z(n1012) );
  AND U1699 ( .A(n1013), .B(n1012), .Z(n1123) );
  OR U1700 ( .A(n1015), .B(n1014), .Z(n1019) );
  OR U1701 ( .A(n1017), .B(n1016), .Z(n1018) );
  NAND U1702 ( .A(n1019), .B(n1018), .Z(n1151) );
  NAND U1703 ( .A(y[644]), .B(x[142]), .Z(n1020) );
  XOR U1704 ( .A(n1021), .B(n1020), .Z(n1138) );
  NAND U1705 ( .A(x[143]), .B(y[643]), .Z(n1137) );
  XOR U1706 ( .A(n1138), .B(n1137), .Z(n1148) );
  NANDN U1707 ( .A(n1022), .B(o[17]), .Z(n1162) );
  AND U1708 ( .A(x[138]), .B(y[648]), .Z(n1024) );
  NAND U1709 ( .A(x[129]), .B(y[657]), .Z(n1023) );
  XNOR U1710 ( .A(n1024), .B(n1023), .Z(n1161) );
  XOR U1711 ( .A(n1148), .B(n1149), .Z(n1150) );
  XNOR U1712 ( .A(n1151), .B(n1150), .Z(n1215) );
  NANDN U1713 ( .A(n1026), .B(n1025), .Z(n1030) );
  NANDN U1714 ( .A(n1028), .B(n1027), .Z(n1029) );
  NAND U1715 ( .A(n1030), .B(n1029), .Z(n1203) );
  NAND U1716 ( .A(x[135]), .B(y[651]), .Z(n1031) );
  XOR U1717 ( .A(n1032), .B(n1031), .Z(n1184) );
  NAND U1718 ( .A(x[132]), .B(y[654]), .Z(n1183) );
  XNOR U1719 ( .A(n1184), .B(n1183), .Z(n1130) );
  AND U1720 ( .A(x[133]), .B(y[653]), .Z(n1297) );
  NAND U1721 ( .A(x[134]), .B(y[652]), .Z(n1129) );
  XNOR U1722 ( .A(n1297), .B(n1129), .Z(n1131) );
  XOR U1723 ( .A(n1203), .B(n1202), .Z(n1205) );
  NAND U1724 ( .A(x[130]), .B(y[656]), .Z(n1145) );
  AND U1725 ( .A(y[647]), .B(x[139]), .Z(n1034) );
  AND U1726 ( .A(x[144]), .B(y[642]), .Z(n1033) );
  XNOR U1727 ( .A(n1034), .B(n1033), .Z(n1144) );
  XOR U1728 ( .A(n1145), .B(n1144), .Z(n1204) );
  XNOR U1729 ( .A(n1205), .B(n1204), .Z(n1214) );
  XOR U1730 ( .A(n1215), .B(n1214), .Z(n1217) );
  OR U1731 ( .A(n1036), .B(n1035), .Z(n1040) );
  OR U1732 ( .A(n1038), .B(n1037), .Z(n1039) );
  NAND U1733 ( .A(n1040), .B(n1039), .Z(n1216) );
  XOR U1734 ( .A(n1217), .B(n1216), .Z(n1220) );
  OR U1735 ( .A(n1042), .B(n1041), .Z(n1046) );
  OR U1736 ( .A(n1044), .B(n1043), .Z(n1045) );
  AND U1737 ( .A(n1046), .B(n1045), .Z(n1192) );
  NANDN U1738 ( .A(n1048), .B(n1047), .Z(n1051) );
  NANDN U1739 ( .A(n1049), .B(n1181), .Z(n1050) );
  NAND U1740 ( .A(n1051), .B(n1050), .Z(n1191) );
  NAND U1741 ( .A(y[655]), .B(x[138]), .Z(n2027) );
  NANDN U1742 ( .A(n2027), .B(n1052), .Z(n1056) );
  OR U1743 ( .A(n1054), .B(n1053), .Z(n1055) );
  AND U1744 ( .A(n1056), .B(n1055), .Z(n1156) );
  NAND U1745 ( .A(x[128]), .B(y[658]), .Z(n1166) );
  NAND U1746 ( .A(x[146]), .B(y[640]), .Z(n1165) );
  XOR U1747 ( .A(n1166), .B(n1165), .Z(n1167) );
  NAND U1748 ( .A(x[145]), .B(y[641]), .Z(n1187) );
  XOR U1749 ( .A(o[18]), .B(n1187), .Z(n1168) );
  XOR U1750 ( .A(n1167), .B(n1168), .Z(n1155) );
  ANDN U1751 ( .B(x[140]), .A(n2618), .Z(n1255) );
  AND U1752 ( .A(y[655]), .B(x[131]), .Z(n1058) );
  NAND U1753 ( .A(x[141]), .B(y[645]), .Z(n1057) );
  XOR U1754 ( .A(n1058), .B(n1057), .Z(n1174) );
  XOR U1755 ( .A(n1255), .B(n1174), .Z(n1154) );
  XNOR U1756 ( .A(n1155), .B(n1154), .Z(n1157) );
  XOR U1757 ( .A(n1156), .B(n1157), .Z(n1208) );
  OR U1758 ( .A(n1060), .B(n1059), .Z(n1064) );
  OR U1759 ( .A(n1062), .B(n1061), .Z(n1063) );
  AND U1760 ( .A(n1064), .B(n1063), .Z(n1209) );
  XNOR U1761 ( .A(n1208), .B(n1209), .Z(n1211) );
  ANDN U1762 ( .B(y[656]), .A(n160), .Z(n2028) );
  NAND U1763 ( .A(n1160), .B(n2028), .Z(n1068) );
  OR U1764 ( .A(n1066), .B(n1065), .Z(n1067) );
  NAND U1765 ( .A(n1068), .B(n1067), .Z(n1210) );
  XNOR U1766 ( .A(n1211), .B(n1210), .Z(n1190) );
  XNOR U1767 ( .A(n1191), .B(n1190), .Z(n1193) );
  XOR U1768 ( .A(n1192), .B(n1193), .Z(n1221) );
  XOR U1769 ( .A(n1220), .B(n1221), .Z(n1223) );
  NANDN U1770 ( .A(n1070), .B(n1069), .Z(n1074) );
  OR U1771 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U1772 ( .A(n1074), .B(n1073), .Z(n1196) );
  NAND U1773 ( .A(n1076), .B(n1075), .Z(n1080) );
  OR U1774 ( .A(n1078), .B(n1077), .Z(n1079) );
  AND U1775 ( .A(n1080), .B(n1079), .Z(n1197) );
  XOR U1776 ( .A(n1196), .B(n1197), .Z(n1198) );
  OR U1777 ( .A(n1082), .B(n1081), .Z(n1086) );
  OR U1778 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U1779 ( .A(n1086), .B(n1085), .Z(n1199) );
  XOR U1780 ( .A(n1223), .B(n1222), .Z(n1229) );
  OR U1781 ( .A(n1088), .B(n1087), .Z(n1092) );
  NAND U1782 ( .A(n1090), .B(n1089), .Z(n1091) );
  NAND U1783 ( .A(n1092), .B(n1091), .Z(n1227) );
  OR U1784 ( .A(n1094), .B(n1093), .Z(n1098) );
  NAND U1785 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1786 ( .A(n1098), .B(n1097), .Z(n1226) );
  XOR U1787 ( .A(n1229), .B(n1228), .Z(n1124) );
  XNOR U1788 ( .A(n1123), .B(n1124), .Z(n1126) );
  OR U1789 ( .A(n1100), .B(n1099), .Z(n1104) );
  NANDN U1790 ( .A(n1102), .B(n1101), .Z(n1103) );
  NAND U1791 ( .A(n1104), .B(n1103), .Z(n1125) );
  XOR U1792 ( .A(n1126), .B(n1125), .Z(n1119) );
  NANDN U1793 ( .A(n1106), .B(n1105), .Z(n1110) );
  NAND U1794 ( .A(n1108), .B(n1107), .Z(n1109) );
  NAND U1795 ( .A(n1110), .B(n1109), .Z(n1117) );
  OR U1796 ( .A(n1112), .B(n1111), .Z(n1116) );
  OR U1797 ( .A(n1114), .B(n1113), .Z(n1115) );
  AND U1798 ( .A(n1116), .B(n1115), .Z(n1118) );
  XNOR U1799 ( .A(n1117), .B(n1118), .Z(n1120) );
  XNOR U1800 ( .A(n1119), .B(n1120), .Z(N51) );
  NANDN U1801 ( .A(n1118), .B(n1117), .Z(n1122) );
  NAND U1802 ( .A(n1120), .B(n1119), .Z(n1121) );
  NAND U1803 ( .A(n1122), .B(n1121), .Z(n1341) );
  OR U1804 ( .A(n1124), .B(n1123), .Z(n1128) );
  OR U1805 ( .A(n1126), .B(n1125), .Z(n1127) );
  AND U1806 ( .A(n1128), .B(n1127), .Z(n1342) );
  XNOR U1807 ( .A(n1341), .B(n1342), .Z(n1343) );
  NANDN U1808 ( .A(n1297), .B(n1129), .Z(n1133) );
  NAND U1809 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U1810 ( .A(n1133), .B(n1132), .Z(n1337) );
  AND U1811 ( .A(x[136]), .B(y[651]), .Z(n1135) );
  NAND U1812 ( .A(x[142]), .B(y[645]), .Z(n1134) );
  XOR U1813 ( .A(n1135), .B(n1134), .Z(n1315) );
  NAND U1814 ( .A(y[658]), .B(x[129]), .Z(n1314) );
  XOR U1815 ( .A(n1315), .B(n1314), .Z(n1281) );
  ANDN U1816 ( .B(x[142]), .A(n2457), .Z(n1815) );
  NAND U1817 ( .A(n1815), .B(n1136), .Z(n1140) );
  OR U1818 ( .A(n1138), .B(n1137), .Z(n1139) );
  NAND U1819 ( .A(n1140), .B(n1139), .Z(n1279) );
  AND U1820 ( .A(y[646]), .B(x[141]), .Z(n1142) );
  NAND U1821 ( .A(y[647]), .B(x[140]), .Z(n1141) );
  XOR U1822 ( .A(n1142), .B(n1141), .Z(n1258) );
  NAND U1823 ( .A(x[130]), .B(y[657]), .Z(n1257) );
  XNOR U1824 ( .A(n1258), .B(n1257), .Z(n1280) );
  XOR U1825 ( .A(n1279), .B(n1280), .Z(n1282) );
  XNOR U1826 ( .A(n1281), .B(n1282), .Z(n1335) );
  AND U1827 ( .A(y[647]), .B(x[144]), .Z(n1627) );
  NANDN U1828 ( .A(n1143), .B(n1627), .Z(n1147) );
  OR U1829 ( .A(n1145), .B(n1144), .Z(n1146) );
  NAND U1830 ( .A(n1147), .B(n1146), .Z(n1336) );
  XNOR U1831 ( .A(n1335), .B(n1336), .Z(n1338) );
  XOR U1832 ( .A(n1337), .B(n1338), .Z(n1244) );
  NANDN U1833 ( .A(n1149), .B(n1148), .Z(n1153) );
  OR U1834 ( .A(n1151), .B(n1150), .Z(n1152) );
  NAND U1835 ( .A(n1153), .B(n1152), .Z(n1330) );
  OR U1836 ( .A(n1155), .B(n1154), .Z(n1159) );
  OR U1837 ( .A(n1157), .B(n1156), .Z(n1158) );
  NAND U1838 ( .A(n1159), .B(n1158), .Z(n1329) );
  XOR U1839 ( .A(n1330), .B(n1329), .Z(n1331) );
  ANDN U1840 ( .B(y[657]), .A(n161), .Z(n2446) );
  NAND U1841 ( .A(n1160), .B(n2446), .Z(n1164) );
  NANDN U1842 ( .A(n1162), .B(n1161), .Z(n1163) );
  NAND U1843 ( .A(n1164), .B(n1163), .Z(n1293) );
  OR U1844 ( .A(n1166), .B(n1165), .Z(n1170) );
  NANDN U1845 ( .A(n1168), .B(n1167), .Z(n1169) );
  NAND U1846 ( .A(n1170), .B(n1169), .Z(n1292) );
  AND U1847 ( .A(y[650]), .B(x[137]), .Z(n1172) );
  NAND U1848 ( .A(x[144]), .B(y[643]), .Z(n1171) );
  XOR U1849 ( .A(n1172), .B(n1171), .Z(n1252) );
  NAND U1850 ( .A(x[143]), .B(y[644]), .Z(n1251) );
  XOR U1851 ( .A(n1252), .B(n1251), .Z(n1291) );
  XNOR U1852 ( .A(n1292), .B(n1291), .Z(n1294) );
  XNOR U1853 ( .A(n1293), .B(n1294), .Z(n1325) );
  ANDN U1854 ( .B(y[655]), .A(n164), .Z(n2580) );
  NAND U1855 ( .A(n1173), .B(n2580), .Z(n1176) );
  NANDN U1856 ( .A(n1174), .B(n1255), .Z(n1175) );
  NAND U1857 ( .A(n1176), .B(n1175), .Z(n1288) );
  AND U1858 ( .A(y[648]), .B(x[139]), .Z(n1178) );
  NAND U1859 ( .A(y[652]), .B(x[135]), .Z(n1177) );
  XOR U1860 ( .A(n1178), .B(n1177), .Z(n1267) );
  NAND U1861 ( .A(y[656]), .B(x[131]), .Z(n1266) );
  XOR U1862 ( .A(n1267), .B(n1266), .Z(n1286) );
  NAND U1863 ( .A(x[146]), .B(y[641]), .Z(n1272) );
  XOR U1864 ( .A(o[19]), .B(n1272), .Z(n1320) );
  AND U1865 ( .A(y[649]), .B(x[138]), .Z(n1180) );
  NAND U1866 ( .A(x[145]), .B(y[642]), .Z(n1179) );
  XNOR U1867 ( .A(n1180), .B(n1179), .Z(n1319) );
  XOR U1868 ( .A(n1288), .B(n1287), .Z(n1323) );
  NANDN U1869 ( .A(n1182), .B(n1181), .Z(n1186) );
  OR U1870 ( .A(n1184), .B(n1183), .Z(n1185) );
  NAND U1871 ( .A(n1186), .B(n1185), .Z(n1273) );
  NANDN U1872 ( .A(n1187), .B(o[18]), .Z(n1304) );
  NAND U1873 ( .A(x[128]), .B(y[659]), .Z(n1302) );
  NAND U1874 ( .A(x[147]), .B(y[640]), .Z(n1301) );
  XOR U1875 ( .A(n1302), .B(n1301), .Z(n1303) );
  XOR U1876 ( .A(n1304), .B(n1303), .Z(n1274) );
  XOR U1877 ( .A(n1273), .B(n1274), .Z(n1276) );
  NAND U1878 ( .A(x[132]), .B(y[655]), .Z(n1418) );
  AND U1879 ( .A(x[134]), .B(y[653]), .Z(n1189) );
  NAND U1880 ( .A(y[654]), .B(x[133]), .Z(n1188) );
  XNOR U1881 ( .A(n1189), .B(n1188), .Z(n1298) );
  XNOR U1882 ( .A(n1276), .B(n1275), .Z(n1324) );
  XNOR U1883 ( .A(n1323), .B(n1324), .Z(n1326) );
  XNOR U1884 ( .A(n1325), .B(n1326), .Z(n1332) );
  XNOR U1885 ( .A(n1331), .B(n1332), .Z(n1245) );
  XNOR U1886 ( .A(n1244), .B(n1245), .Z(n1247) );
  OR U1887 ( .A(n1191), .B(n1190), .Z(n1195) );
  OR U1888 ( .A(n1193), .B(n1192), .Z(n1194) );
  NAND U1889 ( .A(n1195), .B(n1194), .Z(n1246) );
  XOR U1890 ( .A(n1247), .B(n1246), .Z(n1241) );
  OR U1891 ( .A(n1197), .B(n1196), .Z(n1201) );
  NANDN U1892 ( .A(n1199), .B(n1198), .Z(n1200) );
  NAND U1893 ( .A(n1201), .B(n1200), .Z(n1239) );
  NANDN U1894 ( .A(n1203), .B(n1202), .Z(n1207) );
  OR U1895 ( .A(n1205), .B(n1204), .Z(n1206) );
  AND U1896 ( .A(n1207), .B(n1206), .Z(n1235) );
  OR U1897 ( .A(n1209), .B(n1208), .Z(n1213) );
  OR U1898 ( .A(n1211), .B(n1210), .Z(n1212) );
  AND U1899 ( .A(n1213), .B(n1212), .Z(n1232) );
  NANDN U1900 ( .A(n1215), .B(n1214), .Z(n1219) );
  OR U1901 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U1902 ( .A(n1219), .B(n1218), .Z(n1233) );
  XOR U1903 ( .A(n1232), .B(n1233), .Z(n1234) );
  XOR U1904 ( .A(n1239), .B(n1238), .Z(n1240) );
  XNOR U1905 ( .A(n1241), .B(n1240), .Z(n1350) );
  NANDN U1906 ( .A(n1221), .B(n1220), .Z(n1225) );
  OR U1907 ( .A(n1223), .B(n1222), .Z(n1224) );
  NAND U1908 ( .A(n1225), .B(n1224), .Z(n1347) );
  NANDN U1909 ( .A(n1227), .B(n1226), .Z(n1231) );
  NANDN U1910 ( .A(n1229), .B(n1228), .Z(n1230) );
  NAND U1911 ( .A(n1231), .B(n1230), .Z(n1348) );
  XNOR U1912 ( .A(n1350), .B(n1349), .Z(n1344) );
  XOR U1913 ( .A(n1343), .B(n1344), .Z(N52) );
  OR U1914 ( .A(n1233), .B(n1232), .Z(n1237) );
  NANDN U1915 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U1916 ( .A(n1237), .B(n1236), .Z(n1361) );
  OR U1917 ( .A(n1239), .B(n1238), .Z(n1243) );
  NANDN U1918 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U1919 ( .A(n1243), .B(n1242), .Z(n1360) );
  OR U1920 ( .A(n1245), .B(n1244), .Z(n1249) );
  OR U1921 ( .A(n1247), .B(n1246), .Z(n1248) );
  AND U1922 ( .A(n1249), .B(n1248), .Z(n1468) );
  ANDN U1923 ( .B(y[650]), .A(n167), .Z(n2202) );
  NANDN U1924 ( .A(n1250), .B(n2202), .Z(n1254) );
  OR U1925 ( .A(n1252), .B(n1251), .Z(n1253) );
  NAND U1926 ( .A(n1254), .B(n1253), .Z(n1406) );
  AND U1927 ( .A(x[141]), .B(y[647]), .Z(n1256) );
  NAND U1928 ( .A(n1256), .B(n1255), .Z(n1260) );
  OR U1929 ( .A(n1258), .B(n1257), .Z(n1259) );
  NAND U1930 ( .A(n1260), .B(n1259), .Z(n1444) );
  NAND U1931 ( .A(x[130]), .B(y[658]), .Z(n1432) );
  AND U1932 ( .A(y[650]), .B(x[138]), .Z(n1262) );
  NAND U1933 ( .A(x[144]), .B(y[644]), .Z(n1261) );
  XNOR U1934 ( .A(n1262), .B(n1261), .Z(n1431) );
  AND U1935 ( .A(y[645]), .B(x[143]), .Z(n1264) );
  NAND U1936 ( .A(x[137]), .B(y[651]), .Z(n1263) );
  XOR U1937 ( .A(n1264), .B(n1263), .Z(n1391) );
  AND U1938 ( .A(x[142]), .B(y[646]), .Z(n1390) );
  XNOR U1939 ( .A(n1391), .B(n1390), .Z(n1441) );
  XNOR U1940 ( .A(n1444), .B(n1443), .Z(n1407) );
  ANDN U1941 ( .B(y[652]), .A(n162), .Z(n1859) );
  NANDN U1942 ( .A(n1265), .B(n1859), .Z(n1269) );
  OR U1943 ( .A(n1267), .B(n1266), .Z(n1268) );
  AND U1944 ( .A(n1269), .B(n1268), .Z(n1450) );
  AND U1945 ( .A(y[641]), .B(x[147]), .Z(n1394) );
  XNOR U1946 ( .A(o[20]), .B(n1394), .Z(n1397) );
  AND U1947 ( .A(y[649]), .B(x[139]), .Z(n1271) );
  AND U1948 ( .A(y[659]), .B(x[129]), .Z(n1270) );
  XNOR U1949 ( .A(n1271), .B(n1270), .Z(n1396) );
  XNOR U1950 ( .A(n1397), .B(n1396), .Z(n1448) );
  NANDN U1951 ( .A(n1272), .B(o[19]), .Z(n1415) );
  NAND U1952 ( .A(x[148]), .B(y[640]), .Z(n1413) );
  NAND U1953 ( .A(x[128]), .B(y[660]), .Z(n1412) );
  XOR U1954 ( .A(n1413), .B(n1412), .Z(n1414) );
  XNOR U1955 ( .A(n1415), .B(n1414), .Z(n1447) );
  XOR U1956 ( .A(n1448), .B(n1447), .Z(n1449) );
  XOR U1957 ( .A(n1450), .B(n1449), .Z(n1408) );
  NANDN U1958 ( .A(n1274), .B(n1273), .Z(n1278) );
  NANDN U1959 ( .A(n1276), .B(n1275), .Z(n1277) );
  NAND U1960 ( .A(n1278), .B(n1277), .Z(n1365) );
  NANDN U1961 ( .A(n1280), .B(n1279), .Z(n1284) );
  NANDN U1962 ( .A(n1282), .B(n1281), .Z(n1283) );
  AND U1963 ( .A(n1284), .B(n1283), .Z(n1366) );
  XOR U1964 ( .A(n1367), .B(n1368), .Z(n1456) );
  NAND U1965 ( .A(n1286), .B(n1285), .Z(n1290) );
  NAND U1966 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U1967 ( .A(n1290), .B(n1289), .Z(n1454) );
  NAND U1968 ( .A(n1292), .B(n1291), .Z(n1296) );
  NANDN U1969 ( .A(n1294), .B(n1293), .Z(n1295) );
  NAND U1970 ( .A(n1296), .B(n1295), .Z(n1403) );
  ANDN U1971 ( .B(y[654]), .A(n157), .Z(n1377) );
  NAND U1972 ( .A(n1377), .B(n1297), .Z(n1300) );
  NANDN U1973 ( .A(n1418), .B(n1298), .Z(n1299) );
  NAND U1974 ( .A(n1300), .B(n1299), .Z(n1373) );
  OR U1975 ( .A(n1302), .B(n1301), .Z(n1306) );
  NANDN U1976 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1977 ( .A(n1306), .B(n1305), .Z(n1371) );
  AND U1978 ( .A(y[648]), .B(x[140]), .Z(n1308) );
  NAND U1979 ( .A(x[146]), .B(y[642]), .Z(n1307) );
  XOR U1980 ( .A(n1308), .B(n1307), .Z(n1385) );
  NAND U1981 ( .A(x[145]), .B(y[643]), .Z(n1384) );
  XNOR U1982 ( .A(n1385), .B(n1384), .Z(n1372) );
  XOR U1983 ( .A(n1371), .B(n1372), .Z(n1374) );
  NAND U1984 ( .A(x[135]), .B(y[653]), .Z(n1420) );
  AND U1985 ( .A(x[133]), .B(y[655]), .Z(n1310) );
  NAND U1986 ( .A(x[132]), .B(y[656]), .Z(n1309) );
  XOR U1987 ( .A(n1310), .B(n1309), .Z(n1419) );
  XNOR U1988 ( .A(n1420), .B(n1419), .Z(n1378) );
  NAND U1989 ( .A(y[652]), .B(x[136]), .Z(n1427) );
  AND U1990 ( .A(y[657]), .B(x[131]), .Z(n1312) );
  NAND U1991 ( .A(y[647]), .B(x[141]), .Z(n1311) );
  XNOR U1992 ( .A(n1312), .B(n1311), .Z(n1426) );
  XNOR U1993 ( .A(n1380), .B(n1379), .Z(n1438) );
  IV U1994 ( .A(y[651]), .Z(n1388) );
  ANDN U1995 ( .B(x[142]), .A(n1388), .Z(n2057) );
  NAND U1996 ( .A(n2057), .B(n1313), .Z(n1317) );
  OR U1997 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1998 ( .A(n1317), .B(n1316), .Z(n1436) );
  ANDN U1999 ( .B(y[649]), .A(n168), .Z(n2215) );
  NANDN U2000 ( .A(n1318), .B(n2215), .Z(n1322) );
  NANDN U2001 ( .A(n1320), .B(n1319), .Z(n1321) );
  AND U2002 ( .A(n1322), .B(n1321), .Z(n1435) );
  XOR U2003 ( .A(n1438), .B(n1437), .Z(n1401) );
  XNOR U2004 ( .A(n1400), .B(n1401), .Z(n1402) );
  XNOR U2005 ( .A(n1403), .B(n1402), .Z(n1453) );
  XOR U2006 ( .A(n1454), .B(n1453), .Z(n1455) );
  XNOR U2007 ( .A(n1456), .B(n1455), .Z(n1466) );
  OR U2008 ( .A(n1324), .B(n1323), .Z(n1328) );
  OR U2009 ( .A(n1326), .B(n1325), .Z(n1327) );
  NAND U2010 ( .A(n1328), .B(n1327), .Z(n1460) );
  OR U2011 ( .A(n1330), .B(n1329), .Z(n1334) );
  NANDN U2012 ( .A(n1332), .B(n1331), .Z(n1333) );
  NAND U2013 ( .A(n1334), .B(n1333), .Z(n1459) );
  XOR U2014 ( .A(n1460), .B(n1459), .Z(n1461) );
  OR U2015 ( .A(n1336), .B(n1335), .Z(n1340) );
  OR U2016 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U2017 ( .A(n1340), .B(n1339), .Z(n1462) );
  XOR U2018 ( .A(n1466), .B(n1465), .Z(n1467) );
  XOR U2019 ( .A(n1468), .B(n1467), .Z(n1359) );
  XOR U2020 ( .A(n1361), .B(n1362), .Z(n1355) );
  NANDN U2021 ( .A(n1342), .B(n1341), .Z(n1346) );
  NANDN U2022 ( .A(n1344), .B(n1343), .Z(n1345) );
  NAND U2023 ( .A(n1346), .B(n1345), .Z(n1353) );
  NANDN U2024 ( .A(n1348), .B(n1347), .Z(n1352) );
  NANDN U2025 ( .A(n1350), .B(n1349), .Z(n1351) );
  NAND U2026 ( .A(n1352), .B(n1351), .Z(n1354) );
  XNOR U2027 ( .A(n1353), .B(n1354), .Z(n1356) );
  XNOR U2028 ( .A(n1355), .B(n1356), .Z(N53) );
  NANDN U2029 ( .A(n1354), .B(n1353), .Z(n1358) );
  NAND U2030 ( .A(n1356), .B(n1355), .Z(n1357) );
  NAND U2031 ( .A(n1358), .B(n1357), .Z(n1471) );
  NANDN U2032 ( .A(n1360), .B(n1359), .Z(n1364) );
  OR U2033 ( .A(n1362), .B(n1361), .Z(n1363) );
  AND U2034 ( .A(n1364), .B(n1363), .Z(n1472) );
  XNOR U2035 ( .A(n1471), .B(n1472), .Z(n1473) );
  NANDN U2036 ( .A(n1366), .B(n1365), .Z(n1370) );
  NAND U2037 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U2038 ( .A(n1370), .B(n1369), .Z(n1593) );
  NANDN U2039 ( .A(n1372), .B(n1371), .Z(n1376) );
  NANDN U2040 ( .A(n1374), .B(n1373), .Z(n1375) );
  NAND U2041 ( .A(n1376), .B(n1375), .Z(n1503) );
  NANDN U2042 ( .A(n1378), .B(n1377), .Z(n1382) );
  NANDN U2043 ( .A(n1380), .B(n1379), .Z(n1381) );
  NAND U2044 ( .A(n1382), .B(n1381), .Z(n1502) );
  ANDN U2045 ( .B(y[648]), .A(n169), .Z(n2213) );
  NAND U2046 ( .A(n1383), .B(n2213), .Z(n1387) );
  OR U2047 ( .A(n1385), .B(n1384), .Z(n1386) );
  AND U2048 ( .A(n1387), .B(n1386), .Z(n1521) );
  ANDN U2049 ( .B(y[656]), .A(n156), .Z(n1551) );
  AND U2050 ( .A(x[144]), .B(y[645]), .Z(n1550) );
  XOR U2051 ( .A(n1551), .B(n1550), .Z(n1553) );
  ANDN U2052 ( .B(x[143]), .A(n2618), .Z(n1552) );
  XOR U2053 ( .A(n1553), .B(n1552), .Z(n1579) );
  NOR U2054 ( .A(n1388), .B(n166), .Z(n2207) );
  NAND U2055 ( .A(n2207), .B(n1389), .Z(n1393) );
  NANDN U2056 ( .A(n1391), .B(n1390), .Z(n1392) );
  NAND U2057 ( .A(n1393), .B(n1392), .Z(n1580) );
  XNOR U2058 ( .A(n1579), .B(n1580), .Z(n1582) );
  NAND U2059 ( .A(x[128]), .B(y[661]), .Z(n1570) );
  AND U2060 ( .A(n1394), .B(o[20]), .Z(n1568) );
  NAND U2061 ( .A(x[149]), .B(y[640]), .Z(n1567) );
  XNOR U2062 ( .A(n1568), .B(n1567), .Z(n1569) );
  XNOR U2063 ( .A(n1570), .B(n1569), .Z(n1581) );
  XNOR U2064 ( .A(n1582), .B(n1581), .Z(n1519) );
  ANDN U2065 ( .B(y[659]), .A(n162), .Z(n2958) );
  NAND U2066 ( .A(n2958), .B(n1395), .Z(n1399) );
  OR U2067 ( .A(n1397), .B(n1396), .Z(n1398) );
  AND U2068 ( .A(n1399), .B(n1398), .Z(n1520) );
  XOR U2069 ( .A(n1519), .B(n1520), .Z(n1522) );
  XOR U2070 ( .A(n1521), .B(n1522), .Z(n1501) );
  XNOR U2071 ( .A(n1502), .B(n1501), .Z(n1504) );
  XNOR U2072 ( .A(n1503), .B(n1504), .Z(n1591) );
  NANDN U2073 ( .A(n1401), .B(n1400), .Z(n1405) );
  NANDN U2074 ( .A(n1403), .B(n1402), .Z(n1404) );
  NAND U2075 ( .A(n1405), .B(n1404), .Z(n1592) );
  XOR U2076 ( .A(n1591), .B(n1592), .Z(n1594) );
  NANDN U2077 ( .A(n1407), .B(n1406), .Z(n1411) );
  NAND U2078 ( .A(n1409), .B(n1408), .Z(n1410) );
  NAND U2079 ( .A(n1411), .B(n1410), .Z(n1491) );
  OR U2080 ( .A(n1413), .B(n1412), .Z(n1417) );
  NANDN U2081 ( .A(n1415), .B(n1414), .Z(n1416) );
  AND U2082 ( .A(n1417), .B(n1416), .Z(n1507) );
  NANDN U2083 ( .A(n1418), .B(n1551), .Z(n1422) );
  OR U2084 ( .A(n1420), .B(n1419), .Z(n1421) );
  AND U2085 ( .A(n1422), .B(n1421), .Z(n1508) );
  XOR U2086 ( .A(n1507), .B(n1508), .Z(n1510) );
  ANDN U2087 ( .B(y[655]), .A(n157), .Z(n1563) );
  IV U2088 ( .A(y[654]), .Z(n2238) );
  NOR U2089 ( .A(n158), .B(n2238), .Z(n1852) );
  ANDN U2090 ( .B(x[142]), .A(n143), .Z(n1562) );
  XNOR U2091 ( .A(n1852), .B(n1562), .Z(n1564) );
  XNOR U2092 ( .A(n1563), .B(n1564), .Z(n1533) );
  AND U2093 ( .A(x[136]), .B(y[653]), .Z(n1967) );
  XNOR U2094 ( .A(n1531), .B(n1967), .Z(n1532) );
  XNOR U2095 ( .A(n1533), .B(n1532), .Z(n1587) );
  NAND U2096 ( .A(x[132]), .B(y[657]), .Z(n1559) );
  AND U2097 ( .A(x[141]), .B(y[648]), .Z(n1424) );
  AND U2098 ( .A(y[658]), .B(x[131]), .Z(n1423) );
  XNOR U2099 ( .A(n1424), .B(n1423), .Z(n1558) );
  XOR U2100 ( .A(n1559), .B(n1558), .Z(n1585) );
  NAND U2101 ( .A(x[140]), .B(y[649]), .Z(n1538) );
  ANDN U2102 ( .B(y[659]), .A(n153), .Z(n1537) );
  NAND U2103 ( .A(x[145]), .B(y[644]), .Z(n1536) );
  XOR U2104 ( .A(n1537), .B(n1536), .Z(n1539) );
  XNOR U2105 ( .A(n1538), .B(n1539), .Z(n1586) );
  XNOR U2106 ( .A(n1510), .B(n1509), .Z(n1527) );
  IV U2107 ( .A(y[660]), .Z(n2590) );
  ANDN U2108 ( .B(x[129]), .A(n2590), .Z(n1573) );
  ANDN U2109 ( .B(x[146]), .A(n141), .Z(n1574) );
  XNOR U2110 ( .A(n1573), .B(n1574), .Z(n1576) );
  XNOR U2111 ( .A(n1575), .B(n1576), .Z(n1513) );
  NAND U2112 ( .A(y[650]), .B(x[139]), .Z(n1547) );
  AND U2113 ( .A(x[148]), .B(y[641]), .Z(n1556) );
  XNOR U2114 ( .A(o[21]), .B(n1556), .Z(n1545) );
  NAND U2115 ( .A(y[642]), .B(x[147]), .Z(n1544) );
  XOR U2116 ( .A(n1545), .B(n1544), .Z(n1546) );
  XOR U2117 ( .A(n1547), .B(n1546), .Z(n1514) );
  XOR U2118 ( .A(n1513), .B(n1514), .Z(n1516) );
  AND U2119 ( .A(y[657]), .B(x[141]), .Z(n2717) );
  NAND U2120 ( .A(n2717), .B(n1425), .Z(n1429) );
  NANDN U2121 ( .A(n1427), .B(n1426), .Z(n1428) );
  AND U2122 ( .A(n1429), .B(n1428), .Z(n1515) );
  XOR U2123 ( .A(n1516), .B(n1515), .Z(n1526) );
  NAND U2124 ( .A(n1430), .B(n2202), .Z(n1434) );
  NANDN U2125 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U2126 ( .A(n1434), .B(n1433), .Z(n1525) );
  XNOR U2127 ( .A(n1526), .B(n1525), .Z(n1528) );
  XNOR U2128 ( .A(n1527), .B(n1528), .Z(n1490) );
  NANDN U2129 ( .A(n1436), .B(n1435), .Z(n1440) );
  NANDN U2130 ( .A(n1438), .B(n1437), .Z(n1439) );
  AND U2131 ( .A(n1440), .B(n1439), .Z(n1495) );
  NAND U2132 ( .A(n1442), .B(n1441), .Z(n1446) );
  NAND U2133 ( .A(n1444), .B(n1443), .Z(n1445) );
  NAND U2134 ( .A(n1446), .B(n1445), .Z(n1496) );
  XOR U2135 ( .A(n1495), .B(n1496), .Z(n1497) );
  NANDN U2136 ( .A(n1448), .B(n1447), .Z(n1452) );
  OR U2137 ( .A(n1450), .B(n1449), .Z(n1451) );
  NAND U2138 ( .A(n1452), .B(n1451), .Z(n1498) );
  XNOR U2139 ( .A(n1497), .B(n1498), .Z(n1489) );
  XNOR U2140 ( .A(n1490), .B(n1489), .Z(n1492) );
  XOR U2141 ( .A(n1491), .B(n1492), .Z(n1483) );
  NANDN U2142 ( .A(n1454), .B(n1453), .Z(n1458) );
  OR U2143 ( .A(n1456), .B(n1455), .Z(n1457) );
  AND U2144 ( .A(n1458), .B(n1457), .Z(n1484) );
  XOR U2145 ( .A(n1483), .B(n1484), .Z(n1486) );
  XNOR U2146 ( .A(n1485), .B(n1486), .Z(n1479) );
  OR U2147 ( .A(n1460), .B(n1459), .Z(n1464) );
  NANDN U2148 ( .A(n1462), .B(n1461), .Z(n1463) );
  NAND U2149 ( .A(n1464), .B(n1463), .Z(n1478) );
  NAND U2150 ( .A(n1466), .B(n1465), .Z(n1470) );
  NANDN U2151 ( .A(n1468), .B(n1467), .Z(n1469) );
  NAND U2152 ( .A(n1470), .B(n1469), .Z(n1477) );
  XNOR U2153 ( .A(n1478), .B(n1477), .Z(n1480) );
  XOR U2154 ( .A(n1479), .B(n1480), .Z(n1474) );
  XOR U2155 ( .A(n1473), .B(n1474), .Z(N54) );
  NANDN U2156 ( .A(n1472), .B(n1471), .Z(n1476) );
  NANDN U2157 ( .A(n1474), .B(n1473), .Z(n1475) );
  NAND U2158 ( .A(n1476), .B(n1475), .Z(n1597) );
  OR U2159 ( .A(n1478), .B(n1477), .Z(n1482) );
  NANDN U2160 ( .A(n1480), .B(n1479), .Z(n1481) );
  AND U2161 ( .A(n1482), .B(n1481), .Z(n1598) );
  XNOR U2162 ( .A(n1597), .B(n1598), .Z(n1599) );
  NANDN U2163 ( .A(n1484), .B(n1483), .Z(n1488) );
  NANDN U2164 ( .A(n1486), .B(n1485), .Z(n1487) );
  NAND U2165 ( .A(n1488), .B(n1487), .Z(n1606) );
  OR U2166 ( .A(n1490), .B(n1489), .Z(n1494) );
  NANDN U2167 ( .A(n1492), .B(n1491), .Z(n1493) );
  NAND U2168 ( .A(n1494), .B(n1493), .Z(n1726) );
  OR U2169 ( .A(n1496), .B(n1495), .Z(n1500) );
  NANDN U2170 ( .A(n1498), .B(n1497), .Z(n1499) );
  AND U2171 ( .A(n1500), .B(n1499), .Z(n1725) );
  XOR U2172 ( .A(n1726), .B(n1725), .Z(n1727) );
  NAND U2173 ( .A(n1502), .B(n1501), .Z(n1506) );
  NANDN U2174 ( .A(n1504), .B(n1503), .Z(n1505) );
  NAND U2175 ( .A(n1506), .B(n1505), .Z(n1610) );
  OR U2176 ( .A(n1508), .B(n1507), .Z(n1512) );
  NAND U2177 ( .A(n1510), .B(n1509), .Z(n1511) );
  AND U2178 ( .A(n1512), .B(n1511), .Z(n1615) );
  NANDN U2179 ( .A(n1514), .B(n1513), .Z(n1518) );
  OR U2180 ( .A(n1516), .B(n1515), .Z(n1517) );
  AND U2181 ( .A(n1518), .B(n1517), .Z(n1616) );
  XOR U2182 ( .A(n1615), .B(n1616), .Z(n1617) );
  NANDN U2183 ( .A(n1520), .B(n1519), .Z(n1524) );
  OR U2184 ( .A(n1522), .B(n1521), .Z(n1523) );
  AND U2185 ( .A(n1524), .B(n1523), .Z(n1618) );
  XNOR U2186 ( .A(n1617), .B(n1618), .Z(n1609) );
  XNOR U2187 ( .A(n1610), .B(n1609), .Z(n1612) );
  OR U2188 ( .A(n1526), .B(n1525), .Z(n1530) );
  NANDN U2189 ( .A(n1528), .B(n1527), .Z(n1529) );
  NAND U2190 ( .A(n1530), .B(n1529), .Z(n1704) );
  OR U2191 ( .A(n1531), .B(n1967), .Z(n1535) );
  OR U2192 ( .A(n1533), .B(n1532), .Z(n1534) );
  AND U2193 ( .A(n1535), .B(n1534), .Z(n1721) );
  NANDN U2194 ( .A(n1537), .B(n1536), .Z(n1541) );
  NANDN U2195 ( .A(n1539), .B(n1538), .Z(n1540) );
  NAND U2196 ( .A(n1541), .B(n1540), .Z(n1698) );
  NAND U2197 ( .A(x[132]), .B(y[658]), .Z(n1635) );
  AND U2198 ( .A(y[650]), .B(x[140]), .Z(n1543) );
  AND U2199 ( .A(y[644]), .B(x[146]), .Z(n1542) );
  XNOR U2200 ( .A(n1543), .B(n1542), .Z(n1634) );
  XOR U2201 ( .A(n1635), .B(n1634), .Z(n1695) );
  NAND U2202 ( .A(x[144]), .B(y[646]), .Z(n1653) );
  NAND U2203 ( .A(x[145]), .B(y[645]), .Z(n1651) );
  NAND U2204 ( .A(x[133]), .B(y[657]), .Z(n1650) );
  XNOR U2205 ( .A(n1651), .B(n1650), .Z(n1652) );
  XNOR U2206 ( .A(n1653), .B(n1652), .Z(n1696) );
  XNOR U2207 ( .A(n1698), .B(n1697), .Z(n1719) );
  OR U2208 ( .A(n1545), .B(n1544), .Z(n1549) );
  NANDN U2209 ( .A(n1547), .B(n1546), .Z(n1548) );
  NAND U2210 ( .A(n1549), .B(n1548), .Z(n1720) );
  XNOR U2211 ( .A(n1719), .B(n1720), .Z(n1722) );
  XOR U2212 ( .A(n1721), .B(n1722), .Z(n1702) );
  NAND U2213 ( .A(x[148]), .B(y[642]), .Z(n1647) );
  NAND U2214 ( .A(y[649]), .B(x[141]), .Z(n1645) );
  NAND U2215 ( .A(x[130]), .B(y[660]), .Z(n1644) );
  XNOR U2216 ( .A(n1645), .B(n1644), .Z(n1646) );
  XNOR U2217 ( .A(n1647), .B(n1646), .Z(n1624) );
  NAND U2218 ( .A(y[647]), .B(x[143]), .Z(n1660) );
  NAND U2219 ( .A(y[652]), .B(x[138]), .Z(n1658) );
  NAND U2220 ( .A(x[134]), .B(y[656]), .Z(n1657) );
  XNOR U2221 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U2222 ( .A(n1660), .B(n1659), .Z(n1622) );
  NAND U2223 ( .A(n1551), .B(n1550), .Z(n1555) );
  NAND U2224 ( .A(n1553), .B(n1552), .Z(n1554) );
  AND U2225 ( .A(n1555), .B(n1554), .Z(n1621) );
  XNOR U2226 ( .A(n1622), .B(n1621), .Z(n1623) );
  XNOR U2227 ( .A(n1624), .B(n1623), .Z(n1713) );
  NAND U2228 ( .A(y[643]), .B(x[147]), .Z(n1690) );
  NAND U2229 ( .A(x[131]), .B(y[659]), .Z(n1688) );
  NAND U2230 ( .A(x[142]), .B(y[648]), .Z(n1687) );
  XNOR U2231 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U2232 ( .A(n1690), .B(n1689), .Z(n1670) );
  NAND U2233 ( .A(o[21]), .B(n1556), .Z(n1684) );
  AND U2234 ( .A(y[661]), .B(x[129]), .Z(n1681) );
  XNOR U2235 ( .A(n1682), .B(n1681), .Z(n1683) );
  XOR U2236 ( .A(n1684), .B(n1683), .Z(n1669) );
  XOR U2237 ( .A(n1670), .B(n1669), .Z(n1672) );
  IV U2238 ( .A(y[658]), .Z(n2616) );
  ANDN U2239 ( .B(x[141]), .A(n2616), .Z(n2977) );
  NAND U2240 ( .A(n1557), .B(n2977), .Z(n1561) );
  OR U2241 ( .A(n1559), .B(n1558), .Z(n1560) );
  AND U2242 ( .A(n1561), .B(n1560), .Z(n1671) );
  XOR U2243 ( .A(n1672), .B(n1671), .Z(n1714) );
  XOR U2244 ( .A(n1713), .B(n1714), .Z(n1716) );
  AND U2245 ( .A(x[135]), .B(y[655]), .Z(n1565) );
  XNOR U2246 ( .A(n1566), .B(n1565), .Z(n1630) );
  XOR U2247 ( .A(n1629), .B(n1630), .Z(n1664) );
  NAND U2248 ( .A(x[128]), .B(y[662]), .Z(n1639) );
  AND U2249 ( .A(y[640]), .B(x[150]), .Z(n1638) );
  XNOR U2250 ( .A(n1639), .B(n1638), .Z(n1641) );
  NAND U2251 ( .A(y[641]), .B(x[149]), .Z(n1656) );
  XNOR U2252 ( .A(n1656), .B(o[22]), .Z(n1640) );
  XNOR U2253 ( .A(n1641), .B(n1640), .Z(n1663) );
  XOR U2254 ( .A(n1664), .B(n1663), .Z(n1665) );
  NANDN U2255 ( .A(n1568), .B(n1567), .Z(n1572) );
  NAND U2256 ( .A(n1570), .B(n1569), .Z(n1571) );
  AND U2257 ( .A(n1572), .B(n1571), .Z(n1676) );
  OR U2258 ( .A(n1574), .B(n1573), .Z(n1578) );
  OR U2259 ( .A(n1576), .B(n1575), .Z(n1577) );
  AND U2260 ( .A(n1578), .B(n1577), .Z(n1675) );
  XNOR U2261 ( .A(n1676), .B(n1675), .Z(n1677) );
  XNOR U2262 ( .A(n1678), .B(n1677), .Z(n1715) );
  XNOR U2263 ( .A(n1716), .B(n1715), .Z(n1710) );
  OR U2264 ( .A(n1580), .B(n1579), .Z(n1584) );
  OR U2265 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U2266 ( .A(n1584), .B(n1583), .Z(n1707) );
  NANDN U2267 ( .A(n1586), .B(n1585), .Z(n1590) );
  NAND U2268 ( .A(n1588), .B(n1587), .Z(n1589) );
  NAND U2269 ( .A(n1590), .B(n1589), .Z(n1708) );
  XNOR U2270 ( .A(n1707), .B(n1708), .Z(n1709) );
  XNOR U2271 ( .A(n1710), .B(n1709), .Z(n1701) );
  XOR U2272 ( .A(n1702), .B(n1701), .Z(n1703) );
  XOR U2273 ( .A(n1704), .B(n1703), .Z(n1611) );
  XNOR U2274 ( .A(n1612), .B(n1611), .Z(n1728) );
  XNOR U2275 ( .A(n1727), .B(n1728), .Z(n1604) );
  NANDN U2276 ( .A(n1592), .B(n1591), .Z(n1596) );
  NANDN U2277 ( .A(n1594), .B(n1593), .Z(n1595) );
  AND U2278 ( .A(n1596), .B(n1595), .Z(n1603) );
  XOR U2279 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U2280 ( .A(n1606), .B(n1605), .Z(n1600) );
  XOR U2281 ( .A(n1599), .B(n1600), .Z(N55) );
  NANDN U2282 ( .A(n1598), .B(n1597), .Z(n1602) );
  NANDN U2283 ( .A(n1600), .B(n1599), .Z(n1601) );
  NAND U2284 ( .A(n1602), .B(n1601), .Z(n1731) );
  OR U2285 ( .A(n1604), .B(n1603), .Z(n1608) );
  NANDN U2286 ( .A(n1606), .B(n1605), .Z(n1607) );
  NAND U2287 ( .A(n1608), .B(n1607), .Z(n1732) );
  XNOR U2288 ( .A(n1731), .B(n1732), .Z(n1733) );
  OR U2289 ( .A(n1610), .B(n1609), .Z(n1614) );
  OR U2290 ( .A(n1612), .B(n1611), .Z(n1613) );
  AND U2291 ( .A(n1614), .B(n1613), .Z(n1737) );
  OR U2292 ( .A(n1616), .B(n1615), .Z(n1620) );
  NANDN U2293 ( .A(n1618), .B(n1617), .Z(n1619) );
  AND U2294 ( .A(n1620), .B(n1619), .Z(n1757) );
  OR U2295 ( .A(n1622), .B(n1621), .Z(n1626) );
  OR U2296 ( .A(n1624), .B(n1623), .Z(n1625) );
  AND U2297 ( .A(n1626), .B(n1625), .Z(n1827) );
  AND U2298 ( .A(y[641]), .B(x[150]), .Z(n1845) );
  XNOR U2299 ( .A(o[23]), .B(n1845), .Z(n1836) );
  NAND U2300 ( .A(y[640]), .B(x[151]), .Z(n1834) );
  NAND U2301 ( .A(x[128]), .B(y[663]), .Z(n1833) );
  XNOR U2302 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U2303 ( .A(n1836), .B(n1835), .Z(n1775) );
  ANDN U2304 ( .B(x[147]), .A(n2634), .Z(n2100) );
  AND U2305 ( .A(x[148]), .B(y[643]), .Z(n1628) );
  XNOR U2306 ( .A(n1628), .B(n1627), .Z(n1842) );
  XNOR U2307 ( .A(n2100), .B(n1842), .Z(n1773) );
  NAND U2308 ( .A(n1852), .B(n1853), .Z(n1632) );
  NANDN U2309 ( .A(n1630), .B(n1629), .Z(n1631) );
  NAND U2310 ( .A(n1632), .B(n1631), .Z(n1774) );
  XNOR U2311 ( .A(n1773), .B(n1774), .Z(n1776) );
  XOR U2312 ( .A(n1775), .B(n1776), .Z(n1782) );
  ANDN U2313 ( .B(x[146]), .A(n2627), .Z(n2628) );
  NAND U2314 ( .A(n1633), .B(n2628), .Z(n1637) );
  OR U2315 ( .A(n1635), .B(n1634), .Z(n1636) );
  AND U2316 ( .A(n1637), .B(n1636), .Z(n1779) );
  NANDN U2317 ( .A(n1639), .B(n1638), .Z(n1643) );
  NAND U2318 ( .A(n1641), .B(n1640), .Z(n1642) );
  AND U2319 ( .A(n1643), .B(n1642), .Z(n1780) );
  XOR U2320 ( .A(n1779), .B(n1780), .Z(n1781) );
  XOR U2321 ( .A(n1782), .B(n1781), .Z(n1828) );
  XOR U2322 ( .A(n1827), .B(n1828), .Z(n1829) );
  OR U2323 ( .A(n1645), .B(n1644), .Z(n1649) );
  OR U2324 ( .A(n1647), .B(n1646), .Z(n1648) );
  AND U2325 ( .A(n1649), .B(n1648), .Z(n1865) );
  OR U2326 ( .A(n1651), .B(n1650), .Z(n1655) );
  OR U2327 ( .A(n1653), .B(n1652), .Z(n1654) );
  AND U2328 ( .A(n1655), .B(n1654), .Z(n1791) );
  NANDN U2329 ( .A(n1656), .B(o[22]), .Z(n1849) );
  NAND U2330 ( .A(x[129]), .B(y[662]), .Z(n1847) );
  NAND U2331 ( .A(x[140]), .B(y[651]), .Z(n1846) );
  XNOR U2332 ( .A(n1847), .B(n1846), .Z(n1848) );
  XNOR U2333 ( .A(n1849), .B(n1848), .Z(n1792) );
  XOR U2334 ( .A(n1791), .B(n1792), .Z(n1794) );
  NAND U2335 ( .A(x[149]), .B(y[642]), .Z(n1812) );
  NAND U2336 ( .A(x[130]), .B(y[661]), .Z(n1810) );
  AND U2337 ( .A(y[650]), .B(x[141]), .Z(n1809) );
  XNOR U2338 ( .A(n1810), .B(n1809), .Z(n1811) );
  XNOR U2339 ( .A(n1794), .B(n1793), .Z(n1866) );
  XOR U2340 ( .A(n1865), .B(n1866), .Z(n1867) );
  NAND U2341 ( .A(x[132]), .B(y[659]), .Z(n1818) );
  NAND U2342 ( .A(y[660]), .B(x[131]), .Z(n1816) );
  XNOR U2343 ( .A(n1818), .B(n1817), .Z(n1786) );
  NAND U2344 ( .A(x[145]), .B(y[646]), .Z(n1824) );
  NAND U2345 ( .A(x[146]), .B(y[645]), .Z(n1822) );
  AND U2346 ( .A(x[133]), .B(y[658]), .Z(n1821) );
  XNOR U2347 ( .A(n1822), .B(n1821), .Z(n1823) );
  XOR U2348 ( .A(n1786), .B(n1785), .Z(n1788) );
  OR U2349 ( .A(n1658), .B(n1657), .Z(n1662) );
  OR U2350 ( .A(n1660), .B(n1659), .Z(n1661) );
  AND U2351 ( .A(n1662), .B(n1661), .Z(n1787) );
  XNOR U2352 ( .A(n1788), .B(n1787), .Z(n1868) );
  XOR U2353 ( .A(n1867), .B(n1868), .Z(n1830) );
  XOR U2354 ( .A(n1829), .B(n1830), .Z(n1756) );
  OR U2355 ( .A(n1664), .B(n1663), .Z(n1668) );
  NANDN U2356 ( .A(n1666), .B(n1665), .Z(n1667) );
  AND U2357 ( .A(n1668), .B(n1667), .Z(n1767) );
  NANDN U2358 ( .A(n1670), .B(n1669), .Z(n1674) );
  OR U2359 ( .A(n1672), .B(n1671), .Z(n1673) );
  AND U2360 ( .A(n1674), .B(n1673), .Z(n1768) );
  XOR U2361 ( .A(n1767), .B(n1768), .Z(n1769) );
  OR U2362 ( .A(n1676), .B(n1675), .Z(n1680) );
  OR U2363 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U2364 ( .A(n1680), .B(n1679), .Z(n1770) );
  NAND U2365 ( .A(n1682), .B(n1681), .Z(n1686) );
  OR U2366 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U2367 ( .A(n1686), .B(n1685), .Z(n1797) );
  OR U2368 ( .A(n1688), .B(n1687), .Z(n1692) );
  OR U2369 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U2370 ( .A(n1692), .B(n1691), .Z(n1798) );
  XOR U2371 ( .A(n1797), .B(n1798), .Z(n1800) );
  AND U2372 ( .A(x[135]), .B(y[656]), .Z(n1693) );
  XNOR U2373 ( .A(n1694), .B(n1693), .Z(n1854) );
  AND U2374 ( .A(x[138]), .B(y[653]), .Z(n1803) );
  XOR U2375 ( .A(n1804), .B(n1803), .Z(n1806) );
  NAND U2376 ( .A(y[648]), .B(x[143]), .Z(n1858) );
  NAND U2377 ( .A(x[134]), .B(y[657]), .Z(n1857) );
  XNOR U2378 ( .A(n1858), .B(n1857), .Z(n1860) );
  XOR U2379 ( .A(n1806), .B(n1805), .Z(n1799) );
  XNOR U2380 ( .A(n1800), .B(n1799), .Z(n1744) );
  NANDN U2381 ( .A(n1696), .B(n1695), .Z(n1700) );
  NANDN U2382 ( .A(n1698), .B(n1697), .Z(n1699) );
  AND U2383 ( .A(n1700), .B(n1699), .Z(n1743) );
  XOR U2384 ( .A(n1744), .B(n1743), .Z(n1745) );
  XNOR U2385 ( .A(n1756), .B(n1755), .Z(n1758) );
  XOR U2386 ( .A(n1757), .B(n1758), .Z(n1764) );
  NANDN U2387 ( .A(n1702), .B(n1701), .Z(n1706) );
  OR U2388 ( .A(n1704), .B(n1703), .Z(n1705) );
  NAND U2389 ( .A(n1706), .B(n1705), .Z(n1762) );
  OR U2390 ( .A(n1708), .B(n1707), .Z(n1712) );
  OR U2391 ( .A(n1710), .B(n1709), .Z(n1711) );
  AND U2392 ( .A(n1712), .B(n1711), .Z(n1751) );
  NANDN U2393 ( .A(n1714), .B(n1713), .Z(n1718) );
  OR U2394 ( .A(n1716), .B(n1715), .Z(n1717) );
  AND U2395 ( .A(n1718), .B(n1717), .Z(n1750) );
  OR U2396 ( .A(n1720), .B(n1719), .Z(n1724) );
  OR U2397 ( .A(n1722), .B(n1721), .Z(n1723) );
  AND U2398 ( .A(n1724), .B(n1723), .Z(n1749) );
  XNOR U2399 ( .A(n1750), .B(n1749), .Z(n1752) );
  XNOR U2400 ( .A(n1751), .B(n1752), .Z(n1761) );
  XOR U2401 ( .A(n1762), .B(n1761), .Z(n1763) );
  XOR U2402 ( .A(n1764), .B(n1763), .Z(n1738) );
  XOR U2403 ( .A(n1737), .B(n1738), .Z(n1739) );
  OR U2404 ( .A(n1726), .B(n1725), .Z(n1730) );
  NANDN U2405 ( .A(n1728), .B(n1727), .Z(n1729) );
  AND U2406 ( .A(n1730), .B(n1729), .Z(n1740) );
  XOR U2407 ( .A(n1733), .B(n1734), .Z(N56) );
  NANDN U2408 ( .A(n1732), .B(n1731), .Z(n1736) );
  NANDN U2409 ( .A(n1734), .B(n1733), .Z(n1735) );
  NAND U2410 ( .A(n1736), .B(n1735), .Z(n2003) );
  OR U2411 ( .A(n1738), .B(n1737), .Z(n1742) );
  NANDN U2412 ( .A(n1740), .B(n1739), .Z(n1741) );
  AND U2413 ( .A(n1742), .B(n1741), .Z(n2004) );
  XNOR U2414 ( .A(n2003), .B(n2004), .Z(n2005) );
  OR U2415 ( .A(n1744), .B(n1743), .Z(n1748) );
  NANDN U2416 ( .A(n1746), .B(n1745), .Z(n1747) );
  NAND U2417 ( .A(n1748), .B(n1747), .Z(n1872) );
  OR U2418 ( .A(n1750), .B(n1749), .Z(n1754) );
  OR U2419 ( .A(n1752), .B(n1751), .Z(n1753) );
  AND U2420 ( .A(n1754), .B(n1753), .Z(n1871) );
  XOR U2421 ( .A(n1872), .B(n1871), .Z(n1873) );
  OR U2422 ( .A(n1756), .B(n1755), .Z(n1760) );
  OR U2423 ( .A(n1758), .B(n1757), .Z(n1759) );
  NAND U2424 ( .A(n1760), .B(n1759), .Z(n1874) );
  OR U2425 ( .A(n1762), .B(n1761), .Z(n1766) );
  NANDN U2426 ( .A(n1764), .B(n1763), .Z(n1765) );
  AND U2427 ( .A(n1766), .B(n1765), .Z(n2010) );
  OR U2428 ( .A(n1768), .B(n1767), .Z(n1772) );
  NANDN U2429 ( .A(n1770), .B(n1769), .Z(n1771) );
  NAND U2430 ( .A(n1772), .B(n1771), .Z(n1998) );
  OR U2431 ( .A(n1774), .B(n1773), .Z(n1778) );
  OR U2432 ( .A(n1776), .B(n1775), .Z(n1777) );
  NAND U2433 ( .A(n1778), .B(n1777), .Z(n1878) );
  OR U2434 ( .A(n1780), .B(n1779), .Z(n1784) );
  NANDN U2435 ( .A(n1782), .B(n1781), .Z(n1783) );
  AND U2436 ( .A(n1784), .B(n1783), .Z(n1877) );
  XOR U2437 ( .A(n1878), .B(n1877), .Z(n1879) );
  NANDN U2438 ( .A(n1786), .B(n1785), .Z(n1790) );
  OR U2439 ( .A(n1788), .B(n1787), .Z(n1789) );
  AND U2440 ( .A(n1790), .B(n1789), .Z(n1880) );
  OR U2441 ( .A(n1792), .B(n1791), .Z(n1796) );
  NAND U2442 ( .A(n1794), .B(n1793), .Z(n1795) );
  AND U2443 ( .A(n1796), .B(n1795), .Z(n1883) );
  XNOR U2444 ( .A(n1884), .B(n1883), .Z(n1886) );
  OR U2445 ( .A(n1798), .B(n1797), .Z(n1802) );
  NAND U2446 ( .A(n1800), .B(n1799), .Z(n1801) );
  AND U2447 ( .A(n1802), .B(n1801), .Z(n1993) );
  NANDN U2448 ( .A(n1804), .B(n1803), .Z(n1808) );
  OR U2449 ( .A(n1806), .B(n1805), .Z(n1807) );
  AND U2450 ( .A(n1808), .B(n1807), .Z(n1992) );
  NANDN U2451 ( .A(n1810), .B(n1809), .Z(n1814) );
  NANDN U2452 ( .A(n1812), .B(n1811), .Z(n1813) );
  AND U2453 ( .A(n1814), .B(n1813), .Z(n1895) );
  NANDN U2454 ( .A(n1816), .B(n1815), .Z(n1820) );
  OR U2455 ( .A(n1818), .B(n1817), .Z(n1819) );
  AND U2456 ( .A(n1820), .B(n1819), .Z(n1896) );
  XOR U2457 ( .A(n1895), .B(n1896), .Z(n1898) );
  NAND U2458 ( .A(y[646]), .B(x[146]), .Z(n1988) );
  NAND U2459 ( .A(y[647]), .B(x[145]), .Z(n1986) );
  NAND U2460 ( .A(x[135]), .B(y[657]), .Z(n1985) );
  XNOR U2461 ( .A(n1986), .B(n1985), .Z(n1987) );
  XNOR U2462 ( .A(n1988), .B(n1987), .Z(n1914) );
  NANDN U2463 ( .A(n174), .B(y[641]), .Z(n1984) );
  XOR U2464 ( .A(o[24]), .B(n1984), .Z(n1946) );
  NAND U2465 ( .A(x[128]), .B(y[664]), .Z(n1944) );
  AND U2466 ( .A(x[152]), .B(y[640]), .Z(n1943) );
  XNOR U2467 ( .A(n1944), .B(n1943), .Z(n1945) );
  XNOR U2468 ( .A(n1914), .B(n1913), .Z(n1916) );
  NANDN U2469 ( .A(n1822), .B(n1821), .Z(n1826) );
  NANDN U2470 ( .A(n1824), .B(n1823), .Z(n1825) );
  AND U2471 ( .A(n1826), .B(n1825), .Z(n1915) );
  XOR U2472 ( .A(n1916), .B(n1915), .Z(n1897) );
  XOR U2473 ( .A(n1898), .B(n1897), .Z(n1991) );
  XOR U2474 ( .A(n1992), .B(n1991), .Z(n1994) );
  XNOR U2475 ( .A(n1993), .B(n1994), .Z(n1885) );
  XOR U2476 ( .A(n1886), .B(n1885), .Z(n1997) );
  XNOR U2477 ( .A(n1998), .B(n1997), .Z(n2000) );
  OR U2478 ( .A(n1828), .B(n1827), .Z(n1832) );
  NANDN U2479 ( .A(n1830), .B(n1829), .Z(n1831) );
  AND U2480 ( .A(n1832), .B(n1831), .Z(n1934) );
  NAND U2481 ( .A(y[660]), .B(x[132]), .Z(n1952) );
  NAND U2482 ( .A(x[131]), .B(y[661]), .Z(n1950) );
  NAND U2483 ( .A(y[649]), .B(x[143]), .Z(n1949) );
  XNOR U2484 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U2485 ( .A(n1952), .B(n1951), .Z(n1958) );
  OR U2486 ( .A(n1834), .B(n1833), .Z(n1838) );
  OR U2487 ( .A(n1836), .B(n1835), .Z(n1837) );
  AND U2488 ( .A(n1838), .B(n1837), .Z(n1956) );
  NAND U2489 ( .A(x[142]), .B(y[650]), .Z(n1969) );
  AND U2490 ( .A(x[139]), .B(y[653]), .Z(n1840) );
  AND U2491 ( .A(x[136]), .B(y[656]), .Z(n1839) );
  XNOR U2492 ( .A(n1840), .B(n1839), .Z(n1968) );
  XOR U2493 ( .A(n1969), .B(n1968), .Z(n1963) );
  ANDN U2494 ( .B(x[138]), .A(n2238), .Z(n1961) );
  ANDN U2495 ( .B(y[655]), .A(n160), .Z(n1962) );
  XNOR U2496 ( .A(n1961), .B(n1962), .Z(n1964) );
  XNOR U2497 ( .A(n1963), .B(n1964), .Z(n1955) );
  XOR U2498 ( .A(n1956), .B(n1955), .Z(n1957) );
  XOR U2499 ( .A(n1958), .B(n1957), .Z(n1939) );
  NAND U2500 ( .A(x[130]), .B(y[662]), .Z(n1979) );
  NAND U2501 ( .A(y[642]), .B(x[150]), .Z(n1978) );
  XNOR U2502 ( .A(n1979), .B(n1978), .Z(n1981) );
  AND U2503 ( .A(y[643]), .B(x[144]), .Z(n1841) );
  ANDN U2504 ( .B(y[647]), .A(n171), .Z(n2398) );
  NAND U2505 ( .A(n1841), .B(n2398), .Z(n1844) );
  NANDN U2506 ( .A(n1842), .B(n2100), .Z(n1843) );
  AND U2507 ( .A(n1844), .B(n1843), .Z(n1926) );
  NAND U2508 ( .A(n1845), .B(o[23]), .Z(n1975) );
  AND U2509 ( .A(y[663]), .B(x[129]), .Z(n1972) );
  XOR U2510 ( .A(n1973), .B(n1972), .Z(n1974) );
  XNOR U2511 ( .A(n1975), .B(n1974), .Z(n1925) );
  XOR U2512 ( .A(n1926), .B(n1925), .Z(n1927) );
  XNOR U2513 ( .A(n1928), .B(n1927), .Z(n1937) );
  OR U2514 ( .A(n1847), .B(n1846), .Z(n1851) );
  OR U2515 ( .A(n1849), .B(n1848), .Z(n1850) );
  AND U2516 ( .A(n1851), .B(n1850), .Z(n1892) );
  NAND U2517 ( .A(n1852), .B(n2028), .Z(n1856) );
  NANDN U2518 ( .A(n1854), .B(n1853), .Z(n1855) );
  AND U2519 ( .A(n1856), .B(n1855), .Z(n1890) );
  NAND U2520 ( .A(x[133]), .B(y[659]), .Z(n1906) );
  NAND U2521 ( .A(y[643]), .B(x[149]), .Z(n1904) );
  NAND U2522 ( .A(x[144]), .B(y[648]), .Z(n1903) );
  XNOR U2523 ( .A(n1904), .B(n1903), .Z(n1905) );
  XNOR U2524 ( .A(n1906), .B(n1905), .Z(n1922) );
  OR U2525 ( .A(n1858), .B(n1857), .Z(n1862) );
  NANDN U2526 ( .A(n1860), .B(n1859), .Z(n1861) );
  AND U2527 ( .A(n1862), .B(n1861), .Z(n1920) );
  NAND U2528 ( .A(y[658]), .B(x[134]), .Z(n1910) );
  AND U2529 ( .A(x[147]), .B(y[645]), .Z(n1864) );
  AND U2530 ( .A(y[644]), .B(x[148]), .Z(n1863) );
  XNOR U2531 ( .A(n1864), .B(n1863), .Z(n1909) );
  XOR U2532 ( .A(n1910), .B(n1909), .Z(n1919) );
  XOR U2533 ( .A(n1922), .B(n1921), .Z(n1889) );
  XNOR U2534 ( .A(n1890), .B(n1889), .Z(n1891) );
  XNOR U2535 ( .A(n1892), .B(n1891), .Z(n1938) );
  XOR U2536 ( .A(n1937), .B(n1938), .Z(n1940) );
  XNOR U2537 ( .A(n1939), .B(n1940), .Z(n1931) );
  OR U2538 ( .A(n1866), .B(n1865), .Z(n1870) );
  NANDN U2539 ( .A(n1868), .B(n1867), .Z(n1869) );
  AND U2540 ( .A(n1870), .B(n1869), .Z(n1932) );
  XNOR U2541 ( .A(n1931), .B(n1932), .Z(n1933) );
  XNOR U2542 ( .A(n1934), .B(n1933), .Z(n1999) );
  XOR U2543 ( .A(n2000), .B(n1999), .Z(n2009) );
  XOR U2544 ( .A(n2010), .B(n2009), .Z(n2011) );
  XNOR U2545 ( .A(n2012), .B(n2011), .Z(n2006) );
  XOR U2546 ( .A(n2005), .B(n2006), .Z(N57) );
  OR U2547 ( .A(n1872), .B(n1871), .Z(n1876) );
  NANDN U2548 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U2549 ( .A(n1876), .B(n1875), .Z(n2161) );
  OR U2550 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U2551 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2552 ( .A(n1882), .B(n1881), .Z(n2148) );
  OR U2553 ( .A(n1884), .B(n1883), .Z(n1888) );
  OR U2554 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U2555 ( .A(n1888), .B(n1887), .Z(n2147) );
  XOR U2556 ( .A(n2148), .B(n2147), .Z(n2150) );
  NANDN U2557 ( .A(n1890), .B(n1889), .Z(n1894) );
  NANDN U2558 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U2559 ( .A(n1894), .B(n1893), .Z(n2124) );
  OR U2560 ( .A(n1896), .B(n1895), .Z(n1900) );
  NAND U2561 ( .A(n1898), .B(n1897), .Z(n1899) );
  NAND U2562 ( .A(n1900), .B(n1899), .Z(n2123) );
  XOR U2563 ( .A(n2124), .B(n2123), .Z(n2125) );
  AND U2564 ( .A(y[645]), .B(x[148]), .Z(n2101) );
  AND U2565 ( .A(y[646]), .B(x[147]), .Z(n1902) );
  AND U2566 ( .A(y[644]), .B(x[149]), .Z(n1901) );
  XNOR U2567 ( .A(n1902), .B(n1901), .Z(n2102) );
  XOR U2568 ( .A(n2101), .B(n2102), .Z(n2108) );
  ANDN U2569 ( .B(x[150]), .A(n141), .Z(n2084) );
  ANDN U2570 ( .B(x[133]), .A(n2590), .Z(n2082) );
  ANDN U2571 ( .B(y[648]), .A(n168), .Z(n2083) );
  XNOR U2572 ( .A(n2082), .B(n2083), .Z(n2085) );
  XOR U2573 ( .A(n2084), .B(n2085), .Z(n2106) );
  OR U2574 ( .A(n1904), .B(n1903), .Z(n1908) );
  OR U2575 ( .A(n1906), .B(n1905), .Z(n1907) );
  AND U2576 ( .A(n1908), .B(n1907), .Z(n2105) );
  XNOR U2577 ( .A(n2106), .B(n2105), .Z(n2107) );
  XNOR U2578 ( .A(n2108), .B(n2107), .Z(n2046) );
  ANDN U2579 ( .B(x[151]), .A(n140), .Z(n2090) );
  ANDN U2580 ( .B(y[661]), .A(n155), .Z(n2088) );
  ANDN U2581 ( .B(y[649]), .A(n167), .Z(n2089) );
  XNOR U2582 ( .A(n2088), .B(n2089), .Z(n2091) );
  XNOR U2583 ( .A(n2090), .B(n2091), .Z(n2113) );
  ANDN U2584 ( .B(x[143]), .A(n2627), .Z(n2096) );
  ANDN U2585 ( .B(x[146]), .A(n143), .Z(n2094) );
  ANDN U2586 ( .B(y[659]), .A(n157), .Z(n2095) );
  XNOR U2587 ( .A(n2094), .B(n2095), .Z(n2097) );
  XOR U2588 ( .A(n2096), .B(n2097), .Z(n2112) );
  NAND U2589 ( .A(n2100), .B(n2101), .Z(n1912) );
  OR U2590 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2591 ( .A(n1912), .B(n1911), .Z(n2111) );
  XNOR U2592 ( .A(n2112), .B(n2111), .Z(n2114) );
  XOR U2593 ( .A(n2113), .B(n2114), .Z(n2045) );
  XNOR U2594 ( .A(n2046), .B(n2045), .Z(n2048) );
  OR U2595 ( .A(n1914), .B(n1913), .Z(n1918) );
  OR U2596 ( .A(n1916), .B(n1915), .Z(n1917) );
  AND U2597 ( .A(n1918), .B(n1917), .Z(n2047) );
  XOR U2598 ( .A(n2048), .B(n2047), .Z(n2051) );
  NANDN U2599 ( .A(n1920), .B(n1919), .Z(n1924) );
  OR U2600 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U2601 ( .A(n1924), .B(n1923), .Z(n2052) );
  NANDN U2602 ( .A(n1926), .B(n1925), .Z(n1930) );
  OR U2603 ( .A(n1928), .B(n1927), .Z(n1929) );
  AND U2604 ( .A(n1930), .B(n1929), .Z(n2053) );
  XOR U2605 ( .A(n2054), .B(n2053), .Z(n2126) );
  XNOR U2606 ( .A(n2125), .B(n2126), .Z(n2149) );
  NANDN U2607 ( .A(n1932), .B(n1931), .Z(n1936) );
  NANDN U2608 ( .A(n1934), .B(n1933), .Z(n1935) );
  AND U2609 ( .A(n1936), .B(n1935), .Z(n2141) );
  NANDN U2610 ( .A(n1938), .B(n1937), .Z(n1942) );
  OR U2611 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U2612 ( .A(n1942), .B(n1941), .Z(n2135) );
  NAND U2613 ( .A(x[130]), .B(y[663]), .Z(n2060) );
  NAND U2614 ( .A(x[131]), .B(y[662]), .Z(n2058) );
  XNOR U2615 ( .A(n2060), .B(n2059), .Z(n2118) );
  NANDN U2616 ( .A(n1944), .B(n1943), .Z(n1948) );
  NANDN U2617 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2618 ( .A(n1948), .B(n1947), .Z(n2117) );
  XOR U2619 ( .A(n2118), .B(n2117), .Z(n2119) );
  OR U2620 ( .A(n1950), .B(n1949), .Z(n1954) );
  OR U2621 ( .A(n1952), .B(n1951), .Z(n1953) );
  AND U2622 ( .A(n1954), .B(n1953), .Z(n2120) );
  NANDN U2623 ( .A(n1956), .B(n1955), .Z(n1960) );
  OR U2624 ( .A(n1958), .B(n1957), .Z(n1959) );
  AND U2625 ( .A(n1960), .B(n1959), .Z(n2129) );
  XNOR U2626 ( .A(n2130), .B(n2129), .Z(n2132) );
  OR U2627 ( .A(n1962), .B(n1961), .Z(n1966) );
  OR U2628 ( .A(n1964), .B(n1963), .Z(n1965) );
  NAND U2629 ( .A(n1966), .B(n1965), .Z(n2040) );
  NAND U2630 ( .A(n2447), .B(n1967), .Z(n1971) );
  OR U2631 ( .A(n1969), .B(n1968), .Z(n1970) );
  AND U2632 ( .A(n1971), .B(n1970), .Z(n2071) );
  NAND U2633 ( .A(x[129]), .B(y[664]), .Z(n2064) );
  AND U2634 ( .A(y[652]), .B(x[141]), .Z(n2063) );
  XNOR U2635 ( .A(n2064), .B(n2063), .Z(n2066) );
  NAND U2636 ( .A(x[152]), .B(y[641]), .Z(n2075) );
  XNOR U2637 ( .A(n2075), .B(o[25]), .Z(n2065) );
  XNOR U2638 ( .A(n2066), .B(n2065), .Z(n2070) );
  NAND U2639 ( .A(x[139]), .B(y[654]), .Z(n2078) );
  ANDN U2640 ( .B(y[653]), .A(n163), .Z(n2077) );
  NAND U2641 ( .A(y[658]), .B(x[135]), .Z(n2076) );
  XOR U2642 ( .A(n2077), .B(n2076), .Z(n2079) );
  XNOR U2643 ( .A(n2078), .B(n2079), .Z(n2069) );
  XNOR U2644 ( .A(n2070), .B(n2069), .Z(n2072) );
  XNOR U2645 ( .A(n2071), .B(n2072), .Z(n2039) );
  XNOR U2646 ( .A(n2040), .B(n2039), .Z(n2042) );
  NAND U2647 ( .A(n1973), .B(n1972), .Z(n1977) );
  NANDN U2648 ( .A(n1975), .B(n1974), .Z(n1976) );
  AND U2649 ( .A(n1977), .B(n1976), .Z(n2036) );
  OR U2650 ( .A(n1979), .B(n1978), .Z(n1983) );
  NANDN U2651 ( .A(n1981), .B(n1980), .Z(n1982) );
  AND U2652 ( .A(n1983), .B(n1982), .Z(n2034) );
  ANDN U2653 ( .B(y[657]), .A(n159), .Z(n2029) );
  XOR U2654 ( .A(n2028), .B(n2027), .Z(n2030) );
  XOR U2655 ( .A(n2029), .B(n2030), .Z(n2015) );
  ANDN U2656 ( .B(o[24]), .A(n1984), .Z(n2024) );
  IV U2657 ( .A(x[153]), .Z(n14372) );
  ANDN U2658 ( .B(y[640]), .A(n14372), .Z(n2022) );
  NAND U2659 ( .A(x[128]), .B(y[665]), .Z(n2021) );
  XOR U2660 ( .A(n2022), .B(n2021), .Z(n2023) );
  XOR U2661 ( .A(n2024), .B(n2023), .Z(n2016) );
  XNOR U2662 ( .A(n2015), .B(n2016), .Z(n2018) );
  OR U2663 ( .A(n1986), .B(n1985), .Z(n1990) );
  OR U2664 ( .A(n1988), .B(n1987), .Z(n1989) );
  AND U2665 ( .A(n1990), .B(n1989), .Z(n2017) );
  XOR U2666 ( .A(n2018), .B(n2017), .Z(n2033) );
  XNOR U2667 ( .A(n2034), .B(n2033), .Z(n2035) );
  XOR U2668 ( .A(n2036), .B(n2035), .Z(n2041) );
  XNOR U2669 ( .A(n2042), .B(n2041), .Z(n2131) );
  XOR U2670 ( .A(n2132), .B(n2131), .Z(n2136) );
  XOR U2671 ( .A(n2135), .B(n2136), .Z(n2137) );
  NANDN U2672 ( .A(n1992), .B(n1991), .Z(n1996) );
  OR U2673 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2674 ( .A(n1996), .B(n1995), .Z(n2138) );
  XNOR U2675 ( .A(n2137), .B(n2138), .Z(n2142) );
  XNOR U2676 ( .A(n2141), .B(n2142), .Z(n2144) );
  XOR U2677 ( .A(n2143), .B(n2144), .Z(n2159) );
  OR U2678 ( .A(n1998), .B(n1997), .Z(n2002) );
  OR U2679 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2680 ( .A(n2002), .B(n2001), .Z(n2160) );
  XOR U2681 ( .A(n2159), .B(n2160), .Z(n2162) );
  XOR U2682 ( .A(n2161), .B(n2162), .Z(n2155) );
  NANDN U2683 ( .A(n2004), .B(n2003), .Z(n2008) );
  NANDN U2684 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2685 ( .A(n2008), .B(n2007), .Z(n2153) );
  NANDN U2686 ( .A(n2010), .B(n2009), .Z(n2014) );
  OR U2687 ( .A(n2012), .B(n2011), .Z(n2013) );
  AND U2688 ( .A(n2014), .B(n2013), .Z(n2154) );
  XNOR U2689 ( .A(n2153), .B(n2154), .Z(n2156) );
  XNOR U2690 ( .A(n2155), .B(n2156), .Z(N58) );
  OR U2691 ( .A(n2016), .B(n2015), .Z(n2020) );
  OR U2692 ( .A(n2018), .B(n2017), .Z(n2019) );
  AND U2693 ( .A(n2020), .B(n2019), .Z(n2306) );
  NAND U2694 ( .A(x[130]), .B(y[664]), .Z(n2208) );
  AND U2695 ( .A(x[152]), .B(y[642]), .Z(n2209) );
  XNOR U2696 ( .A(n2210), .B(n2209), .Z(n2231) );
  NANDN U2697 ( .A(n2022), .B(n2021), .Z(n2026) );
  OR U2698 ( .A(n2024), .B(n2023), .Z(n2025) );
  NAND U2699 ( .A(n2026), .B(n2025), .Z(n2232) );
  NANDN U2700 ( .A(n2028), .B(n2027), .Z(n2032) );
  OR U2701 ( .A(n2030), .B(n2029), .Z(n2031) );
  NAND U2702 ( .A(n2032), .B(n2031), .Z(n2233) );
  XNOR U2703 ( .A(n2234), .B(n2233), .Z(n2307) );
  XNOR U2704 ( .A(n2306), .B(n2307), .Z(n2309) );
  NANDN U2705 ( .A(n2034), .B(n2033), .Z(n2038) );
  NANDN U2706 ( .A(n2036), .B(n2035), .Z(n2037) );
  AND U2707 ( .A(n2038), .B(n2037), .Z(n2308) );
  XOR U2708 ( .A(n2309), .B(n2308), .Z(n2272) );
  OR U2709 ( .A(n2040), .B(n2039), .Z(n2044) );
  OR U2710 ( .A(n2042), .B(n2041), .Z(n2043) );
  NAND U2711 ( .A(n2044), .B(n2043), .Z(n2270) );
  OR U2712 ( .A(n2046), .B(n2045), .Z(n2050) );
  OR U2713 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U2714 ( .A(n2050), .B(n2049), .Z(n2269) );
  XOR U2715 ( .A(n2270), .B(n2269), .Z(n2271) );
  NANDN U2716 ( .A(n2052), .B(n2051), .Z(n2056) );
  OR U2717 ( .A(n2054), .B(n2053), .Z(n2055) );
  AND U2718 ( .A(n2056), .B(n2055), .Z(n2265) );
  NANDN U2719 ( .A(n2058), .B(n2057), .Z(n2062) );
  OR U2720 ( .A(n2060), .B(n2059), .Z(n2061) );
  NAND U2721 ( .A(n2062), .B(n2061), .Z(n2220) );
  NANDN U2722 ( .A(n2064), .B(n2063), .Z(n2068) );
  NAND U2723 ( .A(n2066), .B(n2065), .Z(n2067) );
  NAND U2724 ( .A(n2068), .B(n2067), .Z(n2219) );
  XOR U2725 ( .A(n2220), .B(n2219), .Z(n2221) );
  ANDN U2726 ( .B(y[657]), .A(n160), .Z(n2302) );
  ANDN U2727 ( .B(x[134]), .A(n2590), .Z(n2300) );
  ANDN U2728 ( .B(x[136]), .A(n2616), .Z(n2301) );
  XNOR U2729 ( .A(n2300), .B(n2301), .Z(n2303) );
  XNOR U2730 ( .A(n2302), .B(n2303), .Z(n2278) );
  ANDN U2731 ( .B(y[659]), .A(n158), .Z(n2275) );
  ANDN U2732 ( .B(y[656]), .A(n161), .Z(n2241) );
  ANDN U2733 ( .B(x[140]), .A(n2238), .Z(n2239) );
  ANDN U2734 ( .B(y[661]), .A(n156), .Z(n2240) );
  XNOR U2735 ( .A(n2239), .B(n2240), .Z(n2242) );
  XNOR U2736 ( .A(n2241), .B(n2242), .Z(n2276) );
  XNOR U2737 ( .A(n2275), .B(n2276), .Z(n2277) );
  XNOR U2738 ( .A(n2278), .B(n2277), .Z(n2222) );
  OR U2739 ( .A(n2070), .B(n2069), .Z(n2074) );
  OR U2740 ( .A(n2072), .B(n2071), .Z(n2073) );
  AND U2741 ( .A(n2074), .B(n2073), .Z(n2258) );
  XNOR U2742 ( .A(n2257), .B(n2258), .Z(n2260) );
  ANDN U2743 ( .B(o[25]), .A(n2075), .Z(n2289) );
  ANDN U2744 ( .B(x[142]), .A(n2617), .Z(n2287) );
  ANDN U2745 ( .B(y[665]), .A(n152), .Z(n2288) );
  XNOR U2746 ( .A(n2287), .B(n2288), .Z(n2290) );
  XOR U2747 ( .A(n2289), .B(n2290), .Z(n2254) );
  NAND U2748 ( .A(y[666]), .B(x[128]), .Z(n2246) );
  AND U2749 ( .A(x[154]), .B(y[640]), .Z(n2245) );
  XNOR U2750 ( .A(n2246), .B(n2245), .Z(n2248) );
  NAND U2751 ( .A(x[153]), .B(y[641]), .Z(n2299) );
  XNOR U2752 ( .A(n2299), .B(o[26]), .Z(n2247) );
  XNOR U2753 ( .A(n2248), .B(n2247), .Z(n2252) );
  NANDN U2754 ( .A(n2077), .B(n2076), .Z(n2081) );
  NANDN U2755 ( .A(n2079), .B(n2078), .Z(n2080) );
  NAND U2756 ( .A(n2081), .B(n2080), .Z(n2251) );
  XOR U2757 ( .A(n2252), .B(n2251), .Z(n2253) );
  OR U2758 ( .A(n2083), .B(n2082), .Z(n2087) );
  OR U2759 ( .A(n2085), .B(n2084), .Z(n2086) );
  AND U2760 ( .A(n2087), .B(n2086), .Z(n2189) );
  OR U2761 ( .A(n2089), .B(n2088), .Z(n2093) );
  OR U2762 ( .A(n2091), .B(n2090), .Z(n2092) );
  AND U2763 ( .A(n2093), .B(n2092), .Z(n2190) );
  XOR U2764 ( .A(n2189), .B(n2190), .Z(n2191) );
  XOR U2765 ( .A(n2192), .B(n2191), .Z(n2227) );
  ANDN U2766 ( .B(y[662]), .A(n155), .Z(n2214) );
  XNOR U2767 ( .A(n2213), .B(n2214), .Z(n2216) );
  XOR U2768 ( .A(n2215), .B(n2216), .Z(n2195) );
  OR U2769 ( .A(n2095), .B(n2094), .Z(n2099) );
  OR U2770 ( .A(n2097), .B(n2096), .Z(n2098) );
  NAND U2771 ( .A(n2099), .B(n2098), .Z(n2196) );
  XNOR U2772 ( .A(n2195), .B(n2196), .Z(n2198) );
  NAND U2773 ( .A(y[647]), .B(x[147]), .Z(n2282) );
  AND U2774 ( .A(y[655]), .B(x[139]), .Z(n2281) );
  XNOR U2775 ( .A(n2282), .B(n2281), .Z(n2283) );
  NAND U2776 ( .A(x[131]), .B(y[663]), .Z(n2284) );
  XOR U2777 ( .A(n2198), .B(n2197), .Z(n2226) );
  ANDN U2778 ( .B(y[646]), .A(n172), .Z(n2384) );
  NAND U2779 ( .A(n2100), .B(n2384), .Z(n2104) );
  NANDN U2780 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U2781 ( .A(n2104), .B(n2103), .Z(n2184) );
  NAND U2782 ( .A(x[150]), .B(y[644]), .Z(n2204) );
  NAND U2783 ( .A(x[151]), .B(y[643]), .Z(n2201) );
  XNOR U2784 ( .A(n2202), .B(n2201), .Z(n2203) );
  XNOR U2785 ( .A(n2204), .B(n2203), .Z(n2183) );
  XNOR U2786 ( .A(n2184), .B(n2183), .Z(n2186) );
  ANDN U2787 ( .B(y[646]), .A(n171), .Z(n2295) );
  ANDN U2788 ( .B(y[645]), .A(n172), .Z(n2294) );
  XNOR U2789 ( .A(n2293), .B(n2294), .Z(n2296) );
  XNOR U2790 ( .A(n2295), .B(n2296), .Z(n2185) );
  XOR U2791 ( .A(n2186), .B(n2185), .Z(n2225) );
  XNOR U2792 ( .A(n2226), .B(n2225), .Z(n2228) );
  XNOR U2793 ( .A(n2227), .B(n2228), .Z(n2259) );
  XOR U2794 ( .A(n2260), .B(n2259), .Z(n2264) );
  OR U2795 ( .A(n2106), .B(n2105), .Z(n2110) );
  OR U2796 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U2797 ( .A(n2110), .B(n2109), .Z(n2312) );
  OR U2798 ( .A(n2112), .B(n2111), .Z(n2116) );
  NANDN U2799 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U2800 ( .A(n2116), .B(n2115), .Z(n2313) );
  XOR U2801 ( .A(n2312), .B(n2313), .Z(n2314) );
  OR U2802 ( .A(n2118), .B(n2117), .Z(n2122) );
  NANDN U2803 ( .A(n2120), .B(n2119), .Z(n2121) );
  AND U2804 ( .A(n2122), .B(n2121), .Z(n2315) );
  XOR U2805 ( .A(n2264), .B(n2263), .Z(n2266) );
  XOR U2806 ( .A(n2265), .B(n2266), .Z(n2177) );
  XOR U2807 ( .A(n2178), .B(n2177), .Z(n2180) );
  OR U2808 ( .A(n2124), .B(n2123), .Z(n2128) );
  NANDN U2809 ( .A(n2126), .B(n2125), .Z(n2127) );
  NAND U2810 ( .A(n2128), .B(n2127), .Z(n2179) );
  XOR U2811 ( .A(n2180), .B(n2179), .Z(n2321) );
  OR U2812 ( .A(n2130), .B(n2129), .Z(n2134) );
  OR U2813 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U2814 ( .A(n2134), .B(n2133), .Z(n2319) );
  OR U2815 ( .A(n2136), .B(n2135), .Z(n2140) );
  NANDN U2816 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U2817 ( .A(n2140), .B(n2139), .Z(n2318) );
  XOR U2818 ( .A(n2319), .B(n2318), .Z(n2320) );
  XOR U2819 ( .A(n2321), .B(n2320), .Z(n2172) );
  OR U2820 ( .A(n2142), .B(n2141), .Z(n2146) );
  NANDN U2821 ( .A(n2144), .B(n2143), .Z(n2145) );
  NAND U2822 ( .A(n2146), .B(n2145), .Z(n2171) );
  XNOR U2823 ( .A(n2172), .B(n2171), .Z(n2173) );
  OR U2824 ( .A(n2148), .B(n2147), .Z(n2152) );
  NAND U2825 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U2826 ( .A(n2152), .B(n2151), .Z(n2174) );
  XOR U2827 ( .A(n2173), .B(n2174), .Z(n2167) );
  NANDN U2828 ( .A(n2154), .B(n2153), .Z(n2158) );
  NAND U2829 ( .A(n2156), .B(n2155), .Z(n2157) );
  NAND U2830 ( .A(n2158), .B(n2157), .Z(n2165) );
  NANDN U2831 ( .A(n2160), .B(n2159), .Z(n2164) );
  OR U2832 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U2833 ( .A(n2164), .B(n2163), .Z(n2166) );
  XNOR U2834 ( .A(n2165), .B(n2166), .Z(n2168) );
  XNOR U2835 ( .A(n2167), .B(n2168), .Z(N59) );
  NANDN U2836 ( .A(n2166), .B(n2165), .Z(n2170) );
  NAND U2837 ( .A(n2168), .B(n2167), .Z(n2169) );
  NAND U2838 ( .A(n2170), .B(n2169), .Z(n2324) );
  OR U2839 ( .A(n2172), .B(n2171), .Z(n2176) );
  OR U2840 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U2841 ( .A(n2176), .B(n2175), .Z(n2325) );
  XNOR U2842 ( .A(n2324), .B(n2325), .Z(n2326) );
  NANDN U2843 ( .A(n2178), .B(n2177), .Z(n2182) );
  OR U2844 ( .A(n2180), .B(n2179), .Z(n2181) );
  NAND U2845 ( .A(n2182), .B(n2181), .Z(n2331) );
  OR U2846 ( .A(n2184), .B(n2183), .Z(n2188) );
  OR U2847 ( .A(n2186), .B(n2185), .Z(n2187) );
  NAND U2848 ( .A(n2188), .B(n2187), .Z(n2349) );
  OR U2849 ( .A(n2190), .B(n2189), .Z(n2194) );
  NANDN U2850 ( .A(n2192), .B(n2191), .Z(n2193) );
  AND U2851 ( .A(n2194), .B(n2193), .Z(n2362) );
  OR U2852 ( .A(n2196), .B(n2195), .Z(n2200) );
  NANDN U2853 ( .A(n2198), .B(n2197), .Z(n2199) );
  NAND U2854 ( .A(n2200), .B(n2199), .Z(n2361) );
  NANDN U2855 ( .A(n2202), .B(n2201), .Z(n2206) );
  NAND U2856 ( .A(n2204), .B(n2203), .Z(n2205) );
  AND U2857 ( .A(n2206), .B(n2205), .Z(n2433) );
  NANDN U2858 ( .A(n2208), .B(n2207), .Z(n2212) );
  NANDN U2859 ( .A(n2210), .B(n2209), .Z(n2211) );
  NAND U2860 ( .A(n2212), .B(n2211), .Z(n2434) );
  XOR U2861 ( .A(n2433), .B(n2434), .Z(n2435) );
  OR U2862 ( .A(n2214), .B(n2213), .Z(n2218) );
  OR U2863 ( .A(n2216), .B(n2215), .Z(n2217) );
  AND U2864 ( .A(n2218), .B(n2217), .Z(n2427) );
  ANDN U2865 ( .B(y[658]), .A(n160), .Z(n2386) );
  ANDN U2866 ( .B(y[649]), .A(n169), .Z(n2385) );
  XNOR U2867 ( .A(n2384), .B(n2385), .Z(n2387) );
  XNOR U2868 ( .A(n2386), .B(n2387), .Z(n2428) );
  XOR U2869 ( .A(n2427), .B(n2428), .Z(n2429) );
  NAND U2870 ( .A(x[128]), .B(y[667]), .Z(n2375) );
  ANDN U2871 ( .B(y[641]), .A(n176), .Z(n2390) );
  XOR U2872 ( .A(o[27]), .B(n2390), .Z(n2373) );
  NAND U2873 ( .A(y[640]), .B(x[155]), .Z(n2372) );
  XNOR U2874 ( .A(n2373), .B(n2372), .Z(n2374) );
  XNOR U2875 ( .A(n2375), .B(n2374), .Z(n2430) );
  XOR U2876 ( .A(n2429), .B(n2430), .Z(n2436) );
  XOR U2877 ( .A(n2361), .B(n2360), .Z(n2363) );
  XOR U2878 ( .A(n2362), .B(n2363), .Z(n2348) );
  XNOR U2879 ( .A(n2349), .B(n2348), .Z(n2351) );
  OR U2880 ( .A(n2220), .B(n2219), .Z(n2224) );
  NANDN U2881 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U2882 ( .A(n2224), .B(n2223), .Z(n2350) );
  XOR U2883 ( .A(n2351), .B(n2350), .Z(n2483) );
  OR U2884 ( .A(n2226), .B(n2225), .Z(n2230) );
  NANDN U2885 ( .A(n2228), .B(n2227), .Z(n2229) );
  AND U2886 ( .A(n2230), .B(n2229), .Z(n2343) );
  NANDN U2887 ( .A(n2232), .B(n2231), .Z(n2236) );
  OR U2888 ( .A(n2234), .B(n2233), .Z(n2235) );
  AND U2889 ( .A(n2236), .B(n2235), .Z(n2368) );
  ANDN U2890 ( .B(x[140]), .A(n2237), .Z(n2464) );
  ANDN U2891 ( .B(x[141]), .A(n2238), .Z(n2465) );
  XNOR U2892 ( .A(n2464), .B(n2465), .Z(n2467) );
  NAND U2893 ( .A(y[651]), .B(x[144]), .Z(n2445) );
  XOR U2894 ( .A(n2446), .B(n2445), .Z(n2448) );
  XNOR U2895 ( .A(n2467), .B(n2466), .Z(n2411) );
  ANDN U2896 ( .B(y[664]), .A(n154), .Z(n2472) );
  ANDN U2897 ( .B(y[665]), .A(n153), .Z(n2470) );
  ANDN U2898 ( .B(x[143]), .A(n2617), .Z(n2471) );
  XNOR U2899 ( .A(n2470), .B(n2471), .Z(n2473) );
  XOR U2900 ( .A(n2472), .B(n2473), .Z(n2409) );
  NAND U2901 ( .A(x[134]), .B(y[661]), .Z(n2393) );
  ANDN U2902 ( .B(y[642]), .A(n14372), .Z(n2392) );
  NAND U2903 ( .A(x[147]), .B(y[648]), .Z(n2391) );
  XOR U2904 ( .A(n2392), .B(n2391), .Z(n2394) );
  XNOR U2905 ( .A(n2393), .B(n2394), .Z(n2410) );
  XNOR U2906 ( .A(n2409), .B(n2410), .Z(n2412) );
  XNOR U2907 ( .A(n2411), .B(n2412), .Z(n2441) );
  OR U2908 ( .A(n2240), .B(n2239), .Z(n2244) );
  OR U2909 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2910 ( .A(n2244), .B(n2243), .Z(n2439) );
  NANDN U2911 ( .A(n2246), .B(n2245), .Z(n2250) );
  NAND U2912 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U2913 ( .A(n2250), .B(n2249), .Z(n2440) );
  XNOR U2914 ( .A(n2439), .B(n2440), .Z(n2442) );
  XOR U2915 ( .A(n2441), .B(n2442), .Z(n2366) );
  OR U2916 ( .A(n2252), .B(n2251), .Z(n2256) );
  NANDN U2917 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2918 ( .A(n2256), .B(n2255), .Z(n2367) );
  XOR U2919 ( .A(n2366), .B(n2367), .Z(n2369) );
  XOR U2920 ( .A(n2368), .B(n2369), .Z(n2342) );
  OR U2921 ( .A(n2258), .B(n2257), .Z(n2262) );
  NANDN U2922 ( .A(n2260), .B(n2259), .Z(n2261) );
  AND U2923 ( .A(n2262), .B(n2261), .Z(n2344) );
  XOR U2924 ( .A(n2345), .B(n2344), .Z(n2482) );
  XNOR U2925 ( .A(n2483), .B(n2482), .Z(n2485) );
  NANDN U2926 ( .A(n2264), .B(n2263), .Z(n2268) );
  OR U2927 ( .A(n2266), .B(n2265), .Z(n2267) );
  AND U2928 ( .A(n2268), .B(n2267), .Z(n2484) );
  XNOR U2929 ( .A(n2485), .B(n2484), .Z(n2478) );
  OR U2930 ( .A(n2270), .B(n2269), .Z(n2274) );
  NANDN U2931 ( .A(n2272), .B(n2271), .Z(n2273) );
  AND U2932 ( .A(n2274), .B(n2273), .Z(n2476) );
  OR U2933 ( .A(n2276), .B(n2275), .Z(n2280) );
  OR U2934 ( .A(n2278), .B(n2277), .Z(n2279) );
  AND U2935 ( .A(n2280), .B(n2279), .Z(n2338) );
  NANDN U2936 ( .A(n2282), .B(n2281), .Z(n2286) );
  NANDN U2937 ( .A(n2284), .B(n2283), .Z(n2285) );
  AND U2938 ( .A(n2286), .B(n2285), .Z(n2417) );
  ANDN U2939 ( .B(x[150]), .A(n142), .Z(n2453) );
  ANDN U2940 ( .B(x[151]), .A(n2634), .Z(n2451) );
  ANDN U2941 ( .B(y[659]), .A(n159), .Z(n2452) );
  XNOR U2942 ( .A(n2451), .B(n2452), .Z(n2454) );
  XOR U2943 ( .A(n2453), .B(n2454), .Z(n2415) );
  NAND U2944 ( .A(y[660]), .B(x[135]), .Z(n2399) );
  NAND U2945 ( .A(y[643]), .B(x[152]), .Z(n2397) );
  XOR U2946 ( .A(n2398), .B(n2397), .Z(n2400) );
  XNOR U2947 ( .A(n2399), .B(n2400), .Z(n2416) );
  XNOR U2948 ( .A(n2415), .B(n2416), .Z(n2418) );
  XOR U2949 ( .A(n2417), .B(n2418), .Z(n2336) );
  OR U2950 ( .A(n2288), .B(n2287), .Z(n2292) );
  OR U2951 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U2952 ( .A(n2292), .B(n2291), .Z(n2404) );
  OR U2953 ( .A(n2294), .B(n2293), .Z(n2298) );
  OR U2954 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2955 ( .A(n2298), .B(n2297), .Z(n2403) );
  XOR U2956 ( .A(n2404), .B(n2403), .Z(n2406) );
  ANDN U2957 ( .B(y[653]), .A(n165), .Z(n2460) );
  ANDN U2958 ( .B(o[26]), .A(n2299), .Z(n2458) );
  IV U2959 ( .A(y[666]), .Z(n2615) );
  ANDN U2960 ( .B(x[129]), .A(n2615), .Z(n2459) );
  XNOR U2961 ( .A(n2458), .B(n2459), .Z(n2461) );
  XOR U2962 ( .A(n2460), .B(n2461), .Z(n2421) );
  NAND U2963 ( .A(x[145]), .B(y[650]), .Z(n2379) );
  AND U2964 ( .A(y[663]), .B(x[132]), .Z(n2378) );
  XOR U2965 ( .A(n2379), .B(n2378), .Z(n2381) );
  AND U2966 ( .A(y[662]), .B(x[133]), .Z(n2380) );
  XOR U2967 ( .A(n2381), .B(n2380), .Z(n2422) );
  XNOR U2968 ( .A(n2421), .B(n2422), .Z(n2424) );
  OR U2969 ( .A(n2301), .B(n2300), .Z(n2305) );
  OR U2970 ( .A(n2303), .B(n2302), .Z(n2304) );
  NAND U2971 ( .A(n2305), .B(n2304), .Z(n2423) );
  XOR U2972 ( .A(n2424), .B(n2423), .Z(n2405) );
  XOR U2973 ( .A(n2406), .B(n2405), .Z(n2337) );
  XNOR U2974 ( .A(n2336), .B(n2337), .Z(n2339) );
  XOR U2975 ( .A(n2338), .B(n2339), .Z(n2354) );
  OR U2976 ( .A(n2307), .B(n2306), .Z(n2311) );
  OR U2977 ( .A(n2309), .B(n2308), .Z(n2310) );
  AND U2978 ( .A(n2311), .B(n2310), .Z(n2355) );
  XNOR U2979 ( .A(n2354), .B(n2355), .Z(n2357) );
  OR U2980 ( .A(n2313), .B(n2312), .Z(n2317) );
  NANDN U2981 ( .A(n2315), .B(n2314), .Z(n2316) );
  AND U2982 ( .A(n2317), .B(n2316), .Z(n2356) );
  XOR U2983 ( .A(n2357), .B(n2356), .Z(n2477) );
  XNOR U2984 ( .A(n2476), .B(n2477), .Z(n2479) );
  XOR U2985 ( .A(n2478), .B(n2479), .Z(n2330) );
  XNOR U2986 ( .A(n2331), .B(n2330), .Z(n2333) );
  OR U2987 ( .A(n2319), .B(n2318), .Z(n2323) );
  NANDN U2988 ( .A(n2321), .B(n2320), .Z(n2322) );
  AND U2989 ( .A(n2323), .B(n2322), .Z(n2332) );
  XOR U2990 ( .A(n2333), .B(n2332), .Z(n2327) );
  XNOR U2991 ( .A(n2326), .B(n2327), .Z(N60) );
  NANDN U2992 ( .A(n2325), .B(n2324), .Z(n2329) );
  NAND U2993 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U2994 ( .A(n2329), .B(n2328), .Z(n2488) );
  OR U2995 ( .A(n2331), .B(n2330), .Z(n2335) );
  OR U2996 ( .A(n2333), .B(n2332), .Z(n2334) );
  AND U2997 ( .A(n2335), .B(n2334), .Z(n2489) );
  XNOR U2998 ( .A(n2488), .B(n2489), .Z(n2490) );
  OR U2999 ( .A(n2337), .B(n2336), .Z(n2341) );
  OR U3000 ( .A(n2339), .B(n2338), .Z(n2340) );
  AND U3001 ( .A(n2341), .B(n2340), .Z(n2656) );
  NANDN U3002 ( .A(n2343), .B(n2342), .Z(n2347) );
  OR U3003 ( .A(n2345), .B(n2344), .Z(n2346) );
  NAND U3004 ( .A(n2347), .B(n2346), .Z(n2654) );
  OR U3005 ( .A(n2349), .B(n2348), .Z(n2353) );
  OR U3006 ( .A(n2351), .B(n2350), .Z(n2352) );
  NAND U3007 ( .A(n2353), .B(n2352), .Z(n2653) );
  XOR U3008 ( .A(n2654), .B(n2653), .Z(n2655) );
  XNOR U3009 ( .A(n2656), .B(n2655), .Z(n2662) );
  OR U3010 ( .A(n2355), .B(n2354), .Z(n2359) );
  OR U3011 ( .A(n2357), .B(n2356), .Z(n2358) );
  AND U3012 ( .A(n2359), .B(n2358), .Z(n2659) );
  NANDN U3013 ( .A(n2361), .B(n2360), .Z(n2365) );
  OR U3014 ( .A(n2363), .B(n2362), .Z(n2364) );
  AND U3015 ( .A(n2365), .B(n2364), .Z(n2641) );
  NANDN U3016 ( .A(n2367), .B(n2366), .Z(n2371) );
  OR U3017 ( .A(n2369), .B(n2368), .Z(n2370) );
  NAND U3018 ( .A(n2371), .B(n2370), .Z(n2642) );
  XOR U3019 ( .A(n2641), .B(n2642), .Z(n2643) );
  NANDN U3020 ( .A(n2373), .B(n2372), .Z(n2377) );
  NAND U3021 ( .A(n2375), .B(n2374), .Z(n2376) );
  AND U3022 ( .A(n2377), .B(n2376), .Z(n2518) );
  NANDN U3023 ( .A(n2379), .B(n2378), .Z(n2383) );
  NANDN U3024 ( .A(n2381), .B(n2380), .Z(n2382) );
  NAND U3025 ( .A(n2383), .B(n2382), .Z(n2519) );
  XOR U3026 ( .A(n2518), .B(n2519), .Z(n2521) );
  OR U3027 ( .A(n2385), .B(n2384), .Z(n2389) );
  OR U3028 ( .A(n2387), .B(n2386), .Z(n2388) );
  AND U3029 ( .A(n2389), .B(n2388), .Z(n2542) );
  ANDN U3030 ( .B(x[138]), .A(n2616), .Z(n2562) );
  ANDN U3031 ( .B(y[659]), .A(n160), .Z(n2560) );
  ANDN U3032 ( .B(x[136]), .A(n2590), .Z(n2561) );
  XNOR U3033 ( .A(n2560), .B(n2561), .Z(n2563) );
  XNOR U3034 ( .A(n2562), .B(n2563), .Z(n2543) );
  XOR U3035 ( .A(n2542), .B(n2543), .Z(n2544) );
  ANDN U3036 ( .B(y[668]), .A(n151), .Z(n2550) );
  AND U3037 ( .A(n2390), .B(o[27]), .Z(n2548) );
  ANDN U3038 ( .B(x[156]), .A(n138), .Z(n2549) );
  XNOR U3039 ( .A(n2548), .B(n2549), .Z(n2551) );
  XNOR U3040 ( .A(n2550), .B(n2551), .Z(n2545) );
  XNOR U3041 ( .A(n2521), .B(n2520), .Z(n2503) );
  ANDN U3042 ( .B(y[645]), .A(n174), .Z(n2578) );
  ANDN U3043 ( .B(y[665]), .A(n154), .Z(n2579) );
  XNOR U3044 ( .A(n2578), .B(n2579), .Z(n2581) );
  XNOR U3045 ( .A(n2580), .B(n2581), .Z(n2526) );
  ANDN U3046 ( .B(y[663]), .A(n156), .Z(n2621) );
  ANDN U3047 ( .B(y[648]), .A(n171), .Z(n2619) );
  ANDN U3048 ( .B(x[149]), .A(n143), .Z(n2620) );
  XNOR U3049 ( .A(n2619), .B(n2620), .Z(n2622) );
  XOR U3050 ( .A(n2621), .B(n2622), .Z(n2524) );
  NANDN U3051 ( .A(n2392), .B(n2391), .Z(n2396) );
  NANDN U3052 ( .A(n2394), .B(n2393), .Z(n2395) );
  NAND U3053 ( .A(n2396), .B(n2395), .Z(n2525) );
  XNOR U3054 ( .A(n2524), .B(n2525), .Z(n2527) );
  XNOR U3055 ( .A(n2526), .B(n2527), .Z(n2501) );
  ANDN U3056 ( .B(y[667]), .A(n152), .Z(n2597) );
  ANDN U3057 ( .B(x[153]), .A(n141), .Z(n2598) );
  XNOR U3058 ( .A(n2597), .B(n2598), .Z(n2600) );
  XOR U3059 ( .A(n2599), .B(n2600), .Z(n2514) );
  ANDN U3060 ( .B(y[652]), .A(n167), .Z(n2605) );
  ANDN U3061 ( .B(y[666]), .A(n153), .Z(n2603) );
  ANDN U3062 ( .B(y[644]), .A(n175), .Z(n2604) );
  XNOR U3063 ( .A(n2603), .B(n2604), .Z(n2606) );
  XOR U3064 ( .A(n2605), .B(n2606), .Z(n2512) );
  NANDN U3065 ( .A(n2398), .B(n2397), .Z(n2402) );
  NANDN U3066 ( .A(n2400), .B(n2399), .Z(n2401) );
  NAND U3067 ( .A(n2402), .B(n2401), .Z(n2513) );
  XNOR U3068 ( .A(n2512), .B(n2513), .Z(n2515) );
  XNOR U3069 ( .A(n2514), .B(n2515), .Z(n2500) );
  XOR U3070 ( .A(n2501), .B(n2500), .Z(n2502) );
  XNOR U3071 ( .A(n2503), .B(n2502), .Z(n2648) );
  OR U3072 ( .A(n2404), .B(n2403), .Z(n2408) );
  NAND U3073 ( .A(n2406), .B(n2405), .Z(n2407) );
  NAND U3074 ( .A(n2408), .B(n2407), .Z(n2539) );
  OR U3075 ( .A(n2410), .B(n2409), .Z(n2414) );
  OR U3076 ( .A(n2412), .B(n2411), .Z(n2413) );
  NAND U3077 ( .A(n2414), .B(n2413), .Z(n2537) );
  OR U3078 ( .A(n2416), .B(n2415), .Z(n2420) );
  OR U3079 ( .A(n2418), .B(n2417), .Z(n2419) );
  NAND U3080 ( .A(n2420), .B(n2419), .Z(n2536) );
  XOR U3081 ( .A(n2537), .B(n2536), .Z(n2538) );
  XOR U3082 ( .A(n2648), .B(n2647), .Z(n2650) );
  OR U3083 ( .A(n2422), .B(n2421), .Z(n2426) );
  OR U3084 ( .A(n2424), .B(n2423), .Z(n2425) );
  AND U3085 ( .A(n2426), .B(n2425), .Z(n2506) );
  OR U3086 ( .A(n2428), .B(n2427), .Z(n2432) );
  NANDN U3087 ( .A(n2430), .B(n2429), .Z(n2431) );
  NAND U3088 ( .A(n2432), .B(n2431), .Z(n2507) );
  XOR U3089 ( .A(n2506), .B(n2507), .Z(n2508) );
  OR U3090 ( .A(n2434), .B(n2433), .Z(n2438) );
  NANDN U3091 ( .A(n2436), .B(n2435), .Z(n2437) );
  NAND U3092 ( .A(n2438), .B(n2437), .Z(n2509) );
  OR U3093 ( .A(n2440), .B(n2439), .Z(n2444) );
  NANDN U3094 ( .A(n2442), .B(n2441), .Z(n2443) );
  AND U3095 ( .A(n2444), .B(n2443), .Z(n2636) );
  ANDN U3096 ( .B(y[661]), .A(n158), .Z(n2611) );
  ANDN U3097 ( .B(y[657]), .A(n162), .Z(n2609) );
  ANDN U3098 ( .B(y[656]), .A(n163), .Z(n2610) );
  XNOR U3099 ( .A(n2609), .B(n2610), .Z(n2612) );
  XOR U3100 ( .A(n2611), .B(n2612), .Z(n2591) );
  NANDN U3101 ( .A(n2446), .B(n2445), .Z(n2450) );
  OR U3102 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U3103 ( .A(n2450), .B(n2449), .Z(n2592) );
  XNOR U3104 ( .A(n2591), .B(n2592), .Z(n2594) );
  NAND U3105 ( .A(x[143]), .B(y[653]), .Z(n2585) );
  AND U3106 ( .A(x[154]), .B(y[642]), .Z(n2584) );
  XNOR U3107 ( .A(n2585), .B(n2584), .Z(n2586) );
  AND U3108 ( .A(y[641]), .B(x[155]), .Z(n2770) );
  XNOR U3109 ( .A(o[28]), .B(n2770), .Z(n2587) );
  XOR U3110 ( .A(n2594), .B(n2593), .Z(n2530) );
  OR U3111 ( .A(n2452), .B(n2451), .Z(n2456) );
  OR U3112 ( .A(n2454), .B(n2453), .Z(n2455) );
  AND U3113 ( .A(n2456), .B(n2455), .Z(n2572) );
  ANDN U3114 ( .B(y[662]), .A(n157), .Z(n2630) );
  ANDN U3115 ( .B(x[147]), .A(n2457), .Z(n2629) );
  XNOR U3116 ( .A(n2628), .B(n2629), .Z(n2631) );
  XNOR U3117 ( .A(n2630), .B(n2631), .Z(n2573) );
  XOR U3118 ( .A(n2572), .B(n2573), .Z(n2575) );
  NAND U3119 ( .A(y[651]), .B(x[145]), .Z(n2556) );
  ANDN U3120 ( .B(y[664]), .A(n155), .Z(n2555) );
  NAND U3121 ( .A(x[150]), .B(y[646]), .Z(n2554) );
  XOR U3122 ( .A(n2555), .B(n2554), .Z(n2557) );
  XNOR U3123 ( .A(n2556), .B(n2557), .Z(n2574) );
  XNOR U3124 ( .A(n2575), .B(n2574), .Z(n2531) );
  XNOR U3125 ( .A(n2530), .B(n2531), .Z(n2533) );
  OR U3126 ( .A(n2459), .B(n2458), .Z(n2463) );
  OR U3127 ( .A(n2461), .B(n2460), .Z(n2462) );
  AND U3128 ( .A(n2463), .B(n2462), .Z(n2569) );
  OR U3129 ( .A(n2465), .B(n2464), .Z(n2469) );
  NANDN U3130 ( .A(n2467), .B(n2466), .Z(n2468) );
  AND U3131 ( .A(n2469), .B(n2468), .Z(n2566) );
  OR U3132 ( .A(n2471), .B(n2470), .Z(n2475) );
  OR U3133 ( .A(n2473), .B(n2472), .Z(n2474) );
  AND U3134 ( .A(n2475), .B(n2474), .Z(n2567) );
  XOR U3135 ( .A(n2566), .B(n2567), .Z(n2568) );
  XOR U3136 ( .A(n2533), .B(n2532), .Z(n2635) );
  XOR U3137 ( .A(n2636), .B(n2635), .Z(n2638) );
  XOR U3138 ( .A(n2637), .B(n2638), .Z(n2649) );
  XNOR U3139 ( .A(n2650), .B(n2649), .Z(n2644) );
  XNOR U3140 ( .A(n2643), .B(n2644), .Z(n2660) );
  XOR U3141 ( .A(n2659), .B(n2660), .Z(n2661) );
  OR U3142 ( .A(n2477), .B(n2476), .Z(n2481) );
  NANDN U3143 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U3144 ( .A(n2481), .B(n2480), .Z(n2495) );
  XNOR U3145 ( .A(n2494), .B(n2495), .Z(n2497) );
  NAND U3146 ( .A(n2483), .B(n2482), .Z(n2487) );
  OR U3147 ( .A(n2485), .B(n2484), .Z(n2486) );
  NAND U3148 ( .A(n2487), .B(n2486), .Z(n2496) );
  XOR U3149 ( .A(n2497), .B(n2496), .Z(n2491) );
  XNOR U3150 ( .A(n2490), .B(n2491), .Z(N61) );
  NANDN U3151 ( .A(n2489), .B(n2488), .Z(n2493) );
  NAND U3152 ( .A(n2491), .B(n2490), .Z(n2492) );
  NAND U3153 ( .A(n2493), .B(n2492), .Z(n2665) );
  OR U3154 ( .A(n2495), .B(n2494), .Z(n2499) );
  OR U3155 ( .A(n2497), .B(n2496), .Z(n2498) );
  AND U3156 ( .A(n2499), .B(n2498), .Z(n2666) );
  XNOR U3157 ( .A(n2665), .B(n2666), .Z(n2667) );
  NANDN U3158 ( .A(n2501), .B(n2500), .Z(n2505) );
  OR U3159 ( .A(n2503), .B(n2502), .Z(n2504) );
  AND U3160 ( .A(n2505), .B(n2504), .Z(n2685) );
  OR U3161 ( .A(n2507), .B(n2506), .Z(n2511) );
  NANDN U3162 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U3163 ( .A(n2511), .B(n2510), .Z(n2679) );
  OR U3164 ( .A(n2513), .B(n2512), .Z(n2517) );
  OR U3165 ( .A(n2515), .B(n2514), .Z(n2516) );
  NAND U3166 ( .A(n2517), .B(n2516), .Z(n2826) );
  OR U3167 ( .A(n2519), .B(n2518), .Z(n2523) );
  NAND U3168 ( .A(n2521), .B(n2520), .Z(n2522) );
  AND U3169 ( .A(n2523), .B(n2522), .Z(n2823) );
  OR U3170 ( .A(n2525), .B(n2524), .Z(n2529) );
  NANDN U3171 ( .A(n2527), .B(n2526), .Z(n2528) );
  NAND U3172 ( .A(n2529), .B(n2528), .Z(n2824) );
  XNOR U3173 ( .A(n2823), .B(n2824), .Z(n2825) );
  XOR U3174 ( .A(n2826), .B(n2825), .Z(n2677) );
  OR U3175 ( .A(n2531), .B(n2530), .Z(n2535) );
  OR U3176 ( .A(n2533), .B(n2532), .Z(n2534) );
  NAND U3177 ( .A(n2535), .B(n2534), .Z(n2678) );
  XNOR U3178 ( .A(n2677), .B(n2678), .Z(n2680) );
  XOR U3179 ( .A(n2679), .B(n2680), .Z(n2683) );
  OR U3180 ( .A(n2537), .B(n2536), .Z(n2541) );
  NANDN U3181 ( .A(n2539), .B(n2538), .Z(n2540) );
  AND U3182 ( .A(n2541), .B(n2540), .Z(n2684) );
  XNOR U3183 ( .A(n2683), .B(n2684), .Z(n2686) );
  XOR U3184 ( .A(n2685), .B(n2686), .Z(n2692) );
  OR U3185 ( .A(n2543), .B(n2542), .Z(n2547) );
  NANDN U3186 ( .A(n2545), .B(n2544), .Z(n2546) );
  AND U3187 ( .A(n2547), .B(n2546), .Z(n2732) );
  OR U3188 ( .A(n2549), .B(n2548), .Z(n2553) );
  OR U3189 ( .A(n2551), .B(n2550), .Z(n2552) );
  AND U3190 ( .A(n2553), .B(n2552), .Z(n2729) );
  NANDN U3191 ( .A(n2555), .B(n2554), .Z(n2559) );
  NANDN U3192 ( .A(n2557), .B(n2556), .Z(n2558) );
  AND U3193 ( .A(n2559), .B(n2558), .Z(n2726) );
  AND U3194 ( .A(y[657]), .B(x[140]), .Z(n2956) );
  ANDN U3195 ( .B(x[150]), .A(n143), .Z(n2806) );
  ANDN U3196 ( .B(y[668]), .A(n152), .Z(n2807) );
  XNOR U3197 ( .A(n2806), .B(n2807), .Z(n2808) );
  XNOR U3198 ( .A(n2956), .B(n2808), .Z(n2704) );
  OR U3199 ( .A(n2561), .B(n2560), .Z(n2565) );
  OR U3200 ( .A(n2563), .B(n2562), .Z(n2564) );
  AND U3201 ( .A(n2565), .B(n2564), .Z(n2701) );
  NAND U3202 ( .A(x[143]), .B(y[654]), .Z(n2810) );
  AND U3203 ( .A(x[149]), .B(y[648]), .Z(n3016) );
  NAND U3204 ( .A(y[649]), .B(x[148]), .Z(n2809) );
  XNOR U3205 ( .A(n3016), .B(n2809), .Z(n2811) );
  XNOR U3206 ( .A(n2701), .B(n2702), .Z(n2703) );
  XNOR U3207 ( .A(n2704), .B(n2703), .Z(n2727) );
  XOR U3208 ( .A(n2726), .B(n2727), .Z(n2728) );
  XNOR U3209 ( .A(n2732), .B(n2733), .Z(n2735) );
  OR U3210 ( .A(n2567), .B(n2566), .Z(n2571) );
  NANDN U3211 ( .A(n2569), .B(n2568), .Z(n2570) );
  AND U3212 ( .A(n2571), .B(n2570), .Z(n2734) );
  XOR U3213 ( .A(n2735), .B(n2734), .Z(n2738) );
  OR U3214 ( .A(n2573), .B(n2572), .Z(n2577) );
  NAND U3215 ( .A(n2575), .B(n2574), .Z(n2576) );
  NAND U3216 ( .A(n2577), .B(n2576), .Z(n2739) );
  XNOR U3217 ( .A(n2738), .B(n2739), .Z(n2741) );
  OR U3218 ( .A(n2579), .B(n2578), .Z(n2583) );
  OR U3219 ( .A(n2581), .B(n2580), .Z(n2582) );
  AND U3220 ( .A(n2583), .B(n2582), .Z(n2744) );
  NANDN U3221 ( .A(n2585), .B(n2584), .Z(n2589) );
  NANDN U3222 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U3223 ( .A(n2589), .B(n2588), .Z(n2745) );
  XOR U3224 ( .A(n2744), .B(n2745), .Z(n2746) );
  ANDN U3225 ( .B(y[663]), .A(n157), .Z(n2788) );
  ANDN U3226 ( .B(y[661]), .A(n159), .Z(n2786) );
  ANDN U3227 ( .B(y[662]), .A(n158), .Z(n2787) );
  XNOR U3228 ( .A(n2786), .B(n2787), .Z(n2789) );
  XNOR U3229 ( .A(n2788), .B(n2789), .Z(n2715) );
  NOR U3230 ( .A(n2590), .B(n160), .Z(n2927) );
  ANDN U3231 ( .B(y[664]), .A(n156), .Z(n2756) );
  ANDN U3232 ( .B(y[659]), .A(n161), .Z(n2757) );
  XNOR U3233 ( .A(n2756), .B(n2757), .Z(n2759) );
  ANDN U3234 ( .B(y[665]), .A(n155), .Z(n2758) );
  XNOR U3235 ( .A(n2759), .B(n2758), .Z(n2713) );
  XNOR U3236 ( .A(n2927), .B(n2713), .Z(n2714) );
  XNOR U3237 ( .A(n2715), .B(n2714), .Z(n2747) );
  XOR U3238 ( .A(n2746), .B(n2747), .Z(n2819) );
  OR U3239 ( .A(n2592), .B(n2591), .Z(n2596) );
  OR U3240 ( .A(n2594), .B(n2593), .Z(n2595) );
  AND U3241 ( .A(n2596), .B(n2595), .Z(n2818) );
  OR U3242 ( .A(n2598), .B(n2597), .Z(n2602) );
  OR U3243 ( .A(n2600), .B(n2599), .Z(n2601) );
  AND U3244 ( .A(n2602), .B(n2601), .Z(n2698) );
  OR U3245 ( .A(n2604), .B(n2603), .Z(n2608) );
  OR U3246 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U3247 ( .A(n2608), .B(n2607), .Z(n2695) );
  OR U3248 ( .A(n2610), .B(n2609), .Z(n2614) );
  OR U3249 ( .A(n2612), .B(n2611), .Z(n2613) );
  AND U3250 ( .A(n2614), .B(n2613), .Z(n2750) );
  ANDN U3251 ( .B(x[131]), .A(n2615), .Z(n2777) );
  ANDN U3252 ( .B(x[139]), .A(n2616), .Z(n2775) );
  ANDN U3253 ( .B(x[145]), .A(n2617), .Z(n2776) );
  XNOR U3254 ( .A(n2775), .B(n2776), .Z(n2778) );
  XNOR U3255 ( .A(n2777), .B(n2778), .Z(n2751) );
  XOR U3256 ( .A(n2750), .B(n2751), .Z(n2752) );
  NAND U3257 ( .A(y[656]), .B(x[141]), .Z(n2783) );
  ANDN U3258 ( .B(x[151]), .A(n2618), .Z(n2781) );
  AND U3259 ( .A(x[152]), .B(y[645]), .Z(n3044) );
  XOR U3260 ( .A(n2781), .B(n3044), .Z(n2782) );
  XNOR U3261 ( .A(n2783), .B(n2782), .Z(n2753) );
  XOR U3262 ( .A(n2752), .B(n2753), .Z(n2696) );
  XOR U3263 ( .A(n2695), .B(n2696), .Z(n2697) );
  OR U3264 ( .A(n2620), .B(n2619), .Z(n2624) );
  OR U3265 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U3266 ( .A(n2624), .B(n2623), .Z(n2794) );
  NAND U3267 ( .A(y[641]), .B(o[28]), .Z(n2625) );
  XNOR U3268 ( .A(y[642]), .B(n2625), .Z(n2626) );
  NAND U3269 ( .A(x[155]), .B(n2626), .Z(n2769) );
  ANDN U3270 ( .B(y[653]), .A(n167), .Z(n2768) );
  XNOR U3271 ( .A(n2769), .B(n2768), .Z(n2795) );
  XOR U3272 ( .A(n2794), .B(n2795), .Z(n2797) );
  ANDN U3273 ( .B(y[651]), .A(n169), .Z(n2762) );
  ANDN U3274 ( .B(x[147]), .A(n2627), .Z(n2763) );
  XNOR U3275 ( .A(n2762), .B(n2763), .Z(n2765) );
  ANDN U3276 ( .B(y[667]), .A(n153), .Z(n2764) );
  XOR U3277 ( .A(n2765), .B(n2764), .Z(n2796) );
  XNOR U3278 ( .A(n2797), .B(n2796), .Z(n2830) );
  OR U3279 ( .A(n2629), .B(n2628), .Z(n2633) );
  OR U3280 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U3281 ( .A(n2633), .B(n2632), .Z(n2710) );
  ANDN U3282 ( .B(x[156]), .A(n139), .Z(n2816) );
  XOR U3283 ( .A(o[29]), .B(n2816), .Z(n2720) );
  ANDN U3284 ( .B(x[157]), .A(n138), .Z(n2721) );
  XNOR U3285 ( .A(n2720), .B(n2721), .Z(n2723) );
  ANDN U3286 ( .B(y[669]), .A(n151), .Z(n2722) );
  XOR U3287 ( .A(n2723), .B(n2722), .Z(n2707) );
  NAND U3288 ( .A(y[655]), .B(x[142]), .Z(n2802) );
  ANDN U3289 ( .B(x[153]), .A(n2634), .Z(n2801) );
  NAND U3290 ( .A(x[154]), .B(y[643]), .Z(n2800) );
  XOR U3291 ( .A(n2801), .B(n2800), .Z(n2803) );
  XNOR U3292 ( .A(n2802), .B(n2803), .Z(n2708) );
  XNOR U3293 ( .A(n2707), .B(n2708), .Z(n2709) );
  XOR U3294 ( .A(n2710), .B(n2709), .Z(n2829) );
  XNOR U3295 ( .A(n2830), .B(n2829), .Z(n2831) );
  XNOR U3296 ( .A(n2832), .B(n2831), .Z(n2817) );
  XOR U3297 ( .A(n2818), .B(n2817), .Z(n2820) );
  XNOR U3298 ( .A(n2819), .B(n2820), .Z(n2740) );
  XOR U3299 ( .A(n2741), .B(n2740), .Z(n2690) );
  NANDN U3300 ( .A(n2636), .B(n2635), .Z(n2640) );
  NANDN U3301 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U3302 ( .A(n2640), .B(n2639), .Z(n2689) );
  XOR U3303 ( .A(n2690), .B(n2689), .Z(n2691) );
  OR U3304 ( .A(n2642), .B(n2641), .Z(n2646) );
  NANDN U3305 ( .A(n2644), .B(n2643), .Z(n2645) );
  AND U3306 ( .A(n2646), .B(n2645), .Z(n2835) );
  NANDN U3307 ( .A(n2648), .B(n2647), .Z(n2652) );
  OR U3308 ( .A(n2650), .B(n2649), .Z(n2651) );
  AND U3309 ( .A(n2652), .B(n2651), .Z(n2836) );
  XOR U3310 ( .A(n2835), .B(n2836), .Z(n2837) );
  XOR U3311 ( .A(n2838), .B(n2837), .Z(n2674) );
  OR U3312 ( .A(n2654), .B(n2653), .Z(n2658) );
  NANDN U3313 ( .A(n2656), .B(n2655), .Z(n2657) );
  AND U3314 ( .A(n2658), .B(n2657), .Z(n2671) );
  OR U3315 ( .A(n2660), .B(n2659), .Z(n2664) );
  NANDN U3316 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U3317 ( .A(n2664), .B(n2663), .Z(n2672) );
  XNOR U3318 ( .A(n2671), .B(n2672), .Z(n2673) );
  XOR U3319 ( .A(n2674), .B(n2673), .Z(n2668) );
  XNOR U3320 ( .A(n2667), .B(n2668), .Z(N62) );
  NANDN U3321 ( .A(n2666), .B(n2665), .Z(n2670) );
  NAND U3322 ( .A(n2668), .B(n2667), .Z(n2669) );
  AND U3323 ( .A(n2670), .B(n2669), .Z(n2843) );
  OR U3324 ( .A(n2672), .B(n2671), .Z(n2676) );
  OR U3325 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U3326 ( .A(n2676), .B(n2675), .Z(n2844) );
  XNOR U3327 ( .A(n2843), .B(n2844), .Z(n2842) );
  OR U3328 ( .A(n2678), .B(n2677), .Z(n2682) );
  OR U3329 ( .A(n2680), .B(n2679), .Z(n2681) );
  NAND U3330 ( .A(n2682), .B(n2681), .Z(n3135) );
  OR U3331 ( .A(n2684), .B(n2683), .Z(n2688) );
  OR U3332 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U3333 ( .A(n2688), .B(n2687), .Z(n3133) );
  OR U3334 ( .A(n2690), .B(n2689), .Z(n2694) );
  NANDN U3335 ( .A(n2692), .B(n2691), .Z(n2693) );
  NAND U3336 ( .A(n2694), .B(n2693), .Z(n3134) );
  XNOR U3337 ( .A(n3133), .B(n3134), .Z(n3136) );
  XOR U3338 ( .A(n3135), .B(n3136), .Z(n3128) );
  OR U3339 ( .A(n2696), .B(n2695), .Z(n2700) );
  NANDN U3340 ( .A(n2698), .B(n2697), .Z(n2699) );
  AND U3341 ( .A(n2700), .B(n2699), .Z(n3095) );
  OR U3342 ( .A(n2702), .B(n2701), .Z(n2706) );
  OR U3343 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U3344 ( .A(n2706), .B(n2705), .Z(n3096) );
  XOR U3345 ( .A(n3095), .B(n3096), .Z(n3093) );
  OR U3346 ( .A(n2708), .B(n2707), .Z(n2712) );
  OR U3347 ( .A(n2710), .B(n2709), .Z(n2711) );
  NAND U3348 ( .A(n2712), .B(n2711), .Z(n3094) );
  XNOR U3349 ( .A(n3093), .B(n3094), .Z(n3090) );
  NAND U3350 ( .A(y[643]), .B(x[155]), .Z(n3050) );
  NAND U3351 ( .A(x[129]), .B(y[669]), .Z(n3049) );
  XNOR U3352 ( .A(n3050), .B(n3049), .Z(n3052) );
  XNOR U3353 ( .A(n3051), .B(n3052), .Z(n2913) );
  AND U3354 ( .A(y[658]), .B(x[140]), .Z(n2716) );
  XNOR U3355 ( .A(n2717), .B(n2716), .Z(n2957) );
  AND U3356 ( .A(y[661]), .B(x[137]), .Z(n2719) );
  AND U3357 ( .A(y[660]), .B(x[138]), .Z(n2718) );
  XNOR U3358 ( .A(n2719), .B(n2718), .Z(n2925) );
  XOR U3359 ( .A(n2926), .B(n2925), .Z(n2915) );
  OR U3360 ( .A(n2721), .B(n2720), .Z(n2725) );
  OR U3361 ( .A(n2723), .B(n2722), .Z(n2724) );
  AND U3362 ( .A(n2725), .B(n2724), .Z(n2916) );
  XNOR U3363 ( .A(n2915), .B(n2916), .Z(n2914) );
  XOR U3364 ( .A(n2913), .B(n2914), .Z(n2869) );
  XNOR U3365 ( .A(n2870), .B(n2869), .Z(n2868) );
  OR U3366 ( .A(n2727), .B(n2726), .Z(n2731) );
  NANDN U3367 ( .A(n2729), .B(n2728), .Z(n2730) );
  NAND U3368 ( .A(n2731), .B(n2730), .Z(n2867) );
  XOR U3369 ( .A(n2868), .B(n2867), .Z(n3089) );
  XOR U3370 ( .A(n3090), .B(n3089), .Z(n3088) );
  OR U3371 ( .A(n2733), .B(n2732), .Z(n2737) );
  OR U3372 ( .A(n2735), .B(n2734), .Z(n2736) );
  NAND U3373 ( .A(n2737), .B(n2736), .Z(n3087) );
  XOR U3374 ( .A(n3088), .B(n3087), .Z(n3117) );
  OR U3375 ( .A(n2739), .B(n2738), .Z(n2743) );
  NANDN U3376 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U3377 ( .A(n2743), .B(n2742), .Z(n3118) );
  OR U3378 ( .A(n2745), .B(n2744), .Z(n2749) );
  NANDN U3379 ( .A(n2747), .B(n2746), .Z(n2748) );
  AND U3380 ( .A(n2749), .B(n2748), .Z(n2859) );
  OR U3381 ( .A(n2751), .B(n2750), .Z(n2755) );
  NANDN U3382 ( .A(n2753), .B(n2752), .Z(n2754) );
  AND U3383 ( .A(n2755), .B(n2754), .Z(n2861) );
  OR U3384 ( .A(n2757), .B(n2756), .Z(n2761) );
  OR U3385 ( .A(n2759), .B(n2758), .Z(n2760) );
  AND U3386 ( .A(n2761), .B(n2760), .Z(n2886) );
  NAND U3387 ( .A(x[134]), .B(y[664]), .Z(n2936) );
  NAND U3388 ( .A(x[133]), .B(y[665]), .Z(n2935) );
  NAND U3389 ( .A(x[147]), .B(y[651]), .Z(n2934) );
  XNOR U3390 ( .A(n2935), .B(n2934), .Z(n2937) );
  XNOR U3391 ( .A(n2936), .B(n2937), .Z(n2905) );
  OR U3392 ( .A(n2763), .B(n2762), .Z(n2767) );
  OR U3393 ( .A(n2765), .B(n2764), .Z(n2766) );
  AND U3394 ( .A(n2767), .B(n2766), .Z(n2907) );
  NAND U3395 ( .A(y[666]), .B(x[132]), .Z(n2951) );
  NAND U3396 ( .A(x[131]), .B(y[667]), .Z(n2952) );
  AND U3397 ( .A(y[652]), .B(x[146]), .Z(n2953) );
  XNOR U3398 ( .A(n2952), .B(n2953), .Z(n2950) );
  XNOR U3399 ( .A(n2951), .B(n2950), .Z(n2908) );
  XOR U3400 ( .A(n2907), .B(n2908), .Z(n2906) );
  XNOR U3401 ( .A(n2905), .B(n2906), .Z(n2885) );
  XOR U3402 ( .A(n2886), .B(n2885), .Z(n2888) );
  OR U3403 ( .A(n2769), .B(n2768), .Z(n2774) );
  NAND U3404 ( .A(o[28]), .B(n2770), .Z(n2772) );
  NAND U3405 ( .A(y[642]), .B(x[155]), .Z(n2771) );
  AND U3406 ( .A(n2772), .B(n2771), .Z(n2773) );
  ANDN U3407 ( .B(n2774), .A(n2773), .Z(n2887) );
  XNOR U3408 ( .A(n2861), .B(n2862), .Z(n2860) );
  XNOR U3409 ( .A(n2859), .B(n2860), .Z(n3112) );
  OR U3410 ( .A(n2776), .B(n2775), .Z(n2780) );
  OR U3411 ( .A(n2778), .B(n2777), .Z(n2779) );
  NAND U3412 ( .A(n2780), .B(n2779), .Z(n2894) );
  NAND U3413 ( .A(x[148]), .B(y[650]), .Z(n3066) );
  AND U3414 ( .A(x[142]), .B(y[656]), .Z(n3065) );
  XOR U3415 ( .A(n3066), .B(n3065), .Z(n3064) );
  AND U3416 ( .A(y[662]), .B(x[136]), .Z(n3063) );
  XOR U3417 ( .A(n3064), .B(n3063), .Z(n2896) );
  NAND U3418 ( .A(y[640]), .B(x[158]), .Z(n2922) );
  NAND U3419 ( .A(y[641]), .B(x[157]), .Z(n2975) );
  XNOR U3420 ( .A(o[30]), .B(n2975), .Z(n2921) );
  XOR U3421 ( .A(n2922), .B(n2921), .Z(n2920) );
  AND U3422 ( .A(y[670]), .B(x[128]), .Z(n2919) );
  XNOR U3423 ( .A(n2920), .B(n2919), .Z(n2895) );
  XOR U3424 ( .A(n2894), .B(n2893), .Z(n2875) );
  OR U3425 ( .A(n2781), .B(n3044), .Z(n2785) );
  NAND U3426 ( .A(n2783), .B(n2782), .Z(n2784) );
  AND U3427 ( .A(n2785), .B(n2784), .Z(n2876) );
  XNOR U3428 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U3429 ( .A(n2787), .B(n2786), .Z(n2791) );
  OR U3430 ( .A(n2789), .B(n2788), .Z(n2790) );
  AND U3431 ( .A(n2791), .B(n2790), .Z(n2970) );
  NAND U3432 ( .A(x[145]), .B(y[653]), .Z(n3021) );
  NAND U3433 ( .A(x[130]), .B(y[668]), .Z(n3023) );
  NAND U3434 ( .A(y[644]), .B(x[154]), .Z(n3022) );
  XNOR U3435 ( .A(n3023), .B(n3022), .Z(n3020) );
  XNOR U3436 ( .A(n3021), .B(n3020), .Z(n2972) );
  NAND U3437 ( .A(x[135]), .B(y[663]), .Z(n3015) );
  AND U3438 ( .A(y[648]), .B(x[150]), .Z(n2793) );
  AND U3439 ( .A(x[149]), .B(y[649]), .Z(n2792) );
  XNOR U3440 ( .A(n2793), .B(n2792), .Z(n3014) );
  XOR U3441 ( .A(n3015), .B(n3014), .Z(n2971) );
  XNOR U3442 ( .A(n2972), .B(n2971), .Z(n2969) );
  XOR U3443 ( .A(n2970), .B(n2969), .Z(n2873) );
  XNOR U3444 ( .A(n2874), .B(n2873), .Z(n2853) );
  OR U3445 ( .A(n2795), .B(n2794), .Z(n2799) );
  NAND U3446 ( .A(n2797), .B(n2796), .Z(n2798) );
  NAND U3447 ( .A(n2799), .B(n2798), .Z(n2856) );
  NANDN U3448 ( .A(n2801), .B(n2800), .Z(n2805) );
  NANDN U3449 ( .A(n2803), .B(n2802), .Z(n2804) );
  AND U3450 ( .A(n2805), .B(n2804), .Z(n2879) );
  NANDN U3451 ( .A(n3016), .B(n2809), .Z(n2813) );
  NAND U3452 ( .A(n2811), .B(n2810), .Z(n2812) );
  AND U3453 ( .A(n2813), .B(n2812), .Z(n2899) );
  NAND U3454 ( .A(y[647]), .B(x[151]), .Z(n3045) );
  AND U3455 ( .A(x[153]), .B(y[645]), .Z(n2815) );
  AND U3456 ( .A(x[152]), .B(y[646]), .Z(n2814) );
  XNOR U3457 ( .A(n2815), .B(n2814), .Z(n3046) );
  XOR U3458 ( .A(n3045), .B(n3046), .Z(n2901) );
  NAND U3459 ( .A(n2816), .B(o[29]), .Z(n3058) );
  NAND U3460 ( .A(x[156]), .B(y[642]), .Z(n3060) );
  AND U3461 ( .A(x[144]), .B(y[654]), .Z(n3059) );
  XNOR U3462 ( .A(n3060), .B(n3059), .Z(n3057) );
  XNOR U3463 ( .A(n3058), .B(n3057), .Z(n2902) );
  XNOR U3464 ( .A(n2901), .B(n2902), .Z(n2900) );
  XOR U3465 ( .A(n2899), .B(n2900), .Z(n2881) );
  XOR U3466 ( .A(n2879), .B(n2880), .Z(n2855) );
  XNOR U3467 ( .A(n2856), .B(n2855), .Z(n2854) );
  XNOR U3468 ( .A(n2853), .B(n2854), .Z(n3111) );
  XNOR U3469 ( .A(n3112), .B(n3111), .Z(n3110) );
  NANDN U3470 ( .A(n2818), .B(n2817), .Z(n2822) );
  NANDN U3471 ( .A(n2820), .B(n2819), .Z(n2821) );
  NAND U3472 ( .A(n2822), .B(n2821), .Z(n3109) );
  XNOR U3473 ( .A(n3110), .B(n3109), .Z(n2847) );
  OR U3474 ( .A(n2824), .B(n2823), .Z(n2828) );
  OR U3475 ( .A(n2826), .B(n2825), .Z(n2827) );
  NAND U3476 ( .A(n2828), .B(n2827), .Z(n2850) );
  OR U3477 ( .A(n2830), .B(n2829), .Z(n2834) );
  OR U3478 ( .A(n2832), .B(n2831), .Z(n2833) );
  NAND U3479 ( .A(n2834), .B(n2833), .Z(n2849) );
  XNOR U3480 ( .A(n2850), .B(n2849), .Z(n2848) );
  XOR U3481 ( .A(n2847), .B(n2848), .Z(n3115) );
  XNOR U3482 ( .A(n3116), .B(n3115), .Z(n3127) );
  XNOR U3483 ( .A(n3128), .B(n3127), .Z(n3130) );
  OR U3484 ( .A(n2836), .B(n2835), .Z(n2840) );
  NANDN U3485 ( .A(n2838), .B(n2837), .Z(n2839) );
  NAND U3486 ( .A(n2840), .B(n2839), .Z(n3129) );
  XOR U3487 ( .A(n3130), .B(n3129), .Z(n2841) );
  XNOR U3488 ( .A(n2842), .B(n2841), .Z(N63) );
  OR U3489 ( .A(n2842), .B(n2841), .Z(n2846) );
  OR U3490 ( .A(n2844), .B(n2843), .Z(n2845) );
  AND U3491 ( .A(n2846), .B(n2845), .Z(n3126) );
  NANDN U3492 ( .A(n2848), .B(n2847), .Z(n2852) );
  NOR U3493 ( .A(n2850), .B(n2849), .Z(n2851) );
  ANDN U3494 ( .B(n2852), .A(n2851), .Z(n3108) );
  NANDN U3495 ( .A(n2854), .B(n2853), .Z(n2858) );
  OR U3496 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U3497 ( .A(n2858), .B(n2857), .Z(n2866) );
  OR U3498 ( .A(n2860), .B(n2859), .Z(n2864) );
  OR U3499 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U3500 ( .A(n2864), .B(n2863), .Z(n2865) );
  XNOR U3501 ( .A(n2866), .B(n2865), .Z(n3106) );
  OR U3502 ( .A(n2868), .B(n2867), .Z(n2872) );
  OR U3503 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3504 ( .A(n2872), .B(n2871), .Z(n3104) );
  OR U3505 ( .A(n2874), .B(n2873), .Z(n2878) );
  OR U3506 ( .A(n2876), .B(n2875), .Z(n2877) );
  AND U3507 ( .A(n2878), .B(n2877), .Z(n3086) );
  OR U3508 ( .A(n2880), .B(n2879), .Z(n2884) );
  NANDN U3509 ( .A(n2882), .B(n2881), .Z(n2883) );
  AND U3510 ( .A(n2884), .B(n2883), .Z(n2892) );
  NOR U3511 ( .A(n2886), .B(n2885), .Z(n2890) );
  ANDN U3512 ( .B(n2888), .A(n2887), .Z(n2889) );
  OR U3513 ( .A(n2890), .B(n2889), .Z(n2891) );
  XNOR U3514 ( .A(n2892), .B(n2891), .Z(n3084) );
  OR U3515 ( .A(n2894), .B(n2893), .Z(n2898) );
  NANDN U3516 ( .A(n2896), .B(n2895), .Z(n2897) );
  AND U3517 ( .A(n2898), .B(n2897), .Z(n3082) );
  OR U3518 ( .A(n2900), .B(n2899), .Z(n2904) );
  OR U3519 ( .A(n2902), .B(n2901), .Z(n2903) );
  AND U3520 ( .A(n2904), .B(n2903), .Z(n2912) );
  NAND U3521 ( .A(n2906), .B(n2905), .Z(n2910) );
  OR U3522 ( .A(n2908), .B(n2907), .Z(n2909) );
  NAND U3523 ( .A(n2910), .B(n2909), .Z(n2911) );
  XNOR U3524 ( .A(n2912), .B(n2911), .Z(n3080) );
  OR U3525 ( .A(n2914), .B(n2913), .Z(n2918) );
  OR U3526 ( .A(n2916), .B(n2915), .Z(n2917) );
  AND U3527 ( .A(n2918), .B(n2917), .Z(n3078) );
  NANDN U3528 ( .A(n2920), .B(n2919), .Z(n2924) );
  NANDN U3529 ( .A(n2922), .B(n2921), .Z(n2923) );
  AND U3530 ( .A(n2924), .B(n2923), .Z(n2931) );
  OR U3531 ( .A(n2926), .B(n2925), .Z(n2929) );
  NAND U3532 ( .A(x[138]), .B(y[661]), .Z(n2976) );
  NANDN U3533 ( .A(n2976), .B(n2927), .Z(n2928) );
  NAND U3534 ( .A(n2929), .B(n2928), .Z(n2930) );
  XNOR U3535 ( .A(n2931), .B(n2930), .Z(n3076) );
  AND U3536 ( .A(y[664]), .B(x[135]), .Z(n2933) );
  NAND U3537 ( .A(y[666]), .B(x[133]), .Z(n2932) );
  XNOR U3538 ( .A(n2933), .B(n2932), .Z(n2949) );
  NOR U3539 ( .A(n2935), .B(n2934), .Z(n2939) );
  NOR U3540 ( .A(n2937), .B(n2936), .Z(n2938) );
  NOR U3541 ( .A(n2939), .B(n2938), .Z(n2947) );
  AND U3542 ( .A(x[159]), .B(y[640]), .Z(n2941) );
  AND U3543 ( .A(y[669]), .B(x[130]), .Z(n2940) );
  XNOR U3544 ( .A(n2941), .B(n2940), .Z(n2945) );
  AND U3545 ( .A(y[654]), .B(x[145]), .Z(n2943) );
  NAND U3546 ( .A(x[142]), .B(y[657]), .Z(n2942) );
  XNOR U3547 ( .A(n2943), .B(n2942), .Z(n2944) );
  XOR U3548 ( .A(n2945), .B(n2944), .Z(n2946) );
  XNOR U3549 ( .A(n2947), .B(n2946), .Z(n2948) );
  XOR U3550 ( .A(n2949), .B(n2948), .Z(n2968) );
  NANDN U3551 ( .A(n2951), .B(n2950), .Z(n2955) );
  ANDN U3552 ( .B(n2953), .A(n2952), .Z(n2954) );
  ANDN U3553 ( .B(n2955), .A(n2954), .Z(n2962) );
  AND U3554 ( .A(n2977), .B(n2956), .Z(n2960) );
  ANDN U3555 ( .B(n2958), .A(n2957), .Z(n2959) );
  OR U3556 ( .A(n2960), .B(n2959), .Z(n2961) );
  XNOR U3557 ( .A(n2962), .B(n2961), .Z(n2966) );
  AND U3558 ( .A(y[648]), .B(x[151]), .Z(n2964) );
  NAND U3559 ( .A(x[132]), .B(y[667]), .Z(n2963) );
  XNOR U3560 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U3561 ( .A(n2966), .B(n2965), .Z(n2967) );
  XNOR U3562 ( .A(n2968), .B(n2967), .Z(n3042) );
  NANDN U3563 ( .A(n2970), .B(n2969), .Z(n2974) );
  ANDN U3564 ( .B(n2972), .A(n2971), .Z(n2973) );
  ANDN U3565 ( .B(n2974), .A(n2973), .Z(n3040) );
  AND U3566 ( .A(y[668]), .B(x[131]), .Z(n2983) );
  ANDN U3567 ( .B(o[30]), .A(n2975), .Z(n2981) );
  NAND U3568 ( .A(y[649]), .B(x[150]), .Z(n3017) );
  XNOR U3569 ( .A(n3017), .B(o[31]), .Z(n2979) );
  XOR U3570 ( .A(n2977), .B(n2976), .Z(n2978) );
  XNOR U3571 ( .A(n2979), .B(n2978), .Z(n2980) );
  XNOR U3572 ( .A(n2981), .B(n2980), .Z(n2982) );
  XNOR U3573 ( .A(n2983), .B(n2982), .Z(n2991) );
  AND U3574 ( .A(y[665]), .B(x[134]), .Z(n2985) );
  NAND U3575 ( .A(y[644]), .B(x[155]), .Z(n2984) );
  XNOR U3576 ( .A(n2985), .B(n2984), .Z(n2989) );
  AND U3577 ( .A(x[146]), .B(y[653]), .Z(n2987) );
  NAND U3578 ( .A(x[152]), .B(y[647]), .Z(n2986) );
  XNOR U3579 ( .A(n2987), .B(n2986), .Z(n2988) );
  XNOR U3580 ( .A(n2989), .B(n2988), .Z(n2990) );
  XNOR U3581 ( .A(n2991), .B(n2990), .Z(n3038) );
  AND U3582 ( .A(y[662]), .B(x[137]), .Z(n2993) );
  NAND U3583 ( .A(x[148]), .B(y[651]), .Z(n2992) );
  XNOR U3584 ( .A(n2993), .B(n2992), .Z(n2997) );
  AND U3585 ( .A(y[652]), .B(x[147]), .Z(n2995) );
  NAND U3586 ( .A(x[144]), .B(y[655]), .Z(n2994) );
  XNOR U3587 ( .A(n2995), .B(n2994), .Z(n2996) );
  XOR U3588 ( .A(n2997), .B(n2996), .Z(n3005) );
  AND U3589 ( .A(y[642]), .B(x[157]), .Z(n2999) );
  NAND U3590 ( .A(y[641]), .B(x[158]), .Z(n2998) );
  XNOR U3591 ( .A(n2999), .B(n2998), .Z(n3003) );
  AND U3592 ( .A(y[663]), .B(x[136]), .Z(n3001) );
  NAND U3593 ( .A(y[650]), .B(x[149]), .Z(n3000) );
  XNOR U3594 ( .A(n3001), .B(n3000), .Z(n3002) );
  XNOR U3595 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U3596 ( .A(n3005), .B(n3004), .Z(n3013) );
  AND U3597 ( .A(y[659]), .B(x[140]), .Z(n3007) );
  NAND U3598 ( .A(y[660]), .B(x[139]), .Z(n3006) );
  XNOR U3599 ( .A(n3007), .B(n3006), .Z(n3011) );
  AND U3600 ( .A(y[671]), .B(x[128]), .Z(n3009) );
  NAND U3601 ( .A(x[154]), .B(y[645]), .Z(n3008) );
  XNOR U3602 ( .A(n3009), .B(n3008), .Z(n3010) );
  XNOR U3603 ( .A(n3011), .B(n3010), .Z(n3012) );
  XNOR U3604 ( .A(n3013), .B(n3012), .Z(n3029) );
  OR U3605 ( .A(n3015), .B(n3014), .Z(n3019) );
  NANDN U3606 ( .A(n3017), .B(n3016), .Z(n3018) );
  AND U3607 ( .A(n3019), .B(n3018), .Z(n3027) );
  OR U3608 ( .A(n3021), .B(n3020), .Z(n3025) );
  OR U3609 ( .A(n3023), .B(n3022), .Z(n3024) );
  NAND U3610 ( .A(n3025), .B(n3024), .Z(n3026) );
  XNOR U3611 ( .A(n3027), .B(n3026), .Z(n3028) );
  XOR U3612 ( .A(n3029), .B(n3028), .Z(n3036) );
  NAND U3613 ( .A(x[153]), .B(y[646]), .Z(n3043) );
  AND U3614 ( .A(y[656]), .B(x[143]), .Z(n3031) );
  NAND U3615 ( .A(x[129]), .B(y[670]), .Z(n3030) );
  XNOR U3616 ( .A(n3031), .B(n3030), .Z(n3033) );
  NAND U3617 ( .A(y[643]), .B(x[156]), .Z(n3032) );
  XNOR U3618 ( .A(n3033), .B(n3032), .Z(n3034) );
  XOR U3619 ( .A(n3043), .B(n3034), .Z(n3035) );
  XNOR U3620 ( .A(n3036), .B(n3035), .Z(n3037) );
  XNOR U3621 ( .A(n3038), .B(n3037), .Z(n3039) );
  XNOR U3622 ( .A(n3040), .B(n3039), .Z(n3041) );
  XOR U3623 ( .A(n3042), .B(n3041), .Z(n3074) );
  ANDN U3624 ( .B(n3044), .A(n3043), .Z(n3048) );
  NOR U3625 ( .A(n3046), .B(n3045), .Z(n3047) );
  NOR U3626 ( .A(n3048), .B(n3047), .Z(n3056) );
  OR U3627 ( .A(n3050), .B(n3049), .Z(n3054) );
  NANDN U3628 ( .A(n3052), .B(n3051), .Z(n3053) );
  AND U3629 ( .A(n3054), .B(n3053), .Z(n3055) );
  XNOR U3630 ( .A(n3056), .B(n3055), .Z(n3072) );
  NANDN U3631 ( .A(n3058), .B(n3057), .Z(n3062) );
  NANDN U3632 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U3633 ( .A(n3062), .B(n3061), .Z(n3070) );
  NANDN U3634 ( .A(n3064), .B(n3063), .Z(n3068) );
  NANDN U3635 ( .A(n3066), .B(n3065), .Z(n3067) );
  NAND U3636 ( .A(n3068), .B(n3067), .Z(n3069) );
  XNOR U3637 ( .A(n3070), .B(n3069), .Z(n3071) );
  XOR U3638 ( .A(n3072), .B(n3071), .Z(n3073) );
  XNOR U3639 ( .A(n3074), .B(n3073), .Z(n3075) );
  XNOR U3640 ( .A(n3076), .B(n3075), .Z(n3077) );
  XNOR U3641 ( .A(n3078), .B(n3077), .Z(n3079) );
  XNOR U3642 ( .A(n3080), .B(n3079), .Z(n3081) );
  XNOR U3643 ( .A(n3082), .B(n3081), .Z(n3083) );
  XNOR U3644 ( .A(n3084), .B(n3083), .Z(n3085) );
  XNOR U3645 ( .A(n3086), .B(n3085), .Z(n3102) );
  OR U3646 ( .A(n3088), .B(n3087), .Z(n3092) );
  NANDN U3647 ( .A(n3090), .B(n3089), .Z(n3091) );
  AND U3648 ( .A(n3092), .B(n3091), .Z(n3100) );
  NANDN U3649 ( .A(n3094), .B(n3093), .Z(n3098) );
  OR U3650 ( .A(n3096), .B(n3095), .Z(n3097) );
  NAND U3651 ( .A(n3098), .B(n3097), .Z(n3099) );
  XNOR U3652 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U3653 ( .A(n3102), .B(n3101), .Z(n3103) );
  XNOR U3654 ( .A(n3104), .B(n3103), .Z(n3105) );
  XNOR U3655 ( .A(n3106), .B(n3105), .Z(n3107) );
  XNOR U3656 ( .A(n3108), .B(n3107), .Z(n3124) );
  OR U3657 ( .A(n3110), .B(n3109), .Z(n3114) );
  OR U3658 ( .A(n3112), .B(n3111), .Z(n3113) );
  AND U3659 ( .A(n3114), .B(n3113), .Z(n3122) );
  OR U3660 ( .A(n3116), .B(n3115), .Z(n3120) );
  NANDN U3661 ( .A(n3118), .B(n3117), .Z(n3119) );
  NAND U3662 ( .A(n3120), .B(n3119), .Z(n3121) );
  XNOR U3663 ( .A(n3122), .B(n3121), .Z(n3123) );
  XNOR U3664 ( .A(n3124), .B(n3123), .Z(n3125) );
  XNOR U3665 ( .A(n3126), .B(n3125), .Z(n3142) );
  NOR U3666 ( .A(n3128), .B(n3127), .Z(n3132) );
  NOR U3667 ( .A(n3130), .B(n3129), .Z(n3131) );
  NOR U3668 ( .A(n3132), .B(n3131), .Z(n3140) );
  OR U3669 ( .A(n3134), .B(n3133), .Z(n3138) );
  NOR U3670 ( .A(n3136), .B(n3135), .Z(n3137) );
  ANDN U3671 ( .B(n3138), .A(n3137), .Z(n3139) );
  XNOR U3672 ( .A(n3140), .B(n3139), .Z(n3141) );
  XNOR U3673 ( .A(n3142), .B(n3141), .Z(N64) );
  AND U3674 ( .A(x[128]), .B(y[672]), .Z(n3852) );
  XOR U3675 ( .A(n3852), .B(o[32]), .Z(N97) );
  AND U3676 ( .A(x[129]), .B(y[672]), .Z(n3143) );
  NAND U3677 ( .A(x[128]), .B(y[673]), .Z(n3149) );
  XNOR U3678 ( .A(n3149), .B(o[33]), .Z(n3144) );
  XOR U3679 ( .A(n3143), .B(n3144), .Z(n3145) );
  AND U3680 ( .A(o[32]), .B(n3852), .Z(n3146) );
  XOR U3681 ( .A(n3145), .B(n3146), .Z(N98) );
  OR U3682 ( .A(n3144), .B(n3143), .Z(n3148) );
  NANDN U3683 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U3684 ( .A(n3148), .B(n3147), .Z(n3151) );
  NAND U3685 ( .A(x[128]), .B(y[674]), .Z(n3162) );
  XOR U3686 ( .A(n3162), .B(o[34]), .Z(n3150) );
  XNOR U3687 ( .A(n3151), .B(n3150), .Z(n3153) );
  ANDN U3688 ( .B(o[33]), .A(n3149), .Z(n3156) );
  ANDN U3689 ( .B(y[672]), .A(n153), .Z(n3157) );
  XNOR U3690 ( .A(n3156), .B(n3157), .Z(n3159) );
  ANDN U3691 ( .B(y[673]), .A(n152), .Z(n3158) );
  XNOR U3692 ( .A(n3159), .B(n3158), .Z(n3152) );
  XNOR U3693 ( .A(n3153), .B(n3152), .Z(N99) );
  NAND U3694 ( .A(n3151), .B(n3150), .Z(n3155) );
  OR U3695 ( .A(n3153), .B(n3152), .Z(n3154) );
  NAND U3696 ( .A(n3155), .B(n3154), .Z(n3166) );
  OR U3697 ( .A(n3157), .B(n3156), .Z(n3161) );
  OR U3698 ( .A(n3159), .B(n3158), .Z(n3160) );
  AND U3699 ( .A(n3161), .B(n3160), .Z(n3167) );
  XNOR U3700 ( .A(n3166), .B(n3167), .Z(n3168) );
  NAND U3701 ( .A(x[130]), .B(y[673]), .Z(n3178) );
  XNOR U3702 ( .A(n3178), .B(o[35]), .Z(n3172) );
  NANDN U3703 ( .A(n3162), .B(o[34]), .Z(n3175) );
  AND U3704 ( .A(x[131]), .B(y[672]), .Z(n3164) );
  NAND U3705 ( .A(x[128]), .B(y[675]), .Z(n3163) );
  XOR U3706 ( .A(n3164), .B(n3163), .Z(n3174) );
  XNOR U3707 ( .A(n3175), .B(n3174), .Z(n3173) );
  ANDN U3708 ( .B(y[674]), .A(n152), .Z(n3202) );
  XOR U3709 ( .A(n3173), .B(n3202), .Z(n3165) );
  XOR U3710 ( .A(n3172), .B(n3165), .Z(n3169) );
  XNOR U3711 ( .A(n3168), .B(n3169), .Z(N100) );
  NANDN U3712 ( .A(n3167), .B(n3166), .Z(n3171) );
  NAND U3713 ( .A(n3169), .B(n3168), .Z(n3170) );
  NAND U3714 ( .A(n3171), .B(n3170), .Z(n3183) );
  XNOR U3715 ( .A(n3183), .B(n3184), .Z(n3185) );
  ANDN U3716 ( .B(y[675]), .A(n154), .Z(n3250) );
  NAND U3717 ( .A(n3852), .B(n3250), .Z(n3177) );
  OR U3718 ( .A(n3175), .B(n3174), .Z(n3176) );
  NAND U3719 ( .A(n3177), .B(n3176), .Z(n3192) );
  NANDN U3720 ( .A(n3178), .B(o[35]), .Z(n3199) );
  AND U3721 ( .A(y[672]), .B(x[132]), .Z(n3180) );
  AND U3722 ( .A(y[676]), .B(x[128]), .Z(n3179) );
  XNOR U3723 ( .A(n3180), .B(n3179), .Z(n3198) );
  XOR U3724 ( .A(n3199), .B(n3198), .Z(n3190) );
  AND U3725 ( .A(x[129]), .B(y[675]), .Z(n3182) );
  NAND U3726 ( .A(x[130]), .B(y[674]), .Z(n3181) );
  XOR U3727 ( .A(n3182), .B(n3181), .Z(n3204) );
  NAND U3728 ( .A(x[131]), .B(y[673]), .Z(n3195) );
  XNOR U3729 ( .A(n3195), .B(o[36]), .Z(n3203) );
  XOR U3730 ( .A(n3192), .B(n3191), .Z(n3186) );
  XOR U3731 ( .A(n3185), .B(n3186), .Z(N101) );
  NANDN U3732 ( .A(n3184), .B(n3183), .Z(n3188) );
  NANDN U3733 ( .A(n3186), .B(n3185), .Z(n3187) );
  NAND U3734 ( .A(n3188), .B(n3187), .Z(n3207) );
  NAND U3735 ( .A(n3190), .B(n3189), .Z(n3194) );
  NAND U3736 ( .A(n3192), .B(n3191), .Z(n3193) );
  NAND U3737 ( .A(n3194), .B(n3193), .Z(n3208) );
  XNOR U3738 ( .A(n3207), .B(n3208), .Z(n3209) );
  NANDN U3739 ( .A(n3195), .B(o[36]), .Z(n3226) );
  AND U3740 ( .A(x[133]), .B(y[672]), .Z(n3197) );
  AND U3741 ( .A(y[677]), .B(x[128]), .Z(n3196) );
  XNOR U3742 ( .A(n3197), .B(n3196), .Z(n3225) );
  XOR U3743 ( .A(n3226), .B(n3225), .Z(n3221) );
  ANDN U3744 ( .B(y[675]), .A(n153), .Z(n3219) );
  ANDN U3745 ( .B(y[676]), .A(n152), .Z(n3234) );
  ANDN U3746 ( .B(y[673]), .A(n155), .Z(n3229) );
  XOR U3747 ( .A(o[37]), .B(n3229), .Z(n3232) );
  ANDN U3748 ( .B(y[674]), .A(n154), .Z(n3233) );
  XNOR U3749 ( .A(n3232), .B(n3233), .Z(n3235) );
  XNOR U3750 ( .A(n3234), .B(n3235), .Z(n3220) );
  XNOR U3751 ( .A(n3219), .B(n3220), .Z(n3222) );
  XNOR U3752 ( .A(n3221), .B(n3222), .Z(n3216) );
  ANDN U3753 ( .B(y[676]), .A(n155), .Z(n3338) );
  NAND U3754 ( .A(n3852), .B(n3338), .Z(n3201) );
  OR U3755 ( .A(n3199), .B(n3198), .Z(n3200) );
  NAND U3756 ( .A(n3201), .B(n3200), .Z(n3214) );
  NAND U3757 ( .A(n3202), .B(n3219), .Z(n3206) );
  NANDN U3758 ( .A(n3204), .B(n3203), .Z(n3205) );
  NAND U3759 ( .A(n3206), .B(n3205), .Z(n3213) );
  XNOR U3760 ( .A(n3214), .B(n3213), .Z(n3215) );
  XNOR U3761 ( .A(n3216), .B(n3215), .Z(n3210) );
  XOR U3762 ( .A(n3209), .B(n3210), .Z(N102) );
  NANDN U3763 ( .A(n3208), .B(n3207), .Z(n3212) );
  NANDN U3764 ( .A(n3210), .B(n3209), .Z(n3211) );
  NAND U3765 ( .A(n3212), .B(n3211), .Z(n3238) );
  OR U3766 ( .A(n3214), .B(n3213), .Z(n3218) );
  OR U3767 ( .A(n3216), .B(n3215), .Z(n3217) );
  AND U3768 ( .A(n3218), .B(n3217), .Z(n3239) );
  XNOR U3769 ( .A(n3238), .B(n3239), .Z(n3240) );
  OR U3770 ( .A(n3220), .B(n3219), .Z(n3224) );
  OR U3771 ( .A(n3222), .B(n3221), .Z(n3223) );
  AND U3772 ( .A(n3224), .B(n3223), .Z(n3244) );
  NAND U3773 ( .A(x[133]), .B(y[677]), .Z(n3602) );
  NANDN U3774 ( .A(n3602), .B(n3852), .Z(n3228) );
  OR U3775 ( .A(n3226), .B(n3225), .Z(n3227) );
  NAND U3776 ( .A(n3228), .B(n3227), .Z(n3266) );
  NAND U3777 ( .A(n3229), .B(o[37]), .Z(n3256) );
  AND U3778 ( .A(x[134]), .B(y[672]), .Z(n3231) );
  AND U3779 ( .A(x[128]), .B(y[678]), .Z(n3230) );
  XNOR U3780 ( .A(n3231), .B(n3230), .Z(n3255) );
  XOR U3781 ( .A(n3256), .B(n3255), .Z(n3265) );
  XNOR U3782 ( .A(n3266), .B(n3265), .Z(n3268) );
  AND U3783 ( .A(y[677]), .B(x[129]), .Z(n3536) );
  NAND U3784 ( .A(x[133]), .B(y[673]), .Z(n3259) );
  XNOR U3785 ( .A(n3259), .B(o[38]), .Z(n3260) );
  XNOR U3786 ( .A(n3536), .B(n3260), .Z(n3262) );
  AND U3787 ( .A(y[674]), .B(x[132]), .Z(n3261) );
  XOR U3788 ( .A(n3262), .B(n3261), .Z(n3251) );
  AND U3789 ( .A(y[676]), .B(x[130]), .Z(n3585) );
  XNOR U3790 ( .A(n3250), .B(n3585), .Z(n3252) );
  XOR U3791 ( .A(n3251), .B(n3252), .Z(n3267) );
  XNOR U3792 ( .A(n3268), .B(n3267), .Z(n3245) );
  XOR U3793 ( .A(n3244), .B(n3245), .Z(n3246) );
  OR U3794 ( .A(n3233), .B(n3232), .Z(n3237) );
  OR U3795 ( .A(n3235), .B(n3234), .Z(n3236) );
  AND U3796 ( .A(n3237), .B(n3236), .Z(n3247) );
  XOR U3797 ( .A(n3240), .B(n3241), .Z(N103) );
  NANDN U3798 ( .A(n3239), .B(n3238), .Z(n3243) );
  NANDN U3799 ( .A(n3241), .B(n3240), .Z(n3242) );
  NAND U3800 ( .A(n3243), .B(n3242), .Z(n3300) );
  OR U3801 ( .A(n3245), .B(n3244), .Z(n3249) );
  NANDN U3802 ( .A(n3247), .B(n3246), .Z(n3248) );
  AND U3803 ( .A(n3249), .B(n3248), .Z(n3301) );
  XNOR U3804 ( .A(n3300), .B(n3301), .Z(n3302) );
  OR U3805 ( .A(n3250), .B(n3585), .Z(n3254) );
  NANDN U3806 ( .A(n3252), .B(n3251), .Z(n3253) );
  NAND U3807 ( .A(n3254), .B(n3253), .Z(n3297) );
  AND U3808 ( .A(y[678]), .B(x[134]), .Z(n3524) );
  NAND U3809 ( .A(n3852), .B(n3524), .Z(n3258) );
  OR U3810 ( .A(n3256), .B(n3255), .Z(n3257) );
  AND U3811 ( .A(n3258), .B(n3257), .Z(n3295) );
  ANDN U3812 ( .B(y[674]), .A(n156), .Z(n3433) );
  AND U3813 ( .A(y[678]), .B(x[129]), .Z(n3652) );
  NAND U3814 ( .A(x[134]), .B(y[673]), .Z(n3283) );
  XNOR U3815 ( .A(o[39]), .B(n3283), .Z(n3284) );
  XNOR U3816 ( .A(n3652), .B(n3284), .Z(n3285) );
  XNOR U3817 ( .A(n3433), .B(n3285), .Z(n3294) );
  XOR U3818 ( .A(n3295), .B(n3294), .Z(n3296) );
  XNOR U3819 ( .A(n3297), .B(n3296), .Z(n3306) );
  ANDN U3820 ( .B(y[677]), .A(n153), .Z(n3730) );
  ANDN U3821 ( .B(y[675]), .A(n155), .Z(n3455) );
  ANDN U3822 ( .B(y[676]), .A(n154), .Z(n3279) );
  XNOR U3823 ( .A(n3455), .B(n3279), .Z(n3280) );
  XOR U3824 ( .A(n3730), .B(n3280), .Z(n3288) );
  NAND U3825 ( .A(x[128]), .B(y[679]), .Z(n3275) );
  ANDN U3826 ( .B(o[38]), .A(n3259), .Z(n3274) );
  NAND U3827 ( .A(y[672]), .B(x[135]), .Z(n3273) );
  XOR U3828 ( .A(n3274), .B(n3273), .Z(n3276) );
  XNOR U3829 ( .A(n3275), .B(n3276), .Z(n3289) );
  XNOR U3830 ( .A(n3288), .B(n3289), .Z(n3291) );
  NAND U3831 ( .A(n3536), .B(n3260), .Z(n3264) );
  NANDN U3832 ( .A(n3262), .B(n3261), .Z(n3263) );
  AND U3833 ( .A(n3264), .B(n3263), .Z(n3290) );
  XOR U3834 ( .A(n3291), .B(n3290), .Z(n3307) );
  XOR U3835 ( .A(n3306), .B(n3307), .Z(n3309) );
  OR U3836 ( .A(n3266), .B(n3265), .Z(n3270) );
  OR U3837 ( .A(n3268), .B(n3267), .Z(n3269) );
  AND U3838 ( .A(n3270), .B(n3269), .Z(n3308) );
  XOR U3839 ( .A(n3309), .B(n3308), .Z(n3303) );
  XNOR U3840 ( .A(n3302), .B(n3303), .Z(N104) );
  AND U3841 ( .A(x[136]), .B(y[672]), .Z(n3272) );
  NAND U3842 ( .A(x[128]), .B(y[680]), .Z(n3271) );
  XOR U3843 ( .A(n3272), .B(n3271), .Z(n3325) );
  NAND U3844 ( .A(x[135]), .B(y[673]), .Z(n3328) );
  XNOR U3845 ( .A(n3328), .B(o[40]), .Z(n3324) );
  XOR U3846 ( .A(n3325), .B(n3324), .Z(n3319) );
  NANDN U3847 ( .A(n3274), .B(n3273), .Z(n3278) );
  NANDN U3848 ( .A(n3276), .B(n3275), .Z(n3277) );
  NAND U3849 ( .A(n3278), .B(n3277), .Z(n3318) );
  XOR U3850 ( .A(n3319), .B(n3318), .Z(n3320) );
  OR U3851 ( .A(n3279), .B(n3455), .Z(n3282) );
  OR U3852 ( .A(n3280), .B(n3730), .Z(n3281) );
  NAND U3853 ( .A(n3282), .B(n3281), .Z(n3321) );
  XNOR U3854 ( .A(n3320), .B(n3321), .Z(n3354) );
  ANDN U3855 ( .B(y[674]), .A(n157), .Z(n3339) );
  XNOR U3856 ( .A(n3338), .B(n3339), .Z(n3340) );
  NOR U3857 ( .A(n153), .B(n146), .Z(n3868) );
  XNOR U3858 ( .A(n3340), .B(n3868), .Z(n3341) );
  ANDN U3859 ( .B(y[677]), .A(n154), .Z(n4144) );
  XNOR U3860 ( .A(n3341), .B(n4144), .Z(n3343) );
  NANDN U3861 ( .A(n3283), .B(o[39]), .Z(n3335) );
  AND U3862 ( .A(x[133]), .B(y[675]), .Z(n3931) );
  AND U3863 ( .A(y[679]), .B(x[129]), .Z(n3847) );
  XNOR U3864 ( .A(n3931), .B(n3847), .Z(n3334) );
  XOR U3865 ( .A(n3335), .B(n3334), .Z(n3342) );
  XNOR U3866 ( .A(n3343), .B(n3342), .Z(n3312) );
  NAND U3867 ( .A(n3652), .B(n3284), .Z(n3287) );
  NANDN U3868 ( .A(n3285), .B(n3433), .Z(n3286) );
  AND U3869 ( .A(n3287), .B(n3286), .Z(n3313) );
  XOR U3870 ( .A(n3312), .B(n3313), .Z(n3315) );
  OR U3871 ( .A(n3289), .B(n3288), .Z(n3293) );
  OR U3872 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3873 ( .A(n3293), .B(n3292), .Z(n3314) );
  XOR U3874 ( .A(n3315), .B(n3314), .Z(n3352) );
  NANDN U3875 ( .A(n3295), .B(n3294), .Z(n3299) );
  OR U3876 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3877 ( .A(n3299), .B(n3298), .Z(n3353) );
  XNOR U3878 ( .A(n3352), .B(n3353), .Z(n3355) );
  XNOR U3879 ( .A(n3354), .B(n3355), .Z(n3349) );
  NANDN U3880 ( .A(n3301), .B(n3300), .Z(n3305) );
  NAND U3881 ( .A(n3303), .B(n3302), .Z(n3304) );
  NAND U3882 ( .A(n3305), .B(n3304), .Z(n3346) );
  NANDN U3883 ( .A(n3307), .B(n3306), .Z(n3311) );
  OR U3884 ( .A(n3309), .B(n3308), .Z(n3310) );
  AND U3885 ( .A(n3311), .B(n3310), .Z(n3347) );
  XNOR U3886 ( .A(n3346), .B(n3347), .Z(n3348) );
  XOR U3887 ( .A(n3349), .B(n3348), .Z(N105) );
  NANDN U3888 ( .A(n3313), .B(n3312), .Z(n3317) );
  OR U3889 ( .A(n3315), .B(n3314), .Z(n3316) );
  NAND U3890 ( .A(n3317), .B(n3316), .Z(n3365) );
  OR U3891 ( .A(n3319), .B(n3318), .Z(n3323) );
  NANDN U3892 ( .A(n3321), .B(n3320), .Z(n3322) );
  NAND U3893 ( .A(n3323), .B(n3322), .Z(n3364) );
  XOR U3894 ( .A(n3365), .B(n3364), .Z(n3366) );
  AND U3895 ( .A(y[680]), .B(x[136]), .Z(n3865) );
  NAND U3896 ( .A(n3852), .B(n3865), .Z(n3327) );
  NANDN U3897 ( .A(n3325), .B(n3324), .Z(n3326) );
  NAND U3898 ( .A(n3327), .B(n3326), .Z(n3373) );
  NANDN U3899 ( .A(n3328), .B(o[40]), .Z(n3404) );
  AND U3900 ( .A(y[676]), .B(x[133]), .Z(n3329) );
  AND U3901 ( .A(y[674]), .B(x[135]), .Z(n3725) );
  XNOR U3902 ( .A(n3329), .B(n3725), .Z(n3403) );
  XOR U3903 ( .A(n3404), .B(n3403), .Z(n3371) );
  AND U3904 ( .A(x[137]), .B(y[672]), .Z(n3331) );
  NAND U3905 ( .A(x[128]), .B(y[681]), .Z(n3330) );
  XOR U3906 ( .A(n3331), .B(n3330), .Z(n3398) );
  NAND U3907 ( .A(x[136]), .B(y[673]), .Z(n3392) );
  XOR U3908 ( .A(n3392), .B(o[41]), .Z(n3397) );
  XNOR U3909 ( .A(n3398), .B(n3397), .Z(n3370) );
  XNOR U3910 ( .A(n3371), .B(n3370), .Z(n3372) );
  XNOR U3911 ( .A(n3373), .B(n3372), .Z(n3382) );
  NAND U3912 ( .A(x[132]), .B(y[677]), .Z(n3857) );
  AND U3913 ( .A(x[134]), .B(y[675]), .Z(n3333) );
  NAND U3914 ( .A(x[129]), .B(y[680]), .Z(n3332) );
  XNOR U3915 ( .A(n3333), .B(n3332), .Z(n3394) );
  XNOR U3916 ( .A(n3857), .B(n3394), .Z(n3376) );
  ANDN U3917 ( .B(y[679]), .A(n153), .Z(n4045) );
  NAND U3918 ( .A(y[678]), .B(x[131]), .Z(n3746) );
  XOR U3919 ( .A(n4045), .B(n3746), .Z(n3377) );
  XNOR U3920 ( .A(n3376), .B(n3377), .Z(n3380) );
  NAND U3921 ( .A(x[129]), .B(y[675]), .Z(n3393) );
  AND U3922 ( .A(y[679]), .B(x[133]), .Z(n3526) );
  NANDN U3923 ( .A(n3393), .B(n3526), .Z(n3337) );
  OR U3924 ( .A(n3335), .B(n3334), .Z(n3336) );
  AND U3925 ( .A(n3337), .B(n3336), .Z(n3381) );
  XOR U3926 ( .A(n3380), .B(n3381), .Z(n3383) );
  XNOR U3927 ( .A(n3382), .B(n3383), .Z(n3388) );
  OR U3928 ( .A(n3341), .B(n4144), .Z(n3345) );
  OR U3929 ( .A(n3343), .B(n3342), .Z(n3344) );
  AND U3930 ( .A(n3345), .B(n3344), .Z(n3386) );
  XNOR U3931 ( .A(n3387), .B(n3386), .Z(n3389) );
  XOR U3932 ( .A(n3388), .B(n3389), .Z(n3367) );
  XOR U3933 ( .A(n3366), .B(n3367), .Z(n3361) );
  NANDN U3934 ( .A(n3347), .B(n3346), .Z(n3351) );
  NANDN U3935 ( .A(n3349), .B(n3348), .Z(n3350) );
  NAND U3936 ( .A(n3351), .B(n3350), .Z(n3358) );
  OR U3937 ( .A(n3353), .B(n3352), .Z(n3357) );
  OR U3938 ( .A(n3355), .B(n3354), .Z(n3356) );
  AND U3939 ( .A(n3357), .B(n3356), .Z(n3359) );
  XNOR U3940 ( .A(n3358), .B(n3359), .Z(n3360) );
  XOR U3941 ( .A(n3361), .B(n3360), .Z(N106) );
  NANDN U3942 ( .A(n3359), .B(n3358), .Z(n3363) );
  NANDN U3943 ( .A(n3361), .B(n3360), .Z(n3362) );
  NAND U3944 ( .A(n3363), .B(n3362), .Z(n3407) );
  OR U3945 ( .A(n3365), .B(n3364), .Z(n3369) );
  NANDN U3946 ( .A(n3367), .B(n3366), .Z(n3368) );
  AND U3947 ( .A(n3369), .B(n3368), .Z(n3408) );
  XNOR U3948 ( .A(n3407), .B(n3408), .Z(n3409) );
  NANDN U3949 ( .A(n3371), .B(n3370), .Z(n3375) );
  NANDN U3950 ( .A(n3373), .B(n3372), .Z(n3374) );
  NAND U3951 ( .A(n3375), .B(n3374), .Z(n3467) );
  NANDN U3952 ( .A(n4045), .B(n3746), .Z(n3379) );
  OR U3953 ( .A(n3377), .B(n3376), .Z(n3378) );
  NAND U3954 ( .A(n3379), .B(n3378), .Z(n3466) );
  XOR U3955 ( .A(n3467), .B(n3466), .Z(n3468) );
  NANDN U3956 ( .A(n3381), .B(n3380), .Z(n3385) );
  OR U3957 ( .A(n3383), .B(n3382), .Z(n3384) );
  AND U3958 ( .A(n3385), .B(n3384), .Z(n3469) );
  XNOR U3959 ( .A(n3468), .B(n3469), .Z(n3416) );
  OR U3960 ( .A(n3387), .B(n3386), .Z(n3391) );
  NANDN U3961 ( .A(n3389), .B(n3388), .Z(n3390) );
  AND U3962 ( .A(n3391), .B(n3390), .Z(n3413) );
  ANDN U3963 ( .B(y[682]), .A(n151), .Z(n3452) );
  NANDN U3964 ( .A(n3392), .B(o[41]), .Z(n3449) );
  ANDN U3965 ( .B(y[672]), .A(n161), .Z(n3450) );
  XNOR U3966 ( .A(n3452), .B(n3451), .Z(n3440) );
  ANDN U3967 ( .B(y[679]), .A(n154), .Z(n4407) );
  IV U3968 ( .A(y[680]), .Z(n4926) );
  NANDN U3969 ( .A(n4926), .B(x[130]), .Z(n3429) );
  XNOR U3970 ( .A(n4407), .B(n3429), .Z(n3430) );
  NAND U3971 ( .A(y[681]), .B(x[129]), .Z(n4365) );
  ANDN U3972 ( .B(y[680]), .A(n157), .Z(n3717) );
  NANDN U3973 ( .A(n3393), .B(n3717), .Z(n3396) );
  NANDN U3974 ( .A(n3857), .B(n3394), .Z(n3395) );
  AND U3975 ( .A(n3396), .B(n3395), .Z(n3439) );
  XOR U3976 ( .A(n3438), .B(n3439), .Z(n3441) );
  XNOR U3977 ( .A(n3440), .B(n3441), .Z(n3460) );
  AND U3978 ( .A(y[681]), .B(x[137]), .Z(n4023) );
  NAND U3979 ( .A(n3852), .B(n4023), .Z(n3400) );
  OR U3980 ( .A(n3398), .B(n3397), .Z(n3399) );
  NAND U3981 ( .A(n3400), .B(n3399), .Z(n3461) );
  XNOR U3982 ( .A(n3460), .B(n3461), .Z(n3463) );
  AND U3983 ( .A(y[674]), .B(x[136]), .Z(n3517) );
  XOR U3984 ( .A(n3517), .B(n3602), .Z(n3435) );
  NAND U3985 ( .A(x[137]), .B(y[673]), .Z(n3444) );
  XOR U3986 ( .A(o[42]), .B(n3444), .Z(n3434) );
  XOR U3987 ( .A(n3435), .B(n3434), .Z(n3419) );
  AND U3988 ( .A(y[676]), .B(x[134]), .Z(n3669) );
  AND U3989 ( .A(x[132]), .B(y[678]), .Z(n3402) );
  NAND U3990 ( .A(x[135]), .B(y[675]), .Z(n3401) );
  XOR U3991 ( .A(n3402), .B(n3401), .Z(n3457) );
  XNOR U3992 ( .A(n3669), .B(n3457), .Z(n3420) );
  XNOR U3993 ( .A(n3419), .B(n3420), .Z(n3422) );
  ANDN U3994 ( .B(y[676]), .A(n158), .Z(n3518) );
  NAND U3995 ( .A(n3433), .B(n3518), .Z(n3406) );
  OR U3996 ( .A(n3404), .B(n3403), .Z(n3405) );
  NAND U3997 ( .A(n3406), .B(n3405), .Z(n3421) );
  XNOR U3998 ( .A(n3422), .B(n3421), .Z(n3462) );
  XNOR U3999 ( .A(n3463), .B(n3462), .Z(n3414) );
  XOR U4000 ( .A(n3413), .B(n3414), .Z(n3415) );
  XOR U4001 ( .A(n3416), .B(n3415), .Z(n3410) );
  XOR U4002 ( .A(n3409), .B(n3410), .Z(N107) );
  NANDN U4003 ( .A(n3408), .B(n3407), .Z(n3412) );
  NANDN U4004 ( .A(n3410), .B(n3409), .Z(n3411) );
  NAND U4005 ( .A(n3412), .B(n3411), .Z(n3472) );
  OR U4006 ( .A(n3414), .B(n3413), .Z(n3418) );
  NANDN U4007 ( .A(n3416), .B(n3415), .Z(n3417) );
  AND U4008 ( .A(n3418), .B(n3417), .Z(n3473) );
  XNOR U4009 ( .A(n3472), .B(n3473), .Z(n3474) );
  OR U4010 ( .A(n3420), .B(n3419), .Z(n3424) );
  OR U4011 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U4012 ( .A(n3424), .B(n3423), .Z(n3487) );
  AND U4013 ( .A(x[136]), .B(y[675]), .Z(n3426) );
  NAND U4014 ( .A(x[137]), .B(y[674]), .Z(n3425) );
  XNOR U4015 ( .A(n3426), .B(n3425), .Z(n3519) );
  XNOR U4016 ( .A(n3518), .B(n3519), .Z(n3498) );
  ANDN U4017 ( .B(y[680]), .A(n154), .Z(n4534) );
  NAND U4018 ( .A(x[132]), .B(y[679]), .Z(n3533) );
  AND U4019 ( .A(x[133]), .B(y[678]), .Z(n3428) );
  NAND U4020 ( .A(x[130]), .B(y[681]), .Z(n3427) );
  XOR U4021 ( .A(n3428), .B(n3427), .Z(n3532) );
  XNOR U4022 ( .A(n3533), .B(n3532), .Z(n3496) );
  XNOR U4023 ( .A(n4534), .B(n3496), .Z(n3497) );
  XNOR U4024 ( .A(n3498), .B(n3497), .Z(n3510) );
  NANDN U4025 ( .A(n4407), .B(n3429), .Z(n3432) );
  NAND U4026 ( .A(n3430), .B(n4365), .Z(n3431) );
  NAND U4027 ( .A(n3432), .B(n3431), .Z(n3507) );
  ANDN U4028 ( .B(y[677]), .A(n159), .Z(n4278) );
  NAND U4029 ( .A(n4278), .B(n3433), .Z(n3437) );
  OR U4030 ( .A(n3435), .B(n3434), .Z(n3436) );
  NAND U4031 ( .A(n3437), .B(n3436), .Z(n3508) );
  XNOR U4032 ( .A(n3510), .B(n3509), .Z(n3485) );
  NANDN U4033 ( .A(n3439), .B(n3438), .Z(n3443) );
  NANDN U4034 ( .A(n3441), .B(n3440), .Z(n3442) );
  NAND U4035 ( .A(n3443), .B(n3442), .Z(n3493) );
  NANDN U4036 ( .A(n3444), .B(o[42]), .Z(n3514) );
  AND U4037 ( .A(x[139]), .B(y[672]), .Z(n3446) );
  NAND U4038 ( .A(x[128]), .B(y[683]), .Z(n3445) );
  XNOR U4039 ( .A(n3446), .B(n3445), .Z(n3513) );
  AND U4040 ( .A(y[677]), .B(x[134]), .Z(n3448) );
  NAND U4041 ( .A(x[129]), .B(y[682]), .Z(n3447) );
  XOR U4042 ( .A(n3448), .B(n3447), .Z(n3538) );
  NAND U4043 ( .A(x[138]), .B(y[673]), .Z(n3522) );
  XOR U4044 ( .A(o[43]), .B(n3522), .Z(n3537) );
  XOR U4045 ( .A(n3538), .B(n3537), .Z(n3501) );
  NANDN U4046 ( .A(n3450), .B(n3449), .Z(n3454) );
  OR U4047 ( .A(n3452), .B(n3451), .Z(n3453) );
  NAND U4048 ( .A(n3454), .B(n3453), .Z(n3504) );
  XOR U4049 ( .A(n3503), .B(n3504), .Z(n3490) );
  AND U4050 ( .A(y[678]), .B(x[135]), .Z(n3456) );
  NAND U4051 ( .A(n3456), .B(n3455), .Z(n3459) );
  NANDN U4052 ( .A(n3457), .B(n3669), .Z(n3458) );
  NAND U4053 ( .A(n3459), .B(n3458), .Z(n3491) );
  XOR U4054 ( .A(n3493), .B(n3492), .Z(n3484) );
  XOR U4055 ( .A(n3485), .B(n3484), .Z(n3486) );
  XOR U4056 ( .A(n3487), .B(n3486), .Z(n3478) );
  OR U4057 ( .A(n3461), .B(n3460), .Z(n3465) );
  OR U4058 ( .A(n3463), .B(n3462), .Z(n3464) );
  AND U4059 ( .A(n3465), .B(n3464), .Z(n3479) );
  XNOR U4060 ( .A(n3478), .B(n3479), .Z(n3481) );
  OR U4061 ( .A(n3467), .B(n3466), .Z(n3471) );
  NANDN U4062 ( .A(n3469), .B(n3468), .Z(n3470) );
  NAND U4063 ( .A(n3471), .B(n3470), .Z(n3480) );
  XOR U4064 ( .A(n3481), .B(n3480), .Z(n3475) );
  XNOR U4065 ( .A(n3474), .B(n3475), .Z(N108) );
  NANDN U4066 ( .A(n3473), .B(n3472), .Z(n3477) );
  NAND U4067 ( .A(n3475), .B(n3474), .Z(n3476) );
  NAND U4068 ( .A(n3477), .B(n3476), .Z(n3541) );
  OR U4069 ( .A(n3479), .B(n3478), .Z(n3483) );
  OR U4070 ( .A(n3481), .B(n3480), .Z(n3482) );
  AND U4071 ( .A(n3483), .B(n3482), .Z(n3542) );
  XNOR U4072 ( .A(n3541), .B(n3542), .Z(n3543) );
  NANDN U4073 ( .A(n3485), .B(n3484), .Z(n3489) );
  OR U4074 ( .A(n3487), .B(n3486), .Z(n3488) );
  NAND U4075 ( .A(n3489), .B(n3488), .Z(n3548) );
  NANDN U4076 ( .A(n3491), .B(n3490), .Z(n3495) );
  NANDN U4077 ( .A(n3493), .B(n3492), .Z(n3494) );
  NAND U4078 ( .A(n3495), .B(n3494), .Z(n3616) );
  NANDN U4079 ( .A(n3496), .B(n4534), .Z(n3500) );
  NANDN U4080 ( .A(n3498), .B(n3497), .Z(n3499) );
  NAND U4081 ( .A(n3500), .B(n3499), .Z(n3614) );
  NAND U4082 ( .A(n3502), .B(n3501), .Z(n3506) );
  NANDN U4083 ( .A(n3504), .B(n3503), .Z(n3505) );
  AND U4084 ( .A(n3506), .B(n3505), .Z(n3613) );
  XNOR U4085 ( .A(n3616), .B(n3615), .Z(n3547) );
  XNOR U4086 ( .A(n3548), .B(n3547), .Z(n3550) );
  NANDN U4087 ( .A(n3508), .B(n3507), .Z(n3512) );
  NANDN U4088 ( .A(n3510), .B(n3509), .Z(n3511) );
  NAND U4089 ( .A(n3512), .B(n3511), .Z(n3609) );
  ANDN U4090 ( .B(y[683]), .A(n162), .Z(n4656) );
  NAND U4091 ( .A(n3852), .B(n4656), .Z(n3516) );
  NANDN U4092 ( .A(n3514), .B(n3513), .Z(n3515) );
  NAND U4093 ( .A(n3516), .B(n3515), .Z(n3555) );
  NAND U4094 ( .A(x[137]), .B(y[675]), .Z(n4233) );
  NANDN U4095 ( .A(n4233), .B(n3517), .Z(n3521) );
  NAND U4096 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U4097 ( .A(n3521), .B(n3520), .Z(n3553) );
  NANDN U4098 ( .A(n3522), .B(o[43]), .Z(n3570) );
  NAND U4099 ( .A(x[129]), .B(y[683]), .Z(n3523) );
  XNOR U4100 ( .A(n3524), .B(n3523), .Z(n3569) );
  XOR U4101 ( .A(n3553), .B(n3554), .Z(n3556) );
  NAND U4102 ( .A(x[135]), .B(y[677]), .Z(n3525) );
  XOR U4103 ( .A(n3526), .B(n3525), .Z(n3604) );
  AND U4104 ( .A(y[674]), .B(x[138]), .Z(n3527) );
  XOR U4105 ( .A(n3527), .B(n4233), .Z(n3562) );
  NAND U4106 ( .A(x[132]), .B(y[680]), .Z(n3561) );
  XNOR U4107 ( .A(n3562), .B(n3561), .Z(n3603) );
  XOR U4108 ( .A(n3604), .B(n3603), .Z(n3597) );
  AND U4109 ( .A(x[140]), .B(y[672]), .Z(n3529) );
  NAND U4110 ( .A(x[128]), .B(y[684]), .Z(n3528) );
  XOR U4111 ( .A(n3529), .B(n3528), .Z(n3574) );
  NAND U4112 ( .A(x[139]), .B(y[673]), .Z(n3592) );
  XOR U4113 ( .A(o[44]), .B(n3592), .Z(n3573) );
  XOR U4114 ( .A(n3574), .B(n3573), .Z(n3595) );
  AND U4115 ( .A(y[676]), .B(x[136]), .Z(n3531) );
  NAND U4116 ( .A(x[130]), .B(y[682]), .Z(n3530) );
  XOR U4117 ( .A(n3531), .B(n3530), .Z(n3587) );
  NAND U4118 ( .A(y[681]), .B(x[131]), .Z(n3586) );
  XNOR U4119 ( .A(n3587), .B(n3586), .Z(n3596) );
  XOR U4120 ( .A(n3595), .B(n3596), .Z(n3598) );
  ANDN U4121 ( .B(y[681]), .A(n156), .Z(n3747) );
  NAND U4122 ( .A(n3868), .B(n3747), .Z(n3535) );
  OR U4123 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U4124 ( .A(n3535), .B(n3534), .Z(n3580) );
  AND U4125 ( .A(y[682]), .B(x[134]), .Z(n3862) );
  NAND U4126 ( .A(n3862), .B(n3536), .Z(n3540) );
  OR U4127 ( .A(n3538), .B(n3537), .Z(n3539) );
  NAND U4128 ( .A(n3540), .B(n3539), .Z(n3579) );
  XOR U4129 ( .A(n3580), .B(n3579), .Z(n3582) );
  XNOR U4130 ( .A(n3581), .B(n3582), .Z(n3608) );
  XOR U4131 ( .A(n3607), .B(n3608), .Z(n3610) );
  XOR U4132 ( .A(n3609), .B(n3610), .Z(n3549) );
  XNOR U4133 ( .A(n3550), .B(n3549), .Z(n3544) );
  XOR U4134 ( .A(n3543), .B(n3544), .Z(N109) );
  NANDN U4135 ( .A(n3542), .B(n3541), .Z(n3546) );
  NANDN U4136 ( .A(n3544), .B(n3543), .Z(n3545) );
  NAND U4137 ( .A(n3546), .B(n3545), .Z(n3684) );
  OR U4138 ( .A(n3548), .B(n3547), .Z(n3552) );
  OR U4139 ( .A(n3550), .B(n3549), .Z(n3551) );
  AND U4140 ( .A(n3552), .B(n3551), .Z(n3685) );
  XNOR U4141 ( .A(n3684), .B(n3685), .Z(n3686) );
  NANDN U4142 ( .A(n3554), .B(n3553), .Z(n3558) );
  NANDN U4143 ( .A(n3556), .B(n3555), .Z(n3557) );
  NAND U4144 ( .A(n3558), .B(n3557), .Z(n3633) );
  AND U4145 ( .A(y[674]), .B(x[137]), .Z(n3560) );
  AND U4146 ( .A(y[675]), .B(x[138]), .Z(n3559) );
  NAND U4147 ( .A(n3560), .B(n3559), .Z(n3564) );
  OR U4148 ( .A(n3562), .B(n3561), .Z(n3563) );
  NAND U4149 ( .A(n3564), .B(n3563), .Z(n3681) );
  AND U4150 ( .A(x[141]), .B(y[672]), .Z(n3566) );
  NAND U4151 ( .A(x[128]), .B(y[685]), .Z(n3565) );
  XOR U4152 ( .A(n3566), .B(n3565), .Z(n3666) );
  NAND U4153 ( .A(x[140]), .B(y[673]), .Z(n3675) );
  XOR U4154 ( .A(o[45]), .B(n3675), .Z(n3665) );
  XOR U4155 ( .A(n3666), .B(n3665), .Z(n3679) );
  AND U4156 ( .A(x[131]), .B(y[682]), .Z(n3568) );
  NAND U4157 ( .A(x[133]), .B(y[680]), .Z(n3567) );
  XOR U4158 ( .A(n3568), .B(n3567), .Z(n3662) );
  NAND U4159 ( .A(y[681]), .B(x[132]), .Z(n3661) );
  XOR U4160 ( .A(n3662), .B(n3661), .Z(n3678) );
  XNOR U4161 ( .A(n3681), .B(n3680), .Z(n3632) );
  ANDN U4162 ( .B(y[683]), .A(n157), .Z(n4053) );
  NAND U4163 ( .A(n3652), .B(n4053), .Z(n3572) );
  NANDN U4164 ( .A(n3570), .B(n3569), .Z(n3571) );
  AND U4165 ( .A(n3572), .B(n3571), .Z(n3640) );
  ANDN U4166 ( .B(y[684]), .A(n163), .Z(n4867) );
  NAND U4167 ( .A(n3852), .B(n4867), .Z(n3576) );
  OR U4168 ( .A(n3574), .B(n3573), .Z(n3575) );
  NAND U4169 ( .A(n3576), .B(n3575), .Z(n3637) );
  AND U4170 ( .A(y[674]), .B(x[139]), .Z(n3578) );
  NAND U4171 ( .A(x[138]), .B(y[675]), .Z(n3577) );
  XNOR U4172 ( .A(n3578), .B(n3577), .Z(n3658) );
  XNOR U4173 ( .A(n4278), .B(n3658), .Z(n3638) );
  XOR U4174 ( .A(n3640), .B(n3639), .Z(n3631) );
  XOR U4175 ( .A(n3632), .B(n3631), .Z(n3634) );
  OR U4176 ( .A(n3580), .B(n3579), .Z(n3584) );
  NAND U4177 ( .A(n3582), .B(n3581), .Z(n3583) );
  AND U4178 ( .A(n3584), .B(n3583), .Z(n3625) );
  AND U4179 ( .A(y[682]), .B(x[136]), .Z(n4010) );
  NAND U4180 ( .A(n4010), .B(n3585), .Z(n3589) );
  OR U4181 ( .A(n3587), .B(n3586), .Z(n3588) );
  NAND U4182 ( .A(n3589), .B(n3588), .Z(n3646) );
  AND U4183 ( .A(y[679]), .B(x[134]), .Z(n3591) );
  NAND U4184 ( .A(x[137]), .B(y[676]), .Z(n3590) );
  XOR U4185 ( .A(n3591), .B(n3590), .Z(n3671) );
  NAND U4186 ( .A(x[130]), .B(y[683]), .Z(n3670) );
  XOR U4187 ( .A(n3671), .B(n3670), .Z(n3644) );
  NANDN U4188 ( .A(n3592), .B(o[44]), .Z(n3655) );
  AND U4189 ( .A(y[684]), .B(x[129]), .Z(n3594) );
  NAND U4190 ( .A(x[135]), .B(y[678]), .Z(n3593) );
  XNOR U4191 ( .A(n3594), .B(n3593), .Z(n3654) );
  XNOR U4192 ( .A(n3646), .B(n3645), .Z(n3622) );
  NANDN U4193 ( .A(n3596), .B(n3595), .Z(n3600) );
  NANDN U4194 ( .A(n3598), .B(n3597), .Z(n3599) );
  AND U4195 ( .A(n3600), .B(n3599), .Z(n3620) );
  AND U4196 ( .A(y[679]), .B(x[135]), .Z(n3601) );
  NANDN U4197 ( .A(n3602), .B(n3601), .Z(n3606) );
  OR U4198 ( .A(n3604), .B(n3603), .Z(n3605) );
  AND U4199 ( .A(n3606), .B(n3605), .Z(n3619) );
  XNOR U4200 ( .A(n3620), .B(n3619), .Z(n3621) );
  XOR U4201 ( .A(n3622), .B(n3621), .Z(n3626) );
  XNOR U4202 ( .A(n3625), .B(n3626), .Z(n3628) );
  XNOR U4203 ( .A(n3627), .B(n3628), .Z(n3693) );
  NANDN U4204 ( .A(n3608), .B(n3607), .Z(n3612) );
  NANDN U4205 ( .A(n3610), .B(n3609), .Z(n3611) );
  NAND U4206 ( .A(n3612), .B(n3611), .Z(n3691) );
  NANDN U4207 ( .A(n3614), .B(n3613), .Z(n3618) );
  NAND U4208 ( .A(n3616), .B(n3615), .Z(n3617) );
  AND U4209 ( .A(n3618), .B(n3617), .Z(n3690) );
  XNOR U4210 ( .A(n3693), .B(n3692), .Z(n3687) );
  XOR U4211 ( .A(n3686), .B(n3687), .Z(N110) );
  OR U4212 ( .A(n3620), .B(n3619), .Z(n3624) );
  OR U4213 ( .A(n3622), .B(n3621), .Z(n3623) );
  NAND U4214 ( .A(n3624), .B(n3623), .Z(n3705) );
  OR U4215 ( .A(n3626), .B(n3625), .Z(n3630) );
  NANDN U4216 ( .A(n3628), .B(n3627), .Z(n3629) );
  AND U4217 ( .A(n3630), .B(n3629), .Z(n3702) );
  NANDN U4218 ( .A(n3632), .B(n3631), .Z(n3636) );
  NANDN U4219 ( .A(n3634), .B(n3633), .Z(n3635) );
  NAND U4220 ( .A(n3636), .B(n3635), .Z(n3782) );
  NANDN U4221 ( .A(n3638), .B(n3637), .Z(n3642) );
  OR U4222 ( .A(n3640), .B(n3639), .Z(n3641) );
  NAND U4223 ( .A(n3642), .B(n3641), .Z(n3710) );
  NAND U4224 ( .A(n3644), .B(n3643), .Z(n3648) );
  NAND U4225 ( .A(n3646), .B(n3645), .Z(n3647) );
  NAND U4226 ( .A(n3648), .B(n3647), .Z(n3708) );
  ANDN U4227 ( .B(y[682]), .A(n155), .Z(n3762) );
  AND U4228 ( .A(y[676]), .B(x[138]), .Z(n4412) );
  AND U4229 ( .A(y[677]), .B(x[137]), .Z(n4359) );
  NAND U4230 ( .A(x[130]), .B(y[684]), .Z(n3649) );
  XOR U4231 ( .A(n4359), .B(n3649), .Z(n3731) );
  XNOR U4232 ( .A(n4412), .B(n3731), .Z(n3761) );
  XOR U4233 ( .A(n3762), .B(n3761), .Z(n3764) );
  AND U4234 ( .A(y[683]), .B(x[131]), .Z(n3651) );
  NAND U4235 ( .A(x[136]), .B(y[678]), .Z(n3650) );
  XOR U4236 ( .A(n3651), .B(n3650), .Z(n3748) );
  XOR U4237 ( .A(n3747), .B(n3748), .Z(n3763) );
  AND U4238 ( .A(y[684]), .B(x[135]), .Z(n3653) );
  NAND U4239 ( .A(n3653), .B(n3652), .Z(n3657) );
  NANDN U4240 ( .A(n3655), .B(n3654), .Z(n3656) );
  NAND U4241 ( .A(n3657), .B(n3656), .Z(n3767) );
  NAND U4242 ( .A(x[138]), .B(y[674]), .Z(n4283) );
  NOR U4243 ( .A(n162), .B(n145), .Z(n3821) );
  NANDN U4244 ( .A(n4283), .B(n3821), .Z(n3660) );
  NAND U4245 ( .A(n3658), .B(n4278), .Z(n3659) );
  AND U4246 ( .A(n3660), .B(n3659), .Z(n3768) );
  XOR U4247 ( .A(n3770), .B(n3769), .Z(n3709) );
  XOR U4248 ( .A(n3710), .B(n3711), .Z(n3779) );
  ANDN U4249 ( .B(y[682]), .A(n156), .Z(n3842) );
  NAND U4250 ( .A(n4534), .B(n3842), .Z(n3664) );
  OR U4251 ( .A(n3662), .B(n3661), .Z(n3663) );
  NAND U4252 ( .A(n3664), .B(n3663), .Z(n3742) );
  IV U4253 ( .A(n3821), .Z(n3715) );
  IV U4254 ( .A(y[685]), .Z(n4890) );
  NANDN U4255 ( .A(n4890), .B(x[129]), .Z(n3714) );
  XNOR U4256 ( .A(n3715), .B(n3714), .Z(n3716) );
  XOR U4257 ( .A(n3717), .B(n3716), .Z(n3741) );
  AND U4258 ( .A(x[141]), .B(y[685]), .Z(n5244) );
  NAND U4259 ( .A(n3852), .B(n5244), .Z(n3668) );
  OR U4260 ( .A(n3666), .B(n3665), .Z(n3667) );
  AND U4261 ( .A(n3668), .B(n3667), .Z(n3740) );
  XNOR U4262 ( .A(n3741), .B(n3740), .Z(n3743) );
  XOR U4263 ( .A(n3742), .B(n3743), .Z(n3775) );
  AND U4264 ( .A(y[679]), .B(x[137]), .Z(n3827) );
  NAND U4265 ( .A(n3827), .B(n3669), .Z(n3673) );
  OR U4266 ( .A(n3671), .B(n3670), .Z(n3672) );
  AND U4267 ( .A(n3673), .B(n3672), .Z(n3737) );
  AND U4268 ( .A(y[674]), .B(x[140]), .Z(n4354) );
  NAND U4269 ( .A(x[135]), .B(y[679]), .Z(n3674) );
  XOR U4270 ( .A(n4354), .B(n3674), .Z(n3727) );
  NAND U4271 ( .A(x[141]), .B(y[673]), .Z(n3720) );
  XOR U4272 ( .A(o[46]), .B(n3720), .Z(n3726) );
  XOR U4273 ( .A(n3727), .B(n3726), .Z(n3735) );
  NANDN U4274 ( .A(n3675), .B(o[45]), .Z(n3752) );
  AND U4275 ( .A(y[686]), .B(x[128]), .Z(n3677) );
  NAND U4276 ( .A(x[142]), .B(y[672]), .Z(n3676) );
  XNOR U4277 ( .A(n3677), .B(n3676), .Z(n3751) );
  XOR U4278 ( .A(n3737), .B(n3736), .Z(n3773) );
  NAND U4279 ( .A(n3679), .B(n3678), .Z(n3683) );
  NAND U4280 ( .A(n3681), .B(n3680), .Z(n3682) );
  NAND U4281 ( .A(n3683), .B(n3682), .Z(n3774) );
  XOR U4282 ( .A(n3773), .B(n3774), .Z(n3776) );
  XNOR U4283 ( .A(n3775), .B(n3776), .Z(n3780) );
  XOR U4284 ( .A(n3782), .B(n3781), .Z(n3703) );
  XNOR U4285 ( .A(n3702), .B(n3703), .Z(n3704) );
  XOR U4286 ( .A(n3705), .B(n3704), .Z(n3698) );
  NANDN U4287 ( .A(n3685), .B(n3684), .Z(n3689) );
  NANDN U4288 ( .A(n3687), .B(n3686), .Z(n3688) );
  NAND U4289 ( .A(n3689), .B(n3688), .Z(n3696) );
  NANDN U4290 ( .A(n3691), .B(n3690), .Z(n3695) );
  NANDN U4291 ( .A(n3693), .B(n3692), .Z(n3694) );
  NAND U4292 ( .A(n3695), .B(n3694), .Z(n3697) );
  XNOR U4293 ( .A(n3696), .B(n3697), .Z(n3699) );
  XNOR U4294 ( .A(n3698), .B(n3699), .Z(N111) );
  NANDN U4295 ( .A(n3697), .B(n3696), .Z(n3701) );
  NAND U4296 ( .A(n3699), .B(n3698), .Z(n3700) );
  NAND U4297 ( .A(n3701), .B(n3700), .Z(n3785) );
  OR U4298 ( .A(n3703), .B(n3702), .Z(n3707) );
  OR U4299 ( .A(n3705), .B(n3704), .Z(n3706) );
  AND U4300 ( .A(n3707), .B(n3706), .Z(n3786) );
  XNOR U4301 ( .A(n3785), .B(n3786), .Z(n3787) );
  NANDN U4302 ( .A(n3709), .B(n3708), .Z(n3713) );
  NANDN U4303 ( .A(n3711), .B(n3710), .Z(n3712) );
  NAND U4304 ( .A(n3713), .B(n3712), .Z(n3876) );
  NAND U4305 ( .A(n3715), .B(n3714), .Z(n3719) );
  OR U4306 ( .A(n3717), .B(n3716), .Z(n3718) );
  AND U4307 ( .A(n3719), .B(n3718), .Z(n3812) );
  NANDN U4308 ( .A(n3720), .B(o[46]), .Z(n3854) );
  AND U4309 ( .A(x[143]), .B(y[672]), .Z(n3722) );
  NAND U4310 ( .A(x[128]), .B(y[687]), .Z(n3721) );
  XOR U4311 ( .A(n3722), .B(n3721), .Z(n3853) );
  XNOR U4312 ( .A(n3854), .B(n3853), .Z(n3815) );
  AND U4313 ( .A(x[140]), .B(y[675]), .Z(n3724) );
  NAND U4314 ( .A(x[139]), .B(y[676]), .Z(n3723) );
  XOR U4315 ( .A(n3724), .B(n3723), .Z(n3823) );
  NAND U4316 ( .A(x[141]), .B(y[674]), .Z(n3822) );
  XOR U4317 ( .A(n3823), .B(n3822), .Z(n3816) );
  AND U4318 ( .A(y[679]), .B(x[140]), .Z(n4112) );
  NAND U4319 ( .A(n3725), .B(n4112), .Z(n3729) );
  OR U4320 ( .A(n3727), .B(n3726), .Z(n3728) );
  AND U4321 ( .A(n3729), .B(n3728), .Z(n3818) );
  XNOR U4322 ( .A(n3817), .B(n3818), .Z(n3810) );
  ANDN U4323 ( .B(y[684]), .A(n160), .Z(n4489) );
  NAND U4324 ( .A(n3730), .B(n4489), .Z(n3733) );
  NANDN U4325 ( .A(n3731), .B(n4412), .Z(n3732) );
  NAND U4326 ( .A(n3733), .B(n3732), .Z(n3809) );
  XOR U4327 ( .A(n3810), .B(n3809), .Z(n3811) );
  XNOR U4328 ( .A(n3812), .B(n3811), .Z(n3797) );
  NAND U4329 ( .A(n3735), .B(n3734), .Z(n3739) );
  NANDN U4330 ( .A(n3737), .B(n3736), .Z(n3738) );
  AND U4331 ( .A(n3739), .B(n3738), .Z(n3798) );
  XNOR U4332 ( .A(n3797), .B(n3798), .Z(n3800) );
  OR U4333 ( .A(n3741), .B(n3740), .Z(n3745) );
  NANDN U4334 ( .A(n3743), .B(n3742), .Z(n3744) );
  AND U4335 ( .A(n3745), .B(n3744), .Z(n3799) );
  XNOR U4336 ( .A(n3800), .B(n3799), .Z(n3873) );
  NAND U4337 ( .A(x[136]), .B(y[683]), .Z(n4153) );
  OR U4338 ( .A(n4153), .B(n3746), .Z(n3750) );
  NANDN U4339 ( .A(n3748), .B(n3747), .Z(n3749) );
  NAND U4340 ( .A(n3750), .B(n3749), .Z(n3837) );
  AND U4341 ( .A(y[686]), .B(x[142]), .Z(n5536) );
  NAND U4342 ( .A(n3852), .B(n5536), .Z(n3754) );
  NANDN U4343 ( .A(n3752), .B(n3751), .Z(n3753) );
  AND U4344 ( .A(n3754), .B(n3753), .Z(n3836) );
  NAND U4345 ( .A(x[142]), .B(y[673]), .Z(n3863) );
  XOR U4346 ( .A(o[47]), .B(n3863), .Z(n3849) );
  AND U4347 ( .A(y[679]), .B(x[136]), .Z(n3756) );
  NAND U4348 ( .A(x[129]), .B(y[686]), .Z(n3755) );
  XOR U4349 ( .A(n3756), .B(n3755), .Z(n3848) );
  XNOR U4350 ( .A(n3849), .B(n3848), .Z(n3830) );
  AND U4351 ( .A(x[137]), .B(y[678]), .Z(n3758) );
  NAND U4352 ( .A(x[130]), .B(y[685]), .Z(n3757) );
  XOR U4353 ( .A(n3758), .B(n3757), .Z(n3870) );
  NAND U4354 ( .A(x[131]), .B(y[684]), .Z(n3869) );
  XOR U4355 ( .A(n3870), .B(n3869), .Z(n3831) );
  ANDN U4356 ( .B(y[680]), .A(n158), .Z(n4215) );
  AND U4357 ( .A(y[677]), .B(x[138]), .Z(n3760) );
  NAND U4358 ( .A(x[132]), .B(y[683]), .Z(n3759) );
  XOR U4359 ( .A(n3760), .B(n3759), .Z(n3858) );
  XOR U4360 ( .A(n4215), .B(n3858), .Z(n3843) );
  AND U4361 ( .A(x[134]), .B(y[681]), .Z(n3938) );
  XNOR U4362 ( .A(n3842), .B(n3938), .Z(n3844) );
  XOR U4363 ( .A(n3838), .B(n3839), .Z(n3803) );
  OR U4364 ( .A(n3762), .B(n3761), .Z(n3766) );
  NAND U4365 ( .A(n3764), .B(n3763), .Z(n3765) );
  NAND U4366 ( .A(n3766), .B(n3765), .Z(n3804) );
  XNOR U4367 ( .A(n3803), .B(n3804), .Z(n3806) );
  NANDN U4368 ( .A(n3768), .B(n3767), .Z(n3772) );
  NANDN U4369 ( .A(n3770), .B(n3769), .Z(n3771) );
  AND U4370 ( .A(n3772), .B(n3771), .Z(n3805) );
  XOR U4371 ( .A(n3806), .B(n3805), .Z(n3874) );
  XNOR U4372 ( .A(n3873), .B(n3874), .Z(n3875) );
  XOR U4373 ( .A(n3876), .B(n3875), .Z(n3791) );
  NANDN U4374 ( .A(n3774), .B(n3773), .Z(n3778) );
  NANDN U4375 ( .A(n3776), .B(n3775), .Z(n3777) );
  NAND U4376 ( .A(n3778), .B(n3777), .Z(n3792) );
  NAND U4377 ( .A(n3780), .B(n3779), .Z(n3784) );
  NANDN U4378 ( .A(n3782), .B(n3781), .Z(n3783) );
  NAND U4379 ( .A(n3784), .B(n3783), .Z(n3794) );
  XNOR U4380 ( .A(n3793), .B(n3794), .Z(n3788) );
  XOR U4381 ( .A(n3787), .B(n3788), .Z(N112) );
  NANDN U4382 ( .A(n3786), .B(n3785), .Z(n3790) );
  NANDN U4383 ( .A(n3788), .B(n3787), .Z(n3789) );
  NAND U4384 ( .A(n3790), .B(n3789), .Z(n3879) );
  NANDN U4385 ( .A(n3792), .B(n3791), .Z(n3796) );
  NANDN U4386 ( .A(n3794), .B(n3793), .Z(n3795) );
  NAND U4387 ( .A(n3796), .B(n3795), .Z(n3880) );
  XNOR U4388 ( .A(n3879), .B(n3880), .Z(n3881) );
  OR U4389 ( .A(n3798), .B(n3797), .Z(n3802) );
  OR U4390 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U4391 ( .A(n3802), .B(n3801), .Z(n3970) );
  OR U4392 ( .A(n3804), .B(n3803), .Z(n3808) );
  OR U4393 ( .A(n3806), .B(n3805), .Z(n3807) );
  NAND U4394 ( .A(n3808), .B(n3807), .Z(n3968) );
  OR U4395 ( .A(n3810), .B(n3809), .Z(n3814) );
  NANDN U4396 ( .A(n3812), .B(n3811), .Z(n3813) );
  AND U4397 ( .A(n3814), .B(n3813), .Z(n3967) );
  XOR U4398 ( .A(n3968), .B(n3967), .Z(n3969) );
  XNOR U4399 ( .A(n3970), .B(n3969), .Z(n3887) );
  NANDN U4400 ( .A(n3816), .B(n3815), .Z(n3820) );
  NAND U4401 ( .A(n3818), .B(n3817), .Z(n3819) );
  NAND U4402 ( .A(n3820), .B(n3819), .Z(n3922) );
  ANDN U4403 ( .B(y[676]), .A(n163), .Z(n4603) );
  NAND U4404 ( .A(n3821), .B(n4603), .Z(n3825) );
  OR U4405 ( .A(n3823), .B(n3822), .Z(n3824) );
  NAND U4406 ( .A(n3825), .B(n3824), .Z(n3905) );
  NAND U4407 ( .A(x[130]), .B(y[686]), .Z(n3826) );
  XOR U4408 ( .A(n3827), .B(n3826), .Z(n3911) );
  NAND U4409 ( .A(y[685]), .B(x[131]), .Z(n3910) );
  XOR U4410 ( .A(n3911), .B(n3910), .Z(n3903) );
  AND U4411 ( .A(x[141]), .B(y[675]), .Z(n3829) );
  NAND U4412 ( .A(x[133]), .B(y[683]), .Z(n3828) );
  XNOR U4413 ( .A(n3829), .B(n3828), .Z(n3932) );
  XNOR U4414 ( .A(n4603), .B(n3932), .Z(n3904) );
  XOR U4415 ( .A(n3903), .B(n3904), .Z(n3906) );
  XOR U4416 ( .A(n3905), .B(n3906), .Z(n3920) );
  NANDN U4417 ( .A(n3831), .B(n3830), .Z(n3835) );
  NAND U4418 ( .A(n3833), .B(n3832), .Z(n3834) );
  AND U4419 ( .A(n3835), .B(n3834), .Z(n3919) );
  XOR U4420 ( .A(n3922), .B(n3921), .Z(n3893) );
  NANDN U4421 ( .A(n3837), .B(n3836), .Z(n3841) );
  NAND U4422 ( .A(n3839), .B(n3838), .Z(n3840) );
  AND U4423 ( .A(n3841), .B(n3840), .Z(n3892) );
  OR U4424 ( .A(n3842), .B(n3938), .Z(n3846) );
  NANDN U4425 ( .A(n3844), .B(n3843), .Z(n3845) );
  NAND U4426 ( .A(n3846), .B(n3845), .Z(n3961) );
  NAND U4427 ( .A(x[136]), .B(y[686]), .Z(n4764) );
  NANDN U4428 ( .A(n4764), .B(n3847), .Z(n3851) );
  OR U4429 ( .A(n3849), .B(n3848), .Z(n3850) );
  NAND U4430 ( .A(n3851), .B(n3850), .Z(n3897) );
  AND U4431 ( .A(y[687]), .B(x[143]), .Z(n5882) );
  NAND U4432 ( .A(n3852), .B(n5882), .Z(n3856) );
  OR U4433 ( .A(n3854), .B(n3853), .Z(n3855) );
  AND U4434 ( .A(n3856), .B(n3855), .Z(n3898) );
  ANDN U4435 ( .B(y[683]), .A(n161), .Z(n4530) );
  NANDN U4436 ( .A(n3857), .B(n4530), .Z(n3860) );
  NANDN U4437 ( .A(n3858), .B(n4215), .Z(n3859) );
  AND U4438 ( .A(n3860), .B(n3859), .Z(n3927) );
  NAND U4439 ( .A(x[128]), .B(y[688]), .Z(n3948) );
  NAND U4440 ( .A(y[672]), .B(x[144]), .Z(n3947) );
  XOR U4441 ( .A(n3948), .B(n3947), .Z(n3949) );
  NAND U4442 ( .A(x[143]), .B(y[673]), .Z(n3935) );
  XOR U4443 ( .A(o[48]), .B(n3935), .Z(n3950) );
  XOR U4444 ( .A(n3949), .B(n3950), .Z(n3926) );
  NAND U4445 ( .A(x[135]), .B(y[681]), .Z(n3861) );
  XOR U4446 ( .A(n3862), .B(n3861), .Z(n3940) );
  NAND U4447 ( .A(x[138]), .B(y[678]), .Z(n3939) );
  XNOR U4448 ( .A(n3940), .B(n3939), .Z(n3925) );
  XNOR U4449 ( .A(n3926), .B(n3925), .Z(n3928) );
  XNOR U4450 ( .A(n3927), .B(n3928), .Z(n3900) );
  XNOR U4451 ( .A(n3899), .B(n3900), .Z(n3962) );
  NANDN U4452 ( .A(n3863), .B(o[47]), .Z(n3944) );
  NAND U4453 ( .A(x[129]), .B(y[687]), .Z(n3864) );
  XOR U4454 ( .A(n3865), .B(n3864), .Z(n3943) );
  XOR U4455 ( .A(n3944), .B(n3943), .Z(n3958) );
  AND U4456 ( .A(y[677]), .B(x[139]), .Z(n3867) );
  NAND U4457 ( .A(x[142]), .B(y[674]), .Z(n3866) );
  XOR U4458 ( .A(n3867), .B(n3866), .Z(n3916) );
  NAND U4459 ( .A(x[132]), .B(y[684]), .Z(n3915) );
  XNOR U4460 ( .A(n3916), .B(n3915), .Z(n3955) );
  ANDN U4461 ( .B(y[685]), .A(n160), .Z(n4599) );
  NAND U4462 ( .A(n3868), .B(n4599), .Z(n3872) );
  OR U4463 ( .A(n3870), .B(n3869), .Z(n3871) );
  NAND U4464 ( .A(n3872), .B(n3871), .Z(n3956) );
  XOR U4465 ( .A(n3958), .B(n3957), .Z(n3963) );
  XOR U4466 ( .A(n3892), .B(n3891), .Z(n3894) );
  NANDN U4467 ( .A(n3874), .B(n3873), .Z(n3878) );
  NANDN U4468 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4469 ( .A(n3878), .B(n3877), .Z(n3886) );
  XOR U4470 ( .A(n3885), .B(n3886), .Z(n3888) );
  XOR U4471 ( .A(n3887), .B(n3888), .Z(n3882) );
  XOR U4472 ( .A(n3881), .B(n3882), .Z(N113) );
  NANDN U4473 ( .A(n3880), .B(n3879), .Z(n3884) );
  NANDN U4474 ( .A(n3882), .B(n3881), .Z(n3883) );
  NAND U4475 ( .A(n3884), .B(n3883), .Z(n3973) );
  NANDN U4476 ( .A(n3886), .B(n3885), .Z(n3890) );
  OR U4477 ( .A(n3888), .B(n3887), .Z(n3889) );
  NAND U4478 ( .A(n3890), .B(n3889), .Z(n3974) );
  XNOR U4479 ( .A(n3973), .B(n3974), .Z(n3975) );
  NANDN U4480 ( .A(n3892), .B(n3891), .Z(n3896) );
  NANDN U4481 ( .A(n3894), .B(n3893), .Z(n3895) );
  NAND U4482 ( .A(n3896), .B(n3895), .Z(n3988) );
  NANDN U4483 ( .A(n3898), .B(n3897), .Z(n3902) );
  NANDN U4484 ( .A(n3900), .B(n3899), .Z(n3901) );
  NAND U4485 ( .A(n3902), .B(n3901), .Z(n3994) );
  NANDN U4486 ( .A(n3904), .B(n3903), .Z(n3908) );
  NANDN U4487 ( .A(n3906), .B(n3905), .Z(n3907) );
  NAND U4488 ( .A(n3908), .B(n3907), .Z(n3992) );
  AND U4489 ( .A(y[682]), .B(x[135]), .Z(n4152) );
  ANDN U4490 ( .B(y[685]), .A(n155), .Z(n4016) );
  ANDN U4491 ( .B(y[678]), .A(n162), .Z(n4014) );
  ANDN U4492 ( .B(y[676]), .A(n164), .Z(n4013) );
  XNOR U4493 ( .A(n4014), .B(n4013), .Z(n4015) );
  XNOR U4494 ( .A(n4016), .B(n4015), .Z(n4036) );
  NAND U4495 ( .A(x[133]), .B(y[684]), .Z(n4055) );
  NAND U4496 ( .A(y[681]), .B(x[136]), .Z(n4052) );
  XNOR U4497 ( .A(n4053), .B(n4052), .Z(n4054) );
  XOR U4498 ( .A(n4055), .B(n4054), .Z(n4037) );
  XNOR U4499 ( .A(n4036), .B(n4037), .Z(n4038) );
  XNOR U4500 ( .A(n4152), .B(n4038), .Z(n4032) );
  AND U4501 ( .A(y[686]), .B(x[137]), .Z(n3909) );
  NAND U4502 ( .A(n3909), .B(n4045), .Z(n3913) );
  OR U4503 ( .A(n3911), .B(n3910), .Z(n3912) );
  NAND U4504 ( .A(n3913), .B(n3912), .Z(n4031) );
  NAND U4505 ( .A(x[139]), .B(y[674]), .Z(n4114) );
  AND U4506 ( .A(y[677]), .B(x[142]), .Z(n3914) );
  NANDN U4507 ( .A(n4114), .B(n3914), .Z(n3918) );
  OR U4508 ( .A(n3916), .B(n3915), .Z(n3917) );
  AND U4509 ( .A(n3918), .B(n3917), .Z(n4030) );
  XNOR U4510 ( .A(n3992), .B(n3991), .Z(n3993) );
  XOR U4511 ( .A(n3994), .B(n3993), .Z(n3985) );
  NANDN U4512 ( .A(n3920), .B(n3919), .Z(n3924) );
  NANDN U4513 ( .A(n3922), .B(n3921), .Z(n3923) );
  AND U4514 ( .A(n3924), .B(n3923), .Z(n3986) );
  XNOR U4515 ( .A(n3988), .B(n3987), .Z(n3979) );
  OR U4516 ( .A(n3926), .B(n3925), .Z(n3930) );
  OR U4517 ( .A(n3928), .B(n3927), .Z(n3929) );
  NAND U4518 ( .A(n3930), .B(n3929), .Z(n4000) );
  ANDN U4519 ( .B(y[683]), .A(n164), .Z(n4878) );
  NAND U4520 ( .A(n3931), .B(n4878), .Z(n3934) );
  NAND U4521 ( .A(n3932), .B(n4603), .Z(n3933) );
  AND U4522 ( .A(n3934), .B(n3933), .Z(n4067) );
  ANDN U4523 ( .B(y[677]), .A(n163), .Z(n4027) );
  ANDN U4524 ( .B(y[675]), .A(n165), .Z(n4025) );
  ANDN U4525 ( .B(y[674]), .A(n166), .Z(n4024) );
  XNOR U4526 ( .A(n4025), .B(n4024), .Z(n4026) );
  XNOR U4527 ( .A(n4027), .B(n4026), .Z(n4064) );
  NANDN U4528 ( .A(n3935), .B(o[48]), .Z(n4042) );
  AND U4529 ( .A(x[137]), .B(y[680]), .Z(n3937) );
  NAND U4530 ( .A(x[129]), .B(y[688]), .Z(n3936) );
  XNOR U4531 ( .A(n3937), .B(n3936), .Z(n4041) );
  XOR U4532 ( .A(n4067), .B(n4066), .Z(n3997) );
  NAND U4533 ( .A(n4152), .B(n3938), .Z(n3942) );
  OR U4534 ( .A(n3940), .B(n3939), .Z(n3941) );
  NAND U4535 ( .A(n3942), .B(n3941), .Z(n4058) );
  NAND U4536 ( .A(x[136]), .B(y[687]), .Z(n4598) );
  ANDN U4537 ( .B(y[680]), .A(n152), .Z(n4131) );
  NANDN U4538 ( .A(n4598), .B(n4131), .Z(n3946) );
  OR U4539 ( .A(n3944), .B(n3943), .Z(n3945) );
  AND U4540 ( .A(n3946), .B(n3945), .Z(n4059) );
  OR U4541 ( .A(n3948), .B(n3947), .Z(n3952) );
  NANDN U4542 ( .A(n3950), .B(n3949), .Z(n3951) );
  NAND U4543 ( .A(n3952), .B(n3951), .Z(n4071) );
  AND U4544 ( .A(y[679]), .B(x[138]), .Z(n3954) );
  NAND U4545 ( .A(x[130]), .B(y[687]), .Z(n3953) );
  XOR U4546 ( .A(n3954), .B(n3953), .Z(n4047) );
  NAND U4547 ( .A(x[131]), .B(y[686]), .Z(n4046) );
  XOR U4548 ( .A(n4047), .B(n4046), .Z(n4070) );
  XNOR U4549 ( .A(n4071), .B(n4070), .Z(n4073) );
  NAND U4550 ( .A(x[144]), .B(y[673]), .Z(n4019) );
  XOR U4551 ( .A(o[49]), .B(n4019), .Z(n4004) );
  NAND U4552 ( .A(y[672]), .B(x[145]), .Z(n4003) );
  XOR U4553 ( .A(n4004), .B(n4003), .Z(n4005) );
  NAND U4554 ( .A(y[689]), .B(x[128]), .Z(n4006) );
  XNOR U4555 ( .A(n4005), .B(n4006), .Z(n4072) );
  XOR U4556 ( .A(n4073), .B(n4072), .Z(n4061) );
  XNOR U4557 ( .A(n4060), .B(n4061), .Z(n3998) );
  XNOR U4558 ( .A(n3997), .B(n3998), .Z(n3999) );
  XOR U4559 ( .A(n4000), .B(n3999), .Z(n4076) );
  NANDN U4560 ( .A(n3956), .B(n3955), .Z(n3960) );
  OR U4561 ( .A(n3958), .B(n3957), .Z(n3959) );
  NAND U4562 ( .A(n3960), .B(n3959), .Z(n4077) );
  NANDN U4563 ( .A(n3962), .B(n3961), .Z(n3966) );
  NAND U4564 ( .A(n3964), .B(n3963), .Z(n3965) );
  NAND U4565 ( .A(n3966), .B(n3965), .Z(n4079) );
  XNOR U4566 ( .A(n4078), .B(n4079), .Z(n3980) );
  XNOR U4567 ( .A(n3979), .B(n3980), .Z(n3982) );
  OR U4568 ( .A(n3968), .B(n3967), .Z(n3972) );
  NANDN U4569 ( .A(n3970), .B(n3969), .Z(n3971) );
  AND U4570 ( .A(n3972), .B(n3971), .Z(n3981) );
  XOR U4571 ( .A(n3982), .B(n3981), .Z(n3976) );
  XNOR U4572 ( .A(n3975), .B(n3976), .Z(N114) );
  NANDN U4573 ( .A(n3974), .B(n3973), .Z(n3978) );
  NAND U4574 ( .A(n3976), .B(n3975), .Z(n3977) );
  NAND U4575 ( .A(n3978), .B(n3977), .Z(n4082) );
  OR U4576 ( .A(n3980), .B(n3979), .Z(n3984) );
  OR U4577 ( .A(n3982), .B(n3981), .Z(n3983) );
  AND U4578 ( .A(n3984), .B(n3983), .Z(n4083) );
  XNOR U4579 ( .A(n4082), .B(n4083), .Z(n4084) );
  NANDN U4580 ( .A(n3986), .B(n3985), .Z(n3990) );
  NANDN U4581 ( .A(n3988), .B(n3987), .Z(n3989) );
  NAND U4582 ( .A(n3990), .B(n3989), .Z(n4091) );
  NANDN U4583 ( .A(n3992), .B(n3991), .Z(n3996) );
  NANDN U4584 ( .A(n3994), .B(n3993), .Z(n3995) );
  AND U4585 ( .A(n3996), .B(n3995), .Z(n4191) );
  NANDN U4586 ( .A(n3998), .B(n3997), .Z(n4002) );
  NANDN U4587 ( .A(n4000), .B(n3999), .Z(n4001) );
  AND U4588 ( .A(n4002), .B(n4001), .Z(n4192) );
  XOR U4589 ( .A(n4191), .B(n4192), .Z(n4193) );
  OR U4590 ( .A(n4004), .B(n4003), .Z(n4008) );
  NANDN U4591 ( .A(n4006), .B(n4005), .Z(n4007) );
  NAND U4592 ( .A(n4008), .B(n4007), .Z(n4174) );
  NAND U4593 ( .A(x[135]), .B(y[683]), .Z(n4009) );
  XOR U4594 ( .A(n4010), .B(n4009), .Z(n4155) );
  NAND U4595 ( .A(x[132]), .B(y[686]), .Z(n4154) );
  XNOR U4596 ( .A(n4155), .B(n4154), .Z(n4100) );
  ANDN U4597 ( .B(y[684]), .A(n157), .Z(n4627) );
  NAND U4598 ( .A(y[685]), .B(x[133]), .Z(n4262) );
  XOR U4599 ( .A(n4627), .B(n4262), .Z(n4101) );
  XNOR U4600 ( .A(n4174), .B(n4173), .Z(n4175) );
  NAND U4601 ( .A(x[130]), .B(y[688]), .Z(n4116) );
  AND U4602 ( .A(y[679]), .B(x[139]), .Z(n4012) );
  NAND U4603 ( .A(x[144]), .B(y[674]), .Z(n4011) );
  XOR U4604 ( .A(n4012), .B(n4011), .Z(n4115) );
  XOR U4605 ( .A(n4116), .B(n4115), .Z(n4176) );
  XOR U4606 ( .A(n4175), .B(n4176), .Z(n4185) );
  OR U4607 ( .A(n4014), .B(n4013), .Z(n4018) );
  OR U4608 ( .A(n4016), .B(n4015), .Z(n4017) );
  NAND U4609 ( .A(n4018), .B(n4017), .Z(n4122) );
  NANDN U4610 ( .A(n4019), .B(o[49]), .Z(n4133) );
  AND U4611 ( .A(x[138]), .B(y[680]), .Z(n4021) );
  NAND U4612 ( .A(x[129]), .B(y[689]), .Z(n4020) );
  XNOR U4613 ( .A(n4021), .B(n4020), .Z(n4132) );
  NAND U4614 ( .A(x[142]), .B(y[676]), .Z(n4022) );
  XOR U4615 ( .A(n4023), .B(n4022), .Z(n4108) );
  NAND U4616 ( .A(y[675]), .B(x[143]), .Z(n4107) );
  XOR U4617 ( .A(n4108), .B(n4107), .Z(n4119) );
  XOR U4618 ( .A(n4122), .B(n4121), .Z(n4186) );
  XOR U4619 ( .A(n4185), .B(n4186), .Z(n4188) );
  OR U4620 ( .A(n4025), .B(n4024), .Z(n4029) );
  OR U4621 ( .A(n4027), .B(n4026), .Z(n4028) );
  AND U4622 ( .A(n4029), .B(n4028), .Z(n4187) );
  NANDN U4623 ( .A(n4031), .B(n4030), .Z(n4035) );
  NAND U4624 ( .A(n4033), .B(n4032), .Z(n4034) );
  NAND U4625 ( .A(n4035), .B(n4034), .Z(n4164) );
  NANDN U4626 ( .A(n4037), .B(n4036), .Z(n4040) );
  NAND U4627 ( .A(n4038), .B(n4152), .Z(n4039) );
  NAND U4628 ( .A(n4040), .B(n4039), .Z(n4162) );
  AND U4629 ( .A(y[688]), .B(x[137]), .Z(n5110) );
  NAND U4630 ( .A(n5110), .B(n4131), .Z(n4044) );
  NANDN U4631 ( .A(n4042), .B(n4041), .Z(n4043) );
  NAND U4632 ( .A(n4044), .B(n4043), .Z(n4182) );
  IV U4633 ( .A(y[687]), .Z(n4750) );
  NOR U4634 ( .A(n161), .B(n4750), .Z(n5109) );
  NAND U4635 ( .A(n5109), .B(n4045), .Z(n4049) );
  OR U4636 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4637 ( .A(n4049), .B(n4048), .Z(n4127) );
  NAND U4638 ( .A(x[128]), .B(y[690]), .Z(n4137) );
  NAND U4639 ( .A(y[672]), .B(x[146]), .Z(n4136) );
  XOR U4640 ( .A(n4137), .B(n4136), .Z(n4138) );
  NAND U4641 ( .A(x[145]), .B(y[673]), .Z(n4160) );
  XOR U4642 ( .A(o[50]), .B(n4160), .Z(n4139) );
  XOR U4643 ( .A(n4138), .B(n4139), .Z(n4126) );
  ANDN U4644 ( .B(y[678]), .A(n163), .Z(n4223) );
  AND U4645 ( .A(x[131]), .B(y[687]), .Z(n4051) );
  NAND U4646 ( .A(x[141]), .B(y[677]), .Z(n4050) );
  XNOR U4647 ( .A(n4051), .B(n4050), .Z(n4145) );
  XOR U4648 ( .A(n4126), .B(n4125), .Z(n4128) );
  XOR U4649 ( .A(n4127), .B(n4128), .Z(n4179) );
  NANDN U4650 ( .A(n4053), .B(n4052), .Z(n4057) );
  NAND U4651 ( .A(n4055), .B(n4054), .Z(n4056) );
  AND U4652 ( .A(n4057), .B(n4056), .Z(n4180) );
  XOR U4653 ( .A(n4179), .B(n4180), .Z(n4181) );
  XNOR U4654 ( .A(n4182), .B(n4181), .Z(n4161) );
  XOR U4655 ( .A(n4162), .B(n4161), .Z(n4163) );
  XOR U4656 ( .A(n4164), .B(n4163), .Z(n4095) );
  XOR U4657 ( .A(n4094), .B(n4095), .Z(n4097) );
  NANDN U4658 ( .A(n4059), .B(n4058), .Z(n4063) );
  NANDN U4659 ( .A(n4061), .B(n4060), .Z(n4062) );
  NAND U4660 ( .A(n4063), .B(n4062), .Z(n4170) );
  NAND U4661 ( .A(n4065), .B(n4064), .Z(n4069) );
  NANDN U4662 ( .A(n4067), .B(n4066), .Z(n4068) );
  NAND U4663 ( .A(n4069), .B(n4068), .Z(n4168) );
  NAND U4664 ( .A(n4071), .B(n4070), .Z(n4075) );
  NANDN U4665 ( .A(n4073), .B(n4072), .Z(n4074) );
  AND U4666 ( .A(n4075), .B(n4074), .Z(n4167) );
  XNOR U4667 ( .A(n4170), .B(n4169), .Z(n4096) );
  XOR U4668 ( .A(n4097), .B(n4096), .Z(n4194) );
  XNOR U4669 ( .A(n4193), .B(n4194), .Z(n4089) );
  NANDN U4670 ( .A(n4077), .B(n4076), .Z(n4081) );
  NANDN U4671 ( .A(n4079), .B(n4078), .Z(n4080) );
  AND U4672 ( .A(n4081), .B(n4080), .Z(n4088) );
  XOR U4673 ( .A(n4089), .B(n4088), .Z(n4090) );
  XOR U4674 ( .A(n4091), .B(n4090), .Z(n4085) );
  XOR U4675 ( .A(n4084), .B(n4085), .Z(N115) );
  NANDN U4676 ( .A(n4083), .B(n4082), .Z(n4087) );
  NANDN U4677 ( .A(n4085), .B(n4084), .Z(n4086) );
  NAND U4678 ( .A(n4087), .B(n4086), .Z(n4197) );
  OR U4679 ( .A(n4089), .B(n4088), .Z(n4093) );
  NAND U4680 ( .A(n4091), .B(n4090), .Z(n4092) );
  NAND U4681 ( .A(n4093), .B(n4092), .Z(n4198) );
  XNOR U4682 ( .A(n4197), .B(n4198), .Z(n4199) );
  NANDN U4683 ( .A(n4095), .B(n4094), .Z(n4099) );
  OR U4684 ( .A(n4097), .B(n4096), .Z(n4098) );
  NAND U4685 ( .A(n4099), .B(n4098), .Z(n4204) );
  NANDN U4686 ( .A(n4627), .B(n4262), .Z(n4103) );
  NANDN U4687 ( .A(n4101), .B(n4100), .Z(n4102) );
  AND U4688 ( .A(n4103), .B(n4102), .Z(n4303) );
  AND U4689 ( .A(y[683]), .B(x[136]), .Z(n4105) );
  NAND U4690 ( .A(x[142]), .B(y[677]), .Z(n4104) );
  XOR U4691 ( .A(n4105), .B(n4104), .Z(n4280) );
  NAND U4692 ( .A(x[129]), .B(y[690]), .Z(n4279) );
  XNOR U4693 ( .A(n4280), .B(n4279), .Z(n4241) );
  AND U4694 ( .A(y[676]), .B(x[137]), .Z(n4106) );
  ANDN U4695 ( .B(y[681]), .A(n165), .Z(n4805) );
  NAND U4696 ( .A(n4106), .B(n4805), .Z(n4110) );
  OR U4697 ( .A(n4108), .B(n4107), .Z(n4109) );
  AND U4698 ( .A(n4110), .B(n4109), .Z(n4239) );
  NAND U4699 ( .A(x[141]), .B(y[678]), .Z(n4111) );
  XOR U4700 ( .A(n4112), .B(n4111), .Z(n4226) );
  AND U4701 ( .A(x[130]), .B(y[689]), .Z(n4225) );
  XOR U4702 ( .A(n4226), .B(n4225), .Z(n4238) );
  XOR U4703 ( .A(n4239), .B(n4238), .Z(n4240) );
  XOR U4704 ( .A(n4241), .B(n4240), .Z(n4300) );
  AND U4705 ( .A(y[679]), .B(x[144]), .Z(n4113) );
  NANDN U4706 ( .A(n4114), .B(n4113), .Z(n4118) );
  OR U4707 ( .A(n4116), .B(n4115), .Z(n4117) );
  NAND U4708 ( .A(n4118), .B(n4117), .Z(n4301) );
  XNOR U4709 ( .A(n4300), .B(n4301), .Z(n4302) );
  XOR U4710 ( .A(n4303), .B(n4302), .Z(n4209) );
  NAND U4711 ( .A(n4120), .B(n4119), .Z(n4124) );
  NANDN U4712 ( .A(n4122), .B(n4121), .Z(n4123) );
  NAND U4713 ( .A(n4124), .B(n4123), .Z(n4295) );
  NANDN U4714 ( .A(n4126), .B(n4125), .Z(n4130) );
  NANDN U4715 ( .A(n4128), .B(n4127), .Z(n4129) );
  NAND U4716 ( .A(n4130), .B(n4129), .Z(n4294) );
  XOR U4717 ( .A(n4295), .B(n4294), .Z(n4296) );
  AND U4718 ( .A(x[138]), .B(y[689]), .Z(n5410) );
  NAND U4719 ( .A(n4131), .B(n5410), .Z(n4135) );
  NANDN U4720 ( .A(n4133), .B(n4132), .Z(n4134) );
  NAND U4721 ( .A(n4135), .B(n4134), .Z(n4258) );
  OR U4722 ( .A(n4137), .B(n4136), .Z(n4141) );
  NANDN U4723 ( .A(n4139), .B(n4138), .Z(n4140) );
  NAND U4724 ( .A(n4141), .B(n4140), .Z(n4257) );
  AND U4725 ( .A(x[137]), .B(y[682]), .Z(n4143) );
  NAND U4726 ( .A(x[144]), .B(y[675]), .Z(n4142) );
  XOR U4727 ( .A(n4143), .B(n4142), .Z(n4235) );
  AND U4728 ( .A(y[676]), .B(x[143]), .Z(n4234) );
  XNOR U4729 ( .A(n4235), .B(n4234), .Z(n4256) );
  XNOR U4730 ( .A(n4257), .B(n4256), .Z(n4259) );
  XNOR U4731 ( .A(n4258), .B(n4259), .Z(n4290) );
  AND U4732 ( .A(x[141]), .B(y[687]), .Z(n5505) );
  NAND U4733 ( .A(n4144), .B(n5505), .Z(n4147) );
  NAND U4734 ( .A(n4145), .B(n4223), .Z(n4146) );
  NAND U4735 ( .A(n4147), .B(n4146), .Z(n4253) );
  AND U4736 ( .A(x[139]), .B(y[680]), .Z(n4149) );
  NAND U4737 ( .A(x[135]), .B(y[684]), .Z(n4148) );
  XOR U4738 ( .A(n4149), .B(n4148), .Z(n4217) );
  NAND U4739 ( .A(x[131]), .B(y[688]), .Z(n4216) );
  XOR U4740 ( .A(n4217), .B(n4216), .Z(n4251) );
  AND U4741 ( .A(y[673]), .B(x[146]), .Z(n4222) );
  XNOR U4742 ( .A(o[51]), .B(n4222), .Z(n4285) );
  AND U4743 ( .A(x[138]), .B(y[681]), .Z(n4151) );
  NAND U4744 ( .A(x[145]), .B(y[674]), .Z(n4150) );
  XOR U4745 ( .A(n4151), .B(n4150), .Z(n4284) );
  XOR U4746 ( .A(n4285), .B(n4284), .Z(n4250) );
  XOR U4747 ( .A(n4253), .B(n4252), .Z(n4288) );
  NANDN U4748 ( .A(n4153), .B(n4152), .Z(n4157) );
  OR U4749 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U4750 ( .A(n4157), .B(n4156), .Z(n4244) );
  ANDN U4751 ( .B(y[687]), .A(n155), .Z(n4400) );
  AND U4752 ( .A(x[134]), .B(y[685]), .Z(n4159) );
  NAND U4753 ( .A(x[133]), .B(y[686]), .Z(n4158) );
  XNOR U4754 ( .A(n4159), .B(n4158), .Z(n4263) );
  XNOR U4755 ( .A(n4400), .B(n4263), .Z(n4245) );
  NANDN U4756 ( .A(n4160), .B(o[50]), .Z(n4269) );
  NAND U4757 ( .A(x[128]), .B(y[691]), .Z(n4267) );
  NAND U4758 ( .A(y[672]), .B(x[147]), .Z(n4266) );
  XOR U4759 ( .A(n4267), .B(n4266), .Z(n4268) );
  XOR U4760 ( .A(n4269), .B(n4268), .Z(n4247) );
  XNOR U4761 ( .A(n4246), .B(n4247), .Z(n4289) );
  XNOR U4762 ( .A(n4288), .B(n4289), .Z(n4291) );
  XNOR U4763 ( .A(n4290), .B(n4291), .Z(n4297) );
  XNOR U4764 ( .A(n4296), .B(n4297), .Z(n4210) );
  XNOR U4765 ( .A(n4209), .B(n4210), .Z(n4211) );
  OR U4766 ( .A(n4162), .B(n4161), .Z(n4166) );
  NAND U4767 ( .A(n4164), .B(n4163), .Z(n4165) );
  NAND U4768 ( .A(n4166), .B(n4165), .Z(n4212) );
  XOR U4769 ( .A(n4211), .B(n4212), .Z(n4308) );
  NANDN U4770 ( .A(n4168), .B(n4167), .Z(n4172) );
  NANDN U4771 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U4772 ( .A(n4172), .B(n4171), .Z(n4306) );
  NANDN U4773 ( .A(n4174), .B(n4173), .Z(n4178) );
  NANDN U4774 ( .A(n4176), .B(n4175), .Z(n4177) );
  AND U4775 ( .A(n4178), .B(n4177), .Z(n4315) );
  NANDN U4776 ( .A(n4180), .B(n4179), .Z(n4184) );
  OR U4777 ( .A(n4182), .B(n4181), .Z(n4183) );
  AND U4778 ( .A(n4184), .B(n4183), .Z(n4312) );
  NANDN U4779 ( .A(n4186), .B(n4185), .Z(n4190) );
  NANDN U4780 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U4781 ( .A(n4190), .B(n4189), .Z(n4313) );
  XOR U4782 ( .A(n4312), .B(n4313), .Z(n4314) );
  XOR U4783 ( .A(n4308), .B(n4309), .Z(n4203) );
  XNOR U4784 ( .A(n4204), .B(n4203), .Z(n4206) );
  OR U4785 ( .A(n4192), .B(n4191), .Z(n4196) );
  NANDN U4786 ( .A(n4194), .B(n4193), .Z(n4195) );
  AND U4787 ( .A(n4196), .B(n4195), .Z(n4205) );
  XOR U4788 ( .A(n4206), .B(n4205), .Z(n4200) );
  XNOR U4789 ( .A(n4199), .B(n4200), .Z(N116) );
  NANDN U4790 ( .A(n4198), .B(n4197), .Z(n4202) );
  NAND U4791 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U4792 ( .A(n4202), .B(n4201), .Z(n4318) );
  OR U4793 ( .A(n4204), .B(n4203), .Z(n4208) );
  OR U4794 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U4795 ( .A(n4208), .B(n4207), .Z(n4319) );
  XNOR U4796 ( .A(n4318), .B(n4319), .Z(n4320) );
  NANDN U4797 ( .A(n4210), .B(n4209), .Z(n4214) );
  NANDN U4798 ( .A(n4212), .B(n4211), .Z(n4213) );
  AND U4799 ( .A(n4214), .B(n4213), .Z(n4425) );
  ANDN U4800 ( .B(y[684]), .A(n162), .Z(n4771) );
  NAND U4801 ( .A(n4771), .B(n4215), .Z(n4219) );
  OR U4802 ( .A(n4217), .B(n4216), .Z(n4218) );
  AND U4803 ( .A(n4219), .B(n4218), .Z(n4390) );
  NAND U4804 ( .A(x[147]), .B(y[673]), .Z(n4364) );
  XOR U4805 ( .A(o[52]), .B(n4364), .Z(n4367) );
  AND U4806 ( .A(x[139]), .B(y[681]), .Z(n4221) );
  NAND U4807 ( .A(x[129]), .B(y[691]), .Z(n4220) );
  XNOR U4808 ( .A(n4221), .B(n4220), .Z(n4366) );
  NAND U4809 ( .A(o[51]), .B(n4222), .Z(n4397) );
  NAND U4810 ( .A(x[148]), .B(y[672]), .Z(n4395) );
  AND U4811 ( .A(x[128]), .B(y[692]), .Z(n4394) );
  XNOR U4812 ( .A(n4395), .B(n4394), .Z(n4396) );
  XNOR U4813 ( .A(n4389), .B(n4388), .Z(n4391) );
  XOR U4814 ( .A(n4390), .B(n4391), .Z(n4373) );
  AND U4815 ( .A(y[679]), .B(x[141]), .Z(n4224) );
  NAND U4816 ( .A(n4224), .B(n4223), .Z(n4228) );
  NANDN U4817 ( .A(n4226), .B(n4225), .Z(n4227) );
  AND U4818 ( .A(n4228), .B(n4227), .Z(n4384) );
  NAND U4819 ( .A(x[130]), .B(y[690]), .Z(n4414) );
  AND U4820 ( .A(y[682]), .B(x[138]), .Z(n4230) );
  AND U4821 ( .A(y[676]), .B(x[144]), .Z(n4229) );
  XNOR U4822 ( .A(n4230), .B(n4229), .Z(n4413) );
  XOR U4823 ( .A(n4414), .B(n4413), .Z(n4382) );
  AND U4824 ( .A(y[677]), .B(x[143]), .Z(n4232) );
  NAND U4825 ( .A(x[137]), .B(y[683]), .Z(n4231) );
  XOR U4826 ( .A(n4232), .B(n4231), .Z(n4361) );
  NAND U4827 ( .A(x[142]), .B(y[678]), .Z(n4360) );
  XNOR U4828 ( .A(n4361), .B(n4360), .Z(n4383) );
  XNOR U4829 ( .A(n4384), .B(n4385), .Z(n4370) );
  AND U4830 ( .A(x[144]), .B(y[682]), .Z(n5168) );
  NANDN U4831 ( .A(n4233), .B(n5168), .Z(n4237) );
  NANDN U4832 ( .A(n4235), .B(n4234), .Z(n4236) );
  NAND U4833 ( .A(n4237), .B(n4236), .Z(n4371) );
  XOR U4834 ( .A(n4370), .B(n4371), .Z(n4372) );
  XOR U4835 ( .A(n4373), .B(n4372), .Z(n4333) );
  OR U4836 ( .A(n4239), .B(n4238), .Z(n4243) );
  NANDN U4837 ( .A(n4241), .B(n4240), .Z(n4242) );
  NAND U4838 ( .A(n4243), .B(n4242), .Z(n4330) );
  NANDN U4839 ( .A(n4245), .B(n4244), .Z(n4249) );
  NANDN U4840 ( .A(n4247), .B(n4246), .Z(n4248) );
  AND U4841 ( .A(n4249), .B(n4248), .Z(n4331) );
  XNOR U4842 ( .A(n4333), .B(n4332), .Z(n4419) );
  NAND U4843 ( .A(n4251), .B(n4250), .Z(n4255) );
  NAND U4844 ( .A(n4253), .B(n4252), .Z(n4254) );
  NAND U4845 ( .A(n4255), .B(n4254), .Z(n4418) );
  NAND U4846 ( .A(n4257), .B(n4256), .Z(n4261) );
  NANDN U4847 ( .A(n4259), .B(n4258), .Z(n4260) );
  NAND U4848 ( .A(n4261), .B(n4260), .Z(n4339) );
  ANDN U4849 ( .B(y[686]), .A(n157), .Z(n4348) );
  NANDN U4850 ( .A(n4262), .B(n4348), .Z(n4265) );
  NAND U4851 ( .A(n4263), .B(n4400), .Z(n4264) );
  AND U4852 ( .A(n4265), .B(n4264), .Z(n4345) );
  OR U4853 ( .A(n4267), .B(n4266), .Z(n4271) );
  NANDN U4854 ( .A(n4269), .B(n4268), .Z(n4270) );
  AND U4855 ( .A(n4271), .B(n4270), .Z(n4343) );
  AND U4856 ( .A(x[140]), .B(y[680]), .Z(n4273) );
  NAND U4857 ( .A(x[146]), .B(y[674]), .Z(n4272) );
  XOR U4858 ( .A(n4273), .B(n4272), .Z(n4356) );
  NAND U4859 ( .A(x[145]), .B(y[675]), .Z(n4355) );
  XOR U4860 ( .A(n4356), .B(n4355), .Z(n4342) );
  XNOR U4861 ( .A(n4343), .B(n4342), .Z(n4344) );
  XOR U4862 ( .A(n4345), .B(n4344), .Z(n4336) );
  NAND U4863 ( .A(x[135]), .B(y[685]), .Z(n4402) );
  AND U4864 ( .A(x[133]), .B(y[687]), .Z(n4275) );
  NAND U4865 ( .A(x[132]), .B(y[688]), .Z(n4274) );
  XOR U4866 ( .A(n4275), .B(n4274), .Z(n4401) );
  XNOR U4867 ( .A(n4402), .B(n4401), .Z(n4349) );
  XOR U4868 ( .A(n4348), .B(n4349), .Z(n4351) );
  NAND U4869 ( .A(x[136]), .B(y[684]), .Z(n4409) );
  AND U4870 ( .A(x[131]), .B(y[689]), .Z(n4277) );
  NAND U4871 ( .A(x[141]), .B(y[679]), .Z(n4276) );
  XOR U4872 ( .A(n4277), .B(n4276), .Z(n4408) );
  XNOR U4873 ( .A(n4409), .B(n4408), .Z(n4350) );
  XNOR U4874 ( .A(n4351), .B(n4350), .Z(n4378) );
  ANDN U4875 ( .B(y[683]), .A(n165), .Z(n5030) );
  NAND U4876 ( .A(n5030), .B(n4278), .Z(n4282) );
  OR U4877 ( .A(n4280), .B(n4279), .Z(n4281) );
  NAND U4878 ( .A(n4282), .B(n4281), .Z(n4377) );
  AND U4879 ( .A(x[145]), .B(y[681]), .Z(n5181) );
  NANDN U4880 ( .A(n4283), .B(n5181), .Z(n4287) );
  OR U4881 ( .A(n4285), .B(n4284), .Z(n4286) );
  NAND U4882 ( .A(n4287), .B(n4286), .Z(n4376) );
  XOR U4883 ( .A(n4377), .B(n4376), .Z(n4379) );
  XNOR U4884 ( .A(n4378), .B(n4379), .Z(n4337) );
  XNOR U4885 ( .A(n4336), .B(n4337), .Z(n4338) );
  XNOR U4886 ( .A(n4339), .B(n4338), .Z(n4417) );
  XOR U4887 ( .A(n4418), .B(n4417), .Z(n4420) );
  XOR U4888 ( .A(n4419), .B(n4420), .Z(n4423) );
  OR U4889 ( .A(n4289), .B(n4288), .Z(n4293) );
  OR U4890 ( .A(n4291), .B(n4290), .Z(n4292) );
  NAND U4891 ( .A(n4293), .B(n4292), .Z(n4430) );
  OR U4892 ( .A(n4295), .B(n4294), .Z(n4299) );
  NANDN U4893 ( .A(n4297), .B(n4296), .Z(n4298) );
  NAND U4894 ( .A(n4299), .B(n4298), .Z(n4429) );
  XOR U4895 ( .A(n4430), .B(n4429), .Z(n4431) );
  NANDN U4896 ( .A(n4301), .B(n4300), .Z(n4305) );
  NANDN U4897 ( .A(n4303), .B(n4302), .Z(n4304) );
  NAND U4898 ( .A(n4305), .B(n4304), .Z(n4432) );
  XNOR U4899 ( .A(n4423), .B(n4424), .Z(n4426) );
  XOR U4900 ( .A(n4425), .B(n4426), .Z(n4324) );
  NANDN U4901 ( .A(n4307), .B(n4306), .Z(n4311) );
  NANDN U4902 ( .A(n4309), .B(n4308), .Z(n4310) );
  AND U4903 ( .A(n4311), .B(n4310), .Z(n4325) );
  XNOR U4904 ( .A(n4324), .B(n4325), .Z(n4327) );
  OR U4905 ( .A(n4313), .B(n4312), .Z(n4317) );
  NANDN U4906 ( .A(n4315), .B(n4314), .Z(n4316) );
  NAND U4907 ( .A(n4317), .B(n4316), .Z(n4326) );
  XOR U4908 ( .A(n4327), .B(n4326), .Z(n4321) );
  XOR U4909 ( .A(n4320), .B(n4321), .Z(N117) );
  NANDN U4910 ( .A(n4319), .B(n4318), .Z(n4323) );
  NANDN U4911 ( .A(n4321), .B(n4320), .Z(n4322) );
  NAND U4912 ( .A(n4323), .B(n4322), .Z(n4435) );
  NAND U4913 ( .A(n4325), .B(n4324), .Z(n4329) );
  OR U4914 ( .A(n4327), .B(n4326), .Z(n4328) );
  NAND U4915 ( .A(n4329), .B(n4328), .Z(n4436) );
  XNOR U4916 ( .A(n4435), .B(n4436), .Z(n4437) );
  NANDN U4917 ( .A(n4331), .B(n4330), .Z(n4335) );
  NANDN U4918 ( .A(n4333), .B(n4332), .Z(n4334) );
  NAND U4919 ( .A(n4335), .B(n4334), .Z(n4456) );
  NANDN U4920 ( .A(n4337), .B(n4336), .Z(n4341) );
  NANDN U4921 ( .A(n4339), .B(n4338), .Z(n4340) );
  NAND U4922 ( .A(n4341), .B(n4340), .Z(n4453) );
  NANDN U4923 ( .A(n4343), .B(n4342), .Z(n4347) );
  NANDN U4924 ( .A(n4345), .B(n4344), .Z(n4346) );
  AND U4925 ( .A(n4347), .B(n4346), .Z(n4462) );
  NANDN U4926 ( .A(n4349), .B(n4348), .Z(n4353) );
  OR U4927 ( .A(n4351), .B(n4350), .Z(n4352) );
  AND U4928 ( .A(n4353), .B(n4352), .Z(n4460) );
  NOR U4929 ( .A(n169), .B(n4926), .Z(n5179) );
  NAND U4930 ( .A(n5179), .B(n4354), .Z(n4358) );
  OR U4931 ( .A(n4356), .B(n4355), .Z(n4357) );
  AND U4932 ( .A(n4358), .B(n4357), .Z(n4468) );
  AND U4933 ( .A(y[688]), .B(x[133]), .Z(n4541) );
  NAND U4934 ( .A(x[144]), .B(y[677]), .Z(n4542) );
  XOR U4935 ( .A(n4541), .B(n4542), .Z(n4544) );
  NAND U4936 ( .A(y[678]), .B(x[143]), .Z(n4543) );
  XOR U4937 ( .A(n4544), .B(n4543), .Z(n4547) );
  ANDN U4938 ( .B(y[683]), .A(n166), .Z(n5173) );
  NAND U4939 ( .A(n4359), .B(n5173), .Z(n4363) );
  OR U4940 ( .A(n4361), .B(n4360), .Z(n4362) );
  NAND U4941 ( .A(n4363), .B(n4362), .Z(n4548) );
  XNOR U4942 ( .A(n4547), .B(n4548), .Z(n4550) );
  NAND U4943 ( .A(y[693]), .B(x[128]), .Z(n4523) );
  NANDN U4944 ( .A(n4364), .B(o[52]), .Z(n4521) );
  NAND U4945 ( .A(y[672]), .B(x[149]), .Z(n4522) );
  XNOR U4946 ( .A(n4521), .B(n4522), .Z(n4524) );
  XOR U4947 ( .A(n4523), .B(n4524), .Z(n4549) );
  XNOR U4948 ( .A(n4550), .B(n4549), .Z(n4465) );
  ANDN U4949 ( .B(y[691]), .A(n162), .Z(n5869) );
  NANDN U4950 ( .A(n4365), .B(n5869), .Z(n4369) );
  NANDN U4951 ( .A(n4367), .B(n4366), .Z(n4368) );
  AND U4952 ( .A(n4369), .B(n4368), .Z(n4466) );
  XNOR U4953 ( .A(n4465), .B(n4466), .Z(n4467) );
  XNOR U4954 ( .A(n4468), .B(n4467), .Z(n4459) );
  XNOR U4955 ( .A(n4460), .B(n4459), .Z(n4461) );
  XNOR U4956 ( .A(n4462), .B(n4461), .Z(n4454) );
  XOR U4957 ( .A(n4453), .B(n4454), .Z(n4455) );
  XNOR U4958 ( .A(n4456), .B(n4455), .Z(n4449) );
  NANDN U4959 ( .A(n4371), .B(n4370), .Z(n4375) );
  OR U4960 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U4961 ( .A(n4375), .B(n4374), .Z(n4555) );
  OR U4962 ( .A(n4377), .B(n4376), .Z(n4381) );
  NAND U4963 ( .A(n4379), .B(n4378), .Z(n4380) );
  AND U4964 ( .A(n4381), .B(n4380), .Z(n4559) );
  NANDN U4965 ( .A(n4383), .B(n4382), .Z(n4387) );
  OR U4966 ( .A(n4385), .B(n4384), .Z(n4386) );
  NAND U4967 ( .A(n4387), .B(n4386), .Z(n4560) );
  XOR U4968 ( .A(n4559), .B(n4560), .Z(n4561) );
  NAND U4969 ( .A(n4389), .B(n4388), .Z(n4393) );
  OR U4970 ( .A(n4391), .B(n4390), .Z(n4392) );
  NAND U4971 ( .A(n4393), .B(n4392), .Z(n4562) );
  NANDN U4972 ( .A(n4395), .B(n4394), .Z(n4399) );
  NANDN U4973 ( .A(n4397), .B(n4396), .Z(n4398) );
  NAND U4974 ( .A(n4399), .B(n4398), .Z(n4471) );
  NAND U4975 ( .A(n4400), .B(n4541), .Z(n4404) );
  OR U4976 ( .A(n4402), .B(n4401), .Z(n4403) );
  AND U4977 ( .A(n4404), .B(n4403), .Z(n4472) );
  ANDN U4978 ( .B(y[687]), .A(n157), .Z(n4515) );
  ANDN U4979 ( .B(y[686]), .A(n158), .Z(n4597) );
  ANDN U4980 ( .B(y[679]), .A(n165), .Z(n4514) );
  XNOR U4981 ( .A(n4597), .B(n4514), .Z(n4516) );
  XNOR U4982 ( .A(n4515), .B(n4516), .Z(n4491) );
  ANDN U4983 ( .B(y[685]), .A(n159), .Z(n4891) );
  XOR U4984 ( .A(n4489), .B(n4891), .Z(n4490) );
  XNOR U4985 ( .A(n4491), .B(n4490), .Z(n4510) );
  NAND U4986 ( .A(x[132]), .B(y[689]), .Z(n4536) );
  AND U4987 ( .A(y[690]), .B(x[131]), .Z(n4406) );
  AND U4988 ( .A(x[141]), .B(y[680]), .Z(n4405) );
  XNOR U4989 ( .A(n4406), .B(n4405), .Z(n4535) );
  XOR U4990 ( .A(n4536), .B(n4535), .Z(n4508) );
  ANDN U4991 ( .B(y[681]), .A(n163), .Z(n4496) );
  ANDN U4992 ( .B(y[691]), .A(n153), .Z(n4494) );
  ANDN U4993 ( .B(y[676]), .A(n168), .Z(n4495) );
  XNOR U4994 ( .A(n4494), .B(n4495), .Z(n4497) );
  XOR U4995 ( .A(n4496), .B(n4497), .Z(n4509) );
  XOR U4996 ( .A(n4508), .B(n4509), .Z(n4511) );
  XNOR U4997 ( .A(n4510), .B(n4511), .Z(n4474) );
  XNOR U4998 ( .A(n4473), .B(n4474), .Z(n4486) );
  NAND U4999 ( .A(x[139]), .B(y[682]), .Z(n4505) );
  NAND U5000 ( .A(x[148]), .B(y[673]), .Z(n4533) );
  XOR U5001 ( .A(o[53]), .B(n4533), .Z(n4503) );
  NAND U5002 ( .A(x[147]), .B(y[674]), .Z(n4502) );
  XNOR U5003 ( .A(n4503), .B(n4502), .Z(n4504) );
  XNOR U5004 ( .A(n4505), .B(n4504), .Z(n4478) );
  ANDN U5005 ( .B(y[692]), .A(n152), .Z(n4528) );
  NAND U5006 ( .A(y[675]), .B(x[146]), .Z(n4527) );
  XOR U5007 ( .A(n4528), .B(n4527), .Z(n4529) );
  XOR U5008 ( .A(n4530), .B(n4529), .Z(n4477) );
  XOR U5009 ( .A(n4478), .B(n4477), .Z(n4479) );
  AND U5010 ( .A(x[141]), .B(y[689]), .Z(n5751) );
  NAND U5011 ( .A(n5751), .B(n4407), .Z(n4411) );
  OR U5012 ( .A(n4409), .B(n4408), .Z(n4410) );
  AND U5013 ( .A(n4411), .B(n4410), .Z(n4480) );
  XOR U5014 ( .A(n4479), .B(n4480), .Z(n4483) );
  NAND U5015 ( .A(n4412), .B(n5168), .Z(n4416) );
  OR U5016 ( .A(n4414), .B(n4413), .Z(n4415) );
  NAND U5017 ( .A(n4416), .B(n4415), .Z(n4484) );
  XOR U5018 ( .A(n4486), .B(n4485), .Z(n4553) );
  XOR U5019 ( .A(n4554), .B(n4553), .Z(n4556) );
  XOR U5020 ( .A(n4555), .B(n4556), .Z(n4447) );
  NANDN U5021 ( .A(n4418), .B(n4417), .Z(n4422) );
  OR U5022 ( .A(n4420), .B(n4419), .Z(n4421) );
  NAND U5023 ( .A(n4422), .B(n4421), .Z(n4448) );
  XOR U5024 ( .A(n4447), .B(n4448), .Z(n4450) );
  XNOR U5025 ( .A(n4449), .B(n4450), .Z(n4444) );
  OR U5026 ( .A(n4424), .B(n4423), .Z(n4428) );
  OR U5027 ( .A(n4426), .B(n4425), .Z(n4427) );
  NAND U5028 ( .A(n4428), .B(n4427), .Z(n4442) );
  OR U5029 ( .A(n4430), .B(n4429), .Z(n4434) );
  NANDN U5030 ( .A(n4432), .B(n4431), .Z(n4433) );
  NAND U5031 ( .A(n4434), .B(n4433), .Z(n4441) );
  XOR U5032 ( .A(n4442), .B(n4441), .Z(n4443) );
  XOR U5033 ( .A(n4444), .B(n4443), .Z(n4438) );
  XOR U5034 ( .A(n4437), .B(n4438), .Z(N118) );
  NANDN U5035 ( .A(n4436), .B(n4435), .Z(n4440) );
  NANDN U5036 ( .A(n4438), .B(n4437), .Z(n4439) );
  NAND U5037 ( .A(n4440), .B(n4439), .Z(n4565) );
  OR U5038 ( .A(n4442), .B(n4441), .Z(n4446) );
  NANDN U5039 ( .A(n4444), .B(n4443), .Z(n4445) );
  AND U5040 ( .A(n4446), .B(n4445), .Z(n4566) );
  XNOR U5041 ( .A(n4565), .B(n4566), .Z(n4567) );
  NANDN U5042 ( .A(n4448), .B(n4447), .Z(n4452) );
  NANDN U5043 ( .A(n4450), .B(n4449), .Z(n4451) );
  NAND U5044 ( .A(n4452), .B(n4451), .Z(n4574) );
  NANDN U5045 ( .A(n4454), .B(n4453), .Z(n4458) );
  OR U5046 ( .A(n4456), .B(n4455), .Z(n4457) );
  NAND U5047 ( .A(n4458), .B(n4457), .Z(n4572) );
  NANDN U5048 ( .A(n4460), .B(n4459), .Z(n4464) );
  NANDN U5049 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U5050 ( .A(n4464), .B(n4463), .Z(n4578) );
  NANDN U5051 ( .A(n4466), .B(n4465), .Z(n4470) );
  NANDN U5052 ( .A(n4468), .B(n4467), .Z(n4469) );
  NAND U5053 ( .A(n4470), .B(n4469), .Z(n4673) );
  NANDN U5054 ( .A(n4472), .B(n4471), .Z(n4476) );
  NANDN U5055 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U5056 ( .A(n4476), .B(n4475), .Z(n4671) );
  OR U5057 ( .A(n4478), .B(n4477), .Z(n4482) );
  NANDN U5058 ( .A(n4480), .B(n4479), .Z(n4481) );
  NAND U5059 ( .A(n4482), .B(n4481), .Z(n4670) );
  XOR U5060 ( .A(n4671), .B(n4670), .Z(n4672) );
  XOR U5061 ( .A(n4578), .B(n4577), .Z(n4580) );
  NANDN U5062 ( .A(n4484), .B(n4483), .Z(n4488) );
  OR U5063 ( .A(n4486), .B(n4485), .Z(n4487) );
  NAND U5064 ( .A(n4488), .B(n4487), .Z(n4679) );
  OR U5065 ( .A(n4891), .B(n4489), .Z(n4493) );
  NANDN U5066 ( .A(n4491), .B(n4490), .Z(n4492) );
  AND U5067 ( .A(n4493), .B(n4492), .Z(n4696) );
  OR U5068 ( .A(n4495), .B(n4494), .Z(n4499) );
  OR U5069 ( .A(n4497), .B(n4496), .Z(n4498) );
  NAND U5070 ( .A(n4499), .B(n4498), .Z(n4667) );
  AND U5071 ( .A(x[140]), .B(y[682]), .Z(n4501) );
  NAND U5072 ( .A(x[146]), .B(y[676]), .Z(n4500) );
  XOR U5073 ( .A(n4501), .B(n4500), .Z(n4605) );
  NAND U5074 ( .A(x[132]), .B(y[690]), .Z(n4604) );
  XOR U5075 ( .A(n4605), .B(n4604), .Z(n4664) );
  NAND U5076 ( .A(x[133]), .B(y[689]), .Z(n4621) );
  NAND U5077 ( .A(x[145]), .B(y[677]), .Z(n4620) );
  XOR U5078 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U5079 ( .A(y[678]), .B(x[144]), .Z(n4623) );
  XOR U5080 ( .A(n4622), .B(n4623), .Z(n4665) );
  XOR U5081 ( .A(n4667), .B(n4666), .Z(n4694) );
  OR U5082 ( .A(n4503), .B(n4502), .Z(n4507) );
  OR U5083 ( .A(n4505), .B(n4504), .Z(n4506) );
  NAND U5084 ( .A(n4507), .B(n4506), .Z(n4695) );
  XNOR U5085 ( .A(n4694), .B(n4695), .Z(n4697) );
  XOR U5086 ( .A(n4696), .B(n4697), .Z(n4677) );
  NANDN U5087 ( .A(n4509), .B(n4508), .Z(n4513) );
  OR U5088 ( .A(n4511), .B(n4510), .Z(n4512) );
  NAND U5089 ( .A(n4513), .B(n4512), .Z(n4683) );
  OR U5090 ( .A(n4514), .B(n4597), .Z(n4518) );
  OR U5091 ( .A(n4516), .B(n4515), .Z(n4517) );
  NAND U5092 ( .A(n4518), .B(n4517), .Z(n4635) );
  AND U5093 ( .A(y[686]), .B(x[136]), .Z(n4520) );
  NAND U5094 ( .A(x[135]), .B(y[687]), .Z(n4519) );
  XNOR U5095 ( .A(n4520), .B(n4519), .Z(n4600) );
  XNOR U5096 ( .A(n4599), .B(n4600), .Z(n4633) );
  NAND U5097 ( .A(x[128]), .B(y[694]), .Z(n4609) );
  NAND U5098 ( .A(y[672]), .B(x[150]), .Z(n4608) );
  XOR U5099 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U5100 ( .A(x[149]), .B(y[673]), .Z(n4626) );
  XOR U5101 ( .A(o[54]), .B(n4626), .Z(n4611) );
  XOR U5102 ( .A(n4610), .B(n4611), .Z(n4632) );
  XOR U5103 ( .A(n4633), .B(n4632), .Z(n4634) );
  XNOR U5104 ( .A(n4635), .B(n4634), .Z(n4647) );
  NAND U5105 ( .A(n4522), .B(n4521), .Z(n4526) );
  NANDN U5106 ( .A(n4524), .B(n4523), .Z(n4525) );
  AND U5107 ( .A(n4526), .B(n4525), .Z(n4644) );
  NANDN U5108 ( .A(n4528), .B(n4527), .Z(n4532) );
  OR U5109 ( .A(n4530), .B(n4529), .Z(n4531) );
  AND U5110 ( .A(n4532), .B(n4531), .Z(n4645) );
  XOR U5111 ( .A(n4644), .B(n4645), .Z(n4646) );
  NAND U5112 ( .A(x[142]), .B(y[680]), .Z(n4651) );
  NAND U5113 ( .A(x[131]), .B(y[691]), .Z(n4650) );
  XOR U5114 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U5115 ( .A(y[675]), .B(x[147]), .Z(n4653) );
  XOR U5116 ( .A(n4652), .B(n4653), .Z(n4639) );
  NANDN U5117 ( .A(n4533), .B(o[53]), .Z(n4659) );
  NAND U5118 ( .A(y[693]), .B(x[129]), .Z(n4657) );
  XOR U5119 ( .A(n4656), .B(n4657), .Z(n4658) );
  XNOR U5120 ( .A(n4659), .B(n4658), .Z(n4638) );
  XNOR U5121 ( .A(n4639), .B(n4638), .Z(n4641) );
  ANDN U5122 ( .B(y[690]), .A(n164), .Z(n5959) );
  NAND U5123 ( .A(n4534), .B(n5959), .Z(n4538) );
  OR U5124 ( .A(n4536), .B(n4535), .Z(n4537) );
  AND U5125 ( .A(n4538), .B(n4537), .Z(n4640) );
  XNOR U5126 ( .A(n4641), .B(n4640), .Z(n4689) );
  NAND U5127 ( .A(x[148]), .B(y[674]), .Z(n4615) );
  NAND U5128 ( .A(y[692]), .B(x[130]), .Z(n4614) );
  XOR U5129 ( .A(n4615), .B(n4614), .Z(n4616) );
  NAND U5130 ( .A(x[141]), .B(y[681]), .Z(n4617) );
  XOR U5131 ( .A(n4616), .B(n4617), .Z(n4592) );
  AND U5132 ( .A(y[688]), .B(x[134]), .Z(n4540) );
  NAND U5133 ( .A(x[138]), .B(y[684]), .Z(n4539) );
  XOR U5134 ( .A(n4540), .B(n4539), .Z(n4629) );
  NAND U5135 ( .A(x[143]), .B(y[679]), .Z(n4628) );
  XNOR U5136 ( .A(n4629), .B(n4628), .Z(n4589) );
  NANDN U5137 ( .A(n4542), .B(n4541), .Z(n4546) );
  OR U5138 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U5139 ( .A(n4546), .B(n4545), .Z(n4590) );
  XOR U5140 ( .A(n4592), .B(n4591), .Z(n4688) );
  XNOR U5141 ( .A(n4689), .B(n4688), .Z(n4691) );
  XOR U5142 ( .A(n4690), .B(n4691), .Z(n4682) );
  XNOR U5143 ( .A(n4683), .B(n4682), .Z(n4685) );
  OR U5144 ( .A(n4548), .B(n4547), .Z(n4552) );
  OR U5145 ( .A(n4550), .B(n4549), .Z(n4551) );
  AND U5146 ( .A(n4552), .B(n4551), .Z(n4684) );
  XNOR U5147 ( .A(n4685), .B(n4684), .Z(n4676) );
  XOR U5148 ( .A(n4677), .B(n4676), .Z(n4678) );
  XOR U5149 ( .A(n4679), .B(n4678), .Z(n4579) );
  XNOR U5150 ( .A(n4580), .B(n4579), .Z(n4585) );
  NANDN U5151 ( .A(n4554), .B(n4553), .Z(n4558) );
  NANDN U5152 ( .A(n4556), .B(n4555), .Z(n4557) );
  NAND U5153 ( .A(n4558), .B(n4557), .Z(n4584) );
  OR U5154 ( .A(n4560), .B(n4559), .Z(n4564) );
  NANDN U5155 ( .A(n4562), .B(n4561), .Z(n4563) );
  NAND U5156 ( .A(n4564), .B(n4563), .Z(n4583) );
  XOR U5157 ( .A(n4584), .B(n4583), .Z(n4586) );
  XNOR U5158 ( .A(n4585), .B(n4586), .Z(n4571) );
  XOR U5159 ( .A(n4572), .B(n4571), .Z(n4573) );
  XOR U5160 ( .A(n4574), .B(n4573), .Z(n4568) );
  XOR U5161 ( .A(n4567), .B(n4568), .Z(N119) );
  NANDN U5162 ( .A(n4566), .B(n4565), .Z(n4570) );
  NANDN U5163 ( .A(n4568), .B(n4567), .Z(n4569) );
  NAND U5164 ( .A(n4570), .B(n4569), .Z(n4700) );
  OR U5165 ( .A(n4572), .B(n4571), .Z(n4576) );
  NAND U5166 ( .A(n4574), .B(n4573), .Z(n4575) );
  NAND U5167 ( .A(n4576), .B(n4575), .Z(n4701) );
  XNOR U5168 ( .A(n4700), .B(n4701), .Z(n4702) );
  NANDN U5169 ( .A(n4578), .B(n4577), .Z(n4582) );
  OR U5170 ( .A(n4580), .B(n4579), .Z(n4581) );
  AND U5171 ( .A(n4582), .B(n4581), .Z(n4706) );
  OR U5172 ( .A(n4584), .B(n4583), .Z(n4588) );
  NAND U5173 ( .A(n4586), .B(n4585), .Z(n4587) );
  NAND U5174 ( .A(n4588), .B(n4587), .Z(n4707) );
  XOR U5175 ( .A(n4706), .B(n4707), .Z(n4709) );
  NANDN U5176 ( .A(n4590), .B(n4589), .Z(n4594) );
  NAND U5177 ( .A(n4592), .B(n4591), .Z(n4593) );
  NAND U5178 ( .A(n4594), .B(n4593), .Z(n4737) );
  NAND U5179 ( .A(x[128]), .B(y[695]), .Z(n4752) );
  NAND U5180 ( .A(y[672]), .B(x[151]), .Z(n4751) );
  XOR U5181 ( .A(n4752), .B(n4751), .Z(n4754) );
  AND U5182 ( .A(y[673]), .B(x[150]), .Z(n4780) );
  XOR U5183 ( .A(o[55]), .B(n4780), .Z(n4753) );
  ANDN U5184 ( .B(y[676]), .A(n170), .Z(n4934) );
  AND U5185 ( .A(x[148]), .B(y[675]), .Z(n4596) );
  NAND U5186 ( .A(x[144]), .B(y[679]), .Z(n4595) );
  XOR U5187 ( .A(n4596), .B(n4595), .Z(n4777) );
  XOR U5188 ( .A(n4934), .B(n4777), .Z(n4835) );
  NANDN U5189 ( .A(n4598), .B(n4597), .Z(n4602) );
  NAND U5190 ( .A(n4600), .B(n4599), .Z(n4601) );
  NAND U5191 ( .A(n4602), .B(n4601), .Z(n4836) );
  NAND U5192 ( .A(n5530), .B(n4603), .Z(n4607) );
  OR U5193 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U5194 ( .A(n4607), .B(n4606), .Z(n4829) );
  OR U5195 ( .A(n4609), .B(n4608), .Z(n4613) );
  NANDN U5196 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U5197 ( .A(n4613), .B(n4612), .Z(n4830) );
  XOR U5198 ( .A(n4737), .B(n4736), .Z(n4739) );
  OR U5199 ( .A(n4615), .B(n4614), .Z(n4619) );
  NANDN U5200 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U5201 ( .A(n4619), .B(n4618), .Z(n4743) );
  NAND U5202 ( .A(x[141]), .B(y[682]), .Z(n4812) );
  NAND U5203 ( .A(y[693]), .B(x[130]), .Z(n4811) );
  XOR U5204 ( .A(n4812), .B(n4811), .Z(n4813) );
  NAND U5205 ( .A(x[149]), .B(y[674]), .Z(n4814) );
  XOR U5206 ( .A(n4813), .B(n4814), .Z(n4820) );
  OR U5207 ( .A(n4621), .B(n4620), .Z(n4625) );
  NANDN U5208 ( .A(n4623), .B(n4622), .Z(n4624) );
  AND U5209 ( .A(n4625), .B(n4624), .Z(n4817) );
  NANDN U5210 ( .A(n4626), .B(o[54]), .Z(n4760) );
  NAND U5211 ( .A(x[140]), .B(y[683]), .Z(n4758) );
  NAND U5212 ( .A(x[129]), .B(y[694]), .Z(n4757) );
  XOR U5213 ( .A(n4758), .B(n4757), .Z(n4759) );
  XOR U5214 ( .A(n4760), .B(n4759), .Z(n4818) );
  XOR U5215 ( .A(n4817), .B(n4818), .Z(n4819) );
  XNOR U5216 ( .A(n4820), .B(n4819), .Z(n4742) );
  XNOR U5217 ( .A(n4743), .B(n4742), .Z(n4745) );
  AND U5218 ( .A(y[688]), .B(x[138]), .Z(n5209) );
  NAND U5219 ( .A(n4627), .B(n5209), .Z(n4631) );
  OR U5220 ( .A(n4629), .B(n4628), .Z(n4630) );
  AND U5221 ( .A(n4631), .B(n4630), .Z(n4826) );
  NAND U5222 ( .A(y[692]), .B(x[131]), .Z(n4806) );
  XOR U5223 ( .A(n4805), .B(n4806), .Z(n4808) );
  NAND U5224 ( .A(x[132]), .B(y[691]), .Z(n4807) );
  XOR U5225 ( .A(n4808), .B(n4807), .Z(n4824) );
  NAND U5226 ( .A(x[133]), .B(y[690]), .Z(n4800) );
  NAND U5227 ( .A(x[146]), .B(y[677]), .Z(n4799) );
  XOR U5228 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U5229 ( .A(y[678]), .B(x[145]), .Z(n4802) );
  XNOR U5230 ( .A(n4801), .B(n4802), .Z(n4823) );
  XNOR U5231 ( .A(n4826), .B(n4825), .Z(n4744) );
  XNOR U5232 ( .A(n4745), .B(n4744), .Z(n4738) );
  XNOR U5233 ( .A(n4739), .B(n4738), .Z(n4724) );
  OR U5234 ( .A(n4633), .B(n4632), .Z(n4637) );
  NANDN U5235 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U5236 ( .A(n4637), .B(n4636), .Z(n4781) );
  OR U5237 ( .A(n4639), .B(n4638), .Z(n4643) );
  OR U5238 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U5239 ( .A(n4643), .B(n4642), .Z(n4782) );
  XOR U5240 ( .A(n4781), .B(n4782), .Z(n4783) );
  OR U5241 ( .A(n4645), .B(n4644), .Z(n4649) );
  NANDN U5242 ( .A(n4647), .B(n4646), .Z(n4648) );
  NAND U5243 ( .A(n4649), .B(n4648), .Z(n4784) );
  OR U5244 ( .A(n4651), .B(n4650), .Z(n4655) );
  NANDN U5245 ( .A(n4653), .B(n4652), .Z(n4654) );
  NAND U5246 ( .A(n4655), .B(n4654), .Z(n4787) );
  NANDN U5247 ( .A(n4657), .B(n4656), .Z(n4661) );
  OR U5248 ( .A(n4659), .B(n4658), .Z(n4660) );
  AND U5249 ( .A(n4661), .B(n4660), .Z(n4788) );
  AND U5250 ( .A(x[136]), .B(y[687]), .Z(n4663) );
  NAND U5251 ( .A(x[137]), .B(y[686]), .Z(n4662) );
  XOR U5252 ( .A(n4663), .B(n4662), .Z(n4766) );
  NAND U5253 ( .A(x[135]), .B(y[688]), .Z(n4765) );
  XOR U5254 ( .A(n4766), .B(n4765), .Z(n4793) );
  NAND U5255 ( .A(y[685]), .B(x[138]), .Z(n4794) );
  XNOR U5256 ( .A(n4793), .B(n4794), .Z(n4795) );
  NAND U5257 ( .A(x[134]), .B(y[689]), .Z(n4770) );
  NAND U5258 ( .A(y[680]), .B(x[143]), .Z(n4769) );
  XOR U5259 ( .A(n4770), .B(n4769), .Z(n4772) );
  XNOR U5260 ( .A(n4771), .B(n4772), .Z(n4796) );
  XNOR U5261 ( .A(n4795), .B(n4796), .Z(n4789) );
  NANDN U5262 ( .A(n4665), .B(n4664), .Z(n4669) );
  OR U5263 ( .A(n4667), .B(n4666), .Z(n4668) );
  AND U5264 ( .A(n4669), .B(n4668), .Z(n4713) );
  XOR U5265 ( .A(n4712), .B(n4713), .Z(n4714) );
  XNOR U5266 ( .A(n4715), .B(n4714), .Z(n4725) );
  XOR U5267 ( .A(n4724), .B(n4725), .Z(n4727) );
  OR U5268 ( .A(n4671), .B(n4670), .Z(n4675) );
  NANDN U5269 ( .A(n4673), .B(n4672), .Z(n4674) );
  NAND U5270 ( .A(n4675), .B(n4674), .Z(n4726) );
  XNOR U5271 ( .A(n4727), .B(n4726), .Z(n4732) );
  NANDN U5272 ( .A(n4677), .B(n4676), .Z(n4681) );
  OR U5273 ( .A(n4679), .B(n4678), .Z(n4680) );
  NAND U5274 ( .A(n4681), .B(n4680), .Z(n4731) );
  OR U5275 ( .A(n4683), .B(n4682), .Z(n4687) );
  OR U5276 ( .A(n4685), .B(n4684), .Z(n4686) );
  AND U5277 ( .A(n4687), .B(n4686), .Z(n4721) );
  OR U5278 ( .A(n4689), .B(n4688), .Z(n4693) );
  OR U5279 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U5280 ( .A(n4693), .B(n4692), .Z(n4719) );
  OR U5281 ( .A(n4695), .B(n4694), .Z(n4699) );
  OR U5282 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U5283 ( .A(n4699), .B(n4698), .Z(n4718) );
  XOR U5284 ( .A(n4719), .B(n4718), .Z(n4720) );
  XOR U5285 ( .A(n4731), .B(n4730), .Z(n4733) );
  XNOR U5286 ( .A(n4709), .B(n4708), .Z(n4703) );
  XOR U5287 ( .A(n4702), .B(n4703), .Z(N120) );
  NANDN U5288 ( .A(n4701), .B(n4700), .Z(n4705) );
  NANDN U5289 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U5290 ( .A(n4705), .B(n4704), .Z(n4841) );
  OR U5291 ( .A(n4707), .B(n4706), .Z(n4711) );
  NAND U5292 ( .A(n4709), .B(n4708), .Z(n4710) );
  AND U5293 ( .A(n4711), .B(n4710), .Z(n4842) );
  XNOR U5294 ( .A(n4841), .B(n4842), .Z(n4843) );
  NANDN U5295 ( .A(n4713), .B(n4712), .Z(n4717) );
  OR U5296 ( .A(n4715), .B(n4714), .Z(n4716) );
  NAND U5297 ( .A(n4717), .B(n4716), .Z(n4977) );
  OR U5298 ( .A(n4719), .B(n4718), .Z(n4723) );
  NANDN U5299 ( .A(n4721), .B(n4720), .Z(n4722) );
  AND U5300 ( .A(n4723), .B(n4722), .Z(n4976) );
  XOR U5301 ( .A(n4977), .B(n4976), .Z(n4978) );
  NANDN U5302 ( .A(n4725), .B(n4724), .Z(n4729) );
  OR U5303 ( .A(n4727), .B(n4726), .Z(n4728) );
  NAND U5304 ( .A(n4729), .B(n4728), .Z(n4979) );
  OR U5305 ( .A(n4731), .B(n4730), .Z(n4735) );
  NAND U5306 ( .A(n4733), .B(n4732), .Z(n4734) );
  AND U5307 ( .A(n4735), .B(n4734), .Z(n4848) );
  NANDN U5308 ( .A(n4737), .B(n4736), .Z(n4741) );
  NANDN U5309 ( .A(n4739), .B(n4738), .Z(n4740) );
  NAND U5310 ( .A(n4741), .B(n4740), .Z(n4855) );
  NAND U5311 ( .A(n4743), .B(n4742), .Z(n4747) );
  NANDN U5312 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U5313 ( .A(n4747), .B(n4746), .Z(n4853) );
  AND U5314 ( .A(x[139]), .B(y[685]), .Z(n4749) );
  NAND U5315 ( .A(x[136]), .B(y[688]), .Z(n4748) );
  XOR U5316 ( .A(n4749), .B(n4748), .Z(n4893) );
  AND U5317 ( .A(x[142]), .B(y[682]), .Z(n4892) );
  XNOR U5318 ( .A(n4893), .B(n4892), .Z(n4887) );
  NOR U5319 ( .A(n160), .B(n4750), .Z(n4763) );
  IV U5320 ( .A(n4763), .Z(n4885) );
  NAND U5321 ( .A(x[138]), .B(y[686]), .Z(n4884) );
  XOR U5322 ( .A(n4885), .B(n4884), .Z(n4886) );
  XNOR U5323 ( .A(n4887), .B(n4886), .Z(n4898) );
  OR U5324 ( .A(n4752), .B(n4751), .Z(n4756) );
  NAND U5325 ( .A(n4754), .B(n4753), .Z(n4755) );
  NAND U5326 ( .A(n4756), .B(n4755), .Z(n4896) );
  NAND U5327 ( .A(x[143]), .B(y[681]), .Z(n4903) );
  NAND U5328 ( .A(y[693]), .B(x[131]), .Z(n4902) );
  XOR U5329 ( .A(n4903), .B(n4902), .Z(n4904) );
  NAND U5330 ( .A(y[692]), .B(x[132]), .Z(n4905) );
  XOR U5331 ( .A(n4904), .B(n4905), .Z(n4897) );
  XOR U5332 ( .A(n4898), .B(n4899), .Z(n4916) );
  OR U5333 ( .A(n4758), .B(n4757), .Z(n4762) );
  NANDN U5334 ( .A(n4760), .B(n4759), .Z(n4761) );
  AND U5335 ( .A(n4762), .B(n4761), .Z(n4961) );
  NANDN U5336 ( .A(n4764), .B(n4763), .Z(n4768) );
  OR U5337 ( .A(n4766), .B(n4765), .Z(n4767) );
  AND U5338 ( .A(n4768), .B(n4767), .Z(n4959) );
  OR U5339 ( .A(n4770), .B(n4769), .Z(n4774) );
  NAND U5340 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U5341 ( .A(n4774), .B(n4773), .Z(n4947) );
  NAND U5342 ( .A(x[134]), .B(y[690]), .Z(n4937) );
  AND U5343 ( .A(y[677]), .B(x[147]), .Z(n4775) );
  AND U5344 ( .A(y[676]), .B(x[148]), .Z(n5074) );
  XNOR U5345 ( .A(n4775), .B(n5074), .Z(n4936) );
  XOR U5346 ( .A(n4937), .B(n4936), .Z(n4946) );
  NAND U5347 ( .A(x[144]), .B(y[680]), .Z(n4931) );
  NAND U5348 ( .A(x[133]), .B(y[691]), .Z(n4929) );
  NAND U5349 ( .A(x[149]), .B(y[675]), .Z(n4928) );
  XNOR U5350 ( .A(n4929), .B(n4928), .Z(n4930) );
  XNOR U5351 ( .A(n4931), .B(n4930), .Z(n4948) );
  XOR U5352 ( .A(n4949), .B(n4948), .Z(n4958) );
  XNOR U5353 ( .A(n4959), .B(n4958), .Z(n4960) );
  XOR U5354 ( .A(n4961), .B(n4960), .Z(n4914) );
  NAND U5355 ( .A(x[130]), .B(y[694]), .Z(n4866) );
  NAND U5356 ( .A(x[150]), .B(y[674]), .Z(n4865) );
  XOR U5357 ( .A(n4866), .B(n4865), .Z(n4868) );
  XNOR U5358 ( .A(n4867), .B(n4868), .Z(n4955) );
  AND U5359 ( .A(y[675]), .B(x[144]), .Z(n4776) );
  AND U5360 ( .A(y[679]), .B(x[148]), .Z(n5342) );
  NAND U5361 ( .A(n4776), .B(n5342), .Z(n4779) );
  NANDN U5362 ( .A(n4777), .B(n4934), .Z(n4778) );
  AND U5363 ( .A(n4779), .B(n4778), .Z(n4953) );
  NAND U5364 ( .A(n4780), .B(o[55]), .Z(n4881) );
  NAND U5365 ( .A(x[129]), .B(y[695]), .Z(n4879) );
  XOR U5366 ( .A(n4878), .B(n4879), .Z(n4880) );
  XOR U5367 ( .A(n4881), .B(n4880), .Z(n4952) );
  XOR U5368 ( .A(n4955), .B(n4954), .Z(n4915) );
  XOR U5369 ( .A(n4914), .B(n4915), .Z(n4917) );
  XOR U5370 ( .A(n4916), .B(n4917), .Z(n4854) );
  XOR U5371 ( .A(n4855), .B(n4856), .Z(n4984) );
  OR U5372 ( .A(n4782), .B(n4781), .Z(n4786) );
  NANDN U5373 ( .A(n4784), .B(n4783), .Z(n4785) );
  NAND U5374 ( .A(n4786), .B(n4785), .Z(n4983) );
  NANDN U5375 ( .A(n4788), .B(n4787), .Z(n4792) );
  NAND U5376 ( .A(n4790), .B(n4789), .Z(n4791) );
  NAND U5377 ( .A(n4792), .B(n4791), .Z(n4861) );
  NANDN U5378 ( .A(n4794), .B(n4793), .Z(n4798) );
  NANDN U5379 ( .A(n4796), .B(n4795), .Z(n4797) );
  NAND U5380 ( .A(n4798), .B(n4797), .Z(n4859) );
  OR U5381 ( .A(n4800), .B(n4799), .Z(n4804) );
  NANDN U5382 ( .A(n4802), .B(n4801), .Z(n4803) );
  AND U5383 ( .A(n4804), .B(n4803), .Z(n4942) );
  NAND U5384 ( .A(x[146]), .B(y[678]), .Z(n4875) );
  NAND U5385 ( .A(x[145]), .B(y[679]), .Z(n4873) );
  NAND U5386 ( .A(y[689]), .B(x[135]), .Z(n4872) );
  XOR U5387 ( .A(n4873), .B(n4872), .Z(n4874) );
  XOR U5388 ( .A(n4875), .B(n4874), .Z(n4941) );
  ANDN U5389 ( .B(y[673]), .A(n174), .Z(n4871) );
  XOR U5390 ( .A(o[56]), .B(n4871), .Z(n4911) );
  NAND U5391 ( .A(x[128]), .B(y[696]), .Z(n4909) );
  NAND U5392 ( .A(y[672]), .B(x[152]), .Z(n4908) );
  XOR U5393 ( .A(n4909), .B(n4908), .Z(n4910) );
  XOR U5394 ( .A(n4941), .B(n4940), .Z(n4943) );
  XNOR U5395 ( .A(n4942), .B(n4943), .Z(n4967) );
  NANDN U5396 ( .A(n4806), .B(n4805), .Z(n4810) );
  OR U5397 ( .A(n4808), .B(n4807), .Z(n4809) );
  AND U5398 ( .A(n4810), .B(n4809), .Z(n4965) );
  OR U5399 ( .A(n4812), .B(n4811), .Z(n4816) );
  NANDN U5400 ( .A(n4814), .B(n4813), .Z(n4815) );
  AND U5401 ( .A(n4816), .B(n4815), .Z(n4964) );
  XNOR U5402 ( .A(n4965), .B(n4964), .Z(n4966) );
  XNOR U5403 ( .A(n4967), .B(n4966), .Z(n4860) );
  XOR U5404 ( .A(n4859), .B(n4860), .Z(n4862) );
  OR U5405 ( .A(n4818), .B(n4817), .Z(n4822) );
  NANDN U5406 ( .A(n4820), .B(n4819), .Z(n4821) );
  NAND U5407 ( .A(n4822), .B(n4821), .Z(n4970) );
  NAND U5408 ( .A(n4824), .B(n4823), .Z(n4828) );
  NANDN U5409 ( .A(n4826), .B(n4825), .Z(n4827) );
  NAND U5410 ( .A(n4828), .B(n4827), .Z(n4923) );
  NANDN U5411 ( .A(n4830), .B(n4829), .Z(n4834) );
  NAND U5412 ( .A(n4832), .B(n4831), .Z(n4833) );
  NAND U5413 ( .A(n4834), .B(n4833), .Z(n4920) );
  NANDN U5414 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U5415 ( .A(n4838), .B(n4837), .Z(n4839) );
  NAND U5416 ( .A(n4840), .B(n4839), .Z(n4921) );
  XNOR U5417 ( .A(n4923), .B(n4922), .Z(n4971) );
  XOR U5418 ( .A(n4972), .B(n4973), .Z(n4982) );
  XNOR U5419 ( .A(n4983), .B(n4982), .Z(n4985) );
  XNOR U5420 ( .A(n4984), .B(n4985), .Z(n4847) );
  XOR U5421 ( .A(n4848), .B(n4847), .Z(n4849) );
  XNOR U5422 ( .A(n4850), .B(n4849), .Z(n4844) );
  XOR U5423 ( .A(n4843), .B(n4844), .Z(N121) );
  NANDN U5424 ( .A(n4842), .B(n4841), .Z(n4846) );
  NANDN U5425 ( .A(n4844), .B(n4843), .Z(n4845) );
  NAND U5426 ( .A(n4846), .B(n4845), .Z(n4988) );
  NANDN U5427 ( .A(n4848), .B(n4847), .Z(n4852) );
  OR U5428 ( .A(n4850), .B(n4849), .Z(n4851) );
  AND U5429 ( .A(n4852), .B(n4851), .Z(n4989) );
  XNOR U5430 ( .A(n4988), .B(n4989), .Z(n4990) );
  NANDN U5431 ( .A(n4854), .B(n4853), .Z(n4858) );
  NANDN U5432 ( .A(n4856), .B(n4855), .Z(n4857) );
  NAND U5433 ( .A(n4858), .B(n4857), .Z(n5136) );
  NANDN U5434 ( .A(n4860), .B(n4859), .Z(n4864) );
  NANDN U5435 ( .A(n4862), .B(n4861), .Z(n4863) );
  NAND U5436 ( .A(n4864), .B(n4863), .Z(n5009) );
  OR U5437 ( .A(n4866), .B(n4865), .Z(n4870) );
  NAND U5438 ( .A(n4868), .B(n4867), .Z(n4869) );
  AND U5439 ( .A(n4870), .B(n4869), .Z(n5116) );
  IV U5440 ( .A(y[689]), .Z(n5570) );
  NANDN U5441 ( .A(n5570), .B(x[136]), .Z(n5111) );
  XNOR U5442 ( .A(n5111), .B(n5112), .Z(n5097) );
  AND U5443 ( .A(n4871), .B(o[56]), .Z(n5106) );
  NAND U5444 ( .A(x[128]), .B(y[697]), .Z(n5104) );
  XNOR U5445 ( .A(n5103), .B(n5104), .Z(n5105) );
  XOR U5446 ( .A(n5106), .B(n5105), .Z(n5098) );
  XNOR U5447 ( .A(n5097), .B(n5098), .Z(n5100) );
  OR U5448 ( .A(n4873), .B(n4872), .Z(n4877) );
  NANDN U5449 ( .A(n4875), .B(n4874), .Z(n4876) );
  AND U5450 ( .A(n4877), .B(n4876), .Z(n5099) );
  XOR U5451 ( .A(n5100), .B(n5099), .Z(n5115) );
  NANDN U5452 ( .A(n4879), .B(n4878), .Z(n4883) );
  OR U5453 ( .A(n4881), .B(n4880), .Z(n4882) );
  AND U5454 ( .A(n4883), .B(n4882), .Z(n5117) );
  XNOR U5455 ( .A(n5118), .B(n5117), .Z(n5123) );
  NAND U5456 ( .A(n4885), .B(n4884), .Z(n4889) );
  NANDN U5457 ( .A(n4887), .B(n4886), .Z(n4888) );
  AND U5458 ( .A(n4889), .B(n4888), .Z(n5121) );
  NANDN U5459 ( .A(n162), .B(y[686]), .Z(n5052) );
  NANDN U5460 ( .A(n4890), .B(x[140]), .Z(n5050) );
  NANDN U5461 ( .A(n158), .B(y[690]), .Z(n5051) );
  XNOR U5462 ( .A(n5050), .B(n5051), .Z(n5053) );
  XNOR U5463 ( .A(n5052), .B(n5053), .Z(n5043) );
  AND U5464 ( .A(y[688]), .B(x[139]), .Z(n5412) );
  NAND U5465 ( .A(n4891), .B(n5412), .Z(n4895) );
  NANDN U5466 ( .A(n4893), .B(n4892), .Z(n4894) );
  AND U5467 ( .A(n4895), .B(n4894), .Z(n5044) );
  XNOR U5468 ( .A(n5043), .B(n5044), .Z(n5046) );
  NAND U5469 ( .A(x[141]), .B(y[684]), .Z(n5037) );
  AND U5470 ( .A(y[696]), .B(x[129]), .Z(n5036) );
  XNOR U5471 ( .A(n5037), .B(n5036), .Z(n5038) );
  ANDN U5472 ( .B(y[673]), .A(n175), .Z(n5049) );
  XNOR U5473 ( .A(o[57]), .B(n5049), .Z(n5039) );
  XOR U5474 ( .A(n5038), .B(n5039), .Z(n5045) );
  XOR U5475 ( .A(n5046), .B(n5045), .Z(n5122) );
  XNOR U5476 ( .A(n5121), .B(n5122), .Z(n5124) );
  XNOR U5477 ( .A(n5123), .B(n5124), .Z(n5014) );
  NANDN U5478 ( .A(n4897), .B(n4896), .Z(n4901) );
  OR U5479 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U5480 ( .A(n4901), .B(n4900), .Z(n5012) );
  OR U5481 ( .A(n4903), .B(n4902), .Z(n4907) );
  NANDN U5482 ( .A(n4905), .B(n4904), .Z(n4906) );
  AND U5483 ( .A(n4907), .B(n4906), .Z(n5094) );
  OR U5484 ( .A(n4909), .B(n4908), .Z(n4913) );
  NAND U5485 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U5486 ( .A(n4913), .B(n4912), .Z(n5091) );
  NAND U5487 ( .A(x[130]), .B(y[695]), .Z(n5033) );
  NAND U5488 ( .A(x[131]), .B(y[694]), .Z(n5031) );
  XOR U5489 ( .A(n5033), .B(n5032), .Z(n5092) );
  XOR U5490 ( .A(n5091), .B(n5092), .Z(n5093) );
  XOR U5491 ( .A(n5014), .B(n5015), .Z(n5007) );
  NANDN U5492 ( .A(n4915), .B(n4914), .Z(n4919) );
  OR U5493 ( .A(n4917), .B(n4916), .Z(n4918) );
  AND U5494 ( .A(n4919), .B(n4918), .Z(n5006) );
  XOR U5495 ( .A(n5007), .B(n5006), .Z(n5008) );
  XOR U5496 ( .A(n5009), .B(n5008), .Z(n5133) );
  NANDN U5497 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U5498 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U5499 ( .A(n4925), .B(n4924), .Z(n5001) );
  NANDN U5500 ( .A(n145), .B(x[150]), .Z(n5058) );
  IV U5501 ( .A(y[692]), .Z(n5515) );
  NANDN U5502 ( .A(n5515), .B(x[133]), .Z(n5056) );
  NANDN U5503 ( .A(n4926), .B(x[145]), .Z(n5057) );
  XNOR U5504 ( .A(n5056), .B(n5057), .Z(n5059) );
  XNOR U5505 ( .A(n5058), .B(n5059), .Z(n5086) );
  NAND U5506 ( .A(x[147]), .B(y[678]), .Z(n5076) );
  AND U5507 ( .A(y[676]), .B(x[149]), .Z(n4927) );
  AND U5508 ( .A(y[677]), .B(x[148]), .Z(n4935) );
  XNOR U5509 ( .A(n4927), .B(n4935), .Z(n5075) );
  XOR U5510 ( .A(n5076), .B(n5075), .Z(n5085) );
  XOR U5511 ( .A(n5086), .B(n5085), .Z(n5088) );
  OR U5512 ( .A(n4929), .B(n4928), .Z(n4933) );
  OR U5513 ( .A(n4931), .B(n4930), .Z(n4932) );
  AND U5514 ( .A(n4933), .B(n4932), .Z(n5087) );
  XOR U5515 ( .A(n5088), .B(n5087), .Z(n5127) );
  AND U5516 ( .A(y[674]), .B(x[151]), .Z(n5064) );
  IV U5517 ( .A(y[693]), .Z(n5042) );
  NANDN U5518 ( .A(n5042), .B(x[132]), .Z(n5062) );
  XNOR U5519 ( .A(n5062), .B(n5063), .Z(n5065) );
  XNOR U5520 ( .A(n5064), .B(n5065), .Z(n5081) );
  AND U5521 ( .A(x[143]), .B(y[682]), .Z(n5070) );
  NANDN U5522 ( .A(n169), .B(y[679]), .Z(n5068) );
  NANDN U5523 ( .A(n157), .B(y[691]), .Z(n5069) );
  XNOR U5524 ( .A(n5068), .B(n5069), .Z(n5071) );
  XOR U5525 ( .A(n5070), .B(n5071), .Z(n5080) );
  NAND U5526 ( .A(n4935), .B(n4934), .Z(n4939) );
  OR U5527 ( .A(n4937), .B(n4936), .Z(n4938) );
  AND U5528 ( .A(n4939), .B(n4938), .Z(n5079) );
  XNOR U5529 ( .A(n5080), .B(n5079), .Z(n5082) );
  XOR U5530 ( .A(n5081), .B(n5082), .Z(n5128) );
  XOR U5531 ( .A(n5127), .B(n5128), .Z(n5130) );
  NANDN U5532 ( .A(n4941), .B(n4940), .Z(n4945) );
  OR U5533 ( .A(n4943), .B(n4942), .Z(n4944) );
  AND U5534 ( .A(n4945), .B(n4944), .Z(n5129) );
  XOR U5535 ( .A(n5130), .B(n5129), .Z(n5024) );
  NANDN U5536 ( .A(n4947), .B(n4946), .Z(n4951) );
  OR U5537 ( .A(n4949), .B(n4948), .Z(n4950) );
  NAND U5538 ( .A(n4951), .B(n4950), .Z(n5025) );
  XNOR U5539 ( .A(n5024), .B(n5025), .Z(n5027) );
  NANDN U5540 ( .A(n4953), .B(n4952), .Z(n4957) );
  OR U5541 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U5542 ( .A(n4957), .B(n4956), .Z(n5026) );
  XOR U5543 ( .A(n5027), .B(n5026), .Z(n5021) );
  NANDN U5544 ( .A(n4959), .B(n4958), .Z(n4963) );
  NANDN U5545 ( .A(n4961), .B(n4960), .Z(n4962) );
  NAND U5546 ( .A(n4963), .B(n4962), .Z(n5019) );
  OR U5547 ( .A(n4965), .B(n4964), .Z(n4969) );
  OR U5548 ( .A(n4967), .B(n4966), .Z(n4968) );
  AND U5549 ( .A(n4969), .B(n4968), .Z(n5018) );
  XNOR U5550 ( .A(n5001), .B(n5000), .Z(n5002) );
  NANDN U5551 ( .A(n4971), .B(n4970), .Z(n4975) );
  NAND U5552 ( .A(n4973), .B(n4972), .Z(n4974) );
  NAND U5553 ( .A(n4975), .B(n4974), .Z(n5003) );
  XNOR U5554 ( .A(n5002), .B(n5003), .Z(n5134) );
  XOR U5555 ( .A(n5136), .B(n5135), .Z(n4997) );
  OR U5556 ( .A(n4977), .B(n4976), .Z(n4981) );
  NANDN U5557 ( .A(n4979), .B(n4978), .Z(n4980) );
  AND U5558 ( .A(n4981), .B(n4980), .Z(n4994) );
  OR U5559 ( .A(n4983), .B(n4982), .Z(n4987) );
  NANDN U5560 ( .A(n4985), .B(n4984), .Z(n4986) );
  AND U5561 ( .A(n4987), .B(n4986), .Z(n4995) );
  XOR U5562 ( .A(n4994), .B(n4995), .Z(n4996) );
  XOR U5563 ( .A(n4997), .B(n4996), .Z(n4991) );
  XOR U5564 ( .A(n4990), .B(n4991), .Z(N122) );
  NANDN U5565 ( .A(n4989), .B(n4988), .Z(n4993) );
  NANDN U5566 ( .A(n4991), .B(n4990), .Z(n4992) );
  NAND U5567 ( .A(n4993), .B(n4992), .Z(n5139) );
  OR U5568 ( .A(n4995), .B(n4994), .Z(n4999) );
  NANDN U5569 ( .A(n4997), .B(n4996), .Z(n4998) );
  AND U5570 ( .A(n4999), .B(n4998), .Z(n5140) );
  XNOR U5571 ( .A(n5139), .B(n5140), .Z(n5141) );
  NANDN U5572 ( .A(n5001), .B(n5000), .Z(n5005) );
  NANDN U5573 ( .A(n5003), .B(n5002), .Z(n5004) );
  NAND U5574 ( .A(n5005), .B(n5004), .Z(n5148) );
  OR U5575 ( .A(n5007), .B(n5006), .Z(n5011) );
  NANDN U5576 ( .A(n5009), .B(n5008), .Z(n5010) );
  NAND U5577 ( .A(n5011), .B(n5010), .Z(n5280) );
  NANDN U5578 ( .A(n5013), .B(n5012), .Z(n5017) );
  OR U5579 ( .A(n5015), .B(n5014), .Z(n5016) );
  NAND U5580 ( .A(n5017), .B(n5016), .Z(n5281) );
  NANDN U5581 ( .A(n5019), .B(n5018), .Z(n5023) );
  NAND U5582 ( .A(n5021), .B(n5020), .Z(n5022) );
  AND U5583 ( .A(n5023), .B(n5022), .Z(n5286) );
  OR U5584 ( .A(n5025), .B(n5024), .Z(n5029) );
  OR U5585 ( .A(n5027), .B(n5026), .Z(n5028) );
  NAND U5586 ( .A(n5029), .B(n5028), .Z(n5192) );
  NANDN U5587 ( .A(n5031), .B(n5030), .Z(n5035) );
  NANDN U5588 ( .A(n5033), .B(n5032), .Z(n5034) );
  NAND U5589 ( .A(n5035), .B(n5034), .Z(n5184) );
  NANDN U5590 ( .A(n5037), .B(n5036), .Z(n5041) );
  NANDN U5591 ( .A(n5039), .B(n5038), .Z(n5040) );
  NAND U5592 ( .A(n5041), .B(n5040), .Z(n5183) );
  XOR U5593 ( .A(n5184), .B(n5183), .Z(n5185) );
  ANDN U5594 ( .B(y[691]), .A(n158), .Z(n5262) );
  NANDN U5595 ( .A(n163), .B(y[686]), .Z(n5207) );
  NANDN U5596 ( .A(n5042), .B(x[133]), .Z(n5208) );
  XNOR U5597 ( .A(n5207), .B(n5208), .Z(n5210) );
  XNOR U5598 ( .A(n5209), .B(n5210), .Z(n5263) );
  XNOR U5599 ( .A(n5262), .B(n5263), .Z(n5265) );
  NANDN U5600 ( .A(n5570), .B(x[137]), .Z(n5252) );
  NANDN U5601 ( .A(n5515), .B(x[134]), .Z(n5250) );
  NANDN U5602 ( .A(n159), .B(y[690]), .Z(n5251) );
  XNOR U5603 ( .A(n5250), .B(n5251), .Z(n5253) );
  XOR U5604 ( .A(n5252), .B(n5253), .Z(n5264) );
  XNOR U5605 ( .A(n5265), .B(n5264), .Z(n5186) );
  OR U5606 ( .A(n5044), .B(n5043), .Z(n5048) );
  OR U5607 ( .A(n5046), .B(n5045), .Z(n5047) );
  AND U5608 ( .A(n5048), .B(n5047), .Z(n5226) );
  XNOR U5609 ( .A(n5225), .B(n5226), .Z(n5228) );
  AND U5610 ( .A(n5049), .B(o[57]), .Z(n5239) );
  ANDN U5611 ( .B(y[684]), .A(n165), .Z(n5237) );
  ANDN U5612 ( .B(y[697]), .A(n152), .Z(n5238) );
  XNOR U5613 ( .A(n5237), .B(n5238), .Z(n5240) );
  XNOR U5614 ( .A(n5239), .B(n5240), .Z(n5219) );
  NAND U5615 ( .A(n5051), .B(n5050), .Z(n5055) );
  NANDN U5616 ( .A(n5053), .B(n5052), .Z(n5054) );
  NAND U5617 ( .A(n5055), .B(n5054), .Z(n5220) );
  XOR U5618 ( .A(n5219), .B(n5220), .Z(n5222) );
  NAND U5619 ( .A(x[128]), .B(y[698]), .Z(n5214) );
  AND U5620 ( .A(x[154]), .B(y[672]), .Z(n5213) );
  XNOR U5621 ( .A(n5214), .B(n5213), .Z(n5215) );
  AND U5622 ( .A(y[673]), .B(x[153]), .Z(n5249) );
  XNOR U5623 ( .A(o[58]), .B(n5249), .Z(n5216) );
  XOR U5624 ( .A(n5222), .B(n5221), .Z(n5160) );
  NAND U5625 ( .A(n5057), .B(n5056), .Z(n5061) );
  NANDN U5626 ( .A(n5059), .B(n5058), .Z(n5060) );
  AND U5627 ( .A(n5061), .B(n5060), .Z(n5157) );
  NAND U5628 ( .A(n5063), .B(n5062), .Z(n5067) );
  OR U5629 ( .A(n5065), .B(n5064), .Z(n5066) );
  AND U5630 ( .A(n5067), .B(n5066), .Z(n5158) );
  XOR U5631 ( .A(n5157), .B(n5158), .Z(n5159) );
  XOR U5632 ( .A(n5160), .B(n5159), .Z(n5197) );
  ANDN U5633 ( .B(y[694]), .A(n155), .Z(n5180) );
  XNOR U5634 ( .A(n5179), .B(n5180), .Z(n5182) );
  XNOR U5635 ( .A(n5181), .B(n5182), .Z(n5161) );
  NAND U5636 ( .A(n5069), .B(n5068), .Z(n5073) );
  OR U5637 ( .A(n5071), .B(n5070), .Z(n5072) );
  NAND U5638 ( .A(n5073), .B(n5072), .Z(n5162) );
  XOR U5639 ( .A(n5161), .B(n5162), .Z(n5164) );
  NAND U5640 ( .A(x[147]), .B(y[679]), .Z(n5257) );
  AND U5641 ( .A(x[139]), .B(y[687]), .Z(n5256) );
  XNOR U5642 ( .A(n5257), .B(n5256), .Z(n5258) );
  NAND U5643 ( .A(x[131]), .B(y[695]), .Z(n5259) );
  XOR U5644 ( .A(n5164), .B(n5163), .Z(n5196) );
  NAND U5645 ( .A(x[149]), .B(y[677]), .Z(n5243) );
  NANDN U5646 ( .A(n5243), .B(n5074), .Z(n5078) );
  OR U5647 ( .A(n5076), .B(n5075), .Z(n5077) );
  NAND U5648 ( .A(n5078), .B(n5077), .Z(n5152) );
  NAND U5649 ( .A(x[150]), .B(y[676]), .Z(n5170) );
  NAND U5650 ( .A(y[675]), .B(x[151]), .Z(n5167) );
  XNOR U5651 ( .A(n5168), .B(n5167), .Z(n5169) );
  XNOR U5652 ( .A(n5170), .B(n5169), .Z(n5151) );
  XNOR U5653 ( .A(n5152), .B(n5151), .Z(n5154) );
  NANDN U5654 ( .A(n146), .B(x[148]), .Z(n5245) );
  XOR U5655 ( .A(n5244), .B(n5243), .Z(n5246) );
  XOR U5656 ( .A(n5245), .B(n5246), .Z(n5153) );
  XOR U5657 ( .A(n5154), .B(n5153), .Z(n5195) );
  XNOR U5658 ( .A(n5196), .B(n5195), .Z(n5198) );
  XNOR U5659 ( .A(n5197), .B(n5198), .Z(n5227) );
  XOR U5660 ( .A(n5228), .B(n5227), .Z(n5190) );
  OR U5661 ( .A(n5080), .B(n5079), .Z(n5084) );
  NANDN U5662 ( .A(n5082), .B(n5081), .Z(n5083) );
  NAND U5663 ( .A(n5084), .B(n5083), .Z(n5275) );
  NANDN U5664 ( .A(n5086), .B(n5085), .Z(n5090) );
  OR U5665 ( .A(n5088), .B(n5087), .Z(n5089) );
  NAND U5666 ( .A(n5090), .B(n5089), .Z(n5274) );
  XOR U5667 ( .A(n5275), .B(n5274), .Z(n5276) );
  OR U5668 ( .A(n5092), .B(n5091), .Z(n5096) );
  NANDN U5669 ( .A(n5094), .B(n5093), .Z(n5095) );
  NAND U5670 ( .A(n5096), .B(n5095), .Z(n5277) );
  XNOR U5671 ( .A(n5276), .B(n5277), .Z(n5189) );
  XNOR U5672 ( .A(n5190), .B(n5189), .Z(n5191) );
  XOR U5673 ( .A(n5192), .B(n5191), .Z(n5287) );
  XOR U5674 ( .A(n5286), .B(n5287), .Z(n5288) );
  OR U5675 ( .A(n5098), .B(n5097), .Z(n5102) );
  OR U5676 ( .A(n5100), .B(n5099), .Z(n5101) );
  AND U5677 ( .A(n5102), .B(n5101), .Z(n5268) );
  NAND U5678 ( .A(x[130]), .B(y[696]), .Z(n5174) );
  XNOR U5679 ( .A(n5174), .B(n5173), .Z(n5176) );
  ANDN U5680 ( .B(y[674]), .A(n175), .Z(n5175) );
  XOR U5681 ( .A(n5176), .B(n5175), .Z(n5201) );
  NAND U5682 ( .A(n5104), .B(n5103), .Z(n5108) );
  OR U5683 ( .A(n5106), .B(n5105), .Z(n5107) );
  AND U5684 ( .A(n5108), .B(n5107), .Z(n5202) );
  XNOR U5685 ( .A(n5201), .B(n5202), .Z(n5204) );
  OR U5686 ( .A(n5110), .B(n5109), .Z(n5114) );
  NANDN U5687 ( .A(n5112), .B(n5111), .Z(n5113) );
  AND U5688 ( .A(n5114), .B(n5113), .Z(n5203) );
  XOR U5689 ( .A(n5204), .B(n5203), .Z(n5269) );
  XNOR U5690 ( .A(n5268), .B(n5269), .Z(n5271) );
  NANDN U5691 ( .A(n5116), .B(n5115), .Z(n5120) );
  OR U5692 ( .A(n5118), .B(n5117), .Z(n5119) );
  AND U5693 ( .A(n5120), .B(n5119), .Z(n5270) );
  XNOR U5694 ( .A(n5271), .B(n5270), .Z(n5233) );
  OR U5695 ( .A(n5122), .B(n5121), .Z(n5126) );
  NANDN U5696 ( .A(n5124), .B(n5123), .Z(n5125) );
  AND U5697 ( .A(n5126), .B(n5125), .Z(n5231) );
  NANDN U5698 ( .A(n5128), .B(n5127), .Z(n5132) );
  OR U5699 ( .A(n5130), .B(n5129), .Z(n5131) );
  NAND U5700 ( .A(n5132), .B(n5131), .Z(n5232) );
  XNOR U5701 ( .A(n5231), .B(n5232), .Z(n5234) );
  XOR U5702 ( .A(n5233), .B(n5234), .Z(n5289) );
  XOR U5703 ( .A(n5288), .B(n5289), .Z(n5283) );
  XOR U5704 ( .A(n5282), .B(n5283), .Z(n5145) );
  NANDN U5705 ( .A(n5134), .B(n5133), .Z(n5138) );
  NAND U5706 ( .A(n5136), .B(n5135), .Z(n5137) );
  AND U5707 ( .A(n5138), .B(n5137), .Z(n5146) );
  XNOR U5708 ( .A(n5148), .B(n5147), .Z(n5142) );
  XOR U5709 ( .A(n5141), .B(n5142), .Z(N123) );
  NANDN U5710 ( .A(n5140), .B(n5139), .Z(n5144) );
  NANDN U5711 ( .A(n5142), .B(n5141), .Z(n5143) );
  NAND U5712 ( .A(n5144), .B(n5143), .Z(n5292) );
  NANDN U5713 ( .A(n5146), .B(n5145), .Z(n5150) );
  NANDN U5714 ( .A(n5148), .B(n5147), .Z(n5149) );
  NAND U5715 ( .A(n5150), .B(n5149), .Z(n5293) );
  XNOR U5716 ( .A(n5292), .B(n5293), .Z(n5294) );
  OR U5717 ( .A(n5152), .B(n5151), .Z(n5156) );
  OR U5718 ( .A(n5154), .B(n5153), .Z(n5155) );
  NAND U5719 ( .A(n5156), .B(n5155), .Z(n5317) );
  NANDN U5720 ( .A(n5162), .B(n5161), .Z(n5166) );
  NANDN U5721 ( .A(n5164), .B(n5163), .Z(n5165) );
  NAND U5722 ( .A(n5166), .B(n5165), .Z(n5426) );
  NANDN U5723 ( .A(n5168), .B(n5167), .Z(n5172) );
  NAND U5724 ( .A(n5170), .B(n5169), .Z(n5171) );
  AND U5725 ( .A(n5172), .B(n5171), .Z(n5379) );
  NANDN U5726 ( .A(n5174), .B(n5173), .Z(n5178) );
  NAND U5727 ( .A(n5176), .B(n5175), .Z(n5177) );
  NAND U5728 ( .A(n5178), .B(n5177), .Z(n5380) );
  XOR U5729 ( .A(n5379), .B(n5380), .Z(n5381) );
  ANDN U5730 ( .B(y[690]), .A(n160), .Z(n5337) );
  ANDN U5731 ( .B(y[681]), .A(n169), .Z(n5335) );
  ANDN U5732 ( .B(y[678]), .A(n172), .Z(n5336) );
  XNOR U5733 ( .A(n5335), .B(n5336), .Z(n5338) );
  XNOR U5734 ( .A(n5337), .B(n5338), .Z(n5374) );
  XOR U5735 ( .A(n5373), .B(n5374), .Z(n5375) );
  NAND U5736 ( .A(x[128]), .B(y[699]), .Z(n5325) );
  ANDN U5737 ( .B(y[673]), .A(n176), .Z(n5334) );
  XOR U5738 ( .A(o[59]), .B(n5334), .Z(n5323) );
  NAND U5739 ( .A(y[672]), .B(x[155]), .Z(n5322) );
  XNOR U5740 ( .A(n5323), .B(n5322), .Z(n5324) );
  XNOR U5741 ( .A(n5325), .B(n5324), .Z(n5376) );
  XOR U5742 ( .A(n5375), .B(n5376), .Z(n5382) );
  XOR U5743 ( .A(n5426), .B(n5425), .Z(n5428) );
  XNOR U5744 ( .A(n5427), .B(n5428), .Z(n5316) );
  XNOR U5745 ( .A(n5317), .B(n5316), .Z(n5319) );
  OR U5746 ( .A(n5184), .B(n5183), .Z(n5188) );
  NANDN U5747 ( .A(n5186), .B(n5185), .Z(n5187) );
  NAND U5748 ( .A(n5188), .B(n5187), .Z(n5318) );
  XOR U5749 ( .A(n5319), .B(n5318), .Z(n5443) );
  OR U5750 ( .A(n5190), .B(n5189), .Z(n5194) );
  OR U5751 ( .A(n5192), .B(n5191), .Z(n5193) );
  AND U5752 ( .A(n5194), .B(n5193), .Z(n5444) );
  OR U5753 ( .A(n5196), .B(n5195), .Z(n5200) );
  NANDN U5754 ( .A(n5198), .B(n5197), .Z(n5199) );
  AND U5755 ( .A(n5200), .B(n5199), .Z(n5311) );
  NAND U5756 ( .A(n5202), .B(n5201), .Z(n5206) );
  NANDN U5757 ( .A(n5204), .B(n5203), .Z(n5205) );
  AND U5758 ( .A(n5206), .B(n5205), .Z(n5423) );
  ANDN U5759 ( .B(y[687]), .A(n163), .Z(n5397) );
  ANDN U5760 ( .B(y[686]), .A(n164), .Z(n5398) );
  XNOR U5761 ( .A(n5397), .B(n5398), .Z(n5400) );
  NAND U5762 ( .A(x[144]), .B(y[683]), .Z(n5409) );
  XOR U5763 ( .A(n5410), .B(n5409), .Z(n5411) );
  XOR U5764 ( .A(n5412), .B(n5411), .Z(n5399) );
  XNOR U5765 ( .A(n5400), .B(n5399), .Z(n5359) );
  ANDN U5766 ( .B(y[696]), .A(n154), .Z(n5405) );
  ANDN U5767 ( .B(y[697]), .A(n153), .Z(n5403) );
  ANDN U5768 ( .B(y[684]), .A(n166), .Z(n5404) );
  XNOR U5769 ( .A(n5403), .B(n5404), .Z(n5406) );
  XOR U5770 ( .A(n5405), .B(n5406), .Z(n5357) );
  NAND U5771 ( .A(y[693]), .B(x[134]), .Z(n5349) );
  ANDN U5772 ( .B(y[674]), .A(n14372), .Z(n5348) );
  NAND U5773 ( .A(y[680]), .B(x[147]), .Z(n5347) );
  XOR U5774 ( .A(n5348), .B(n5347), .Z(n5350) );
  XNOR U5775 ( .A(n5349), .B(n5350), .Z(n5358) );
  XNOR U5776 ( .A(n5357), .B(n5358), .Z(n5360) );
  XNOR U5777 ( .A(n5359), .B(n5360), .Z(n5387) );
  NAND U5778 ( .A(n5208), .B(n5207), .Z(n5212) );
  OR U5779 ( .A(n5210), .B(n5209), .Z(n5211) );
  AND U5780 ( .A(n5212), .B(n5211), .Z(n5385) );
  NANDN U5781 ( .A(n5214), .B(n5213), .Z(n5218) );
  NANDN U5782 ( .A(n5216), .B(n5215), .Z(n5217) );
  NAND U5783 ( .A(n5218), .B(n5217), .Z(n5386) );
  XNOR U5784 ( .A(n5385), .B(n5386), .Z(n5388) );
  XOR U5785 ( .A(n5387), .B(n5388), .Z(n5421) );
  NANDN U5786 ( .A(n5220), .B(n5219), .Z(n5224) );
  OR U5787 ( .A(n5222), .B(n5221), .Z(n5223) );
  AND U5788 ( .A(n5224), .B(n5223), .Z(n5422) );
  XOR U5789 ( .A(n5421), .B(n5422), .Z(n5424) );
  XOR U5790 ( .A(n5423), .B(n5424), .Z(n5310) );
  OR U5791 ( .A(n5226), .B(n5225), .Z(n5230) );
  NANDN U5792 ( .A(n5228), .B(n5227), .Z(n5229) );
  AND U5793 ( .A(n5230), .B(n5229), .Z(n5312) );
  XOR U5794 ( .A(n5313), .B(n5312), .Z(n5445) );
  XOR U5795 ( .A(n5446), .B(n5445), .Z(n5439) );
  OR U5796 ( .A(n5232), .B(n5231), .Z(n5236) );
  NANDN U5797 ( .A(n5234), .B(n5233), .Z(n5235) );
  AND U5798 ( .A(n5236), .B(n5235), .Z(n5437) );
  OR U5799 ( .A(n5238), .B(n5237), .Z(n5242) );
  OR U5800 ( .A(n5240), .B(n5239), .Z(n5241) );
  NAND U5801 ( .A(n5242), .B(n5241), .Z(n5354) );
  NANDN U5802 ( .A(n5244), .B(n5243), .Z(n5248) );
  NANDN U5803 ( .A(n5246), .B(n5245), .Z(n5247) );
  NAND U5804 ( .A(n5248), .B(n5247), .Z(n5353) );
  XOR U5805 ( .A(n5354), .B(n5353), .Z(n5355) );
  ANDN U5806 ( .B(y[685]), .A(n165), .Z(n5393) );
  AND U5807 ( .A(n5249), .B(o[58]), .Z(n5391) );
  ANDN U5808 ( .B(y[698]), .A(n152), .Z(n5392) );
  XNOR U5809 ( .A(n5391), .B(n5392), .Z(n5394) );
  XOR U5810 ( .A(n5393), .B(n5394), .Z(n5368) );
  NAND U5811 ( .A(x[145]), .B(y[682]), .Z(n5329) );
  ANDN U5812 ( .B(y[695]), .A(n155), .Z(n5328) );
  XNOR U5813 ( .A(n5329), .B(n5328), .Z(n5331) );
  ANDN U5814 ( .B(y[694]), .A(n156), .Z(n5330) );
  XOR U5815 ( .A(n5331), .B(n5330), .Z(n5367) );
  XOR U5816 ( .A(n5368), .B(n5367), .Z(n5370) );
  NAND U5817 ( .A(n5251), .B(n5250), .Z(n5255) );
  NANDN U5818 ( .A(n5253), .B(n5252), .Z(n5254) );
  NAND U5819 ( .A(n5255), .B(n5254), .Z(n5369) );
  XNOR U5820 ( .A(n5370), .B(n5369), .Z(n5356) );
  XOR U5821 ( .A(n5355), .B(n5356), .Z(n5304) );
  NANDN U5822 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U5823 ( .A(n5259), .B(n5258), .Z(n5260) );
  AND U5824 ( .A(n5261), .B(n5260), .Z(n5365) );
  ANDN U5825 ( .B(y[677]), .A(n173), .Z(n5417) );
  ANDN U5826 ( .B(y[676]), .A(n174), .Z(n5415) );
  ANDN U5827 ( .B(y[691]), .A(n159), .Z(n5416) );
  XNOR U5828 ( .A(n5415), .B(n5416), .Z(n5418) );
  XOR U5829 ( .A(n5417), .B(n5418), .Z(n5363) );
  AND U5830 ( .A(x[135]), .B(y[692]), .Z(n5343) );
  NANDN U5831 ( .A(n145), .B(x[152]), .Z(n5341) );
  XOR U5832 ( .A(n5342), .B(n5341), .Z(n5344) );
  XOR U5833 ( .A(n5343), .B(n5344), .Z(n5364) );
  XOR U5834 ( .A(n5363), .B(n5364), .Z(n5366) );
  XOR U5835 ( .A(n5365), .B(n5366), .Z(n5305) );
  XNOR U5836 ( .A(n5304), .B(n5305), .Z(n5307) );
  OR U5837 ( .A(n5263), .B(n5262), .Z(n5267) );
  OR U5838 ( .A(n5265), .B(n5264), .Z(n5266) );
  AND U5839 ( .A(n5267), .B(n5266), .Z(n5306) );
  XOR U5840 ( .A(n5307), .B(n5306), .Z(n5431) );
  OR U5841 ( .A(n5269), .B(n5268), .Z(n5273) );
  OR U5842 ( .A(n5271), .B(n5270), .Z(n5272) );
  AND U5843 ( .A(n5273), .B(n5272), .Z(n5432) );
  XNOR U5844 ( .A(n5431), .B(n5432), .Z(n5434) );
  OR U5845 ( .A(n5275), .B(n5274), .Z(n5279) );
  NANDN U5846 ( .A(n5277), .B(n5276), .Z(n5278) );
  NAND U5847 ( .A(n5279), .B(n5278), .Z(n5433) );
  XOR U5848 ( .A(n5434), .B(n5433), .Z(n5438) );
  XNOR U5849 ( .A(n5437), .B(n5438), .Z(n5440) );
  XNOR U5850 ( .A(n5439), .B(n5440), .Z(n5301) );
  NANDN U5851 ( .A(n5281), .B(n5280), .Z(n5285) );
  NANDN U5852 ( .A(n5283), .B(n5282), .Z(n5284) );
  NAND U5853 ( .A(n5285), .B(n5284), .Z(n5299) );
  OR U5854 ( .A(n5287), .B(n5286), .Z(n5291) );
  NANDN U5855 ( .A(n5289), .B(n5288), .Z(n5290) );
  AND U5856 ( .A(n5291), .B(n5290), .Z(n5298) );
  XNOR U5857 ( .A(n5301), .B(n5300), .Z(n5295) );
  XOR U5858 ( .A(n5294), .B(n5295), .Z(N124) );
  NANDN U5859 ( .A(n5293), .B(n5292), .Z(n5297) );
  NANDN U5860 ( .A(n5295), .B(n5294), .Z(n5296) );
  NAND U5861 ( .A(n5297), .B(n5296), .Z(n5605) );
  NANDN U5862 ( .A(n5299), .B(n5298), .Z(n5303) );
  NANDN U5863 ( .A(n5301), .B(n5300), .Z(n5302) );
  NAND U5864 ( .A(n5303), .B(n5302), .Z(n5606) );
  XNOR U5865 ( .A(n5605), .B(n5606), .Z(n5607) );
  NAND U5866 ( .A(n5305), .B(n5304), .Z(n5309) );
  OR U5867 ( .A(n5307), .B(n5306), .Z(n5308) );
  AND U5868 ( .A(n5309), .B(n5308), .Z(n5458) );
  NANDN U5869 ( .A(n5311), .B(n5310), .Z(n5315) );
  OR U5870 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U5871 ( .A(n5315), .B(n5314), .Z(n5456) );
  OR U5872 ( .A(n5317), .B(n5316), .Z(n5321) );
  OR U5873 ( .A(n5319), .B(n5318), .Z(n5320) );
  NAND U5874 ( .A(n5321), .B(n5320), .Z(n5455) );
  XOR U5875 ( .A(n5456), .B(n5455), .Z(n5457) );
  XNOR U5876 ( .A(n5458), .B(n5457), .Z(n5452) );
  NANDN U5877 ( .A(n5323), .B(n5322), .Z(n5327) );
  NAND U5878 ( .A(n5325), .B(n5324), .Z(n5326) );
  AND U5879 ( .A(n5327), .B(n5326), .Z(n5479) );
  NANDN U5880 ( .A(n5329), .B(n5328), .Z(n5333) );
  NAND U5881 ( .A(n5331), .B(n5330), .Z(n5332) );
  NAND U5882 ( .A(n5333), .B(n5332), .Z(n5480) );
  XOR U5883 ( .A(n5479), .B(n5480), .Z(n5482) );
  AND U5884 ( .A(n5334), .B(o[59]), .Z(n5577) );
  IV U5885 ( .A(x[156]), .Z(n14373) );
  ANDN U5886 ( .B(y[672]), .A(n14373), .Z(n5578) );
  XNOR U5887 ( .A(n5577), .B(n5578), .Z(n5580) );
  ANDN U5888 ( .B(y[700]), .A(n151), .Z(n5579) );
  XNOR U5889 ( .A(n5580), .B(n5579), .Z(n5561) );
  OR U5890 ( .A(n5336), .B(n5335), .Z(n5340) );
  OR U5891 ( .A(n5338), .B(n5337), .Z(n5339) );
  AND U5892 ( .A(n5340), .B(n5339), .Z(n5558) );
  ANDN U5893 ( .B(y[691]), .A(n160), .Z(n5571) );
  ANDN U5894 ( .B(y[692]), .A(n159), .Z(n5572) );
  XNOR U5895 ( .A(n5571), .B(n5572), .Z(n5574) );
  ANDN U5896 ( .B(y[690]), .A(n161), .Z(n5573) );
  XNOR U5897 ( .A(n5574), .B(n5573), .Z(n5559) );
  XOR U5898 ( .A(n5558), .B(n5559), .Z(n5560) );
  XNOR U5899 ( .A(n5482), .B(n5481), .Z(n5464) );
  ANDN U5900 ( .B(y[699]), .A(n152), .Z(n5534) );
  ANDN U5901 ( .B(y[675]), .A(n14372), .Z(n5535) );
  XNOR U5902 ( .A(n5534), .B(n5535), .Z(n5537) );
  XNOR U5903 ( .A(n5536), .B(n5537), .Z(n5475) );
  ANDN U5904 ( .B(y[684]), .A(n167), .Z(n5542) );
  ANDN U5905 ( .B(y[698]), .A(n153), .Z(n5540) );
  ANDN U5906 ( .B(y[676]), .A(n175), .Z(n5541) );
  XNOR U5907 ( .A(n5540), .B(n5541), .Z(n5543) );
  XOR U5908 ( .A(n5542), .B(n5543), .Z(n5473) );
  NANDN U5909 ( .A(n5342), .B(n5341), .Z(n5346) );
  OR U5910 ( .A(n5344), .B(n5343), .Z(n5345) );
  NAND U5911 ( .A(n5346), .B(n5345), .Z(n5474) );
  XNOR U5912 ( .A(n5473), .B(n5474), .Z(n5476) );
  XNOR U5913 ( .A(n5475), .B(n5476), .Z(n5462) );
  ANDN U5914 ( .B(y[677]), .A(n174), .Z(n5503) );
  ANDN U5915 ( .B(y[697]), .A(n154), .Z(n5504) );
  XNOR U5916 ( .A(n5503), .B(n5504), .Z(n5506) );
  XOR U5917 ( .A(n5505), .B(n5506), .Z(n5487) );
  ANDN U5918 ( .B(y[695]), .A(n156), .Z(n5524) );
  ANDN U5919 ( .B(y[680]), .A(n171), .Z(n5522) );
  ANDN U5920 ( .B(y[679]), .A(n172), .Z(n5523) );
  XNOR U5921 ( .A(n5522), .B(n5523), .Z(n5525) );
  XOR U5922 ( .A(n5524), .B(n5525), .Z(n5485) );
  NANDN U5923 ( .A(n5348), .B(n5347), .Z(n5352) );
  NANDN U5924 ( .A(n5350), .B(n5349), .Z(n5351) );
  NAND U5925 ( .A(n5352), .B(n5351), .Z(n5486) );
  XNOR U5926 ( .A(n5485), .B(n5486), .Z(n5488) );
  XNOR U5927 ( .A(n5487), .B(n5488), .Z(n5461) );
  XOR U5928 ( .A(n5462), .B(n5461), .Z(n5463) );
  XNOR U5929 ( .A(n5464), .B(n5463), .Z(n5596) );
  OR U5930 ( .A(n5358), .B(n5357), .Z(n5362) );
  OR U5931 ( .A(n5360), .B(n5359), .Z(n5361) );
  NAND U5932 ( .A(n5362), .B(n5361), .Z(n5498) );
  XOR U5933 ( .A(n5498), .B(n5497), .Z(n5499) );
  XOR U5934 ( .A(n5596), .B(n5595), .Z(n5598) );
  NANDN U5935 ( .A(n5368), .B(n5367), .Z(n5372) );
  OR U5936 ( .A(n5370), .B(n5369), .Z(n5371) );
  AND U5937 ( .A(n5372), .B(n5371), .Z(n5491) );
  OR U5938 ( .A(n5374), .B(n5373), .Z(n5378) );
  NANDN U5939 ( .A(n5376), .B(n5375), .Z(n5377) );
  NAND U5940 ( .A(n5378), .B(n5377), .Z(n5492) );
  XOR U5941 ( .A(n5491), .B(n5492), .Z(n5493) );
  OR U5942 ( .A(n5380), .B(n5379), .Z(n5384) );
  NANDN U5943 ( .A(n5382), .B(n5381), .Z(n5383) );
  NAND U5944 ( .A(n5384), .B(n5383), .Z(n5494) );
  OR U5945 ( .A(n5386), .B(n5385), .Z(n5390) );
  NANDN U5946 ( .A(n5388), .B(n5387), .Z(n5389) );
  AND U5947 ( .A(n5390), .B(n5389), .Z(n5590) );
  OR U5948 ( .A(n5392), .B(n5391), .Z(n5396) );
  OR U5949 ( .A(n5394), .B(n5393), .Z(n5395) );
  AND U5950 ( .A(n5396), .B(n5395), .Z(n5586) );
  OR U5951 ( .A(n5398), .B(n5397), .Z(n5402) );
  NANDN U5952 ( .A(n5400), .B(n5399), .Z(n5401) );
  AND U5953 ( .A(n5402), .B(n5401), .Z(n5583) );
  OR U5954 ( .A(n5404), .B(n5403), .Z(n5408) );
  OR U5955 ( .A(n5406), .B(n5405), .Z(n5407) );
  AND U5956 ( .A(n5408), .B(n5407), .Z(n5584) );
  XOR U5957 ( .A(n5583), .B(n5584), .Z(n5585) );
  ANDN U5958 ( .B(y[693]), .A(n158), .Z(n5548) );
  ANDN U5959 ( .B(y[689]), .A(n162), .Z(n5546) );
  ANDN U5960 ( .B(y[688]), .A(n163), .Z(n5547) );
  XNOR U5961 ( .A(n5546), .B(n5547), .Z(n5549) );
  XOR U5962 ( .A(n5548), .B(n5549), .Z(n5516) );
  NANDN U5963 ( .A(n5410), .B(n5409), .Z(n5414) );
  OR U5964 ( .A(n5412), .B(n5411), .Z(n5413) );
  NAND U5965 ( .A(n5414), .B(n5413), .Z(n5517) );
  XNOR U5966 ( .A(n5516), .B(n5517), .Z(n5519) );
  NAND U5967 ( .A(x[143]), .B(y[685]), .Z(n5510) );
  AND U5968 ( .A(y[674]), .B(x[154]), .Z(n5509) );
  XNOR U5969 ( .A(n5510), .B(n5509), .Z(n5511) );
  AND U5970 ( .A(y[673]), .B(x[155]), .Z(n5659) );
  XNOR U5971 ( .A(o[60]), .B(n5659), .Z(n5512) );
  XOR U5972 ( .A(n5519), .B(n5518), .Z(n5467) );
  OR U5973 ( .A(n5416), .B(n5415), .Z(n5420) );
  OR U5974 ( .A(n5418), .B(n5417), .Z(n5419) );
  AND U5975 ( .A(n5420), .B(n5419), .Z(n5552) );
  ANDN U5976 ( .B(y[694]), .A(n157), .Z(n5532) );
  ANDN U5977 ( .B(y[681]), .A(n170), .Z(n5531) );
  XNOR U5978 ( .A(n5530), .B(n5531), .Z(n5533) );
  XNOR U5979 ( .A(n5532), .B(n5533), .Z(n5553) );
  XOR U5980 ( .A(n5552), .B(n5553), .Z(n5555) );
  NAND U5981 ( .A(x[145]), .B(y[683]), .Z(n5566) );
  ANDN U5982 ( .B(y[696]), .A(n155), .Z(n5565) );
  NAND U5983 ( .A(y[678]), .B(x[150]), .Z(n5564) );
  XOR U5984 ( .A(n5565), .B(n5564), .Z(n5567) );
  XNOR U5985 ( .A(n5566), .B(n5567), .Z(n5554) );
  XNOR U5986 ( .A(n5555), .B(n5554), .Z(n5468) );
  XNOR U5987 ( .A(n5467), .B(n5468), .Z(n5469) );
  XOR U5988 ( .A(n5470), .B(n5469), .Z(n5589) );
  XOR U5989 ( .A(n5590), .B(n5589), .Z(n5592) );
  XOR U5990 ( .A(n5591), .B(n5592), .Z(n5597) );
  XOR U5991 ( .A(n5598), .B(n5597), .Z(n5604) );
  NANDN U5992 ( .A(n5426), .B(n5425), .Z(n5430) );
  NANDN U5993 ( .A(n5428), .B(n5427), .Z(n5429) );
  NAND U5994 ( .A(n5430), .B(n5429), .Z(n5602) );
  XOR U5995 ( .A(n5601), .B(n5602), .Z(n5603) );
  XOR U5996 ( .A(n5604), .B(n5603), .Z(n5450) );
  OR U5997 ( .A(n5432), .B(n5431), .Z(n5436) );
  OR U5998 ( .A(n5434), .B(n5433), .Z(n5435) );
  AND U5999 ( .A(n5436), .B(n5435), .Z(n5449) );
  XOR U6000 ( .A(n5450), .B(n5449), .Z(n5451) );
  OR U6001 ( .A(n5438), .B(n5437), .Z(n5442) );
  NANDN U6002 ( .A(n5440), .B(n5439), .Z(n5441) );
  AND U6003 ( .A(n5442), .B(n5441), .Z(n5612) );
  XNOR U6004 ( .A(n5611), .B(n5612), .Z(n5614) );
  NANDN U6005 ( .A(n5444), .B(n5443), .Z(n5448) );
  NANDN U6006 ( .A(n5446), .B(n5445), .Z(n5447) );
  NAND U6007 ( .A(n5448), .B(n5447), .Z(n5613) );
  XOR U6008 ( .A(n5614), .B(n5613), .Z(n5608) );
  XNOR U6009 ( .A(n5607), .B(n5608), .Z(N125) );
  OR U6010 ( .A(n5450), .B(n5449), .Z(n5454) );
  NANDN U6011 ( .A(n5452), .B(n5451), .Z(n5453) );
  NAND U6012 ( .A(n5454), .B(n5453), .Z(n5626) );
  OR U6013 ( .A(n5456), .B(n5455), .Z(n5460) );
  NANDN U6014 ( .A(n5458), .B(n5457), .Z(n5459) );
  AND U6015 ( .A(n5460), .B(n5459), .Z(n5623) );
  NANDN U6016 ( .A(n5462), .B(n5461), .Z(n5466) );
  OR U6017 ( .A(n5464), .B(n5463), .Z(n5465) );
  AND U6018 ( .A(n5466), .B(n5465), .Z(n5787) );
  OR U6019 ( .A(n5468), .B(n5467), .Z(n5472) );
  OR U6020 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U6021 ( .A(n5472), .B(n5471), .Z(n5780) );
  OR U6022 ( .A(n5474), .B(n5473), .Z(n5478) );
  NANDN U6023 ( .A(n5476), .B(n5475), .Z(n5477) );
  NAND U6024 ( .A(n5478), .B(n5477), .Z(n5715) );
  OR U6025 ( .A(n5480), .B(n5479), .Z(n5484) );
  NAND U6026 ( .A(n5482), .B(n5481), .Z(n5483) );
  AND U6027 ( .A(n5484), .B(n5483), .Z(n5712) );
  OR U6028 ( .A(n5486), .B(n5485), .Z(n5490) );
  OR U6029 ( .A(n5488), .B(n5487), .Z(n5489) );
  NAND U6030 ( .A(n5490), .B(n5489), .Z(n5713) );
  XNOR U6031 ( .A(n5712), .B(n5713), .Z(n5714) );
  XOR U6032 ( .A(n5715), .B(n5714), .Z(n5779) );
  XNOR U6033 ( .A(n5780), .B(n5779), .Z(n5782) );
  OR U6034 ( .A(n5492), .B(n5491), .Z(n5496) );
  NANDN U6035 ( .A(n5494), .B(n5493), .Z(n5495) );
  AND U6036 ( .A(n5496), .B(n5495), .Z(n5781) );
  XOR U6037 ( .A(n5782), .B(n5781), .Z(n5785) );
  OR U6038 ( .A(n5498), .B(n5497), .Z(n5502) );
  NANDN U6039 ( .A(n5500), .B(n5499), .Z(n5501) );
  AND U6040 ( .A(n5502), .B(n5501), .Z(n5786) );
  XNOR U6041 ( .A(n5785), .B(n5786), .Z(n5788) );
  XOR U6042 ( .A(n5787), .B(n5788), .Z(n5775) );
  OR U6043 ( .A(n5504), .B(n5503), .Z(n5508) );
  OR U6044 ( .A(n5506), .B(n5505), .Z(n5507) );
  AND U6045 ( .A(n5508), .B(n5507), .Z(n5633) );
  NANDN U6046 ( .A(n5510), .B(n5509), .Z(n5514) );
  NANDN U6047 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U6048 ( .A(n5514), .B(n5513), .Z(n5634) );
  XOR U6049 ( .A(n5633), .B(n5634), .Z(n5635) );
  ANDN U6050 ( .B(y[693]), .A(n159), .Z(n5675) );
  ANDN U6051 ( .B(y[694]), .A(n158), .Z(n5676) );
  XNOR U6052 ( .A(n5675), .B(n5676), .Z(n5678) );
  ANDN U6053 ( .B(y[695]), .A(n157), .Z(n5677) );
  XNOR U6054 ( .A(n5678), .B(n5677), .Z(n5750) );
  NOR U6055 ( .A(n160), .B(n5515), .Z(n5921) );
  ANDN U6056 ( .B(y[696]), .A(n156), .Z(n5645) );
  ANDN U6057 ( .B(y[691]), .A(n161), .Z(n5646) );
  XNOR U6058 ( .A(n5645), .B(n5646), .Z(n5648) );
  ANDN U6059 ( .B(y[697]), .A(n155), .Z(n5647) );
  XNOR U6060 ( .A(n5648), .B(n5647), .Z(n5748) );
  XNOR U6061 ( .A(n5921), .B(n5748), .Z(n5749) );
  XNOR U6062 ( .A(n5750), .B(n5749), .Z(n5636) );
  OR U6063 ( .A(n5517), .B(n5516), .Z(n5521) );
  OR U6064 ( .A(n5519), .B(n5518), .Z(n5520) );
  AND U6065 ( .A(n5521), .B(n5520), .Z(n5706) );
  OR U6066 ( .A(n5523), .B(n5522), .Z(n5527) );
  OR U6067 ( .A(n5525), .B(n5524), .Z(n5526) );
  AND U6068 ( .A(n5527), .B(n5526), .Z(n5683) );
  ANDN U6069 ( .B(y[685]), .A(n167), .Z(n5657) );
  NAND U6070 ( .A(y[673]), .B(o[60]), .Z(n5528) );
  XNOR U6071 ( .A(y[674]), .B(n5528), .Z(n5529) );
  NAND U6072 ( .A(x[155]), .B(n5529), .Z(n5658) );
  XNOR U6073 ( .A(n5657), .B(n5658), .Z(n5684) );
  XOR U6074 ( .A(n5683), .B(n5684), .Z(n5686) );
  NAND U6075 ( .A(x[130]), .B(y[699]), .Z(n5653) );
  ANDN U6076 ( .B(y[683]), .A(n169), .Z(n5652) );
  NAND U6077 ( .A(y[682]), .B(x[147]), .Z(n5651) );
  XOR U6078 ( .A(n5652), .B(n5651), .Z(n5654) );
  XNOR U6079 ( .A(n5653), .B(n5654), .Z(n5685) );
  XNOR U6080 ( .A(n5686), .B(n5685), .Z(n5719) );
  ANDN U6081 ( .B(y[673]), .A(n14373), .Z(n5705) );
  XOR U6082 ( .A(o[61]), .B(n5705), .Z(n5755) );
  IV U6083 ( .A(x[157]), .Z(n11441) );
  ANDN U6084 ( .B(y[672]), .A(n11441), .Z(n5756) );
  XNOR U6085 ( .A(n5755), .B(n5756), .Z(n5758) );
  ANDN U6086 ( .B(y[701]), .A(n151), .Z(n5757) );
  XOR U6087 ( .A(n5758), .B(n5757), .Z(n5743) );
  ANDN U6088 ( .B(y[687]), .A(n165), .Z(n5691) );
  ANDN U6089 ( .B(y[676]), .A(n14372), .Z(n5689) );
  ANDN U6090 ( .B(y[675]), .A(n176), .Z(n5690) );
  XNOR U6091 ( .A(n5689), .B(n5690), .Z(n5692) );
  XNOR U6092 ( .A(n5691), .B(n5692), .Z(n5742) );
  XOR U6093 ( .A(n5743), .B(n5742), .Z(n5744) );
  XOR U6094 ( .A(n5745), .B(n5744), .Z(n5718) );
  XNOR U6095 ( .A(n5719), .B(n5718), .Z(n5721) );
  OR U6096 ( .A(n5535), .B(n5534), .Z(n5539) );
  OR U6097 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U6098 ( .A(n5539), .B(n5538), .Z(n5733) );
  OR U6099 ( .A(n5541), .B(n5540), .Z(n5545) );
  OR U6100 ( .A(n5543), .B(n5542), .Z(n5544) );
  AND U6101 ( .A(n5545), .B(n5544), .Z(n5730) );
  OR U6102 ( .A(n5547), .B(n5546), .Z(n5551) );
  OR U6103 ( .A(n5549), .B(n5548), .Z(n5550) );
  AND U6104 ( .A(n5551), .B(n5550), .Z(n5639) );
  ANDN U6105 ( .B(y[690]), .A(n162), .Z(n5664) );
  ANDN U6106 ( .B(y[684]), .A(n168), .Z(n5665) );
  XNOR U6107 ( .A(n5664), .B(n5665), .Z(n5667) );
  ANDN U6108 ( .B(y[698]), .A(n154), .Z(n5666) );
  XNOR U6109 ( .A(n5667), .B(n5666), .Z(n5640) );
  XOR U6110 ( .A(n5639), .B(n5640), .Z(n5642) );
  ANDN U6111 ( .B(y[678]), .A(n174), .Z(n5670) );
  ANDN U6112 ( .B(y[677]), .A(n175), .Z(n5890) );
  XNOR U6113 ( .A(n5670), .B(n5890), .Z(n5672) );
  ANDN U6114 ( .B(y[688]), .A(n164), .Z(n5671) );
  XOR U6115 ( .A(n5672), .B(n5671), .Z(n5641) );
  XNOR U6116 ( .A(n5642), .B(n5641), .Z(n5731) );
  XOR U6117 ( .A(n5730), .B(n5731), .Z(n5732) );
  XOR U6118 ( .A(n5721), .B(n5720), .Z(n5707) );
  XOR U6119 ( .A(n5706), .B(n5707), .Z(n5708) );
  OR U6120 ( .A(n5553), .B(n5552), .Z(n5557) );
  NAND U6121 ( .A(n5555), .B(n5554), .Z(n5556) );
  AND U6122 ( .A(n5557), .B(n5556), .Z(n5724) );
  OR U6123 ( .A(n5559), .B(n5558), .Z(n5563) );
  NANDN U6124 ( .A(n5561), .B(n5560), .Z(n5562) );
  AND U6125 ( .A(n5563), .B(n5562), .Z(n5767) );
  NANDN U6126 ( .A(n5565), .B(n5564), .Z(n5569) );
  NANDN U6127 ( .A(n5567), .B(n5566), .Z(n5568) );
  AND U6128 ( .A(n5569), .B(n5568), .Z(n5761) );
  NOR U6129 ( .A(n163), .B(n5570), .Z(n5871) );
  ANDN U6130 ( .B(y[679]), .A(n173), .Z(n5695) );
  ANDN U6131 ( .B(y[700]), .A(n152), .Z(n5696) );
  XNOR U6132 ( .A(n5695), .B(n5696), .Z(n5697) );
  XNOR U6133 ( .A(n5871), .B(n5697), .Z(n5739) );
  OR U6134 ( .A(n5572), .B(n5571), .Z(n5576) );
  OR U6135 ( .A(n5574), .B(n5573), .Z(n5575) );
  AND U6136 ( .A(n5576), .B(n5575), .Z(n5736) );
  NAND U6137 ( .A(x[143]), .B(y[686]), .Z(n5699) );
  AND U6138 ( .A(x[149]), .B(y[680]), .Z(n5999) );
  NAND U6139 ( .A(y[681]), .B(x[148]), .Z(n5698) );
  XNOR U6140 ( .A(n5999), .B(n5698), .Z(n5700) );
  XNOR U6141 ( .A(n5736), .B(n5737), .Z(n5738) );
  XNOR U6142 ( .A(n5739), .B(n5738), .Z(n5762) );
  XOR U6143 ( .A(n5761), .B(n5762), .Z(n5763) );
  OR U6144 ( .A(n5578), .B(n5577), .Z(n5582) );
  OR U6145 ( .A(n5580), .B(n5579), .Z(n5581) );
  AND U6146 ( .A(n5582), .B(n5581), .Z(n5764) );
  XNOR U6147 ( .A(n5767), .B(n5768), .Z(n5770) );
  OR U6148 ( .A(n5584), .B(n5583), .Z(n5588) );
  NANDN U6149 ( .A(n5586), .B(n5585), .Z(n5587) );
  AND U6150 ( .A(n5588), .B(n5587), .Z(n5769) );
  XNOR U6151 ( .A(n5770), .B(n5769), .Z(n5725) );
  XNOR U6152 ( .A(n5724), .B(n5725), .Z(n5727) );
  XOR U6153 ( .A(n5726), .B(n5727), .Z(n5773) );
  NANDN U6154 ( .A(n5590), .B(n5589), .Z(n5594) );
  NANDN U6155 ( .A(n5592), .B(n5591), .Z(n5593) );
  NAND U6156 ( .A(n5594), .B(n5593), .Z(n5774) );
  XOR U6157 ( .A(n5773), .B(n5774), .Z(n5776) );
  XNOR U6158 ( .A(n5775), .B(n5776), .Z(n5631) );
  NANDN U6159 ( .A(n5596), .B(n5595), .Z(n5600) );
  OR U6160 ( .A(n5598), .B(n5597), .Z(n5599) );
  NAND U6161 ( .A(n5600), .B(n5599), .Z(n5630) );
  XOR U6162 ( .A(n5630), .B(n5629), .Z(n5632) );
  XOR U6163 ( .A(n5631), .B(n5632), .Z(n5624) );
  XNOR U6164 ( .A(n5623), .B(n5624), .Z(n5625) );
  XNOR U6165 ( .A(n5626), .B(n5625), .Z(n5620) );
  NANDN U6166 ( .A(n5606), .B(n5605), .Z(n5610) );
  NAND U6167 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U6168 ( .A(n5610), .B(n5609), .Z(n5617) );
  OR U6169 ( .A(n5612), .B(n5611), .Z(n5616) );
  OR U6170 ( .A(n5614), .B(n5613), .Z(n5615) );
  AND U6171 ( .A(n5616), .B(n5615), .Z(n5618) );
  XNOR U6172 ( .A(n5617), .B(n5618), .Z(n5619) );
  XOR U6173 ( .A(n5620), .B(n5619), .Z(N126) );
  NANDN U6174 ( .A(n5618), .B(n5617), .Z(n5622) );
  NANDN U6175 ( .A(n5620), .B(n5619), .Z(n5621) );
  AND U6176 ( .A(n5622), .B(n5621), .Z(n5793) );
  OR U6177 ( .A(n5624), .B(n5623), .Z(n5628) );
  OR U6178 ( .A(n5626), .B(n5625), .Z(n5627) );
  AND U6179 ( .A(n5628), .B(n5627), .Z(n5794) );
  XNOR U6180 ( .A(n5793), .B(n5794), .Z(n5792) );
  OR U6181 ( .A(n5634), .B(n5633), .Z(n5638) );
  NANDN U6182 ( .A(n5636), .B(n5635), .Z(n5637) );
  AND U6183 ( .A(n5638), .B(n5637), .Z(n5809) );
  OR U6184 ( .A(n5640), .B(n5639), .Z(n5644) );
  NAND U6185 ( .A(n5642), .B(n5641), .Z(n5643) );
  AND U6186 ( .A(n5644), .B(n5643), .Z(n5811) );
  OR U6187 ( .A(n5646), .B(n5645), .Z(n5650) );
  OR U6188 ( .A(n5648), .B(n5647), .Z(n5649) );
  AND U6189 ( .A(n5650), .B(n5649), .Z(n5836) );
  NAND U6190 ( .A(x[134]), .B(y[696]), .Z(n5894) );
  NAND U6191 ( .A(x[133]), .B(y[697]), .Z(n5896) );
  NAND U6192 ( .A(x[147]), .B(y[683]), .Z(n5895) );
  XNOR U6193 ( .A(n5896), .B(n5895), .Z(n5893) );
  XNOR U6194 ( .A(n5894), .B(n5893), .Z(n5952) );
  NANDN U6195 ( .A(n5652), .B(n5651), .Z(n5656) );
  NANDN U6196 ( .A(n5654), .B(n5653), .Z(n5655) );
  AND U6197 ( .A(n5656), .B(n5655), .Z(n5954) );
  NAND U6198 ( .A(x[132]), .B(y[698]), .Z(n6004) );
  NAND U6199 ( .A(x[131]), .B(y[699]), .Z(n6006) );
  AND U6200 ( .A(y[684]), .B(x[146]), .Z(n6005) );
  XNOR U6201 ( .A(n6006), .B(n6005), .Z(n6003) );
  XNOR U6202 ( .A(n6004), .B(n6003), .Z(n5955) );
  XOR U6203 ( .A(n5954), .B(n5955), .Z(n5953) );
  XNOR U6204 ( .A(n5952), .B(n5953), .Z(n5835) );
  XOR U6205 ( .A(n5836), .B(n5835), .Z(n5838) );
  OR U6206 ( .A(n5658), .B(n5657), .Z(n5663) );
  NAND U6207 ( .A(o[60]), .B(n5659), .Z(n5661) );
  NAND U6208 ( .A(x[155]), .B(y[674]), .Z(n5660) );
  AND U6209 ( .A(n5661), .B(n5660), .Z(n5662) );
  ANDN U6210 ( .B(n5663), .A(n5662), .Z(n5837) );
  XNOR U6211 ( .A(n5811), .B(n5812), .Z(n5810) );
  XNOR U6212 ( .A(n5809), .B(n5810), .Z(n5800) );
  OR U6213 ( .A(n5665), .B(n5664), .Z(n5669) );
  OR U6214 ( .A(n5667), .B(n5666), .Z(n5668) );
  NAND U6215 ( .A(n5669), .B(n5668), .Z(n5864) );
  NAND U6216 ( .A(x[148]), .B(y[682]), .Z(n5943) );
  AND U6217 ( .A(y[688]), .B(x[142]), .Z(n5942) );
  XOR U6218 ( .A(n5943), .B(n5942), .Z(n5941) );
  AND U6219 ( .A(y[694]), .B(x[136]), .Z(n5940) );
  XOR U6220 ( .A(n5941), .B(n5940), .Z(n5866) );
  NAND U6221 ( .A(y[672]), .B(x[158]), .Z(n5927) );
  NAND U6222 ( .A(x[157]), .B(y[673]), .Z(n5958) );
  XNOR U6223 ( .A(o[62]), .B(n5958), .Z(n5926) );
  XOR U6224 ( .A(n5927), .B(n5926), .Z(n5929) );
  AND U6225 ( .A(y[702]), .B(x[128]), .Z(n5928) );
  XNOR U6226 ( .A(n5929), .B(n5928), .Z(n5865) );
  XOR U6227 ( .A(n5864), .B(n5863), .Z(n5819) );
  OR U6228 ( .A(n5890), .B(n5670), .Z(n5674) );
  OR U6229 ( .A(n5672), .B(n5671), .Z(n5673) );
  AND U6230 ( .A(n5674), .B(n5673), .Z(n5820) );
  XNOR U6231 ( .A(n5819), .B(n5820), .Z(n5818) );
  OR U6232 ( .A(n5676), .B(n5675), .Z(n5680) );
  OR U6233 ( .A(n5678), .B(n5677), .Z(n5679) );
  AND U6234 ( .A(n5680), .B(n5679), .Z(n5856) );
  NAND U6235 ( .A(x[145]), .B(y[685]), .Z(n5935) );
  NAND U6236 ( .A(x[130]), .B(y[700]), .Z(n5937) );
  NAND U6237 ( .A(x[154]), .B(y[676]), .Z(n5936) );
  XNOR U6238 ( .A(n5937), .B(n5936), .Z(n5934) );
  XNOR U6239 ( .A(n5935), .B(n5934), .Z(n5857) );
  NAND U6240 ( .A(x[135]), .B(y[695]), .Z(n5998) );
  AND U6241 ( .A(x[150]), .B(y[680]), .Z(n5682) );
  AND U6242 ( .A(x[149]), .B(y[681]), .Z(n5681) );
  XNOR U6243 ( .A(n5682), .B(n5681), .Z(n5997) );
  XOR U6244 ( .A(n5998), .B(n5997), .Z(n5858) );
  XNOR U6245 ( .A(n5857), .B(n5858), .Z(n5855) );
  XOR U6246 ( .A(n5856), .B(n5855), .Z(n5817) );
  XNOR U6247 ( .A(n5818), .B(n5817), .Z(n5803) );
  OR U6248 ( .A(n5684), .B(n5683), .Z(n5688) );
  NAND U6249 ( .A(n5686), .B(n5685), .Z(n5687) );
  NAND U6250 ( .A(n5688), .B(n5687), .Z(n5806) );
  OR U6251 ( .A(n5690), .B(n5689), .Z(n5694) );
  OR U6252 ( .A(n5692), .B(n5691), .Z(n5693) );
  AND U6253 ( .A(n5694), .B(n5693), .Z(n5829) );
  NANDN U6254 ( .A(n5999), .B(n5698), .Z(n5702) );
  NAND U6255 ( .A(n5700), .B(n5699), .Z(n5701) );
  AND U6256 ( .A(n5702), .B(n5701), .Z(n5849) );
  NAND U6257 ( .A(x[151]), .B(y[679]), .Z(n5889) );
  AND U6258 ( .A(y[677]), .B(x[153]), .Z(n5704) );
  AND U6259 ( .A(x[152]), .B(y[678]), .Z(n5703) );
  XNOR U6260 ( .A(n5704), .B(n5703), .Z(n5888) );
  XOR U6261 ( .A(n5889), .B(n5888), .Z(n5851) );
  NAND U6262 ( .A(n5705), .B(o[61]), .Z(n5875) );
  NAND U6263 ( .A(x[156]), .B(y[674]), .Z(n5877) );
  AND U6264 ( .A(y[686]), .B(x[144]), .Z(n5876) );
  XNOR U6265 ( .A(n5877), .B(n5876), .Z(n5874) );
  XNOR U6266 ( .A(n5875), .B(n5874), .Z(n5852) );
  XNOR U6267 ( .A(n5851), .B(n5852), .Z(n5850) );
  XOR U6268 ( .A(n5849), .B(n5850), .Z(n5831) );
  XOR U6269 ( .A(n5829), .B(n5830), .Z(n5805) );
  XNOR U6270 ( .A(n5806), .B(n5805), .Z(n5804) );
  XNOR U6271 ( .A(n5803), .B(n5804), .Z(n5799) );
  XNOR U6272 ( .A(n5800), .B(n5799), .Z(n5798) );
  OR U6273 ( .A(n5707), .B(n5706), .Z(n5711) );
  NANDN U6274 ( .A(n5709), .B(n5708), .Z(n5710) );
  NAND U6275 ( .A(n5711), .B(n5710), .Z(n5797) );
  XOR U6276 ( .A(n5798), .B(n5797), .Z(n6066) );
  OR U6277 ( .A(n5713), .B(n5712), .Z(n5717) );
  OR U6278 ( .A(n5715), .B(n5714), .Z(n5716) );
  NAND U6279 ( .A(n5717), .B(n5716), .Z(n6068) );
  OR U6280 ( .A(n5719), .B(n5718), .Z(n5723) );
  OR U6281 ( .A(n5721), .B(n5720), .Z(n5722) );
  NAND U6282 ( .A(n5723), .B(n5722), .Z(n6067) );
  XOR U6283 ( .A(n6068), .B(n6067), .Z(n6065) );
  XOR U6284 ( .A(n6066), .B(n6065), .Z(n6060) );
  OR U6285 ( .A(n5725), .B(n5724), .Z(n5729) );
  NANDN U6286 ( .A(n5727), .B(n5726), .Z(n5728) );
  NAND U6287 ( .A(n5729), .B(n5728), .Z(n6062) );
  OR U6288 ( .A(n5731), .B(n5730), .Z(n5735) );
  NANDN U6289 ( .A(n5733), .B(n5732), .Z(n5734) );
  AND U6290 ( .A(n5735), .B(n5734), .Z(n6045) );
  OR U6291 ( .A(n5737), .B(n5736), .Z(n5741) );
  OR U6292 ( .A(n5739), .B(n5738), .Z(n5740) );
  AND U6293 ( .A(n5741), .B(n5740), .Z(n6046) );
  XOR U6294 ( .A(n6045), .B(n6046), .Z(n6043) );
  NANDN U6295 ( .A(n5743), .B(n5742), .Z(n5747) );
  OR U6296 ( .A(n5745), .B(n5744), .Z(n5746) );
  NAND U6297 ( .A(n5747), .B(n5746), .Z(n6044) );
  XNOR U6298 ( .A(n6043), .B(n6044), .Z(n6040) );
  NAND U6299 ( .A(x[155]), .B(y[675]), .Z(n5885) );
  NAND U6300 ( .A(x[129]), .B(y[701]), .Z(n5884) );
  XNOR U6301 ( .A(n5885), .B(n5884), .Z(n5883) );
  XNOR U6302 ( .A(n5882), .B(n5883), .Z(n5843) );
  AND U6303 ( .A(y[690]), .B(x[140]), .Z(n5752) );
  XNOR U6304 ( .A(n5752), .B(n5751), .Z(n5870) );
  XNOR U6305 ( .A(n5869), .B(n5870), .Z(n5923) );
  AND U6306 ( .A(x[138]), .B(y[692]), .Z(n5754) );
  AND U6307 ( .A(x[137]), .B(y[693]), .Z(n5753) );
  XNOR U6308 ( .A(n5754), .B(n5753), .Z(n5922) );
  XNOR U6309 ( .A(n5923), .B(n5922), .Z(n5845) );
  OR U6310 ( .A(n5756), .B(n5755), .Z(n5760) );
  OR U6311 ( .A(n5758), .B(n5757), .Z(n5759) );
  AND U6312 ( .A(n5760), .B(n5759), .Z(n5846) );
  XNOR U6313 ( .A(n5845), .B(n5846), .Z(n5844) );
  XOR U6314 ( .A(n5843), .B(n5844), .Z(n5825) );
  XNOR U6315 ( .A(n5826), .B(n5825), .Z(n5824) );
  OR U6316 ( .A(n5762), .B(n5761), .Z(n5766) );
  NANDN U6317 ( .A(n5764), .B(n5763), .Z(n5765) );
  NAND U6318 ( .A(n5766), .B(n5765), .Z(n5823) );
  XOR U6319 ( .A(n5824), .B(n5823), .Z(n6039) );
  XOR U6320 ( .A(n6040), .B(n6039), .Z(n6038) );
  OR U6321 ( .A(n5768), .B(n5767), .Z(n5772) );
  OR U6322 ( .A(n5770), .B(n5769), .Z(n5771) );
  NAND U6323 ( .A(n5772), .B(n5771), .Z(n6037) );
  XOR U6324 ( .A(n6038), .B(n6037), .Z(n6061) );
  XNOR U6325 ( .A(n6060), .B(n6059), .Z(n6078) );
  NANDN U6326 ( .A(n5774), .B(n5773), .Z(n5778) );
  OR U6327 ( .A(n5776), .B(n5775), .Z(n5777) );
  AND U6328 ( .A(n5778), .B(n5777), .Z(n6085) );
  OR U6329 ( .A(n5780), .B(n5779), .Z(n5784) );
  OR U6330 ( .A(n5782), .B(n5781), .Z(n5783) );
  AND U6331 ( .A(n5784), .B(n5783), .Z(n6083) );
  OR U6332 ( .A(n5786), .B(n5785), .Z(n5790) );
  OR U6333 ( .A(n5788), .B(n5787), .Z(n5789) );
  NAND U6334 ( .A(n5790), .B(n5789), .Z(n6084) );
  XNOR U6335 ( .A(n6083), .B(n6084), .Z(n6086) );
  XOR U6336 ( .A(n6085), .B(n6086), .Z(n6077) );
  XNOR U6337 ( .A(n6078), .B(n6077), .Z(n6079) );
  XOR U6338 ( .A(n6080), .B(n6079), .Z(n5791) );
  XOR U6339 ( .A(n5792), .B(n5791), .Z(N127) );
  NANDN U6340 ( .A(n5792), .B(n5791), .Z(n5796) );
  OR U6341 ( .A(n5794), .B(n5793), .Z(n5795) );
  AND U6342 ( .A(n5796), .B(n5795), .Z(n6076) );
  OR U6343 ( .A(n5798), .B(n5797), .Z(n5802) );
  OR U6344 ( .A(n5800), .B(n5799), .Z(n5801) );
  AND U6345 ( .A(n5802), .B(n5801), .Z(n6058) );
  NANDN U6346 ( .A(n5804), .B(n5803), .Z(n5808) );
  OR U6347 ( .A(n5806), .B(n5805), .Z(n5807) );
  AND U6348 ( .A(n5808), .B(n5807), .Z(n5816) );
  OR U6349 ( .A(n5810), .B(n5809), .Z(n5814) );
  OR U6350 ( .A(n5812), .B(n5811), .Z(n5813) );
  NAND U6351 ( .A(n5814), .B(n5813), .Z(n5815) );
  XNOR U6352 ( .A(n5816), .B(n5815), .Z(n6056) );
  OR U6353 ( .A(n5818), .B(n5817), .Z(n5822) );
  OR U6354 ( .A(n5820), .B(n5819), .Z(n5821) );
  AND U6355 ( .A(n5822), .B(n5821), .Z(n6054) );
  OR U6356 ( .A(n5824), .B(n5823), .Z(n5828) );
  OR U6357 ( .A(n5826), .B(n5825), .Z(n5827) );
  AND U6358 ( .A(n5828), .B(n5827), .Z(n6036) );
  OR U6359 ( .A(n5830), .B(n5829), .Z(n5834) );
  NANDN U6360 ( .A(n5832), .B(n5831), .Z(n5833) );
  AND U6361 ( .A(n5834), .B(n5833), .Z(n5842) );
  NOR U6362 ( .A(n5836), .B(n5835), .Z(n5840) );
  ANDN U6363 ( .B(n5838), .A(n5837), .Z(n5839) );
  OR U6364 ( .A(n5840), .B(n5839), .Z(n5841) );
  XNOR U6365 ( .A(n5842), .B(n5841), .Z(n6034) );
  OR U6366 ( .A(n5844), .B(n5843), .Z(n5848) );
  OR U6367 ( .A(n5846), .B(n5845), .Z(n5847) );
  AND U6368 ( .A(n5848), .B(n5847), .Z(n6032) );
  OR U6369 ( .A(n5850), .B(n5849), .Z(n5854) );
  OR U6370 ( .A(n5852), .B(n5851), .Z(n5853) );
  AND U6371 ( .A(n5854), .B(n5853), .Z(n5862) );
  NANDN U6372 ( .A(n5856), .B(n5855), .Z(n5860) );
  NANDN U6373 ( .A(n5858), .B(n5857), .Z(n5859) );
  NAND U6374 ( .A(n5860), .B(n5859), .Z(n5861) );
  XNOR U6375 ( .A(n5862), .B(n5861), .Z(n6030) );
  OR U6376 ( .A(n5864), .B(n5863), .Z(n5868) );
  NANDN U6377 ( .A(n5866), .B(n5865), .Z(n5867) );
  AND U6378 ( .A(n5868), .B(n5867), .Z(n6028) );
  NANDN U6379 ( .A(n5870), .B(n5869), .Z(n5873) );
  NAND U6380 ( .A(n5871), .B(n5959), .Z(n5872) );
  AND U6381 ( .A(n5873), .B(n5872), .Z(n5881) );
  NANDN U6382 ( .A(n5875), .B(n5874), .Z(n5879) );
  NANDN U6383 ( .A(n5877), .B(n5876), .Z(n5878) );
  NAND U6384 ( .A(n5879), .B(n5878), .Z(n5880) );
  XNOR U6385 ( .A(n5881), .B(n5880), .Z(n5920) );
  NANDN U6386 ( .A(n5883), .B(n5882), .Z(n5887) );
  OR U6387 ( .A(n5885), .B(n5884), .Z(n5886) );
  AND U6388 ( .A(n5887), .B(n5886), .Z(n5918) );
  OR U6389 ( .A(n5889), .B(n5888), .Z(n5892) );
  NAND U6390 ( .A(x[153]), .B(y[678]), .Z(n5960) );
  NANDN U6391 ( .A(n5960), .B(n5890), .Z(n5891) );
  AND U6392 ( .A(n5892), .B(n5891), .Z(n5900) );
  OR U6393 ( .A(n5894), .B(n5893), .Z(n5898) );
  OR U6394 ( .A(n5896), .B(n5895), .Z(n5897) );
  NAND U6395 ( .A(n5898), .B(n5897), .Z(n5899) );
  XNOR U6396 ( .A(n5900), .B(n5899), .Z(n5916) );
  AND U6397 ( .A(x[158]), .B(y[673]), .Z(n5902) );
  NAND U6398 ( .A(x[157]), .B(y[674]), .Z(n5901) );
  XNOR U6399 ( .A(n5902), .B(n5901), .Z(n5906) );
  AND U6400 ( .A(x[151]), .B(y[680]), .Z(n5904) );
  NAND U6401 ( .A(x[155]), .B(y[676]), .Z(n5903) );
  XNOR U6402 ( .A(n5904), .B(n5903), .Z(n5905) );
  XOR U6403 ( .A(n5906), .B(n5905), .Z(n5914) );
  AND U6404 ( .A(y[691]), .B(x[140]), .Z(n5908) );
  NAND U6405 ( .A(x[139]), .B(y[692]), .Z(n5907) );
  XNOR U6406 ( .A(n5908), .B(n5907), .Z(n5912) );
  AND U6407 ( .A(x[156]), .B(y[675]), .Z(n5910) );
  NAND U6408 ( .A(x[154]), .B(y[677]), .Z(n5909) );
  XNOR U6409 ( .A(n5910), .B(n5909), .Z(n5911) );
  XNOR U6410 ( .A(n5912), .B(n5911), .Z(n5913) );
  XNOR U6411 ( .A(n5914), .B(n5913), .Z(n5915) );
  XNOR U6412 ( .A(n5916), .B(n5915), .Z(n5917) );
  XNOR U6413 ( .A(n5918), .B(n5917), .Z(n5919) );
  XOR U6414 ( .A(n5920), .B(n5919), .Z(n5951) );
  NAND U6415 ( .A(x[138]), .B(y[693]), .Z(n6018) );
  ANDN U6416 ( .B(n5921), .A(n6018), .Z(n5925) );
  ANDN U6417 ( .B(n5923), .A(n5922), .Z(n5924) );
  NOR U6418 ( .A(n5925), .B(n5924), .Z(n5933) );
  NANDN U6419 ( .A(n5927), .B(n5926), .Z(n5931) );
  NANDN U6420 ( .A(n5929), .B(n5928), .Z(n5930) );
  AND U6421 ( .A(n5931), .B(n5930), .Z(n5932) );
  XNOR U6422 ( .A(n5933), .B(n5932), .Z(n5949) );
  OR U6423 ( .A(n5935), .B(n5934), .Z(n5939) );
  OR U6424 ( .A(n5937), .B(n5936), .Z(n5938) );
  AND U6425 ( .A(n5939), .B(n5938), .Z(n5947) );
  NANDN U6426 ( .A(n5941), .B(n5940), .Z(n5945) );
  NANDN U6427 ( .A(n5943), .B(n5942), .Z(n5944) );
  NAND U6428 ( .A(n5945), .B(n5944), .Z(n5946) );
  XNOR U6429 ( .A(n5947), .B(n5946), .Z(n5948) );
  XOR U6430 ( .A(n5949), .B(n5948), .Z(n5950) );
  XNOR U6431 ( .A(n5951), .B(n5950), .Z(n6026) );
  NAND U6432 ( .A(n5953), .B(n5952), .Z(n5957) );
  OR U6433 ( .A(n5955), .B(n5954), .Z(n5956) );
  AND U6434 ( .A(n5957), .B(n5956), .Z(n6024) );
  AND U6435 ( .A(y[703]), .B(x[128]), .Z(n5966) );
  ANDN U6436 ( .B(o[62]), .A(n5958), .Z(n5964) );
  XOR U6437 ( .A(n5959), .B(o[63]), .Z(n5962) );
  NAND U6438 ( .A(x[150]), .B(y[681]), .Z(n6000) );
  XNOR U6439 ( .A(n6000), .B(n5960), .Z(n5961) );
  XNOR U6440 ( .A(n5962), .B(n5961), .Z(n5963) );
  XNOR U6441 ( .A(n5964), .B(n5963), .Z(n5965) );
  XNOR U6442 ( .A(n5966), .B(n5965), .Z(n5974) );
  AND U6443 ( .A(y[694]), .B(x[137]), .Z(n5968) );
  NAND U6444 ( .A(x[142]), .B(y[689]), .Z(n5967) );
  XNOR U6445 ( .A(n5968), .B(n5967), .Z(n5972) );
  AND U6446 ( .A(y[688]), .B(x[143]), .Z(n5970) );
  NAND U6447 ( .A(x[129]), .B(y[702]), .Z(n5969) );
  XNOR U6448 ( .A(n5970), .B(n5969), .Z(n5971) );
  XNOR U6449 ( .A(n5972), .B(n5971), .Z(n5973) );
  XNOR U6450 ( .A(n5974), .B(n5973), .Z(n6022) );
  AND U6451 ( .A(y[686]), .B(x[145]), .Z(n5976) );
  NAND U6452 ( .A(x[130]), .B(y[701]), .Z(n5975) );
  XNOR U6453 ( .A(n5976), .B(n5975), .Z(n5980) );
  AND U6454 ( .A(y[695]), .B(x[136]), .Z(n5978) );
  NAND U6455 ( .A(x[149]), .B(y[682]), .Z(n5977) );
  XNOR U6456 ( .A(n5978), .B(n5977), .Z(n5979) );
  XOR U6457 ( .A(n5980), .B(n5979), .Z(n5988) );
  AND U6458 ( .A(y[698]), .B(x[133]), .Z(n5982) );
  NAND U6459 ( .A(x[135]), .B(y[696]), .Z(n5981) );
  XNOR U6460 ( .A(n5982), .B(n5981), .Z(n5986) );
  AND U6461 ( .A(x[159]), .B(y[672]), .Z(n5984) );
  NAND U6462 ( .A(x[147]), .B(y[684]), .Z(n5983) );
  XNOR U6463 ( .A(n5984), .B(n5983), .Z(n5985) );
  XNOR U6464 ( .A(n5986), .B(n5985), .Z(n5987) );
  XNOR U6465 ( .A(n5988), .B(n5987), .Z(n5996) );
  AND U6466 ( .A(y[699]), .B(x[132]), .Z(n5990) );
  NAND U6467 ( .A(x[152]), .B(y[679]), .Z(n5989) );
  XNOR U6468 ( .A(n5990), .B(n5989), .Z(n5994) );
  AND U6469 ( .A(y[700]), .B(x[131]), .Z(n5992) );
  NAND U6470 ( .A(x[134]), .B(y[697]), .Z(n5991) );
  XNOR U6471 ( .A(n5992), .B(n5991), .Z(n5993) );
  XNOR U6472 ( .A(n5994), .B(n5993), .Z(n5995) );
  XNOR U6473 ( .A(n5996), .B(n5995), .Z(n6012) );
  OR U6474 ( .A(n5998), .B(n5997), .Z(n6002) );
  NANDN U6475 ( .A(n6000), .B(n5999), .Z(n6001) );
  AND U6476 ( .A(n6002), .B(n6001), .Z(n6010) );
  NANDN U6477 ( .A(n6004), .B(n6003), .Z(n6008) );
  NANDN U6478 ( .A(n6006), .B(n6005), .Z(n6007) );
  NAND U6479 ( .A(n6008), .B(n6007), .Z(n6009) );
  XNOR U6480 ( .A(n6010), .B(n6009), .Z(n6011) );
  XOR U6481 ( .A(n6012), .B(n6011), .Z(n6020) );
  AND U6482 ( .A(x[146]), .B(y[685]), .Z(n6014) );
  NAND U6483 ( .A(x[148]), .B(y[683]), .Z(n6013) );
  XNOR U6484 ( .A(n6014), .B(n6013), .Z(n6016) );
  NAND U6485 ( .A(x[144]), .B(y[687]), .Z(n6015) );
  XNOR U6486 ( .A(n6016), .B(n6015), .Z(n6017) );
  XOR U6487 ( .A(n6018), .B(n6017), .Z(n6019) );
  XNOR U6488 ( .A(n6020), .B(n6019), .Z(n6021) );
  XNOR U6489 ( .A(n6022), .B(n6021), .Z(n6023) );
  XNOR U6490 ( .A(n6024), .B(n6023), .Z(n6025) );
  XNOR U6491 ( .A(n6026), .B(n6025), .Z(n6027) );
  XNOR U6492 ( .A(n6028), .B(n6027), .Z(n6029) );
  XNOR U6493 ( .A(n6030), .B(n6029), .Z(n6031) );
  XNOR U6494 ( .A(n6032), .B(n6031), .Z(n6033) );
  XNOR U6495 ( .A(n6034), .B(n6033), .Z(n6035) );
  XNOR U6496 ( .A(n6036), .B(n6035), .Z(n6052) );
  OR U6497 ( .A(n6038), .B(n6037), .Z(n6042) );
  NANDN U6498 ( .A(n6040), .B(n6039), .Z(n6041) );
  AND U6499 ( .A(n6042), .B(n6041), .Z(n6050) );
  NANDN U6500 ( .A(n6044), .B(n6043), .Z(n6048) );
  OR U6501 ( .A(n6046), .B(n6045), .Z(n6047) );
  NAND U6502 ( .A(n6048), .B(n6047), .Z(n6049) );
  XNOR U6503 ( .A(n6050), .B(n6049), .Z(n6051) );
  XNOR U6504 ( .A(n6052), .B(n6051), .Z(n6053) );
  XNOR U6505 ( .A(n6054), .B(n6053), .Z(n6055) );
  XNOR U6506 ( .A(n6056), .B(n6055), .Z(n6057) );
  XNOR U6507 ( .A(n6058), .B(n6057), .Z(n6074) );
  NANDN U6508 ( .A(n6060), .B(n6059), .Z(n6064) );
  NANDN U6509 ( .A(n6062), .B(n6061), .Z(n6063) );
  AND U6510 ( .A(n6064), .B(n6063), .Z(n6072) );
  NANDN U6511 ( .A(n6066), .B(n6065), .Z(n6070) );
  OR U6512 ( .A(n6068), .B(n6067), .Z(n6069) );
  NAND U6513 ( .A(n6070), .B(n6069), .Z(n6071) );
  XNOR U6514 ( .A(n6072), .B(n6071), .Z(n6073) );
  XNOR U6515 ( .A(n6074), .B(n6073), .Z(n6075) );
  XNOR U6516 ( .A(n6076), .B(n6075), .Z(n6092) );
  NOR U6517 ( .A(n6078), .B(n6077), .Z(n6082) );
  NOR U6518 ( .A(n6080), .B(n6079), .Z(n6081) );
  NOR U6519 ( .A(n6082), .B(n6081), .Z(n6090) );
  OR U6520 ( .A(n6084), .B(n6083), .Z(n6088) );
  OR U6521 ( .A(n6086), .B(n6085), .Z(n6087) );
  AND U6522 ( .A(n6088), .B(n6087), .Z(n6089) );
  XNOR U6523 ( .A(n6090), .B(n6089), .Z(n6091) );
  XNOR U6524 ( .A(n6092), .B(n6091), .Z(N128) );
  AND U6525 ( .A(y[704]), .B(x[128]), .Z(n6773) );
  XOR U6526 ( .A(n6773), .B(o[64]), .Z(N161) );
  AND U6527 ( .A(y[704]), .B(x[129]), .Z(n6093) );
  NAND U6528 ( .A(x[128]), .B(y[705]), .Z(n6099) );
  XNOR U6529 ( .A(n6099), .B(o[65]), .Z(n6094) );
  XOR U6530 ( .A(n6093), .B(n6094), .Z(n6095) );
  AND U6531 ( .A(o[64]), .B(n6773), .Z(n6096) );
  XOR U6532 ( .A(n6095), .B(n6096), .Z(N162) );
  OR U6533 ( .A(n6094), .B(n6093), .Z(n6098) );
  NANDN U6534 ( .A(n6096), .B(n6095), .Z(n6097) );
  NAND U6535 ( .A(n6098), .B(n6097), .Z(n6101) );
  NAND U6536 ( .A(x[128]), .B(y[706]), .Z(n6112) );
  XOR U6537 ( .A(n6112), .B(o[66]), .Z(n6100) );
  XNOR U6538 ( .A(n6101), .B(n6100), .Z(n6103) );
  ANDN U6539 ( .B(o[65]), .A(n6099), .Z(n6106) );
  ANDN U6540 ( .B(y[704]), .A(n153), .Z(n6107) );
  XNOR U6541 ( .A(n6106), .B(n6107), .Z(n6109) );
  ANDN U6542 ( .B(y[705]), .A(n152), .Z(n6108) );
  XNOR U6543 ( .A(n6109), .B(n6108), .Z(n6102) );
  XNOR U6544 ( .A(n6103), .B(n6102), .Z(N163) );
  NAND U6545 ( .A(n6101), .B(n6100), .Z(n6105) );
  OR U6546 ( .A(n6103), .B(n6102), .Z(n6104) );
  NAND U6547 ( .A(n6105), .B(n6104), .Z(n6115) );
  OR U6548 ( .A(n6107), .B(n6106), .Z(n6111) );
  OR U6549 ( .A(n6109), .B(n6108), .Z(n6110) );
  AND U6550 ( .A(n6111), .B(n6110), .Z(n6116) );
  XNOR U6551 ( .A(n6115), .B(n6116), .Z(n6117) );
  AND U6552 ( .A(y[706]), .B(x[129]), .Z(n6154) );
  NAND U6553 ( .A(x[130]), .B(y[705]), .Z(n6130) );
  XOR U6554 ( .A(o[67]), .B(n6130), .Z(n6121) );
  XOR U6555 ( .A(n6154), .B(n6121), .Z(n6123) );
  NANDN U6556 ( .A(n6112), .B(o[66]), .Z(n6127) );
  AND U6557 ( .A(y[704]), .B(x[131]), .Z(n6114) );
  NAND U6558 ( .A(x[128]), .B(y[707]), .Z(n6113) );
  XNOR U6559 ( .A(n6114), .B(n6113), .Z(n6126) );
  XNOR U6560 ( .A(n6123), .B(n6122), .Z(n6118) );
  XOR U6561 ( .A(n6117), .B(n6118), .Z(N164) );
  NANDN U6562 ( .A(n6116), .B(n6115), .Z(n6120) );
  NANDN U6563 ( .A(n6118), .B(n6117), .Z(n6119) );
  NAND U6564 ( .A(n6120), .B(n6119), .Z(n6135) );
  NANDN U6565 ( .A(n6121), .B(n6154), .Z(n6125) );
  NANDN U6566 ( .A(n6123), .B(n6122), .Z(n6124) );
  NAND U6567 ( .A(n6125), .B(n6124), .Z(n6136) );
  XNOR U6568 ( .A(n6135), .B(n6136), .Z(n6137) );
  ANDN U6569 ( .B(y[707]), .A(n154), .Z(n6202) );
  NAND U6570 ( .A(n6773), .B(n6202), .Z(n6129) );
  NANDN U6571 ( .A(n6127), .B(n6126), .Z(n6128) );
  NAND U6572 ( .A(n6129), .B(n6128), .Z(n6144) );
  NANDN U6573 ( .A(n6130), .B(o[67]), .Z(n6151) );
  AND U6574 ( .A(y[704]), .B(x[132]), .Z(n6132) );
  AND U6575 ( .A(y[708]), .B(x[128]), .Z(n6131) );
  XNOR U6576 ( .A(n6132), .B(n6131), .Z(n6150) );
  XOR U6577 ( .A(n6151), .B(n6150), .Z(n6142) );
  AND U6578 ( .A(x[129]), .B(y[707]), .Z(n6134) );
  NAND U6579 ( .A(x[130]), .B(y[706]), .Z(n6133) );
  XOR U6580 ( .A(n6134), .B(n6133), .Z(n6156) );
  NAND U6581 ( .A(x[131]), .B(y[705]), .Z(n6147) );
  XNOR U6582 ( .A(n6147), .B(o[68]), .Z(n6155) );
  XOR U6583 ( .A(n6144), .B(n6143), .Z(n6138) );
  XOR U6584 ( .A(n6137), .B(n6138), .Z(N165) );
  NANDN U6585 ( .A(n6136), .B(n6135), .Z(n6140) );
  NANDN U6586 ( .A(n6138), .B(n6137), .Z(n6139) );
  NAND U6587 ( .A(n6140), .B(n6139), .Z(n6159) );
  NAND U6588 ( .A(n6142), .B(n6141), .Z(n6146) );
  NAND U6589 ( .A(n6144), .B(n6143), .Z(n6145) );
  NAND U6590 ( .A(n6146), .B(n6145), .Z(n6160) );
  XNOR U6591 ( .A(n6159), .B(n6160), .Z(n6161) );
  NANDN U6592 ( .A(n6147), .B(o[68]), .Z(n6178) );
  AND U6593 ( .A(y[704]), .B(x[133]), .Z(n6149) );
  AND U6594 ( .A(y[709]), .B(x[128]), .Z(n6148) );
  XNOR U6595 ( .A(n6149), .B(n6148), .Z(n6177) );
  XOR U6596 ( .A(n6178), .B(n6177), .Z(n6173) );
  ANDN U6597 ( .B(y[707]), .A(n153), .Z(n6171) );
  ANDN U6598 ( .B(y[708]), .A(n152), .Z(n6186) );
  ANDN U6599 ( .B(y[705]), .A(n155), .Z(n6181) );
  XOR U6600 ( .A(o[69]), .B(n6181), .Z(n6184) );
  ANDN U6601 ( .B(y[706]), .A(n154), .Z(n6185) );
  XNOR U6602 ( .A(n6184), .B(n6185), .Z(n6187) );
  XNOR U6603 ( .A(n6186), .B(n6187), .Z(n6172) );
  XNOR U6604 ( .A(n6171), .B(n6172), .Z(n6174) );
  XNOR U6605 ( .A(n6173), .B(n6174), .Z(n6168) );
  ANDN U6606 ( .B(y[708]), .A(n155), .Z(n6290) );
  NAND U6607 ( .A(n6773), .B(n6290), .Z(n6153) );
  OR U6608 ( .A(n6151), .B(n6150), .Z(n6152) );
  NAND U6609 ( .A(n6153), .B(n6152), .Z(n6166) );
  NAND U6610 ( .A(n6154), .B(n6171), .Z(n6158) );
  NANDN U6611 ( .A(n6156), .B(n6155), .Z(n6157) );
  NAND U6612 ( .A(n6158), .B(n6157), .Z(n6165) );
  XNOR U6613 ( .A(n6166), .B(n6165), .Z(n6167) );
  XNOR U6614 ( .A(n6168), .B(n6167), .Z(n6162) );
  XOR U6615 ( .A(n6161), .B(n6162), .Z(N166) );
  NANDN U6616 ( .A(n6160), .B(n6159), .Z(n6164) );
  NANDN U6617 ( .A(n6162), .B(n6161), .Z(n6163) );
  NAND U6618 ( .A(n6164), .B(n6163), .Z(n6190) );
  OR U6619 ( .A(n6166), .B(n6165), .Z(n6170) );
  OR U6620 ( .A(n6168), .B(n6167), .Z(n6169) );
  AND U6621 ( .A(n6170), .B(n6169), .Z(n6191) );
  XNOR U6622 ( .A(n6190), .B(n6191), .Z(n6192) );
  OR U6623 ( .A(n6172), .B(n6171), .Z(n6176) );
  OR U6624 ( .A(n6174), .B(n6173), .Z(n6175) );
  AND U6625 ( .A(n6176), .B(n6175), .Z(n6196) );
  NAND U6626 ( .A(x[133]), .B(y[709]), .Z(n6520) );
  NANDN U6627 ( .A(n6520), .B(n6773), .Z(n6180) );
  OR U6628 ( .A(n6178), .B(n6177), .Z(n6179) );
  NAND U6629 ( .A(n6180), .B(n6179), .Z(n6218) );
  NAND U6630 ( .A(n6181), .B(o[69]), .Z(n6208) );
  AND U6631 ( .A(y[704]), .B(x[134]), .Z(n6183) );
  AND U6632 ( .A(x[128]), .B(y[710]), .Z(n6182) );
  XNOR U6633 ( .A(n6183), .B(n6182), .Z(n6207) );
  XOR U6634 ( .A(n6208), .B(n6207), .Z(n6217) );
  XNOR U6635 ( .A(n6218), .B(n6217), .Z(n6220) );
  AND U6636 ( .A(y[709]), .B(x[129]), .Z(n6468) );
  NAND U6637 ( .A(x[133]), .B(y[705]), .Z(n6211) );
  XNOR U6638 ( .A(n6211), .B(o[70]), .Z(n6212) );
  XNOR U6639 ( .A(n6468), .B(n6212), .Z(n6214) );
  AND U6640 ( .A(y[706]), .B(x[132]), .Z(n6213) );
  XOR U6641 ( .A(n6214), .B(n6213), .Z(n6203) );
  AND U6642 ( .A(y[708]), .B(x[130]), .Z(n6509) );
  XNOR U6643 ( .A(n6202), .B(n6509), .Z(n6204) );
  XOR U6644 ( .A(n6203), .B(n6204), .Z(n6219) );
  XNOR U6645 ( .A(n6220), .B(n6219), .Z(n6197) );
  XOR U6646 ( .A(n6196), .B(n6197), .Z(n6198) );
  OR U6647 ( .A(n6185), .B(n6184), .Z(n6189) );
  OR U6648 ( .A(n6187), .B(n6186), .Z(n6188) );
  AND U6649 ( .A(n6189), .B(n6188), .Z(n6199) );
  XOR U6650 ( .A(n6192), .B(n6193), .Z(N167) );
  NANDN U6651 ( .A(n6191), .B(n6190), .Z(n6195) );
  NANDN U6652 ( .A(n6193), .B(n6192), .Z(n6194) );
  NAND U6653 ( .A(n6195), .B(n6194), .Z(n6252) );
  OR U6654 ( .A(n6197), .B(n6196), .Z(n6201) );
  NANDN U6655 ( .A(n6199), .B(n6198), .Z(n6200) );
  AND U6656 ( .A(n6201), .B(n6200), .Z(n6253) );
  XNOR U6657 ( .A(n6252), .B(n6253), .Z(n6254) );
  OR U6658 ( .A(n6202), .B(n6509), .Z(n6206) );
  NANDN U6659 ( .A(n6204), .B(n6203), .Z(n6205) );
  NAND U6660 ( .A(n6206), .B(n6205), .Z(n6249) );
  AND U6661 ( .A(y[710]), .B(x[134]), .Z(n6484) );
  NAND U6662 ( .A(n6773), .B(n6484), .Z(n6210) );
  OR U6663 ( .A(n6208), .B(n6207), .Z(n6209) );
  AND U6664 ( .A(n6210), .B(n6209), .Z(n6247) );
  ANDN U6665 ( .B(y[706]), .A(n156), .Z(n6383) );
  ANDN U6666 ( .B(y[710]), .A(n152), .Z(n6602) );
  NAND U6667 ( .A(x[134]), .B(y[705]), .Z(n6241) );
  XNOR U6668 ( .A(o[71]), .B(n6241), .Z(n6242) );
  XNOR U6669 ( .A(n6602), .B(n6242), .Z(n6243) );
  XNOR U6670 ( .A(n6383), .B(n6243), .Z(n6246) );
  XOR U6671 ( .A(n6247), .B(n6246), .Z(n6248) );
  XNOR U6672 ( .A(n6249), .B(n6248), .Z(n6258) );
  ANDN U6673 ( .B(y[709]), .A(n153), .Z(n6697) );
  ANDN U6674 ( .B(y[707]), .A(n155), .Z(n6405) );
  ANDN U6675 ( .B(y[708]), .A(n154), .Z(n6231) );
  XNOR U6676 ( .A(n6405), .B(n6231), .Z(n6232) );
  XOR U6677 ( .A(n6697), .B(n6232), .Z(n6235) );
  NAND U6678 ( .A(x[128]), .B(y[711]), .Z(n6227) );
  ANDN U6679 ( .B(o[70]), .A(n6211), .Z(n6226) );
  NAND U6680 ( .A(x[135]), .B(y[704]), .Z(n6225) );
  XOR U6681 ( .A(n6226), .B(n6225), .Z(n6228) );
  XNOR U6682 ( .A(n6227), .B(n6228), .Z(n6236) );
  XNOR U6683 ( .A(n6235), .B(n6236), .Z(n6238) );
  NAND U6684 ( .A(n6468), .B(n6212), .Z(n6216) );
  NANDN U6685 ( .A(n6214), .B(n6213), .Z(n6215) );
  AND U6686 ( .A(n6216), .B(n6215), .Z(n6237) );
  XOR U6687 ( .A(n6238), .B(n6237), .Z(n6259) );
  XOR U6688 ( .A(n6258), .B(n6259), .Z(n6261) );
  OR U6689 ( .A(n6218), .B(n6217), .Z(n6222) );
  OR U6690 ( .A(n6220), .B(n6219), .Z(n6221) );
  AND U6691 ( .A(n6222), .B(n6221), .Z(n6260) );
  XOR U6692 ( .A(n6261), .B(n6260), .Z(n6255) );
  XNOR U6693 ( .A(n6254), .B(n6255), .Z(N168) );
  AND U6694 ( .A(y[704]), .B(x[136]), .Z(n6224) );
  NAND U6695 ( .A(x[128]), .B(y[712]), .Z(n6223) );
  XOR U6696 ( .A(n6224), .B(n6223), .Z(n6277) );
  NAND U6697 ( .A(x[135]), .B(y[705]), .Z(n6280) );
  XNOR U6698 ( .A(n6280), .B(o[72]), .Z(n6276) );
  XOR U6699 ( .A(n6277), .B(n6276), .Z(n6271) );
  NANDN U6700 ( .A(n6226), .B(n6225), .Z(n6230) );
  NANDN U6701 ( .A(n6228), .B(n6227), .Z(n6229) );
  NAND U6702 ( .A(n6230), .B(n6229), .Z(n6270) );
  XOR U6703 ( .A(n6271), .B(n6270), .Z(n6272) );
  OR U6704 ( .A(n6231), .B(n6405), .Z(n6234) );
  OR U6705 ( .A(n6232), .B(n6697), .Z(n6233) );
  NAND U6706 ( .A(n6234), .B(n6233), .Z(n6273) );
  XNOR U6707 ( .A(n6272), .B(n6273), .Z(n6306) );
  OR U6708 ( .A(n6236), .B(n6235), .Z(n6240) );
  OR U6709 ( .A(n6238), .B(n6237), .Z(n6239) );
  AND U6710 ( .A(n6240), .B(n6239), .Z(n6266) );
  ANDN U6711 ( .B(y[706]), .A(n157), .Z(n6291) );
  XNOR U6712 ( .A(n6290), .B(n6291), .Z(n6292) );
  NOR U6713 ( .A(n153), .B(n148), .Z(n6789) );
  XNOR U6714 ( .A(n6292), .B(n6789), .Z(n6293) );
  ANDN U6715 ( .B(y[709]), .A(n154), .Z(n7106) );
  XNOR U6716 ( .A(n6293), .B(n7106), .Z(n6295) );
  NANDN U6717 ( .A(n6241), .B(o[71]), .Z(n6287) );
  AND U6718 ( .A(y[707]), .B(x[133]), .Z(n6907) );
  AND U6719 ( .A(y[711]), .B(x[129]), .Z(n6768) );
  XNOR U6720 ( .A(n6907), .B(n6768), .Z(n6286) );
  XOR U6721 ( .A(n6287), .B(n6286), .Z(n6294) );
  XNOR U6722 ( .A(n6295), .B(n6294), .Z(n6264) );
  NAND U6723 ( .A(n6602), .B(n6242), .Z(n6245) );
  NANDN U6724 ( .A(n6243), .B(n6383), .Z(n6244) );
  AND U6725 ( .A(n6245), .B(n6244), .Z(n6265) );
  XOR U6726 ( .A(n6264), .B(n6265), .Z(n6267) );
  XOR U6727 ( .A(n6266), .B(n6267), .Z(n6304) );
  NANDN U6728 ( .A(n6247), .B(n6246), .Z(n6251) );
  OR U6729 ( .A(n6249), .B(n6248), .Z(n6250) );
  NAND U6730 ( .A(n6251), .B(n6250), .Z(n6305) );
  XNOR U6731 ( .A(n6304), .B(n6305), .Z(n6307) );
  XNOR U6732 ( .A(n6306), .B(n6307), .Z(n6301) );
  NANDN U6733 ( .A(n6253), .B(n6252), .Z(n6257) );
  NAND U6734 ( .A(n6255), .B(n6254), .Z(n6256) );
  NAND U6735 ( .A(n6257), .B(n6256), .Z(n6298) );
  NANDN U6736 ( .A(n6259), .B(n6258), .Z(n6263) );
  OR U6737 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U6738 ( .A(n6263), .B(n6262), .Z(n6299) );
  XNOR U6739 ( .A(n6298), .B(n6299), .Z(n6300) );
  XOR U6740 ( .A(n6301), .B(n6300), .Z(N169) );
  NANDN U6741 ( .A(n6265), .B(n6264), .Z(n6269) );
  OR U6742 ( .A(n6267), .B(n6266), .Z(n6268) );
  NAND U6743 ( .A(n6269), .B(n6268), .Z(n6317) );
  OR U6744 ( .A(n6271), .B(n6270), .Z(n6275) );
  NANDN U6745 ( .A(n6273), .B(n6272), .Z(n6274) );
  NAND U6746 ( .A(n6275), .B(n6274), .Z(n6316) );
  XOR U6747 ( .A(n6317), .B(n6316), .Z(n6318) );
  AND U6748 ( .A(y[712]), .B(x[136]), .Z(n6786) );
  NAND U6749 ( .A(n6773), .B(n6786), .Z(n6279) );
  NANDN U6750 ( .A(n6277), .B(n6276), .Z(n6278) );
  NAND U6751 ( .A(n6279), .B(n6278), .Z(n6325) );
  NANDN U6752 ( .A(n6280), .B(o[72]), .Z(n6354) );
  AND U6753 ( .A(y[708]), .B(x[133]), .Z(n6281) );
  AND U6754 ( .A(y[706]), .B(x[135]), .Z(n6701) );
  XNOR U6755 ( .A(n6281), .B(n6701), .Z(n6353) );
  XOR U6756 ( .A(n6354), .B(n6353), .Z(n6323) );
  AND U6757 ( .A(y[704]), .B(x[137]), .Z(n6283) );
  NAND U6758 ( .A(x[128]), .B(y[713]), .Z(n6282) );
  XOR U6759 ( .A(n6283), .B(n6282), .Z(n6348) );
  NAND U6760 ( .A(x[136]), .B(y[705]), .Z(n6342) );
  XOR U6761 ( .A(n6342), .B(o[73]), .Z(n6347) );
  XNOR U6762 ( .A(n6348), .B(n6347), .Z(n6322) );
  XNOR U6763 ( .A(n6323), .B(n6322), .Z(n6324) );
  XNOR U6764 ( .A(n6325), .B(n6324), .Z(n6332) );
  NAND U6765 ( .A(x[132]), .B(y[709]), .Z(n6780) );
  AND U6766 ( .A(x[134]), .B(y[707]), .Z(n6285) );
  NAND U6767 ( .A(x[129]), .B(y[712]), .Z(n6284) );
  XNOR U6768 ( .A(n6285), .B(n6284), .Z(n6344) );
  XNOR U6769 ( .A(n6780), .B(n6344), .Z(n6328) );
  NOR U6770 ( .A(n154), .B(n148), .Z(n6670) );
  ANDN U6771 ( .B(y[711]), .A(n153), .Z(n6995) );
  XNOR U6772 ( .A(n6670), .B(n6995), .Z(n6329) );
  XNOR U6773 ( .A(n6328), .B(n6329), .Z(n6330) );
  NAND U6774 ( .A(x[129]), .B(y[707]), .Z(n6343) );
  AND U6775 ( .A(y[711]), .B(x[133]), .Z(n6458) );
  NANDN U6776 ( .A(n6343), .B(n6458), .Z(n6289) );
  OR U6777 ( .A(n6287), .B(n6286), .Z(n6288) );
  AND U6778 ( .A(n6289), .B(n6288), .Z(n6331) );
  XOR U6779 ( .A(n6330), .B(n6331), .Z(n6333) );
  XNOR U6780 ( .A(n6332), .B(n6333), .Z(n6338) );
  OR U6781 ( .A(n6293), .B(n7106), .Z(n6297) );
  OR U6782 ( .A(n6295), .B(n6294), .Z(n6296) );
  AND U6783 ( .A(n6297), .B(n6296), .Z(n6336) );
  XNOR U6784 ( .A(n6337), .B(n6336), .Z(n6339) );
  XOR U6785 ( .A(n6338), .B(n6339), .Z(n6319) );
  XOR U6786 ( .A(n6318), .B(n6319), .Z(n6313) );
  NANDN U6787 ( .A(n6299), .B(n6298), .Z(n6303) );
  NANDN U6788 ( .A(n6301), .B(n6300), .Z(n6302) );
  NAND U6789 ( .A(n6303), .B(n6302), .Z(n6310) );
  OR U6790 ( .A(n6305), .B(n6304), .Z(n6309) );
  OR U6791 ( .A(n6307), .B(n6306), .Z(n6308) );
  AND U6792 ( .A(n6309), .B(n6308), .Z(n6311) );
  XNOR U6793 ( .A(n6310), .B(n6311), .Z(n6312) );
  XOR U6794 ( .A(n6313), .B(n6312), .Z(N170) );
  NANDN U6795 ( .A(n6311), .B(n6310), .Z(n6315) );
  NANDN U6796 ( .A(n6313), .B(n6312), .Z(n6314) );
  NAND U6797 ( .A(n6315), .B(n6314), .Z(n6357) );
  OR U6798 ( .A(n6317), .B(n6316), .Z(n6321) );
  NANDN U6799 ( .A(n6319), .B(n6318), .Z(n6320) );
  AND U6800 ( .A(n6321), .B(n6320), .Z(n6358) );
  XNOR U6801 ( .A(n6357), .B(n6358), .Z(n6359) );
  NANDN U6802 ( .A(n6323), .B(n6322), .Z(n6327) );
  NANDN U6803 ( .A(n6325), .B(n6324), .Z(n6326) );
  NAND U6804 ( .A(n6327), .B(n6326), .Z(n6417) );
  XOR U6805 ( .A(n6417), .B(n6416), .Z(n6418) );
  NANDN U6806 ( .A(n6331), .B(n6330), .Z(n6335) );
  OR U6807 ( .A(n6333), .B(n6332), .Z(n6334) );
  AND U6808 ( .A(n6335), .B(n6334), .Z(n6419) );
  XNOR U6809 ( .A(n6418), .B(n6419), .Z(n6366) );
  OR U6810 ( .A(n6337), .B(n6336), .Z(n6341) );
  NANDN U6811 ( .A(n6339), .B(n6338), .Z(n6340) );
  AND U6812 ( .A(n6341), .B(n6340), .Z(n6363) );
  ANDN U6813 ( .B(y[714]), .A(n151), .Z(n6402) );
  NANDN U6814 ( .A(n6342), .B(o[73]), .Z(n6399) );
  ANDN U6815 ( .B(y[704]), .A(n161), .Z(n6400) );
  XNOR U6816 ( .A(n6402), .B(n6401), .Z(n6391) );
  ANDN U6817 ( .B(y[713]), .A(n152), .Z(n7302) );
  ANDN U6818 ( .B(y[711]), .A(n154), .Z(n7338) );
  XNOR U6819 ( .A(n7338), .B(n6379), .Z(n6380) );
  XNOR U6820 ( .A(n7302), .B(n6380), .Z(n6389) );
  ANDN U6821 ( .B(y[712]), .A(n157), .Z(n6714) );
  NANDN U6822 ( .A(n6343), .B(n6714), .Z(n6346) );
  NANDN U6823 ( .A(n6780), .B(n6344), .Z(n6345) );
  AND U6824 ( .A(n6346), .B(n6345), .Z(n6388) );
  XOR U6825 ( .A(n6389), .B(n6388), .Z(n6390) );
  XOR U6826 ( .A(n6391), .B(n6390), .Z(n6410) );
  AND U6827 ( .A(y[713]), .B(x[137]), .Z(n6972) );
  NAND U6828 ( .A(n6773), .B(n6972), .Z(n6350) );
  OR U6829 ( .A(n6348), .B(n6347), .Z(n6349) );
  NAND U6830 ( .A(n6350), .B(n6349), .Z(n6411) );
  XNOR U6831 ( .A(n6410), .B(n6411), .Z(n6413) );
  AND U6832 ( .A(y[706]), .B(x[136]), .Z(n6477) );
  XOR U6833 ( .A(n6477), .B(n6520), .Z(n6385) );
  NAND U6834 ( .A(x[137]), .B(y[705]), .Z(n6394) );
  XOR U6835 ( .A(o[74]), .B(n6394), .Z(n6384) );
  XOR U6836 ( .A(n6385), .B(n6384), .Z(n6369) );
  AND U6837 ( .A(y[708]), .B(x[134]), .Z(n6617) );
  AND U6838 ( .A(x[132]), .B(y[710]), .Z(n6352) );
  NAND U6839 ( .A(x[135]), .B(y[707]), .Z(n6351) );
  XOR U6840 ( .A(n6352), .B(n6351), .Z(n6407) );
  XNOR U6841 ( .A(n6617), .B(n6407), .Z(n6370) );
  XNOR U6842 ( .A(n6369), .B(n6370), .Z(n6372) );
  ANDN U6843 ( .B(y[708]), .A(n158), .Z(n6478) );
  NAND U6844 ( .A(n6383), .B(n6478), .Z(n6356) );
  OR U6845 ( .A(n6354), .B(n6353), .Z(n6355) );
  NAND U6846 ( .A(n6356), .B(n6355), .Z(n6371) );
  XNOR U6847 ( .A(n6372), .B(n6371), .Z(n6412) );
  XNOR U6848 ( .A(n6413), .B(n6412), .Z(n6364) );
  XOR U6849 ( .A(n6363), .B(n6364), .Z(n6365) );
  XOR U6850 ( .A(n6366), .B(n6365), .Z(n6360) );
  XOR U6851 ( .A(n6359), .B(n6360), .Z(N171) );
  NANDN U6852 ( .A(n6358), .B(n6357), .Z(n6362) );
  NANDN U6853 ( .A(n6360), .B(n6359), .Z(n6361) );
  NAND U6854 ( .A(n6362), .B(n6361), .Z(n6422) );
  OR U6855 ( .A(n6364), .B(n6363), .Z(n6368) );
  NANDN U6856 ( .A(n6366), .B(n6365), .Z(n6367) );
  AND U6857 ( .A(n6368), .B(n6367), .Z(n6423) );
  XNOR U6858 ( .A(n6422), .B(n6423), .Z(n6424) );
  OR U6859 ( .A(n6370), .B(n6369), .Z(n6374) );
  OR U6860 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U6861 ( .A(n6374), .B(n6373), .Z(n6454) );
  ANDN U6862 ( .B(y[712]), .A(n154), .Z(n7481) );
  AND U6863 ( .A(x[133]), .B(y[710]), .Z(n6376) );
  NAND U6864 ( .A(x[130]), .B(y[713]), .Z(n6375) );
  XOR U6865 ( .A(n6376), .B(n6375), .Z(n6465) );
  NAND U6866 ( .A(x[132]), .B(y[711]), .Z(n6464) );
  XNOR U6867 ( .A(n6465), .B(n6464), .Z(n6440) );
  XNOR U6868 ( .A(n7481), .B(n6440), .Z(n6441) );
  AND U6869 ( .A(x[136]), .B(y[707]), .Z(n6378) );
  NAND U6870 ( .A(x[137]), .B(y[706]), .Z(n6377) );
  XNOR U6871 ( .A(n6378), .B(n6377), .Z(n6479) );
  XNOR U6872 ( .A(n6478), .B(n6479), .Z(n6442) );
  XNOR U6873 ( .A(n6441), .B(n6442), .Z(n6488) );
  NANDN U6874 ( .A(n7338), .B(n6379), .Z(n6382) );
  NANDN U6875 ( .A(n7302), .B(n6380), .Z(n6381) );
  NAND U6876 ( .A(n6382), .B(n6381), .Z(n6485) );
  ANDN U6877 ( .B(y[709]), .A(n159), .Z(n7221) );
  NAND U6878 ( .A(n7221), .B(n6383), .Z(n6387) );
  OR U6879 ( .A(n6385), .B(n6384), .Z(n6386) );
  NAND U6880 ( .A(n6387), .B(n6386), .Z(n6486) );
  XNOR U6881 ( .A(n6488), .B(n6487), .Z(n6452) );
  OR U6882 ( .A(n6389), .B(n6388), .Z(n6393) );
  NAND U6883 ( .A(n6391), .B(n6390), .Z(n6392) );
  NAND U6884 ( .A(n6393), .B(n6392), .Z(n6437) );
  NANDN U6885 ( .A(n6394), .B(o[74]), .Z(n6474) );
  AND U6886 ( .A(y[704]), .B(x[139]), .Z(n6396) );
  NAND U6887 ( .A(x[128]), .B(y[715]), .Z(n6395) );
  XNOR U6888 ( .A(n6396), .B(n6395), .Z(n6473) );
  AND U6889 ( .A(y[709]), .B(x[134]), .Z(n6398) );
  NAND U6890 ( .A(x[129]), .B(y[714]), .Z(n6397) );
  XOR U6891 ( .A(n6398), .B(n6397), .Z(n6470) );
  NAND U6892 ( .A(x[138]), .B(y[705]), .Z(n6482) );
  XOR U6893 ( .A(o[75]), .B(n6482), .Z(n6469) );
  XOR U6894 ( .A(n6470), .B(n6469), .Z(n6445) );
  NANDN U6895 ( .A(n6400), .B(n6399), .Z(n6404) );
  OR U6896 ( .A(n6402), .B(n6401), .Z(n6403) );
  NAND U6897 ( .A(n6404), .B(n6403), .Z(n6448) );
  XOR U6898 ( .A(n6447), .B(n6448), .Z(n6434) );
  AND U6899 ( .A(y[710]), .B(x[135]), .Z(n6406) );
  NAND U6900 ( .A(n6406), .B(n6405), .Z(n6409) );
  NANDN U6901 ( .A(n6407), .B(n6617), .Z(n6408) );
  NAND U6902 ( .A(n6409), .B(n6408), .Z(n6435) );
  XOR U6903 ( .A(n6437), .B(n6436), .Z(n6451) );
  XOR U6904 ( .A(n6452), .B(n6451), .Z(n6453) );
  XOR U6905 ( .A(n6454), .B(n6453), .Z(n6428) );
  OR U6906 ( .A(n6411), .B(n6410), .Z(n6415) );
  OR U6907 ( .A(n6413), .B(n6412), .Z(n6414) );
  AND U6908 ( .A(n6415), .B(n6414), .Z(n6429) );
  XNOR U6909 ( .A(n6428), .B(n6429), .Z(n6431) );
  OR U6910 ( .A(n6417), .B(n6416), .Z(n6421) );
  NANDN U6911 ( .A(n6419), .B(n6418), .Z(n6420) );
  NAND U6912 ( .A(n6421), .B(n6420), .Z(n6430) );
  XOR U6913 ( .A(n6431), .B(n6430), .Z(n6425) );
  XNOR U6914 ( .A(n6424), .B(n6425), .Z(N172) );
  NANDN U6915 ( .A(n6423), .B(n6422), .Z(n6427) );
  NAND U6916 ( .A(n6425), .B(n6424), .Z(n6426) );
  NAND U6917 ( .A(n6427), .B(n6426), .Z(n6491) );
  OR U6918 ( .A(n6429), .B(n6428), .Z(n6433) );
  OR U6919 ( .A(n6431), .B(n6430), .Z(n6432) );
  AND U6920 ( .A(n6433), .B(n6432), .Z(n6492) );
  XNOR U6921 ( .A(n6491), .B(n6492), .Z(n6493) );
  NANDN U6922 ( .A(n6435), .B(n6434), .Z(n6439) );
  NANDN U6923 ( .A(n6437), .B(n6436), .Z(n6438) );
  NAND U6924 ( .A(n6439), .B(n6438), .Z(n6566) );
  NANDN U6925 ( .A(n6440), .B(n7481), .Z(n6444) );
  NANDN U6926 ( .A(n6442), .B(n6441), .Z(n6443) );
  NAND U6927 ( .A(n6444), .B(n6443), .Z(n6563) );
  NAND U6928 ( .A(n6446), .B(n6445), .Z(n6450) );
  NANDN U6929 ( .A(n6448), .B(n6447), .Z(n6449) );
  AND U6930 ( .A(n6450), .B(n6449), .Z(n6564) );
  XNOR U6931 ( .A(n6566), .B(n6565), .Z(n6497) );
  NANDN U6932 ( .A(n6452), .B(n6451), .Z(n6456) );
  OR U6933 ( .A(n6454), .B(n6453), .Z(n6455) );
  NAND U6934 ( .A(n6456), .B(n6455), .Z(n6498) );
  XNOR U6935 ( .A(n6497), .B(n6498), .Z(n6500) );
  NAND U6936 ( .A(x[135]), .B(y[709]), .Z(n6457) );
  XOR U6937 ( .A(n6458), .B(n6457), .Z(n6522) );
  AND U6938 ( .A(y[706]), .B(x[138]), .Z(n6459) );
  NAND U6939 ( .A(x[137]), .B(y[707]), .Z(n7170) );
  XOR U6940 ( .A(n6459), .B(n7170), .Z(n6550) );
  NAND U6941 ( .A(x[132]), .B(y[712]), .Z(n6549) );
  XNOR U6942 ( .A(n6550), .B(n6549), .Z(n6521) );
  XOR U6943 ( .A(n6522), .B(n6521), .Z(n6527) );
  AND U6944 ( .A(y[704]), .B(x[140]), .Z(n6461) );
  NAND U6945 ( .A(x[128]), .B(y[716]), .Z(n6460) );
  XOR U6946 ( .A(n6461), .B(n6460), .Z(n6542) );
  NAND U6947 ( .A(x[139]), .B(y[705]), .Z(n6516) );
  XOR U6948 ( .A(o[76]), .B(n6516), .Z(n6541) );
  XOR U6949 ( .A(n6542), .B(n6541), .Z(n6525) );
  AND U6950 ( .A(y[708]), .B(x[136]), .Z(n6463) );
  NAND U6951 ( .A(x[130]), .B(y[714]), .Z(n6462) );
  XOR U6952 ( .A(n6463), .B(n6462), .Z(n6511) );
  NAND U6953 ( .A(y[713]), .B(x[131]), .Z(n6510) );
  XNOR U6954 ( .A(n6511), .B(n6510), .Z(n6526) );
  XOR U6955 ( .A(n6525), .B(n6526), .Z(n6528) );
  XOR U6956 ( .A(n6527), .B(n6528), .Z(n6505) );
  ANDN U6957 ( .B(y[713]), .A(n156), .Z(n6671) );
  NAND U6958 ( .A(n6789), .B(n6671), .Z(n6467) );
  OR U6959 ( .A(n6465), .B(n6464), .Z(n6466) );
  NAND U6960 ( .A(n6467), .B(n6466), .Z(n6504) );
  AND U6961 ( .A(y[714]), .B(x[134]), .Z(n6779) );
  NAND U6962 ( .A(n6779), .B(n6468), .Z(n6472) );
  OR U6963 ( .A(n6470), .B(n6469), .Z(n6471) );
  NAND U6964 ( .A(n6472), .B(n6471), .Z(n6503) );
  XNOR U6965 ( .A(n6504), .B(n6503), .Z(n6506) );
  XNOR U6966 ( .A(n6505), .B(n6506), .Z(n6558) );
  AND U6967 ( .A(y[715]), .B(x[139]), .Z(n7603) );
  NAND U6968 ( .A(n6773), .B(n7603), .Z(n6476) );
  NANDN U6969 ( .A(n6474), .B(n6473), .Z(n6475) );
  NAND U6970 ( .A(n6476), .B(n6475), .Z(n6533) );
  NANDN U6971 ( .A(n7170), .B(n6477), .Z(n6481) );
  NAND U6972 ( .A(n6479), .B(n6478), .Z(n6480) );
  NAND U6973 ( .A(n6481), .B(n6480), .Z(n6532) );
  NANDN U6974 ( .A(n6482), .B(o[75]), .Z(n6538) );
  NAND U6975 ( .A(x[129]), .B(y[715]), .Z(n6483) );
  XNOR U6976 ( .A(n6484), .B(n6483), .Z(n6537) );
  XNOR U6977 ( .A(n6532), .B(n6531), .Z(n6534) );
  XOR U6978 ( .A(n6558), .B(n6557), .Z(n6560) );
  NANDN U6979 ( .A(n6486), .B(n6485), .Z(n6490) );
  NANDN U6980 ( .A(n6488), .B(n6487), .Z(n6489) );
  AND U6981 ( .A(n6490), .B(n6489), .Z(n6559) );
  XNOR U6982 ( .A(n6560), .B(n6559), .Z(n6499) );
  XNOR U6983 ( .A(n6500), .B(n6499), .Z(n6494) );
  XOR U6984 ( .A(n6493), .B(n6494), .Z(N173) );
  NANDN U6985 ( .A(n6492), .B(n6491), .Z(n6496) );
  NANDN U6986 ( .A(n6494), .B(n6493), .Z(n6495) );
  NAND U6987 ( .A(n6496), .B(n6495), .Z(n6634) );
  OR U6988 ( .A(n6498), .B(n6497), .Z(n6502) );
  OR U6989 ( .A(n6500), .B(n6499), .Z(n6501) );
  AND U6990 ( .A(n6502), .B(n6501), .Z(n6635) );
  XNOR U6991 ( .A(n6634), .B(n6635), .Z(n6636) );
  OR U6992 ( .A(n6504), .B(n6503), .Z(n6508) );
  NANDN U6993 ( .A(n6506), .B(n6505), .Z(n6507) );
  AND U6994 ( .A(n6508), .B(n6507), .Z(n6575) );
  AND U6995 ( .A(y[714]), .B(x[136]), .Z(n6980) );
  NAND U6996 ( .A(n6980), .B(n6509), .Z(n6513) );
  OR U6997 ( .A(n6511), .B(n6510), .Z(n6512) );
  NAND U6998 ( .A(n6513), .B(n6512), .Z(n6596) );
  AND U6999 ( .A(y[711]), .B(x[134]), .Z(n6515) );
  NAND U7000 ( .A(x[137]), .B(y[708]), .Z(n6514) );
  XOR U7001 ( .A(n6515), .B(n6514), .Z(n6619) );
  NAND U7002 ( .A(x[130]), .B(y[715]), .Z(n6618) );
  XOR U7003 ( .A(n6619), .B(n6618), .Z(n6594) );
  NANDN U7004 ( .A(n6516), .B(o[76]), .Z(n6605) );
  AND U7005 ( .A(y[716]), .B(x[129]), .Z(n6518) );
  NAND U7006 ( .A(x[135]), .B(y[710]), .Z(n6517) );
  XNOR U7007 ( .A(n6518), .B(n6517), .Z(n6604) );
  XNOR U7008 ( .A(n6596), .B(n6595), .Z(n6570) );
  AND U7009 ( .A(y[711]), .B(x[135]), .Z(n6519) );
  NANDN U7010 ( .A(n6520), .B(n6519), .Z(n6524) );
  OR U7011 ( .A(n6522), .B(n6521), .Z(n6523) );
  AND U7012 ( .A(n6524), .B(n6523), .Z(n6569) );
  XOR U7013 ( .A(n6570), .B(n6569), .Z(n6571) );
  NANDN U7014 ( .A(n6526), .B(n6525), .Z(n6530) );
  NANDN U7015 ( .A(n6528), .B(n6527), .Z(n6529) );
  AND U7016 ( .A(n6530), .B(n6529), .Z(n6572) );
  XNOR U7017 ( .A(n6571), .B(n6572), .Z(n6576) );
  XOR U7018 ( .A(n6575), .B(n6576), .Z(n6577) );
  NAND U7019 ( .A(n6532), .B(n6531), .Z(n6536) );
  NANDN U7020 ( .A(n6534), .B(n6533), .Z(n6535) );
  NAND U7021 ( .A(n6536), .B(n6535), .Z(n6584) );
  ANDN U7022 ( .B(y[715]), .A(n157), .Z(n7002) );
  NAND U7023 ( .A(n7002), .B(n6602), .Z(n6540) );
  NANDN U7024 ( .A(n6538), .B(n6537), .Z(n6539) );
  NAND U7025 ( .A(n6540), .B(n6539), .Z(n6589) );
  ANDN U7026 ( .B(y[716]), .A(n163), .Z(n7814) );
  NAND U7027 ( .A(n6773), .B(n7814), .Z(n6544) );
  OR U7028 ( .A(n6542), .B(n6541), .Z(n6543) );
  NAND U7029 ( .A(n6544), .B(n6543), .Z(n6587) );
  AND U7030 ( .A(y[706]), .B(x[139]), .Z(n6546) );
  NAND U7031 ( .A(x[138]), .B(y[707]), .Z(n6545) );
  XNOR U7032 ( .A(n6546), .B(n6545), .Z(n6608) );
  XNOR U7033 ( .A(n7221), .B(n6608), .Z(n6588) );
  XOR U7034 ( .A(n6589), .B(n6590), .Z(n6581) );
  AND U7035 ( .A(y[706]), .B(x[137]), .Z(n6548) );
  AND U7036 ( .A(y[707]), .B(x[138]), .Z(n6547) );
  NAND U7037 ( .A(n6548), .B(n6547), .Z(n6552) );
  OR U7038 ( .A(n6550), .B(n6549), .Z(n6551) );
  NAND U7039 ( .A(n6552), .B(n6551), .Z(n6614) );
  AND U7040 ( .A(y[704]), .B(x[141]), .Z(n6554) );
  NAND U7041 ( .A(x[128]), .B(y[717]), .Z(n6553) );
  XOR U7042 ( .A(n6554), .B(n6553), .Z(n6631) );
  NAND U7043 ( .A(x[140]), .B(y[705]), .Z(n6623) );
  XOR U7044 ( .A(o[77]), .B(n6623), .Z(n6630) );
  XOR U7045 ( .A(n6631), .B(n6630), .Z(n6612) );
  AND U7046 ( .A(x[131]), .B(y[714]), .Z(n6556) );
  NAND U7047 ( .A(x[133]), .B(y[712]), .Z(n6555) );
  XOR U7048 ( .A(n6556), .B(n6555), .Z(n6627) );
  NAND U7049 ( .A(y[713]), .B(x[132]), .Z(n6626) );
  XOR U7050 ( .A(n6627), .B(n6626), .Z(n6611) );
  XOR U7051 ( .A(n6614), .B(n6613), .Z(n6582) );
  XNOR U7052 ( .A(n6581), .B(n6582), .Z(n6583) );
  XOR U7053 ( .A(n6584), .B(n6583), .Z(n6578) );
  XNOR U7054 ( .A(n6577), .B(n6578), .Z(n6643) );
  NANDN U7055 ( .A(n6558), .B(n6557), .Z(n6562) );
  NANDN U7056 ( .A(n6560), .B(n6559), .Z(n6561) );
  NAND U7057 ( .A(n6562), .B(n6561), .Z(n6640) );
  NANDN U7058 ( .A(n6564), .B(n6563), .Z(n6568) );
  NANDN U7059 ( .A(n6566), .B(n6565), .Z(n6567) );
  AND U7060 ( .A(n6568), .B(n6567), .Z(n6641) );
  XNOR U7061 ( .A(n6643), .B(n6642), .Z(n6637) );
  XOR U7062 ( .A(n6636), .B(n6637), .Z(N174) );
  OR U7063 ( .A(n6570), .B(n6569), .Z(n6574) );
  NANDN U7064 ( .A(n6572), .B(n6571), .Z(n6573) );
  NAND U7065 ( .A(n6574), .B(n6573), .Z(n6655) );
  OR U7066 ( .A(n6576), .B(n6575), .Z(n6580) );
  NANDN U7067 ( .A(n6578), .B(n6577), .Z(n6579) );
  AND U7068 ( .A(n6580), .B(n6579), .Z(n6652) );
  NANDN U7069 ( .A(n6582), .B(n6581), .Z(n6586) );
  NANDN U7070 ( .A(n6584), .B(n6583), .Z(n6585) );
  NAND U7071 ( .A(n6586), .B(n6585), .Z(n6660) );
  NANDN U7072 ( .A(n6588), .B(n6587), .Z(n6592) );
  NANDN U7073 ( .A(n6590), .B(n6589), .Z(n6591) );
  NAND U7074 ( .A(n6592), .B(n6591), .Z(n6666) );
  NAND U7075 ( .A(n6594), .B(n6593), .Z(n6598) );
  NAND U7076 ( .A(n6596), .B(n6595), .Z(n6597) );
  NAND U7077 ( .A(n6598), .B(n6597), .Z(n6664) );
  ANDN U7078 ( .B(y[714]), .A(n155), .Z(n6686) );
  AND U7079 ( .A(y[708]), .B(x[138]), .Z(n7343) );
  AND U7080 ( .A(y[709]), .B(x[137]), .Z(n7307) );
  NAND U7081 ( .A(x[130]), .B(y[716]), .Z(n6599) );
  XOR U7082 ( .A(n7307), .B(n6599), .Z(n6698) );
  XNOR U7083 ( .A(n7343), .B(n6698), .Z(n6685) );
  XOR U7084 ( .A(n6686), .B(n6685), .Z(n6688) );
  AND U7085 ( .A(y[715]), .B(x[131]), .Z(n6601) );
  NAND U7086 ( .A(x[136]), .B(y[710]), .Z(n6600) );
  XOR U7087 ( .A(n6601), .B(n6600), .Z(n6672) );
  XOR U7088 ( .A(n6671), .B(n6672), .Z(n6687) );
  AND U7089 ( .A(y[716]), .B(x[135]), .Z(n6603) );
  NAND U7090 ( .A(n6603), .B(n6602), .Z(n6607) );
  NANDN U7091 ( .A(n6605), .B(n6604), .Z(n6606) );
  NAND U7092 ( .A(n6607), .B(n6606), .Z(n6691) );
  NAND U7093 ( .A(x[138]), .B(y[706]), .Z(n7226) );
  NOR U7094 ( .A(n162), .B(n147), .Z(n6810) );
  NANDN U7095 ( .A(n7226), .B(n6810), .Z(n6610) );
  NAND U7096 ( .A(n6608), .B(n7221), .Z(n6609) );
  AND U7097 ( .A(n6610), .B(n6609), .Z(n6692) );
  XOR U7098 ( .A(n6694), .B(n6693), .Z(n6665) );
  XOR U7099 ( .A(n6666), .B(n6667), .Z(n6658) );
  NAND U7100 ( .A(n6612), .B(n6611), .Z(n6616) );
  NAND U7101 ( .A(n6614), .B(n6613), .Z(n6615) );
  NAND U7102 ( .A(n6616), .B(n6615), .Z(n6732) );
  AND U7103 ( .A(y[711]), .B(x[137]), .Z(n6807) );
  NAND U7104 ( .A(n6807), .B(n6617), .Z(n6621) );
  OR U7105 ( .A(n6619), .B(n6618), .Z(n6620) );
  AND U7106 ( .A(n6621), .B(n6620), .Z(n6720) );
  AND U7107 ( .A(y[706]), .B(x[140]), .Z(n7297) );
  NAND U7108 ( .A(x[135]), .B(y[711]), .Z(n6622) );
  XOR U7109 ( .A(n7297), .B(n6622), .Z(n6703) );
  NAND U7110 ( .A(x[141]), .B(y[705]), .Z(n6706) );
  XOR U7111 ( .A(o[78]), .B(n6706), .Z(n6702) );
  XOR U7112 ( .A(n6703), .B(n6702), .Z(n6718) );
  NANDN U7113 ( .A(n6623), .B(o[77]), .Z(n6676) );
  AND U7114 ( .A(x[128]), .B(y[718]), .Z(n6625) );
  NAND U7115 ( .A(x[142]), .B(y[704]), .Z(n6624) );
  XNOR U7116 ( .A(n6625), .B(n6624), .Z(n6675) );
  XOR U7117 ( .A(n6720), .B(n6719), .Z(n6729) );
  ANDN U7118 ( .B(y[714]), .A(n156), .Z(n6765) );
  NAND U7119 ( .A(n7481), .B(n6765), .Z(n6629) );
  OR U7120 ( .A(n6627), .B(n6626), .Z(n6628) );
  NAND U7121 ( .A(n6629), .B(n6628), .Z(n6726) );
  IV U7122 ( .A(n6810), .Z(n6712) );
  XNOR U7123 ( .A(n6712), .B(n6711), .Z(n6713) );
  XOR U7124 ( .A(n6714), .B(n6713), .Z(n6724) );
  AND U7125 ( .A(x[141]), .B(y[717]), .Z(n8209) );
  NAND U7126 ( .A(n6773), .B(n8209), .Z(n6633) );
  OR U7127 ( .A(n6631), .B(n6630), .Z(n6632) );
  AND U7128 ( .A(n6633), .B(n6632), .Z(n6723) );
  XOR U7129 ( .A(n6724), .B(n6723), .Z(n6725) );
  XOR U7130 ( .A(n6726), .B(n6725), .Z(n6730) );
  XNOR U7131 ( .A(n6729), .B(n6730), .Z(n6731) );
  XOR U7132 ( .A(n6732), .B(n6731), .Z(n6659) );
  XOR U7133 ( .A(n6658), .B(n6659), .Z(n6661) );
  XOR U7134 ( .A(n6660), .B(n6661), .Z(n6653) );
  XNOR U7135 ( .A(n6652), .B(n6653), .Z(n6654) );
  XNOR U7136 ( .A(n6655), .B(n6654), .Z(n6649) );
  NANDN U7137 ( .A(n6635), .B(n6634), .Z(n6639) );
  NANDN U7138 ( .A(n6637), .B(n6636), .Z(n6638) );
  NAND U7139 ( .A(n6639), .B(n6638), .Z(n6646) );
  NANDN U7140 ( .A(n6641), .B(n6640), .Z(n6645) );
  NANDN U7141 ( .A(n6643), .B(n6642), .Z(n6644) );
  NAND U7142 ( .A(n6645), .B(n6644), .Z(n6647) );
  XNOR U7143 ( .A(n6646), .B(n6647), .Z(n6648) );
  XOR U7144 ( .A(n6649), .B(n6648), .Z(N175) );
  NANDN U7145 ( .A(n6647), .B(n6646), .Z(n6651) );
  NANDN U7146 ( .A(n6649), .B(n6648), .Z(n6650) );
  NAND U7147 ( .A(n6651), .B(n6650), .Z(n6735) );
  OR U7148 ( .A(n6653), .B(n6652), .Z(n6657) );
  OR U7149 ( .A(n6655), .B(n6654), .Z(n6656) );
  AND U7150 ( .A(n6657), .B(n6656), .Z(n6736) );
  XNOR U7151 ( .A(n6735), .B(n6736), .Z(n6737) );
  NANDN U7152 ( .A(n6659), .B(n6658), .Z(n6663) );
  NANDN U7153 ( .A(n6661), .B(n6660), .Z(n6662) );
  NAND U7154 ( .A(n6663), .B(n6662), .Z(n6744) );
  NANDN U7155 ( .A(n6665), .B(n6664), .Z(n6669) );
  NANDN U7156 ( .A(n6667), .B(n6666), .Z(n6668) );
  NAND U7157 ( .A(n6669), .B(n6668), .Z(n6824) );
  NAND U7158 ( .A(x[136]), .B(y[715]), .Z(n7094) );
  NANDN U7159 ( .A(n7094), .B(n6670), .Z(n6674) );
  NANDN U7160 ( .A(n6672), .B(n6671), .Z(n6673) );
  NAND U7161 ( .A(n6674), .B(n6673), .Z(n6795) );
  AND U7162 ( .A(x[142]), .B(y[718]), .Z(n8399) );
  NAND U7163 ( .A(n6773), .B(n8399), .Z(n6678) );
  NANDN U7164 ( .A(n6676), .B(n6675), .Z(n6677) );
  AND U7165 ( .A(n6678), .B(n6677), .Z(n6794) );
  ANDN U7166 ( .B(y[712]), .A(n158), .Z(n7185) );
  AND U7167 ( .A(y[709]), .B(x[138]), .Z(n6680) );
  NAND U7168 ( .A(x[132]), .B(y[715]), .Z(n6679) );
  XOR U7169 ( .A(n6680), .B(n6679), .Z(n6781) );
  XNOR U7170 ( .A(n7185), .B(n6781), .Z(n6767) );
  IV U7171 ( .A(y[713]), .Z(n7055) );
  NOR U7172 ( .A(n157), .B(n7055), .Z(n6902) );
  XOR U7173 ( .A(n6765), .B(n6902), .Z(n6766) );
  XOR U7174 ( .A(n6767), .B(n6766), .Z(n6803) );
  AND U7175 ( .A(y[705]), .B(x[142]), .Z(n6784) );
  XNOR U7176 ( .A(o[79]), .B(n6784), .Z(n6770) );
  AND U7177 ( .A(y[711]), .B(x[136]), .Z(n6682) );
  NAND U7178 ( .A(x[129]), .B(y[718]), .Z(n6681) );
  XNOR U7179 ( .A(n6682), .B(n6681), .Z(n6769) );
  XNOR U7180 ( .A(n6770), .B(n6769), .Z(n6801) );
  NAND U7181 ( .A(x[131]), .B(y[716]), .Z(n6791) );
  AND U7182 ( .A(x[137]), .B(y[710]), .Z(n6684) );
  NAND U7183 ( .A(x[130]), .B(y[717]), .Z(n6683) );
  XOR U7184 ( .A(n6684), .B(n6683), .Z(n6790) );
  XNOR U7185 ( .A(n6791), .B(n6790), .Z(n6800) );
  XOR U7186 ( .A(n6801), .B(n6800), .Z(n6802) );
  XNOR U7187 ( .A(n6803), .B(n6802), .Z(n6797) );
  XNOR U7188 ( .A(n6796), .B(n6797), .Z(n6759) );
  OR U7189 ( .A(n6686), .B(n6685), .Z(n6690) );
  NAND U7190 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U7191 ( .A(n6690), .B(n6689), .Z(n6760) );
  XNOR U7192 ( .A(n6759), .B(n6760), .Z(n6762) );
  NANDN U7193 ( .A(n6692), .B(n6691), .Z(n6696) );
  NANDN U7194 ( .A(n6694), .B(n6693), .Z(n6695) );
  AND U7195 ( .A(n6696), .B(n6695), .Z(n6761) );
  XOR U7196 ( .A(n6762), .B(n6761), .Z(n6822) );
  ANDN U7197 ( .B(y[716]), .A(n160), .Z(n7438) );
  NAND U7198 ( .A(n6697), .B(n7438), .Z(n6700) );
  NANDN U7199 ( .A(n6698), .B(n7343), .Z(n6699) );
  AND U7200 ( .A(n6700), .B(n6699), .Z(n6753) );
  AND U7201 ( .A(y[711]), .B(x[140]), .Z(n7062) );
  NAND U7202 ( .A(n6701), .B(n7062), .Z(n6705) );
  OR U7203 ( .A(n6703), .B(n6702), .Z(n6704) );
  NAND U7204 ( .A(n6705), .B(n6704), .Z(n6818) );
  NANDN U7205 ( .A(n6706), .B(o[78]), .Z(n6775) );
  AND U7206 ( .A(y[704]), .B(x[143]), .Z(n6708) );
  NAND U7207 ( .A(x[128]), .B(y[719]), .Z(n6707) );
  XOR U7208 ( .A(n6708), .B(n6707), .Z(n6774) );
  XNOR U7209 ( .A(n6775), .B(n6774), .Z(n6815) );
  NAND U7210 ( .A(x[141]), .B(y[706]), .Z(n6812) );
  AND U7211 ( .A(x[140]), .B(y[707]), .Z(n6710) );
  NAND U7212 ( .A(x[139]), .B(y[708]), .Z(n6709) );
  XOR U7213 ( .A(n6710), .B(n6709), .Z(n6811) );
  XOR U7214 ( .A(n6812), .B(n6811), .Z(n6816) );
  XNOR U7215 ( .A(n6818), .B(n6817), .Z(n6754) );
  XOR U7216 ( .A(n6753), .B(n6754), .Z(n6755) );
  NAND U7217 ( .A(n6712), .B(n6711), .Z(n6716) );
  OR U7218 ( .A(n6714), .B(n6713), .Z(n6715) );
  NAND U7219 ( .A(n6716), .B(n6715), .Z(n6756) );
  NAND U7220 ( .A(n6718), .B(n6717), .Z(n6722) );
  NANDN U7221 ( .A(n6720), .B(n6719), .Z(n6721) );
  AND U7222 ( .A(n6722), .B(n6721), .Z(n6747) );
  XNOR U7223 ( .A(n6748), .B(n6747), .Z(n6750) );
  OR U7224 ( .A(n6724), .B(n6723), .Z(n6728) );
  NAND U7225 ( .A(n6726), .B(n6725), .Z(n6727) );
  AND U7226 ( .A(n6728), .B(n6727), .Z(n6749) );
  XOR U7227 ( .A(n6750), .B(n6749), .Z(n6821) );
  XNOR U7228 ( .A(n6824), .B(n6823), .Z(n6742) );
  NANDN U7229 ( .A(n6730), .B(n6729), .Z(n6734) );
  NANDN U7230 ( .A(n6732), .B(n6731), .Z(n6733) );
  AND U7231 ( .A(n6734), .B(n6733), .Z(n6741) );
  XNOR U7232 ( .A(n6744), .B(n6743), .Z(n6738) );
  XOR U7233 ( .A(n6737), .B(n6738), .Z(N176) );
  NANDN U7234 ( .A(n6736), .B(n6735), .Z(n6740) );
  NANDN U7235 ( .A(n6738), .B(n6737), .Z(n6739) );
  NAND U7236 ( .A(n6740), .B(n6739), .Z(n6827) );
  NANDN U7237 ( .A(n6742), .B(n6741), .Z(n6746) );
  NANDN U7238 ( .A(n6744), .B(n6743), .Z(n6745) );
  NAND U7239 ( .A(n6746), .B(n6745), .Z(n6828) );
  XNOR U7240 ( .A(n6827), .B(n6828), .Z(n6829) );
  OR U7241 ( .A(n6748), .B(n6747), .Z(n6752) );
  OR U7242 ( .A(n6750), .B(n6749), .Z(n6751) );
  NAND U7243 ( .A(n6752), .B(n6751), .Z(n6917) );
  OR U7244 ( .A(n6754), .B(n6753), .Z(n6758) );
  NANDN U7245 ( .A(n6756), .B(n6755), .Z(n6757) );
  NAND U7246 ( .A(n6758), .B(n6757), .Z(n6915) );
  OR U7247 ( .A(n6760), .B(n6759), .Z(n6764) );
  OR U7248 ( .A(n6762), .B(n6761), .Z(n6763) );
  NAND U7249 ( .A(n6764), .B(n6763), .Z(n6914) );
  XOR U7250 ( .A(n6915), .B(n6914), .Z(n6916) );
  XNOR U7251 ( .A(n6917), .B(n6916), .Z(n6836) );
  AND U7252 ( .A(y[718]), .B(x[136]), .Z(n7467) );
  NAND U7253 ( .A(n6768), .B(n7467), .Z(n6772) );
  NANDN U7254 ( .A(n6770), .B(n6769), .Z(n6771) );
  AND U7255 ( .A(n6772), .B(n6771), .Z(n6854) );
  AND U7256 ( .A(y[719]), .B(x[143]), .Z(n8949) );
  NAND U7257 ( .A(n6773), .B(n8949), .Z(n6777) );
  OR U7258 ( .A(n6775), .B(n6774), .Z(n6776) );
  AND U7259 ( .A(n6777), .B(n6776), .Z(n6855) );
  XOR U7260 ( .A(n6854), .B(n6855), .Z(n6857) );
  NAND U7261 ( .A(x[144]), .B(y[704]), .Z(n6893) );
  AND U7262 ( .A(y[720]), .B(x[128]), .Z(n6892) );
  XNOR U7263 ( .A(n6893), .B(n6892), .Z(n6895) );
  NAND U7264 ( .A(x[143]), .B(y[705]), .Z(n6911) );
  XNOR U7265 ( .A(n6911), .B(o[80]), .Z(n6894) );
  XNOR U7266 ( .A(n6895), .B(n6894), .Z(n6885) );
  NAND U7267 ( .A(x[138]), .B(y[710]), .Z(n6904) );
  NAND U7268 ( .A(x[135]), .B(y[713]), .Z(n6778) );
  XOR U7269 ( .A(n6779), .B(n6778), .Z(n6903) );
  XNOR U7270 ( .A(n6904), .B(n6903), .Z(n6884) );
  XNOR U7271 ( .A(n6885), .B(n6884), .Z(n6887) );
  ANDN U7272 ( .B(y[715]), .A(n161), .Z(n7477) );
  NANDN U7273 ( .A(n6780), .B(n7477), .Z(n6783) );
  NANDN U7274 ( .A(n6781), .B(n7185), .Z(n6782) );
  AND U7275 ( .A(n6783), .B(n6782), .Z(n6886) );
  XOR U7276 ( .A(n6887), .B(n6886), .Z(n6856) );
  XOR U7277 ( .A(n6857), .B(n6856), .Z(n6873) );
  XOR U7278 ( .A(n6872), .B(n6873), .Z(n6874) );
  NAND U7279 ( .A(o[79]), .B(n6784), .Z(n6899) );
  AND U7280 ( .A(x[129]), .B(y[719]), .Z(n6785) );
  XNOR U7281 ( .A(n6786), .B(n6785), .Z(n6898) );
  XNOR U7282 ( .A(n6899), .B(n6898), .Z(n6880) );
  NAND U7283 ( .A(x[132]), .B(y[716]), .Z(n6845) );
  AND U7284 ( .A(y[709]), .B(x[139]), .Z(n6788) );
  AND U7285 ( .A(y[706]), .B(x[142]), .Z(n6787) );
  XNOR U7286 ( .A(n6788), .B(n6787), .Z(n6844) );
  XOR U7287 ( .A(n6845), .B(n6844), .Z(n6879) );
  AND U7288 ( .A(y[717]), .B(x[137]), .Z(n7561) );
  NAND U7289 ( .A(n6789), .B(n7561), .Z(n6793) );
  OR U7290 ( .A(n6791), .B(n6790), .Z(n6792) );
  NAND U7291 ( .A(n6793), .B(n6792), .Z(n6878) );
  XNOR U7292 ( .A(n6879), .B(n6878), .Z(n6881) );
  XOR U7293 ( .A(n6880), .B(n6881), .Z(n6875) );
  XOR U7294 ( .A(n6874), .B(n6875), .Z(n6867) );
  NANDN U7295 ( .A(n6795), .B(n6794), .Z(n6799) );
  NANDN U7296 ( .A(n6797), .B(n6796), .Z(n6798) );
  AND U7297 ( .A(n6799), .B(n6798), .Z(n6866) );
  XOR U7298 ( .A(n6867), .B(n6866), .Z(n6868) );
  NANDN U7299 ( .A(n6801), .B(n6800), .Z(n6805) );
  OR U7300 ( .A(n6803), .B(n6802), .Z(n6804) );
  AND U7301 ( .A(n6805), .B(n6804), .Z(n6860) );
  NAND U7302 ( .A(x[131]), .B(y[717]), .Z(n6840) );
  AND U7303 ( .A(x[130]), .B(y[718]), .Z(n6806) );
  XNOR U7304 ( .A(n6807), .B(n6806), .Z(n6839) );
  XOR U7305 ( .A(n6840), .B(n6839), .Z(n6849) );
  AND U7306 ( .A(y[708]), .B(x[140]), .Z(n7565) );
  AND U7307 ( .A(x[141]), .B(y[707]), .Z(n6809) );
  NAND U7308 ( .A(x[133]), .B(y[715]), .Z(n6808) );
  XOR U7309 ( .A(n6809), .B(n6808), .Z(n6908) );
  XNOR U7310 ( .A(n7565), .B(n6908), .Z(n6848) );
  XNOR U7311 ( .A(n6849), .B(n6848), .Z(n6851) );
  NAND U7312 ( .A(n6810), .B(n7565), .Z(n6814) );
  OR U7313 ( .A(n6812), .B(n6811), .Z(n6813) );
  AND U7314 ( .A(n6814), .B(n6813), .Z(n6850) );
  XOR U7315 ( .A(n6851), .B(n6850), .Z(n6861) );
  XOR U7316 ( .A(n6860), .B(n6861), .Z(n6862) );
  NANDN U7317 ( .A(n6816), .B(n6815), .Z(n6820) );
  NANDN U7318 ( .A(n6818), .B(n6817), .Z(n6819) );
  AND U7319 ( .A(n6820), .B(n6819), .Z(n6863) );
  XNOR U7320 ( .A(n6868), .B(n6869), .Z(n6834) );
  NAND U7321 ( .A(n6822), .B(n6821), .Z(n6826) );
  NAND U7322 ( .A(n6824), .B(n6823), .Z(n6825) );
  AND U7323 ( .A(n6826), .B(n6825), .Z(n6833) );
  XOR U7324 ( .A(n6834), .B(n6833), .Z(n6835) );
  XNOR U7325 ( .A(n6836), .B(n6835), .Z(n6830) );
  XOR U7326 ( .A(n6829), .B(n6830), .Z(N177) );
  NANDN U7327 ( .A(n6828), .B(n6827), .Z(n6832) );
  NANDN U7328 ( .A(n6830), .B(n6829), .Z(n6831) );
  NAND U7329 ( .A(n6832), .B(n6831), .Z(n6920) );
  OR U7330 ( .A(n6834), .B(n6833), .Z(n6838) );
  NANDN U7331 ( .A(n6836), .B(n6835), .Z(n6837) );
  NAND U7332 ( .A(n6838), .B(n6837), .Z(n6921) );
  XNOR U7333 ( .A(n6920), .B(n6921), .Z(n6922) );
  AND U7334 ( .A(y[714]), .B(x[135]), .Z(n7093) );
  ANDN U7335 ( .B(y[713]), .A(n159), .Z(n7003) );
  XNOR U7336 ( .A(n7002), .B(n7003), .Z(n7005) );
  ANDN U7337 ( .B(y[716]), .A(n156), .Z(n7004) );
  XOR U7338 ( .A(n7005), .B(n7004), .Z(n6990) );
  ANDN U7339 ( .B(y[717]), .A(n155), .Z(n6964) );
  ANDN U7340 ( .B(y[710]), .A(n162), .Z(n6962) );
  ANDN U7341 ( .B(y[708]), .A(n164), .Z(n6963) );
  XNOR U7342 ( .A(n6962), .B(n6963), .Z(n6965) );
  XNOR U7343 ( .A(n6964), .B(n6965), .Z(n6989) );
  XOR U7344 ( .A(n6990), .B(n6989), .Z(n6991) );
  XOR U7345 ( .A(n7093), .B(n6991), .Z(n7014) );
  AND U7346 ( .A(y[718]), .B(x[137]), .Z(n7601) );
  NAND U7347 ( .A(n7601), .B(n6995), .Z(n6842) );
  OR U7348 ( .A(n6840), .B(n6839), .Z(n6841) );
  NAND U7349 ( .A(n6842), .B(n6841), .Z(n7013) );
  NAND U7350 ( .A(x[139]), .B(y[706]), .Z(n7063) );
  AND U7351 ( .A(y[709]), .B(x[142]), .Z(n6843) );
  NANDN U7352 ( .A(n7063), .B(n6843), .Z(n6847) );
  OR U7353 ( .A(n6845), .B(n6844), .Z(n6846) );
  NAND U7354 ( .A(n6847), .B(n6846), .Z(n7012) );
  XOR U7355 ( .A(n7013), .B(n7012), .Z(n7015) );
  XNOR U7356 ( .A(n7014), .B(n7015), .Z(n6939) );
  NAND U7357 ( .A(n6849), .B(n6848), .Z(n6853) );
  OR U7358 ( .A(n6851), .B(n6850), .Z(n6852) );
  NAND U7359 ( .A(n6853), .B(n6852), .Z(n6938) );
  XOR U7360 ( .A(n6939), .B(n6938), .Z(n6940) );
  OR U7361 ( .A(n6855), .B(n6854), .Z(n6859) );
  NAND U7362 ( .A(n6857), .B(n6856), .Z(n6858) );
  NAND U7363 ( .A(n6859), .B(n6858), .Z(n6941) );
  XNOR U7364 ( .A(n6940), .B(n6941), .Z(n7018) );
  OR U7365 ( .A(n6861), .B(n6860), .Z(n6865) );
  NANDN U7366 ( .A(n6863), .B(n6862), .Z(n6864) );
  NAND U7367 ( .A(n6865), .B(n6864), .Z(n7019) );
  XNOR U7368 ( .A(n7018), .B(n7019), .Z(n7021) );
  OR U7369 ( .A(n6867), .B(n6866), .Z(n6871) );
  NANDN U7370 ( .A(n6869), .B(n6868), .Z(n6870) );
  NAND U7371 ( .A(n6871), .B(n6870), .Z(n7020) );
  XOR U7372 ( .A(n7021), .B(n7020), .Z(n6928) );
  OR U7373 ( .A(n6873), .B(n6872), .Z(n6877) );
  NANDN U7374 ( .A(n6875), .B(n6874), .Z(n6876) );
  NAND U7375 ( .A(n6877), .B(n6876), .Z(n7027) );
  OR U7376 ( .A(n6879), .B(n6878), .Z(n6883) );
  NANDN U7377 ( .A(n6881), .B(n6880), .Z(n6882) );
  NAND U7378 ( .A(n6883), .B(n6882), .Z(n7025) );
  OR U7379 ( .A(n6885), .B(n6884), .Z(n6889) );
  OR U7380 ( .A(n6887), .B(n6886), .Z(n6888) );
  NAND U7381 ( .A(n6889), .B(n6888), .Z(n6935) );
  NAND U7382 ( .A(x[128]), .B(y[721]), .Z(n6976) );
  NAND U7383 ( .A(x[144]), .B(y[705]), .Z(n6968) );
  XOR U7384 ( .A(o[81]), .B(n6968), .Z(n6974) );
  NAND U7385 ( .A(x[145]), .B(y[704]), .Z(n6973) );
  XNOR U7386 ( .A(n6974), .B(n6973), .Z(n6975) );
  XNOR U7387 ( .A(n6976), .B(n6975), .Z(n6953) );
  NAND U7388 ( .A(x[131]), .B(y[718]), .Z(n6997) );
  AND U7389 ( .A(y[711]), .B(x[138]), .Z(n6891) );
  AND U7390 ( .A(x[130]), .B(y[719]), .Z(n6890) );
  XNOR U7391 ( .A(n6891), .B(n6890), .Z(n6996) );
  XOR U7392 ( .A(n6997), .B(n6996), .Z(n6950) );
  NANDN U7393 ( .A(n6893), .B(n6892), .Z(n6897) );
  NAND U7394 ( .A(n6895), .B(n6894), .Z(n6896) );
  AND U7395 ( .A(n6897), .B(n6896), .Z(n6951) );
  XOR U7396 ( .A(n6953), .B(n6952), .Z(n6959) );
  IV U7397 ( .A(y[719]), .Z(n6994) );
  ANDN U7398 ( .B(x[136]), .A(n6994), .Z(n7744) );
  ANDN U7399 ( .B(y[712]), .A(n152), .Z(n7080) );
  NAND U7400 ( .A(n7744), .B(n7080), .Z(n6901) );
  OR U7401 ( .A(n6899), .B(n6898), .Z(n6900) );
  AND U7402 ( .A(n6901), .B(n6900), .Z(n6957) );
  NAND U7403 ( .A(n6902), .B(n7093), .Z(n6906) );
  OR U7404 ( .A(n6904), .B(n6903), .Z(n6905) );
  AND U7405 ( .A(n6906), .B(n6905), .Z(n6956) );
  XNOR U7406 ( .A(n6957), .B(n6956), .Z(n6958) );
  XOR U7407 ( .A(n6959), .B(n6958), .Z(n6933) );
  ANDN U7408 ( .B(y[715]), .A(n164), .Z(n7807) );
  NAND U7409 ( .A(n6907), .B(n7807), .Z(n6910) );
  NANDN U7410 ( .A(n6908), .B(n7565), .Z(n6909) );
  AND U7411 ( .A(n6910), .B(n6909), .Z(n6947) );
  ANDN U7412 ( .B(y[709]), .A(n163), .Z(n6985) );
  ANDN U7413 ( .B(y[707]), .A(n165), .Z(n6983) );
  ANDN U7414 ( .B(y[706]), .A(n166), .Z(n6984) );
  XNOR U7415 ( .A(n6983), .B(n6984), .Z(n6986) );
  XOR U7416 ( .A(n6985), .B(n6986), .Z(n6945) );
  NANDN U7417 ( .A(n6911), .B(o[80]), .Z(n7009) );
  AND U7418 ( .A(x[137]), .B(y[712]), .Z(n6913) );
  NAND U7419 ( .A(x[129]), .B(y[720]), .Z(n6912) );
  XOR U7420 ( .A(n6913), .B(n6912), .Z(n7008) );
  XNOR U7421 ( .A(n7009), .B(n7008), .Z(n6944) );
  XOR U7422 ( .A(n6945), .B(n6944), .Z(n6946) );
  XOR U7423 ( .A(n6947), .B(n6946), .Z(n6932) );
  XOR U7424 ( .A(n6933), .B(n6932), .Z(n6934) );
  XOR U7425 ( .A(n6935), .B(n6934), .Z(n7024) );
  XNOR U7426 ( .A(n7025), .B(n7024), .Z(n7026) );
  XNOR U7427 ( .A(n7027), .B(n7026), .Z(n6926) );
  OR U7428 ( .A(n6915), .B(n6914), .Z(n6919) );
  NANDN U7429 ( .A(n6917), .B(n6916), .Z(n6918) );
  AND U7430 ( .A(n6919), .B(n6918), .Z(n6927) );
  XOR U7431 ( .A(n6926), .B(n6927), .Z(n6929) );
  XNOR U7432 ( .A(n6928), .B(n6929), .Z(n6923) );
  XOR U7433 ( .A(n6922), .B(n6923), .Z(N178) );
  NANDN U7434 ( .A(n6921), .B(n6920), .Z(n6925) );
  NANDN U7435 ( .A(n6923), .B(n6922), .Z(n6924) );
  NAND U7436 ( .A(n6925), .B(n6924), .Z(n7030) );
  NANDN U7437 ( .A(n6927), .B(n6926), .Z(n6931) );
  OR U7438 ( .A(n6929), .B(n6928), .Z(n6930) );
  AND U7439 ( .A(n6931), .B(n6930), .Z(n7031) );
  XNOR U7440 ( .A(n7030), .B(n7031), .Z(n7032) );
  NANDN U7441 ( .A(n6933), .B(n6932), .Z(n6937) );
  OR U7442 ( .A(n6935), .B(n6934), .Z(n6936) );
  AND U7443 ( .A(n6937), .B(n6936), .Z(n7140) );
  OR U7444 ( .A(n6939), .B(n6938), .Z(n6943) );
  NANDN U7445 ( .A(n6941), .B(n6940), .Z(n6942) );
  AND U7446 ( .A(n6943), .B(n6942), .Z(n7141) );
  XOR U7447 ( .A(n7140), .B(n7141), .Z(n7143) );
  OR U7448 ( .A(n6945), .B(n6944), .Z(n6949) );
  NANDN U7449 ( .A(n6947), .B(n6946), .Z(n6948) );
  AND U7450 ( .A(n6949), .B(n6948), .Z(n7116) );
  NANDN U7451 ( .A(n6951), .B(n6950), .Z(n6955) );
  NANDN U7452 ( .A(n6953), .B(n6952), .Z(n6954) );
  AND U7453 ( .A(n6955), .B(n6954), .Z(n7117) );
  XOR U7454 ( .A(n7116), .B(n7117), .Z(n7118) );
  OR U7455 ( .A(n6957), .B(n6956), .Z(n6961) );
  OR U7456 ( .A(n6959), .B(n6958), .Z(n6960) );
  AND U7457 ( .A(n6961), .B(n6960), .Z(n7119) );
  OR U7458 ( .A(n6963), .B(n6962), .Z(n6967) );
  OR U7459 ( .A(n6965), .B(n6964), .Z(n6966) );
  NAND U7460 ( .A(n6967), .B(n6966), .Z(n7071) );
  NANDN U7461 ( .A(n6968), .B(o[81]), .Z(n7082) );
  AND U7462 ( .A(x[138]), .B(y[712]), .Z(n6970) );
  NAND U7463 ( .A(x[129]), .B(y[721]), .Z(n6969) );
  XNOR U7464 ( .A(n6970), .B(n6969), .Z(n7081) );
  XNOR U7465 ( .A(n7082), .B(n7081), .Z(n7068) );
  NAND U7466 ( .A(x[142]), .B(y[708]), .Z(n6971) );
  XOR U7467 ( .A(n6972), .B(n6971), .Z(n7058) );
  NAND U7468 ( .A(y[707]), .B(x[143]), .Z(n7057) );
  XNOR U7469 ( .A(n7058), .B(n7057), .Z(n7069) );
  XOR U7470 ( .A(n7068), .B(n7069), .Z(n7070) );
  XNOR U7471 ( .A(n7071), .B(n7070), .Z(n7135) );
  OR U7472 ( .A(n6974), .B(n6973), .Z(n6978) );
  OR U7473 ( .A(n6976), .B(n6975), .Z(n6977) );
  NAND U7474 ( .A(n6978), .B(n6977), .Z(n7123) );
  NAND U7475 ( .A(x[135]), .B(y[715]), .Z(n6979) );
  XOR U7476 ( .A(n6980), .B(n6979), .Z(n7096) );
  NAND U7477 ( .A(y[718]), .B(x[132]), .Z(n7095) );
  XNOR U7478 ( .A(n7096), .B(n7095), .Z(n7049) );
  AND U7479 ( .A(x[133]), .B(y[717]), .Z(n7211) );
  NAND U7480 ( .A(x[134]), .B(y[716]), .Z(n7048) );
  XNOR U7481 ( .A(n7211), .B(n7048), .Z(n7050) );
  XOR U7482 ( .A(n7123), .B(n7122), .Z(n7125) );
  NAND U7483 ( .A(x[130]), .B(y[720]), .Z(n7065) );
  AND U7484 ( .A(y[711]), .B(x[139]), .Z(n6982) );
  AND U7485 ( .A(y[706]), .B(x[144]), .Z(n6981) );
  XNOR U7486 ( .A(n6982), .B(n6981), .Z(n7064) );
  XOR U7487 ( .A(n7065), .B(n7064), .Z(n7124) );
  XNOR U7488 ( .A(n7125), .B(n7124), .Z(n7134) );
  XOR U7489 ( .A(n7135), .B(n7134), .Z(n7137) );
  OR U7490 ( .A(n6984), .B(n6983), .Z(n6988) );
  OR U7491 ( .A(n6986), .B(n6985), .Z(n6987) );
  NAND U7492 ( .A(n6988), .B(n6987), .Z(n7136) );
  XNOR U7493 ( .A(n7137), .B(n7136), .Z(n7042) );
  NANDN U7494 ( .A(n6990), .B(n6989), .Z(n6993) );
  NANDN U7495 ( .A(n6991), .B(n7093), .Z(n6992) );
  NAND U7496 ( .A(n6993), .B(n6992), .Z(n7111) );
  NOR U7497 ( .A(n161), .B(n6994), .Z(n7962) );
  NAND U7498 ( .A(n7962), .B(n6995), .Z(n6999) );
  OR U7499 ( .A(n6997), .B(n6996), .Z(n6998) );
  AND U7500 ( .A(n6999), .B(n6998), .Z(n7076) );
  NAND U7501 ( .A(x[128]), .B(y[722]), .Z(n7086) );
  NAND U7502 ( .A(x[146]), .B(y[704]), .Z(n7085) );
  XOR U7503 ( .A(n7086), .B(n7085), .Z(n7087) );
  NAND U7504 ( .A(x[145]), .B(y[705]), .Z(n7099) );
  XOR U7505 ( .A(o[82]), .B(n7099), .Z(n7088) );
  XOR U7506 ( .A(n7087), .B(n7088), .Z(n7075) );
  ANDN U7507 ( .B(y[710]), .A(n163), .Z(n7175) );
  AND U7508 ( .A(x[131]), .B(y[719]), .Z(n7001) );
  NAND U7509 ( .A(x[141]), .B(y[709]), .Z(n7000) );
  XOR U7510 ( .A(n7001), .B(n7000), .Z(n7107) );
  XOR U7511 ( .A(n7175), .B(n7107), .Z(n7074) );
  XNOR U7512 ( .A(n7075), .B(n7074), .Z(n7077) );
  XOR U7513 ( .A(n7076), .B(n7077), .Z(n7128) );
  OR U7514 ( .A(n7003), .B(n7002), .Z(n7007) );
  OR U7515 ( .A(n7005), .B(n7004), .Z(n7006) );
  AND U7516 ( .A(n7007), .B(n7006), .Z(n7129) );
  XNOR U7517 ( .A(n7128), .B(n7129), .Z(n7131) );
  AND U7518 ( .A(y[720]), .B(x[137]), .Z(n7963) );
  NAND U7519 ( .A(n7080), .B(n7963), .Z(n7011) );
  OR U7520 ( .A(n7009), .B(n7008), .Z(n7010) );
  NAND U7521 ( .A(n7011), .B(n7010), .Z(n7130) );
  XNOR U7522 ( .A(n7131), .B(n7130), .Z(n7110) );
  XNOR U7523 ( .A(n7111), .B(n7110), .Z(n7113) );
  OR U7524 ( .A(n7013), .B(n7012), .Z(n7017) );
  NAND U7525 ( .A(n7015), .B(n7014), .Z(n7016) );
  AND U7526 ( .A(n7017), .B(n7016), .Z(n7112) );
  XNOR U7527 ( .A(n7113), .B(n7112), .Z(n7043) );
  XOR U7528 ( .A(n7042), .B(n7043), .Z(n7045) );
  XNOR U7529 ( .A(n7044), .B(n7045), .Z(n7142) );
  XNOR U7530 ( .A(n7143), .B(n7142), .Z(n7039) );
  OR U7531 ( .A(n7019), .B(n7018), .Z(n7023) );
  OR U7532 ( .A(n7021), .B(n7020), .Z(n7022) );
  NAND U7533 ( .A(n7023), .B(n7022), .Z(n7037) );
  OR U7534 ( .A(n7025), .B(n7024), .Z(n7029) );
  OR U7535 ( .A(n7027), .B(n7026), .Z(n7028) );
  NAND U7536 ( .A(n7029), .B(n7028), .Z(n7036) );
  XNOR U7537 ( .A(n7037), .B(n7036), .Z(n7038) );
  XNOR U7538 ( .A(n7039), .B(n7038), .Z(n7033) );
  XOR U7539 ( .A(n7032), .B(n7033), .Z(N179) );
  NANDN U7540 ( .A(n7031), .B(n7030), .Z(n7035) );
  NANDN U7541 ( .A(n7033), .B(n7032), .Z(n7034) );
  NAND U7542 ( .A(n7035), .B(n7034), .Z(n7255) );
  OR U7543 ( .A(n7037), .B(n7036), .Z(n7041) );
  OR U7544 ( .A(n7039), .B(n7038), .Z(n7040) );
  AND U7545 ( .A(n7041), .B(n7040), .Z(n7256) );
  XNOR U7546 ( .A(n7255), .B(n7256), .Z(n7257) );
  NANDN U7547 ( .A(n7043), .B(n7042), .Z(n7047) );
  NANDN U7548 ( .A(n7045), .B(n7044), .Z(n7046) );
  AND U7549 ( .A(n7047), .B(n7046), .Z(n7261) );
  NANDN U7550 ( .A(n7211), .B(n7048), .Z(n7052) );
  NAND U7551 ( .A(n7050), .B(n7049), .Z(n7051) );
  AND U7552 ( .A(n7052), .B(n7051), .Z(n7245) );
  AND U7553 ( .A(y[715]), .B(x[136]), .Z(n7054) );
  NAND U7554 ( .A(x[142]), .B(y[709]), .Z(n7053) );
  XOR U7555 ( .A(n7054), .B(n7053), .Z(n7223) );
  NAND U7556 ( .A(y[722]), .B(x[129]), .Z(n7222) );
  XOR U7557 ( .A(n7223), .B(n7222), .Z(n7160) );
  ANDN U7558 ( .B(x[142]), .A(n7055), .Z(n7704) );
  AND U7559 ( .A(y[708]), .B(x[137]), .Z(n7056) );
  NAND U7560 ( .A(n7704), .B(n7056), .Z(n7060) );
  OR U7561 ( .A(n7058), .B(n7057), .Z(n7059) );
  NAND U7562 ( .A(n7060), .B(n7059), .Z(n7158) );
  NAND U7563 ( .A(x[141]), .B(y[710]), .Z(n7061) );
  XOR U7564 ( .A(n7062), .B(n7061), .Z(n7178) );
  NAND U7565 ( .A(y[721]), .B(x[130]), .Z(n7177) );
  XNOR U7566 ( .A(n7178), .B(n7177), .Z(n7159) );
  XOR U7567 ( .A(n7158), .B(n7159), .Z(n7161) );
  XNOR U7568 ( .A(n7160), .B(n7161), .Z(n7243) );
  AND U7569 ( .A(y[711]), .B(x[144]), .Z(n7559) );
  NANDN U7570 ( .A(n7063), .B(n7559), .Z(n7067) );
  OR U7571 ( .A(n7065), .B(n7064), .Z(n7066) );
  NAND U7572 ( .A(n7067), .B(n7066), .Z(n7244) );
  XNOR U7573 ( .A(n7243), .B(n7244), .Z(n7246) );
  XOR U7574 ( .A(n7245), .B(n7246), .Z(n7249) );
  NANDN U7575 ( .A(n7069), .B(n7068), .Z(n7073) );
  OR U7576 ( .A(n7071), .B(n7070), .Z(n7072) );
  NAND U7577 ( .A(n7073), .B(n7072), .Z(n7238) );
  OR U7578 ( .A(n7075), .B(n7074), .Z(n7079) );
  OR U7579 ( .A(n7077), .B(n7076), .Z(n7078) );
  NAND U7580 ( .A(n7079), .B(n7078), .Z(n7237) );
  XOR U7581 ( .A(n7238), .B(n7237), .Z(n7239) );
  AND U7582 ( .A(x[138]), .B(y[721]), .Z(n8328) );
  NAND U7583 ( .A(n7080), .B(n8328), .Z(n7084) );
  NANDN U7584 ( .A(n7082), .B(n7081), .Z(n7083) );
  NAND U7585 ( .A(n7084), .B(n7083), .Z(n7201) );
  OR U7586 ( .A(n7086), .B(n7085), .Z(n7090) );
  NANDN U7587 ( .A(n7088), .B(n7087), .Z(n7089) );
  NAND U7588 ( .A(n7090), .B(n7089), .Z(n7200) );
  AND U7589 ( .A(x[137]), .B(y[714]), .Z(n7092) );
  NAND U7590 ( .A(x[144]), .B(y[707]), .Z(n7091) );
  XOR U7591 ( .A(n7092), .B(n7091), .Z(n7172) );
  NAND U7592 ( .A(x[143]), .B(y[708]), .Z(n7171) );
  XOR U7593 ( .A(n7172), .B(n7171), .Z(n7199) );
  XNOR U7594 ( .A(n7200), .B(n7199), .Z(n7202) );
  XNOR U7595 ( .A(n7201), .B(n7202), .Z(n7233) );
  NANDN U7596 ( .A(n7094), .B(n7093), .Z(n7098) );
  OR U7597 ( .A(n7096), .B(n7095), .Z(n7097) );
  NAND U7598 ( .A(n7098), .B(n7097), .Z(n7164) );
  NANDN U7599 ( .A(n7099), .B(o[82]), .Z(n7208) );
  NAND U7600 ( .A(x[128]), .B(y[723]), .Z(n7206) );
  NAND U7601 ( .A(x[147]), .B(y[704]), .Z(n7205) );
  XOR U7602 ( .A(n7206), .B(n7205), .Z(n7207) );
  XOR U7603 ( .A(n7208), .B(n7207), .Z(n7165) );
  XOR U7604 ( .A(n7164), .B(n7165), .Z(n7167) );
  NAND U7605 ( .A(x[132]), .B(y[719]), .Z(n7331) );
  AND U7606 ( .A(x[134]), .B(y[717]), .Z(n7101) );
  NAND U7607 ( .A(x[133]), .B(y[718]), .Z(n7100) );
  XNOR U7608 ( .A(n7101), .B(n7100), .Z(n7212) );
  XNOR U7609 ( .A(n7167), .B(n7166), .Z(n7231) );
  AND U7610 ( .A(x[139]), .B(y[712]), .Z(n7103) );
  NAND U7611 ( .A(x[135]), .B(y[716]), .Z(n7102) );
  XOR U7612 ( .A(n7103), .B(n7102), .Z(n7187) );
  NAND U7613 ( .A(x[131]), .B(y[720]), .Z(n7186) );
  XNOR U7614 ( .A(n7187), .B(n7186), .Z(n7196) );
  NAND U7615 ( .A(x[146]), .B(y[705]), .Z(n7192) );
  XOR U7616 ( .A(o[83]), .B(n7192), .Z(n7228) );
  AND U7617 ( .A(x[138]), .B(y[713]), .Z(n7105) );
  NAND U7618 ( .A(x[145]), .B(y[706]), .Z(n7104) );
  XOR U7619 ( .A(n7105), .B(n7104), .Z(n7227) );
  XNOR U7620 ( .A(n7228), .B(n7227), .Z(n7193) );
  AND U7621 ( .A(x[141]), .B(y[719]), .Z(n8435) );
  NAND U7622 ( .A(n7106), .B(n8435), .Z(n7109) );
  NANDN U7623 ( .A(n7107), .B(n7175), .Z(n7108) );
  NAND U7624 ( .A(n7109), .B(n7108), .Z(n7194) );
  XNOR U7625 ( .A(n7196), .B(n7195), .Z(n7232) );
  XNOR U7626 ( .A(n7231), .B(n7232), .Z(n7234) );
  XNOR U7627 ( .A(n7233), .B(n7234), .Z(n7240) );
  XNOR U7628 ( .A(n7239), .B(n7240), .Z(n7250) );
  XNOR U7629 ( .A(n7249), .B(n7250), .Z(n7252) );
  OR U7630 ( .A(n7111), .B(n7110), .Z(n7115) );
  OR U7631 ( .A(n7113), .B(n7112), .Z(n7114) );
  NAND U7632 ( .A(n7115), .B(n7114), .Z(n7251) );
  XOR U7633 ( .A(n7252), .B(n7251), .Z(n7155) );
  OR U7634 ( .A(n7117), .B(n7116), .Z(n7121) );
  NANDN U7635 ( .A(n7119), .B(n7118), .Z(n7120) );
  NAND U7636 ( .A(n7121), .B(n7120), .Z(n7153) );
  NANDN U7637 ( .A(n7123), .B(n7122), .Z(n7127) );
  OR U7638 ( .A(n7125), .B(n7124), .Z(n7126) );
  AND U7639 ( .A(n7127), .B(n7126), .Z(n7148) );
  OR U7640 ( .A(n7129), .B(n7128), .Z(n7133) );
  OR U7641 ( .A(n7131), .B(n7130), .Z(n7132) );
  AND U7642 ( .A(n7133), .B(n7132), .Z(n7146) );
  NANDN U7643 ( .A(n7135), .B(n7134), .Z(n7139) );
  OR U7644 ( .A(n7137), .B(n7136), .Z(n7138) );
  NAND U7645 ( .A(n7139), .B(n7138), .Z(n7147) );
  XNOR U7646 ( .A(n7146), .B(n7147), .Z(n7149) );
  XNOR U7647 ( .A(n7148), .B(n7149), .Z(n7152) );
  XOR U7648 ( .A(n7153), .B(n7152), .Z(n7154) );
  XOR U7649 ( .A(n7155), .B(n7154), .Z(n7262) );
  XOR U7650 ( .A(n7261), .B(n7262), .Z(n7263) );
  OR U7651 ( .A(n7141), .B(n7140), .Z(n7145) );
  NAND U7652 ( .A(n7143), .B(n7142), .Z(n7144) );
  AND U7653 ( .A(n7145), .B(n7144), .Z(n7264) );
  XOR U7654 ( .A(n7257), .B(n7258), .Z(N180) );
  OR U7655 ( .A(n7147), .B(n7146), .Z(n7151) );
  OR U7656 ( .A(n7149), .B(n7148), .Z(n7150) );
  AND U7657 ( .A(n7151), .B(n7150), .Z(n7276) );
  OR U7658 ( .A(n7153), .B(n7152), .Z(n7157) );
  NANDN U7659 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U7660 ( .A(n7157), .B(n7156), .Z(n7273) );
  NANDN U7661 ( .A(n7159), .B(n7158), .Z(n7163) );
  NANDN U7662 ( .A(n7161), .B(n7160), .Z(n7162) );
  NAND U7663 ( .A(n7163), .B(n7162), .Z(n7279) );
  NANDN U7664 ( .A(n7165), .B(n7164), .Z(n7169) );
  NANDN U7665 ( .A(n7167), .B(n7166), .Z(n7168) );
  AND U7666 ( .A(n7169), .B(n7168), .Z(n7280) );
  AND U7667 ( .A(x[144]), .B(y[714]), .Z(n8127) );
  NANDN U7668 ( .A(n7170), .B(n8127), .Z(n7174) );
  OR U7669 ( .A(n7172), .B(n7171), .Z(n7173) );
  NAND U7670 ( .A(n7174), .B(n7173), .Z(n7319) );
  AND U7671 ( .A(y[711]), .B(x[141]), .Z(n7176) );
  NAND U7672 ( .A(n7176), .B(n7175), .Z(n7180) );
  OR U7673 ( .A(n7178), .B(n7177), .Z(n7179) );
  NAND U7674 ( .A(n7180), .B(n7179), .Z(n7357) );
  NAND U7675 ( .A(x[130]), .B(y[722]), .Z(n7345) );
  AND U7676 ( .A(x[138]), .B(y[714]), .Z(n7182) );
  NAND U7677 ( .A(x[144]), .B(y[708]), .Z(n7181) );
  XNOR U7678 ( .A(n7182), .B(n7181), .Z(n7344) );
  AND U7679 ( .A(y[709]), .B(x[143]), .Z(n7184) );
  NAND U7680 ( .A(x[137]), .B(y[715]), .Z(n7183) );
  XOR U7681 ( .A(n7184), .B(n7183), .Z(n7309) );
  NAND U7682 ( .A(y[710]), .B(x[142]), .Z(n7308) );
  XOR U7683 ( .A(n7309), .B(n7308), .Z(n7354) );
  XNOR U7684 ( .A(n7357), .B(n7356), .Z(n7320) );
  ANDN U7685 ( .B(y[716]), .A(n162), .Z(n7739) );
  NAND U7686 ( .A(n7739), .B(n7185), .Z(n7189) );
  OR U7687 ( .A(n7187), .B(n7186), .Z(n7188) );
  AND U7688 ( .A(n7189), .B(n7188), .Z(n7362) );
  AND U7689 ( .A(y[705]), .B(x[147]), .Z(n7312) );
  XNOR U7690 ( .A(o[84]), .B(n7312), .Z(n7304) );
  AND U7691 ( .A(x[139]), .B(y[713]), .Z(n7191) );
  NAND U7692 ( .A(x[129]), .B(y[723]), .Z(n7190) );
  XNOR U7693 ( .A(n7191), .B(n7190), .Z(n7303) );
  XOR U7694 ( .A(n7304), .B(n7303), .Z(n7361) );
  NANDN U7695 ( .A(n7192), .B(o[83]), .Z(n7328) );
  NAND U7696 ( .A(x[148]), .B(y[704]), .Z(n7326) );
  NAND U7697 ( .A(y[724]), .B(x[128]), .Z(n7325) );
  XOR U7698 ( .A(n7326), .B(n7325), .Z(n7327) );
  XNOR U7699 ( .A(n7328), .B(n7327), .Z(n7360) );
  XOR U7700 ( .A(n7361), .B(n7360), .Z(n7363) );
  XOR U7701 ( .A(n7362), .B(n7363), .Z(n7321) );
  NANDN U7702 ( .A(n7194), .B(n7193), .Z(n7198) );
  NAND U7703 ( .A(n7196), .B(n7195), .Z(n7197) );
  NAND U7704 ( .A(n7198), .B(n7197), .Z(n7366) );
  NAND U7705 ( .A(n7200), .B(n7199), .Z(n7204) );
  NANDN U7706 ( .A(n7202), .B(n7201), .Z(n7203) );
  NAND U7707 ( .A(n7204), .B(n7203), .Z(n7316) );
  OR U7708 ( .A(n7206), .B(n7205), .Z(n7210) );
  NANDN U7709 ( .A(n7208), .B(n7207), .Z(n7209) );
  NAND U7710 ( .A(n7210), .B(n7209), .Z(n7287) );
  ANDN U7711 ( .B(y[718]), .A(n157), .Z(n7291) );
  NAND U7712 ( .A(n7291), .B(n7211), .Z(n7214) );
  NANDN U7713 ( .A(n7331), .B(n7212), .Z(n7213) );
  NAND U7714 ( .A(n7214), .B(n7213), .Z(n7285) );
  AND U7715 ( .A(x[140]), .B(y[712]), .Z(n7216) );
  NAND U7716 ( .A(x[146]), .B(y[706]), .Z(n7215) );
  XOR U7717 ( .A(n7216), .B(n7215), .Z(n7299) );
  NAND U7718 ( .A(y[707]), .B(x[145]), .Z(n7298) );
  XNOR U7719 ( .A(n7299), .B(n7298), .Z(n7286) );
  XOR U7720 ( .A(n7285), .B(n7286), .Z(n7288) );
  NAND U7721 ( .A(x[135]), .B(y[717]), .Z(n7333) );
  AND U7722 ( .A(x[133]), .B(y[719]), .Z(n7218) );
  NAND U7723 ( .A(x[132]), .B(y[720]), .Z(n7217) );
  XNOR U7724 ( .A(n7218), .B(n7217), .Z(n7332) );
  XNOR U7725 ( .A(n7291), .B(n7292), .Z(n7294) );
  NAND U7726 ( .A(x[136]), .B(y[716]), .Z(n7340) );
  AND U7727 ( .A(x[131]), .B(y[721]), .Z(n7220) );
  NAND U7728 ( .A(x[141]), .B(y[711]), .Z(n7219) );
  XNOR U7729 ( .A(n7220), .B(n7219), .Z(n7339) );
  XOR U7730 ( .A(n7294), .B(n7293), .Z(n7351) );
  ANDN U7731 ( .B(y[715]), .A(n165), .Z(n8013) );
  NAND U7732 ( .A(n8013), .B(n7221), .Z(n7225) );
  OR U7733 ( .A(n7223), .B(n7222), .Z(n7224) );
  NAND U7734 ( .A(n7225), .B(n7224), .Z(n7349) );
  ANDN U7735 ( .B(y[713]), .A(n168), .Z(n8140) );
  NANDN U7736 ( .A(n7226), .B(n8140), .Z(n7230) );
  OR U7737 ( .A(n7228), .B(n7227), .Z(n7229) );
  AND U7738 ( .A(n7230), .B(n7229), .Z(n7348) );
  XNOR U7739 ( .A(n7351), .B(n7350), .Z(n7314) );
  XNOR U7740 ( .A(n7313), .B(n7314), .Z(n7315) );
  XOR U7741 ( .A(n7316), .B(n7315), .Z(n7367) );
  XOR U7742 ( .A(n7366), .B(n7367), .Z(n7368) );
  XOR U7743 ( .A(n7369), .B(n7368), .Z(n7372) );
  OR U7744 ( .A(n7232), .B(n7231), .Z(n7236) );
  OR U7745 ( .A(n7234), .B(n7233), .Z(n7235) );
  NAND U7746 ( .A(n7236), .B(n7235), .Z(n7379) );
  OR U7747 ( .A(n7238), .B(n7237), .Z(n7242) );
  NANDN U7748 ( .A(n7240), .B(n7239), .Z(n7241) );
  NAND U7749 ( .A(n7242), .B(n7241), .Z(n7378) );
  XOR U7750 ( .A(n7379), .B(n7378), .Z(n7380) );
  OR U7751 ( .A(n7244), .B(n7243), .Z(n7248) );
  OR U7752 ( .A(n7246), .B(n7245), .Z(n7247) );
  NAND U7753 ( .A(n7248), .B(n7247), .Z(n7381) );
  XNOR U7754 ( .A(n7372), .B(n7373), .Z(n7375) );
  OR U7755 ( .A(n7250), .B(n7249), .Z(n7254) );
  OR U7756 ( .A(n7252), .B(n7251), .Z(n7253) );
  AND U7757 ( .A(n7254), .B(n7253), .Z(n7374) );
  XOR U7758 ( .A(n7375), .B(n7374), .Z(n7274) );
  XNOR U7759 ( .A(n7273), .B(n7274), .Z(n7275) );
  XOR U7760 ( .A(n7276), .B(n7275), .Z(n7269) );
  NANDN U7761 ( .A(n7256), .B(n7255), .Z(n7260) );
  NANDN U7762 ( .A(n7258), .B(n7257), .Z(n7259) );
  NAND U7763 ( .A(n7260), .B(n7259), .Z(n7267) );
  OR U7764 ( .A(n7262), .B(n7261), .Z(n7266) );
  NANDN U7765 ( .A(n7264), .B(n7263), .Z(n7265) );
  AND U7766 ( .A(n7266), .B(n7265), .Z(n7268) );
  XNOR U7767 ( .A(n7267), .B(n7268), .Z(n7270) );
  XNOR U7768 ( .A(n7269), .B(n7270), .Z(N181) );
  NANDN U7769 ( .A(n7268), .B(n7267), .Z(n7272) );
  NAND U7770 ( .A(n7270), .B(n7269), .Z(n7271) );
  NAND U7771 ( .A(n7272), .B(n7271), .Z(n7384) );
  OR U7772 ( .A(n7274), .B(n7273), .Z(n7278) );
  OR U7773 ( .A(n7276), .B(n7275), .Z(n7277) );
  AND U7774 ( .A(n7278), .B(n7277), .Z(n7385) );
  XNOR U7775 ( .A(n7384), .B(n7385), .Z(n7386) );
  NANDN U7776 ( .A(n7280), .B(n7279), .Z(n7284) );
  NAND U7777 ( .A(n7282), .B(n7281), .Z(n7283) );
  NAND U7778 ( .A(n7284), .B(n7283), .Z(n7405) );
  NANDN U7779 ( .A(n7286), .B(n7285), .Z(n7290) );
  NANDN U7780 ( .A(n7288), .B(n7287), .Z(n7289) );
  NAND U7781 ( .A(n7290), .B(n7289), .Z(n7429) );
  NAND U7782 ( .A(n7292), .B(n7291), .Z(n7296) );
  NANDN U7783 ( .A(n7294), .B(n7293), .Z(n7295) );
  NAND U7784 ( .A(n7296), .B(n7295), .Z(n7426) );
  ANDN U7785 ( .B(y[712]), .A(n169), .Z(n8138) );
  NAND U7786 ( .A(n7297), .B(n8138), .Z(n7301) );
  OR U7787 ( .A(n7299), .B(n7298), .Z(n7300) );
  NAND U7788 ( .A(n7301), .B(n7300), .Z(n7423) );
  AND U7789 ( .A(y[723]), .B(x[139]), .Z(n8943) );
  NAND U7790 ( .A(n7302), .B(n8943), .Z(n7306) );
  NANDN U7791 ( .A(n7304), .B(n7303), .Z(n7305) );
  NAND U7792 ( .A(n7306), .B(n7305), .Z(n7420) );
  ANDN U7793 ( .B(y[720]), .A(n156), .Z(n7487) );
  AND U7794 ( .A(y[709]), .B(x[144]), .Z(n7486) );
  XOR U7795 ( .A(n7487), .B(n7486), .Z(n7489) );
  ANDN U7796 ( .B(y[710]), .A(n166), .Z(n7488) );
  XOR U7797 ( .A(n7489), .B(n7488), .Z(n7492) );
  ANDN U7798 ( .B(y[715]), .A(n166), .Z(n8132) );
  NAND U7799 ( .A(n7307), .B(n8132), .Z(n7311) );
  OR U7800 ( .A(n7309), .B(n7308), .Z(n7310) );
  NAND U7801 ( .A(n7311), .B(n7310), .Z(n7493) );
  XNOR U7802 ( .A(n7492), .B(n7493), .Z(n7495) );
  ANDN U7803 ( .B(y[725]), .A(n151), .Z(n7470) );
  AND U7804 ( .A(n7312), .B(o[84]), .Z(n7468) );
  ANDN U7805 ( .B(y[704]), .A(n172), .Z(n7469) );
  XNOR U7806 ( .A(n7468), .B(n7469), .Z(n7471) );
  XNOR U7807 ( .A(n7470), .B(n7471), .Z(n7494) );
  XOR U7808 ( .A(n7495), .B(n7494), .Z(n7421) );
  XNOR U7809 ( .A(n7423), .B(n7422), .Z(n7427) );
  XNOR U7810 ( .A(n7429), .B(n7428), .Z(n7403) );
  NANDN U7811 ( .A(n7314), .B(n7313), .Z(n7318) );
  NANDN U7812 ( .A(n7316), .B(n7315), .Z(n7317) );
  AND U7813 ( .A(n7318), .B(n7317), .Z(n7402) );
  XNOR U7814 ( .A(n7405), .B(n7404), .Z(n7399) );
  NANDN U7815 ( .A(n7320), .B(n7319), .Z(n7324) );
  NAND U7816 ( .A(n7322), .B(n7321), .Z(n7323) );
  NAND U7817 ( .A(n7324), .B(n7323), .Z(n7500) );
  OR U7818 ( .A(n7326), .B(n7325), .Z(n7330) );
  NANDN U7819 ( .A(n7328), .B(n7327), .Z(n7329) );
  NAND U7820 ( .A(n7330), .B(n7329), .Z(n7408) );
  NANDN U7821 ( .A(n7331), .B(n7487), .Z(n7335) );
  NANDN U7822 ( .A(n7333), .B(n7332), .Z(n7334) );
  AND U7823 ( .A(n7335), .B(n7334), .Z(n7409) );
  ANDN U7824 ( .B(y[719]), .A(n157), .Z(n7464) );
  ANDN U7825 ( .B(y[711]), .A(n165), .Z(n7463) );
  XNOR U7826 ( .A(n7743), .B(n7463), .Z(n7465) );
  XNOR U7827 ( .A(n7464), .B(n7465), .Z(n7440) );
  AND U7828 ( .A(x[136]), .B(y[717]), .Z(n7801) );
  XNOR U7829 ( .A(n7438), .B(n7801), .Z(n7439) );
  XOR U7830 ( .A(n7440), .B(n7439), .Z(n7459) );
  NAND U7831 ( .A(x[132]), .B(y[721]), .Z(n7483) );
  AND U7832 ( .A(y[722]), .B(x[131]), .Z(n7337) );
  AND U7833 ( .A(x[141]), .B(y[712]), .Z(n7336) );
  XNOR U7834 ( .A(n7337), .B(n7336), .Z(n7482) );
  XOR U7835 ( .A(n7483), .B(n7482), .Z(n7457) );
  ANDN U7836 ( .B(y[713]), .A(n163), .Z(n7445) );
  ANDN U7837 ( .B(y[723]), .A(n153), .Z(n7443) );
  ANDN U7838 ( .B(y[708]), .A(n168), .Z(n7444) );
  XNOR U7839 ( .A(n7443), .B(n7444), .Z(n7446) );
  XOR U7840 ( .A(n7445), .B(n7446), .Z(n7458) );
  XOR U7841 ( .A(n7457), .B(n7458), .Z(n7460) );
  XNOR U7842 ( .A(n7459), .B(n7460), .Z(n7411) );
  XOR U7843 ( .A(n7410), .B(n7411), .Z(n7434) );
  ANDN U7844 ( .B(y[724]), .A(n152), .Z(n7475) );
  NAND U7845 ( .A(y[707]), .B(x[146]), .Z(n7474) );
  XOR U7846 ( .A(n7475), .B(n7474), .Z(n7476) );
  XOR U7847 ( .A(n7477), .B(n7476), .Z(n7414) );
  NAND U7848 ( .A(x[139]), .B(y[714]), .Z(n7454) );
  AND U7849 ( .A(y[705]), .B(x[148]), .Z(n7480) );
  XNOR U7850 ( .A(o[85]), .B(n7480), .Z(n7452) );
  NAND U7851 ( .A(x[147]), .B(y[706]), .Z(n7451) );
  XOR U7852 ( .A(n7452), .B(n7451), .Z(n7453) );
  XOR U7853 ( .A(n7454), .B(n7453), .Z(n7415) );
  XOR U7854 ( .A(n7414), .B(n7415), .Z(n7416) );
  AND U7855 ( .A(x[141]), .B(y[721]), .Z(n8590) );
  NAND U7856 ( .A(n8590), .B(n7338), .Z(n7342) );
  NANDN U7857 ( .A(n7340), .B(n7339), .Z(n7341) );
  AND U7858 ( .A(n7342), .B(n7341), .Z(n7417) );
  XOR U7859 ( .A(n7416), .B(n7417), .Z(n7432) );
  NAND U7860 ( .A(n7343), .B(n8127), .Z(n7347) );
  NANDN U7861 ( .A(n7345), .B(n7344), .Z(n7346) );
  NAND U7862 ( .A(n7347), .B(n7346), .Z(n7433) );
  XOR U7863 ( .A(n7434), .B(n7435), .Z(n7498) );
  NANDN U7864 ( .A(n7349), .B(n7348), .Z(n7353) );
  NAND U7865 ( .A(n7351), .B(n7350), .Z(n7352) );
  AND U7866 ( .A(n7353), .B(n7352), .Z(n7504) );
  NAND U7867 ( .A(n7355), .B(n7354), .Z(n7359) );
  NAND U7868 ( .A(n7357), .B(n7356), .Z(n7358) );
  NAND U7869 ( .A(n7359), .B(n7358), .Z(n7505) );
  XOR U7870 ( .A(n7504), .B(n7505), .Z(n7506) );
  NANDN U7871 ( .A(n7361), .B(n7360), .Z(n7365) );
  OR U7872 ( .A(n7363), .B(n7362), .Z(n7364) );
  NAND U7873 ( .A(n7365), .B(n7364), .Z(n7507) );
  XNOR U7874 ( .A(n7506), .B(n7507), .Z(n7499) );
  XOR U7875 ( .A(n7498), .B(n7499), .Z(n7501) );
  XOR U7876 ( .A(n7500), .B(n7501), .Z(n7397) );
  NANDN U7877 ( .A(n7367), .B(n7366), .Z(n7371) );
  OR U7878 ( .A(n7369), .B(n7368), .Z(n7370) );
  AND U7879 ( .A(n7371), .B(n7370), .Z(n7396) );
  XNOR U7880 ( .A(n7399), .B(n7398), .Z(n7393) );
  OR U7881 ( .A(n7373), .B(n7372), .Z(n7377) );
  OR U7882 ( .A(n7375), .B(n7374), .Z(n7376) );
  NAND U7883 ( .A(n7377), .B(n7376), .Z(n7391) );
  OR U7884 ( .A(n7379), .B(n7378), .Z(n7383) );
  NANDN U7885 ( .A(n7381), .B(n7380), .Z(n7382) );
  NAND U7886 ( .A(n7383), .B(n7382), .Z(n7390) );
  XOR U7887 ( .A(n7391), .B(n7390), .Z(n7392) );
  XOR U7888 ( .A(n7393), .B(n7392), .Z(n7387) );
  XOR U7889 ( .A(n7386), .B(n7387), .Z(N182) );
  NANDN U7890 ( .A(n7385), .B(n7384), .Z(n7389) );
  NANDN U7891 ( .A(n7387), .B(n7386), .Z(n7388) );
  NAND U7892 ( .A(n7389), .B(n7388), .Z(n7510) );
  OR U7893 ( .A(n7391), .B(n7390), .Z(n7395) );
  NANDN U7894 ( .A(n7393), .B(n7392), .Z(n7394) );
  AND U7895 ( .A(n7395), .B(n7394), .Z(n7511) );
  XNOR U7896 ( .A(n7510), .B(n7511), .Z(n7512) );
  NANDN U7897 ( .A(n7397), .B(n7396), .Z(n7401) );
  NANDN U7898 ( .A(n7399), .B(n7398), .Z(n7400) );
  NAND U7899 ( .A(n7401), .B(n7400), .Z(n7519) );
  NANDN U7900 ( .A(n7403), .B(n7402), .Z(n7407) );
  NAND U7901 ( .A(n7405), .B(n7404), .Z(n7406) );
  NAND U7902 ( .A(n7407), .B(n7406), .Z(n7516) );
  NANDN U7903 ( .A(n7409), .B(n7408), .Z(n7413) );
  NANDN U7904 ( .A(n7411), .B(n7410), .Z(n7412) );
  AND U7905 ( .A(n7413), .B(n7412), .Z(n7534) );
  OR U7906 ( .A(n7415), .B(n7414), .Z(n7419) );
  NANDN U7907 ( .A(n7417), .B(n7416), .Z(n7418) );
  AND U7908 ( .A(n7419), .B(n7418), .Z(n7535) );
  XOR U7909 ( .A(n7534), .B(n7535), .Z(n7536) );
  NANDN U7910 ( .A(n7421), .B(n7420), .Z(n7425) );
  NAND U7911 ( .A(n7423), .B(n7422), .Z(n7424) );
  AND U7912 ( .A(n7425), .B(n7424), .Z(n7537) );
  XNOR U7913 ( .A(n7536), .B(n7537), .Z(n7522) );
  NANDN U7914 ( .A(n7427), .B(n7426), .Z(n7431) );
  NAND U7915 ( .A(n7429), .B(n7428), .Z(n7430) );
  NAND U7916 ( .A(n7431), .B(n7430), .Z(n7523) );
  XNOR U7917 ( .A(n7522), .B(n7523), .Z(n7525) );
  NANDN U7918 ( .A(n7433), .B(n7432), .Z(n7437) );
  NANDN U7919 ( .A(n7435), .B(n7434), .Z(n7436) );
  NAND U7920 ( .A(n7437), .B(n7436), .Z(n7623) );
  OR U7921 ( .A(n7438), .B(n7801), .Z(n7442) );
  OR U7922 ( .A(n7440), .B(n7439), .Z(n7441) );
  AND U7923 ( .A(n7442), .B(n7441), .Z(n7640) );
  OR U7924 ( .A(n7444), .B(n7443), .Z(n7448) );
  OR U7925 ( .A(n7446), .B(n7445), .Z(n7447) );
  NAND U7926 ( .A(n7448), .B(n7447), .Z(n7617) );
  NAND U7927 ( .A(x[132]), .B(y[722]), .Z(n7567) );
  AND U7928 ( .A(x[140]), .B(y[714]), .Z(n7450) );
  AND U7929 ( .A(y[708]), .B(x[146]), .Z(n7449) );
  XNOR U7930 ( .A(n7450), .B(n7449), .Z(n7566) );
  XOR U7931 ( .A(n7567), .B(n7566), .Z(n7614) );
  NAND U7932 ( .A(x[144]), .B(y[710]), .Z(n7543) );
  NAND U7933 ( .A(x[145]), .B(y[709]), .Z(n7541) );
  NAND U7934 ( .A(x[133]), .B(y[721]), .Z(n7540) );
  XNOR U7935 ( .A(n7541), .B(n7540), .Z(n7542) );
  XNOR U7936 ( .A(n7543), .B(n7542), .Z(n7615) );
  XNOR U7937 ( .A(n7617), .B(n7616), .Z(n7638) );
  OR U7938 ( .A(n7452), .B(n7451), .Z(n7456) );
  NANDN U7939 ( .A(n7454), .B(n7453), .Z(n7455) );
  NAND U7940 ( .A(n7456), .B(n7455), .Z(n7639) );
  XNOR U7941 ( .A(n7638), .B(n7639), .Z(n7641) );
  XOR U7942 ( .A(n7640), .B(n7641), .Z(n7621) );
  NANDN U7943 ( .A(n7458), .B(n7457), .Z(n7462) );
  OR U7944 ( .A(n7460), .B(n7459), .Z(n7461) );
  NAND U7945 ( .A(n7462), .B(n7461), .Z(n7627) );
  AND U7946 ( .A(x[135]), .B(y[719]), .Z(n7466) );
  XNOR U7947 ( .A(n7467), .B(n7466), .Z(n7562) );
  XOR U7948 ( .A(n7561), .B(n7562), .Z(n7583) );
  NAND U7949 ( .A(x[128]), .B(y[726]), .Z(n7571) );
  AND U7950 ( .A(y[704]), .B(x[150]), .Z(n7570) );
  XNOR U7951 ( .A(n7571), .B(n7570), .Z(n7573) );
  NAND U7952 ( .A(x[149]), .B(y[705]), .Z(n7546) );
  XNOR U7953 ( .A(n7546), .B(o[86]), .Z(n7572) );
  XNOR U7954 ( .A(n7573), .B(n7572), .Z(n7582) );
  XOR U7955 ( .A(n7583), .B(n7582), .Z(n7584) );
  XNOR U7956 ( .A(n7585), .B(n7584), .Z(n7597) );
  OR U7957 ( .A(n7469), .B(n7468), .Z(n7473) );
  OR U7958 ( .A(n7471), .B(n7470), .Z(n7472) );
  AND U7959 ( .A(n7473), .B(n7472), .Z(n7594) );
  NANDN U7960 ( .A(n7475), .B(n7474), .Z(n7479) );
  OR U7961 ( .A(n7477), .B(n7476), .Z(n7478) );
  AND U7962 ( .A(n7479), .B(n7478), .Z(n7595) );
  XOR U7963 ( .A(n7594), .B(n7595), .Z(n7596) );
  XOR U7964 ( .A(n7597), .B(n7596), .Z(n7635) );
  NAND U7965 ( .A(x[147]), .B(y[707]), .Z(n7611) );
  NAND U7966 ( .A(x[131]), .B(y[723]), .Z(n7609) );
  NAND U7967 ( .A(x[142]), .B(y[712]), .Z(n7608) );
  XNOR U7968 ( .A(n7609), .B(n7608), .Z(n7610) );
  XNOR U7969 ( .A(n7611), .B(n7610), .Z(n7589) );
  NAND U7970 ( .A(o[85]), .B(n7480), .Z(n7605) );
  AND U7971 ( .A(y[725]), .B(x[129]), .Z(n7602) );
  XNOR U7972 ( .A(n7603), .B(n7602), .Z(n7604) );
  XOR U7973 ( .A(n7605), .B(n7604), .Z(n7588) );
  XOR U7974 ( .A(n7589), .B(n7588), .Z(n7591) );
  ANDN U7975 ( .B(y[722]), .A(n164), .Z(n8945) );
  NAND U7976 ( .A(n7481), .B(n8945), .Z(n7485) );
  OR U7977 ( .A(n7483), .B(n7482), .Z(n7484) );
  AND U7978 ( .A(n7485), .B(n7484), .Z(n7590) );
  XOR U7979 ( .A(n7591), .B(n7590), .Z(n7632) );
  NAND U7980 ( .A(x[141]), .B(y[713]), .Z(n7556) );
  NAND U7981 ( .A(x[130]), .B(y[724]), .Z(n7554) );
  NAND U7982 ( .A(x[148]), .B(y[706]), .Z(n7553) );
  XNOR U7983 ( .A(n7554), .B(n7553), .Z(n7555) );
  XNOR U7984 ( .A(n7556), .B(n7555), .Z(n7579) );
  NAND U7985 ( .A(x[138]), .B(y[716]), .Z(n7548) );
  AND U7986 ( .A(y[720]), .B(x[134]), .Z(n7547) );
  XOR U7987 ( .A(n7548), .B(n7547), .Z(n7550) );
  AND U7988 ( .A(y[711]), .B(x[143]), .Z(n7549) );
  XOR U7989 ( .A(n7550), .B(n7549), .Z(n7577) );
  NAND U7990 ( .A(n7487), .B(n7486), .Z(n7491) );
  NAND U7991 ( .A(n7489), .B(n7488), .Z(n7490) );
  AND U7992 ( .A(n7491), .B(n7490), .Z(n7576) );
  XNOR U7993 ( .A(n7577), .B(n7576), .Z(n7578) );
  XOR U7994 ( .A(n7579), .B(n7578), .Z(n7633) );
  XNOR U7995 ( .A(n7632), .B(n7633), .Z(n7634) );
  XNOR U7996 ( .A(n7635), .B(n7634), .Z(n7626) );
  XNOR U7997 ( .A(n7627), .B(n7626), .Z(n7629) );
  OR U7998 ( .A(n7493), .B(n7492), .Z(n7497) );
  OR U7999 ( .A(n7495), .B(n7494), .Z(n7496) );
  AND U8000 ( .A(n7497), .B(n7496), .Z(n7628) );
  XNOR U8001 ( .A(n7629), .B(n7628), .Z(n7620) );
  XOR U8002 ( .A(n7621), .B(n7620), .Z(n7622) );
  XOR U8003 ( .A(n7623), .B(n7622), .Z(n7524) );
  XNOR U8004 ( .A(n7525), .B(n7524), .Z(n7530) );
  NANDN U8005 ( .A(n7499), .B(n7498), .Z(n7503) );
  NANDN U8006 ( .A(n7501), .B(n7500), .Z(n7502) );
  AND U8007 ( .A(n7503), .B(n7502), .Z(n7528) );
  OR U8008 ( .A(n7505), .B(n7504), .Z(n7509) );
  NANDN U8009 ( .A(n7507), .B(n7506), .Z(n7508) );
  NAND U8010 ( .A(n7509), .B(n7508), .Z(n7529) );
  XOR U8011 ( .A(n7528), .B(n7529), .Z(n7531) );
  XNOR U8012 ( .A(n7530), .B(n7531), .Z(n7517) );
  XOR U8013 ( .A(n7519), .B(n7518), .Z(n7513) );
  XOR U8014 ( .A(n7512), .B(n7513), .Z(N183) );
  NANDN U8015 ( .A(n7511), .B(n7510), .Z(n7515) );
  NANDN U8016 ( .A(n7513), .B(n7512), .Z(n7514) );
  NAND U8017 ( .A(n7515), .B(n7514), .Z(n7644) );
  NANDN U8018 ( .A(n7517), .B(n7516), .Z(n7521) );
  NAND U8019 ( .A(n7519), .B(n7518), .Z(n7520) );
  NAND U8020 ( .A(n7521), .B(n7520), .Z(n7645) );
  XNOR U8021 ( .A(n7644), .B(n7645), .Z(n7646) );
  OR U8022 ( .A(n7523), .B(n7522), .Z(n7527) );
  OR U8023 ( .A(n7525), .B(n7524), .Z(n7526) );
  AND U8024 ( .A(n7527), .B(n7526), .Z(n7650) );
  OR U8025 ( .A(n7529), .B(n7528), .Z(n7533) );
  NAND U8026 ( .A(n7531), .B(n7530), .Z(n7532) );
  NAND U8027 ( .A(n7533), .B(n7532), .Z(n7651) );
  XOR U8028 ( .A(n7650), .B(n7651), .Z(n7653) );
  OR U8029 ( .A(n7535), .B(n7534), .Z(n7539) );
  NANDN U8030 ( .A(n7537), .B(n7536), .Z(n7538) );
  AND U8031 ( .A(n7539), .B(n7538), .Z(n7779) );
  OR U8032 ( .A(n7541), .B(n7540), .Z(n7545) );
  OR U8033 ( .A(n7543), .B(n7542), .Z(n7544) );
  AND U8034 ( .A(n7545), .B(n7544), .Z(n7668) );
  NANDN U8035 ( .A(n7546), .B(o[86]), .Z(n7751) );
  NAND U8036 ( .A(x[129]), .B(y[726]), .Z(n7749) );
  NAND U8037 ( .A(x[140]), .B(y[715]), .Z(n7748) );
  XNOR U8038 ( .A(n7749), .B(n7748), .Z(n7750) );
  XNOR U8039 ( .A(n7751), .B(n7750), .Z(n7669) );
  XOR U8040 ( .A(n7668), .B(n7669), .Z(n7670) );
  NAND U8041 ( .A(x[149]), .B(y[706]), .Z(n7701) );
  NAND U8042 ( .A(x[130]), .B(y[725]), .Z(n7699) );
  AND U8043 ( .A(x[141]), .B(y[714]), .Z(n7698) );
  XNOR U8044 ( .A(n7699), .B(n7698), .Z(n7700) );
  XOR U8045 ( .A(n7670), .B(n7671), .Z(n7725) );
  NAND U8046 ( .A(x[132]), .B(y[723]), .Z(n7707) );
  NAND U8047 ( .A(x[131]), .B(y[724]), .Z(n7705) );
  XNOR U8048 ( .A(n7707), .B(n7706), .Z(n7677) );
  NANDN U8049 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U8050 ( .A(n7550), .B(n7549), .Z(n7551) );
  AND U8051 ( .A(n7552), .B(n7551), .Z(n7675) );
  ANDN U8052 ( .B(y[710]), .A(n168), .Z(n7818) );
  NAND U8053 ( .A(x[146]), .B(y[709]), .Z(n7711) );
  AND U8054 ( .A(x[133]), .B(y[722]), .Z(n7710) );
  XNOR U8055 ( .A(n7711), .B(n7710), .Z(n7712) );
  XOR U8056 ( .A(n7818), .B(n7712), .Z(n7674) );
  XOR U8057 ( .A(n7675), .B(n7674), .Z(n7676) );
  XNOR U8058 ( .A(n7677), .B(n7676), .Z(n7723) );
  OR U8059 ( .A(n7554), .B(n7553), .Z(n7558) );
  OR U8060 ( .A(n7556), .B(n7555), .Z(n7557) );
  NAND U8061 ( .A(n7558), .B(n7557), .Z(n7724) );
  XOR U8062 ( .A(n7723), .B(n7724), .Z(n7726) );
  XNOR U8063 ( .A(n7725), .B(n7726), .Z(n7762) );
  AND U8064 ( .A(y[705]), .B(x[150]), .Z(n7758) );
  XNOR U8065 ( .A(o[87]), .B(n7758), .Z(n7732) );
  NAND U8066 ( .A(x[128]), .B(y[727]), .Z(n7730) );
  NAND U8067 ( .A(x[151]), .B(y[704]), .Z(n7729) );
  XNOR U8068 ( .A(n7730), .B(n7729), .Z(n7731) );
  XOR U8069 ( .A(n7732), .B(n7731), .Z(n7682) );
  ANDN U8070 ( .B(y[708]), .A(n170), .Z(n7992) );
  AND U8071 ( .A(y[707]), .B(x[148]), .Z(n7560) );
  XNOR U8072 ( .A(n7560), .B(n7559), .Z(n7755) );
  XNOR U8073 ( .A(n7992), .B(n7755), .Z(n7680) );
  NAND U8074 ( .A(n7743), .B(n7744), .Z(n7564) );
  NANDN U8075 ( .A(n7562), .B(n7561), .Z(n7563) );
  NAND U8076 ( .A(n7564), .B(n7563), .Z(n7681) );
  XNOR U8077 ( .A(n7680), .B(n7681), .Z(n7683) );
  XOR U8078 ( .A(n7682), .B(n7683), .Z(n7689) );
  NAND U8079 ( .A(n8423), .B(n7565), .Z(n7569) );
  OR U8080 ( .A(n7567), .B(n7566), .Z(n7568) );
  AND U8081 ( .A(n7569), .B(n7568), .Z(n7686) );
  NANDN U8082 ( .A(n7571), .B(n7570), .Z(n7575) );
  NAND U8083 ( .A(n7573), .B(n7572), .Z(n7574) );
  AND U8084 ( .A(n7575), .B(n7574), .Z(n7687) );
  XOR U8085 ( .A(n7686), .B(n7687), .Z(n7688) );
  XOR U8086 ( .A(n7689), .B(n7688), .Z(n7760) );
  OR U8087 ( .A(n7577), .B(n7576), .Z(n7581) );
  OR U8088 ( .A(n7579), .B(n7578), .Z(n7580) );
  AND U8089 ( .A(n7581), .B(n7580), .Z(n7759) );
  XOR U8090 ( .A(n7760), .B(n7759), .Z(n7761) );
  XOR U8091 ( .A(n7762), .B(n7761), .Z(n7778) );
  OR U8092 ( .A(n7583), .B(n7582), .Z(n7587) );
  NANDN U8093 ( .A(n7585), .B(n7584), .Z(n7586) );
  AND U8094 ( .A(n7587), .B(n7586), .Z(n7662) );
  NANDN U8095 ( .A(n7589), .B(n7588), .Z(n7593) );
  OR U8096 ( .A(n7591), .B(n7590), .Z(n7592) );
  AND U8097 ( .A(n7593), .B(n7592), .Z(n7663) );
  XOR U8098 ( .A(n7662), .B(n7663), .Z(n7664) );
  OR U8099 ( .A(n7595), .B(n7594), .Z(n7599) );
  NANDN U8100 ( .A(n7597), .B(n7596), .Z(n7598) );
  NAND U8101 ( .A(n7599), .B(n7598), .Z(n7665) );
  AND U8102 ( .A(y[720]), .B(x[135]), .Z(n7600) );
  XNOR U8103 ( .A(n7601), .B(n7600), .Z(n7745) );
  AND U8104 ( .A(x[138]), .B(y[717]), .Z(n7692) );
  XOR U8105 ( .A(n7693), .B(n7692), .Z(n7695) );
  NAND U8106 ( .A(x[143]), .B(y[712]), .Z(n7738) );
  AND U8107 ( .A(x[134]), .B(y[721]), .Z(n7737) );
  XNOR U8108 ( .A(n7738), .B(n7737), .Z(n7740) );
  XOR U8109 ( .A(n7695), .B(n7694), .Z(n7719) );
  NAND U8110 ( .A(n7603), .B(n7602), .Z(n7607) );
  OR U8111 ( .A(n7605), .B(n7604), .Z(n7606) );
  NAND U8112 ( .A(n7607), .B(n7606), .Z(n7718) );
  OR U8113 ( .A(n7609), .B(n7608), .Z(n7613) );
  OR U8114 ( .A(n7611), .B(n7610), .Z(n7612) );
  NAND U8115 ( .A(n7613), .B(n7612), .Z(n7717) );
  XNOR U8116 ( .A(n7718), .B(n7717), .Z(n7720) );
  XOR U8117 ( .A(n7719), .B(n7720), .Z(n7765) );
  NANDN U8118 ( .A(n7615), .B(n7614), .Z(n7619) );
  NANDN U8119 ( .A(n7617), .B(n7616), .Z(n7618) );
  AND U8120 ( .A(n7619), .B(n7618), .Z(n7766) );
  XOR U8121 ( .A(n7765), .B(n7766), .Z(n7767) );
  XOR U8122 ( .A(n7768), .B(n7767), .Z(n7777) );
  XOR U8123 ( .A(n7778), .B(n7777), .Z(n7780) );
  XNOR U8124 ( .A(n7779), .B(n7780), .Z(n7658) );
  NANDN U8125 ( .A(n7621), .B(n7620), .Z(n7625) );
  OR U8126 ( .A(n7623), .B(n7622), .Z(n7624) );
  NAND U8127 ( .A(n7625), .B(n7624), .Z(n7657) );
  OR U8128 ( .A(n7627), .B(n7626), .Z(n7631) );
  OR U8129 ( .A(n7629), .B(n7628), .Z(n7630) );
  AND U8130 ( .A(n7631), .B(n7630), .Z(n7774) );
  OR U8131 ( .A(n7633), .B(n7632), .Z(n7637) );
  OR U8132 ( .A(n7635), .B(n7634), .Z(n7636) );
  AND U8133 ( .A(n7637), .B(n7636), .Z(n7771) );
  OR U8134 ( .A(n7639), .B(n7638), .Z(n7643) );
  OR U8135 ( .A(n7641), .B(n7640), .Z(n7642) );
  AND U8136 ( .A(n7643), .B(n7642), .Z(n7772) );
  XOR U8137 ( .A(n7771), .B(n7772), .Z(n7773) );
  XOR U8138 ( .A(n7657), .B(n7656), .Z(n7659) );
  XNOR U8139 ( .A(n7653), .B(n7652), .Z(n7647) );
  XOR U8140 ( .A(n7646), .B(n7647), .Z(N184) );
  NANDN U8141 ( .A(n7645), .B(n7644), .Z(n7649) );
  NANDN U8142 ( .A(n7647), .B(n7646), .Z(n7648) );
  NAND U8143 ( .A(n7649), .B(n7648), .Z(n7916) );
  OR U8144 ( .A(n7651), .B(n7650), .Z(n7655) );
  NAND U8145 ( .A(n7653), .B(n7652), .Z(n7654) );
  AND U8146 ( .A(n7655), .B(n7654), .Z(n7917) );
  XNOR U8147 ( .A(n7916), .B(n7917), .Z(n7918) );
  OR U8148 ( .A(n7657), .B(n7656), .Z(n7661) );
  NAND U8149 ( .A(n7659), .B(n7658), .Z(n7660) );
  AND U8150 ( .A(n7661), .B(n7660), .Z(n7922) );
  OR U8151 ( .A(n7663), .B(n7662), .Z(n7667) );
  NANDN U8152 ( .A(n7665), .B(n7664), .Z(n7666) );
  NAND U8153 ( .A(n7667), .B(n7666), .Z(n7911) );
  OR U8154 ( .A(n7669), .B(n7668), .Z(n7673) );
  NANDN U8155 ( .A(n7671), .B(n7670), .Z(n7672) );
  AND U8156 ( .A(n7673), .B(n7672), .Z(n7898) );
  NANDN U8157 ( .A(n7675), .B(n7674), .Z(n7679) );
  OR U8158 ( .A(n7677), .B(n7676), .Z(n7678) );
  NAND U8159 ( .A(n7679), .B(n7678), .Z(n7851) );
  OR U8160 ( .A(n7681), .B(n7680), .Z(n7685) );
  OR U8161 ( .A(n7683), .B(n7682), .Z(n7684) );
  AND U8162 ( .A(n7685), .B(n7684), .Z(n7848) );
  OR U8163 ( .A(n7687), .B(n7686), .Z(n7691) );
  NANDN U8164 ( .A(n7689), .B(n7688), .Z(n7690) );
  NAND U8165 ( .A(n7691), .B(n7690), .Z(n7849) );
  XOR U8166 ( .A(n7848), .B(n7849), .Z(n7850) );
  XNOR U8167 ( .A(n7851), .B(n7850), .Z(n7899) );
  XOR U8168 ( .A(n7898), .B(n7899), .Z(n7900) );
  NANDN U8169 ( .A(n7693), .B(n7692), .Z(n7697) );
  NANDN U8170 ( .A(n7695), .B(n7694), .Z(n7696) );
  NAND U8171 ( .A(n7697), .B(n7696), .Z(n7843) );
  NANDN U8172 ( .A(n7699), .B(n7698), .Z(n7703) );
  NANDN U8173 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U8174 ( .A(n7703), .B(n7702), .Z(n7886) );
  NANDN U8175 ( .A(n7705), .B(n7704), .Z(n7709) );
  OR U8176 ( .A(n7707), .B(n7706), .Z(n7708) );
  AND U8177 ( .A(n7709), .B(n7708), .Z(n7887) );
  XOR U8178 ( .A(n7886), .B(n7887), .Z(n7888) );
  NAND U8179 ( .A(x[128]), .B(y[728]), .Z(n7831) );
  AND U8180 ( .A(y[704]), .B(x[152]), .Z(n7830) );
  XNOR U8181 ( .A(n7831), .B(n7830), .Z(n7832) );
  ANDN U8182 ( .B(y[705]), .A(n174), .Z(n7823) );
  XNOR U8183 ( .A(o[88]), .B(n7823), .Z(n7833) );
  NANDN U8184 ( .A(n7711), .B(n7710), .Z(n7714) );
  NAND U8185 ( .A(n7712), .B(n7818), .Z(n7713) );
  AND U8186 ( .A(n7714), .B(n7713), .Z(n7869) );
  AND U8187 ( .A(x[146]), .B(y[710]), .Z(n7716) );
  NAND U8188 ( .A(x[145]), .B(y[711]), .Z(n7715) );
  XOR U8189 ( .A(n7716), .B(n7715), .Z(n7820) );
  AND U8190 ( .A(x[135]), .B(y[721]), .Z(n7819) );
  XNOR U8191 ( .A(n7820), .B(n7819), .Z(n7868) );
  XNOR U8192 ( .A(n7871), .B(n7870), .Z(n7889) );
  XOR U8193 ( .A(n7843), .B(n7842), .Z(n7845) );
  OR U8194 ( .A(n7718), .B(n7717), .Z(n7722) );
  NANDN U8195 ( .A(n7720), .B(n7719), .Z(n7721) );
  AND U8196 ( .A(n7722), .B(n7721), .Z(n7844) );
  XOR U8197 ( .A(n7845), .B(n7844), .Z(n7901) );
  XNOR U8198 ( .A(n7911), .B(n7910), .Z(n7913) );
  NANDN U8199 ( .A(n7724), .B(n7723), .Z(n7728) );
  NANDN U8200 ( .A(n7726), .B(n7725), .Z(n7727) );
  NAND U8201 ( .A(n7728), .B(n7727), .Z(n7905) );
  OR U8202 ( .A(n7730), .B(n7729), .Z(n7734) );
  OR U8203 ( .A(n7732), .B(n7731), .Z(n7733) );
  AND U8204 ( .A(n7734), .B(n7733), .Z(n7836) );
  NAND U8205 ( .A(x[143]), .B(y[713]), .Z(n7825) );
  AND U8206 ( .A(y[725]), .B(x[131]), .Z(n7824) );
  XOR U8207 ( .A(n7825), .B(n7824), .Z(n7827) );
  AND U8208 ( .A(x[132]), .B(y[724]), .Z(n7826) );
  XOR U8209 ( .A(n7827), .B(n7826), .Z(n7837) );
  XNOR U8210 ( .A(n7836), .B(n7837), .Z(n7839) );
  AND U8211 ( .A(x[139]), .B(y[717]), .Z(n7736) );
  NAND U8212 ( .A(x[136]), .B(y[720]), .Z(n7735) );
  XOR U8213 ( .A(n7736), .B(n7735), .Z(n7803) );
  ANDN U8214 ( .B(y[714]), .A(n165), .Z(n7802) );
  XNOR U8215 ( .A(n7803), .B(n7802), .Z(n7797) );
  ANDN U8216 ( .B(y[718]), .A(n161), .Z(n7795) );
  ANDN U8217 ( .B(y[719]), .A(n160), .Z(n7796) );
  XNOR U8218 ( .A(n7795), .B(n7796), .Z(n7798) );
  XNOR U8219 ( .A(n7797), .B(n7798), .Z(n7838) );
  XOR U8220 ( .A(n7839), .B(n7838), .Z(n7792) );
  NAND U8221 ( .A(x[134]), .B(y[722]), .Z(n7863) );
  AND U8222 ( .A(y[709]), .B(x[147]), .Z(n7862) );
  XOR U8223 ( .A(n7863), .B(n7862), .Z(n7865) );
  AND U8224 ( .A(y[708]), .B(x[148]), .Z(n7864) );
  XOR U8225 ( .A(n7865), .B(n7864), .Z(n7875) );
  NAND U8226 ( .A(x[149]), .B(y[707]), .Z(n7855) );
  AND U8227 ( .A(y[723]), .B(x[133]), .Z(n7854) );
  XNOR U8228 ( .A(n7855), .B(n7854), .Z(n7856) );
  NAND U8229 ( .A(x[144]), .B(y[712]), .Z(n7857) );
  XOR U8230 ( .A(n7875), .B(n7874), .Z(n7877) );
  NANDN U8231 ( .A(n7738), .B(n7737), .Z(n7742) );
  NAND U8232 ( .A(n7740), .B(n7739), .Z(n7741) );
  AND U8233 ( .A(n7742), .B(n7741), .Z(n7876) );
  XOR U8234 ( .A(n7877), .B(n7876), .Z(n7892) );
  NAND U8235 ( .A(n7743), .B(n7963), .Z(n7747) );
  NANDN U8236 ( .A(n7745), .B(n7744), .Z(n7746) );
  AND U8237 ( .A(n7747), .B(n7746), .Z(n7893) );
  OR U8238 ( .A(n7749), .B(n7748), .Z(n7753) );
  OR U8239 ( .A(n7751), .B(n7750), .Z(n7752) );
  AND U8240 ( .A(n7753), .B(n7752), .Z(n7894) );
  XNOR U8241 ( .A(n7895), .B(n7894), .Z(n7790) );
  AND U8242 ( .A(y[707]), .B(x[144]), .Z(n7754) );
  AND U8243 ( .A(y[711]), .B(x[148]), .Z(n8278) );
  NAND U8244 ( .A(n7754), .B(n8278), .Z(n7757) );
  NANDN U8245 ( .A(n7755), .B(n7992), .Z(n7756) );
  AND U8246 ( .A(n7757), .B(n7756), .Z(n7881) );
  NAND U8247 ( .A(n7758), .B(o[87]), .Z(n7809) );
  AND U8248 ( .A(y[727]), .B(x[129]), .Z(n7806) );
  XOR U8249 ( .A(n7807), .B(n7806), .Z(n7808) );
  XNOR U8250 ( .A(n7809), .B(n7808), .Z(n7880) );
  NAND U8251 ( .A(x[150]), .B(y[706]), .Z(n7813) );
  AND U8252 ( .A(y[726]), .B(x[130]), .Z(n7812) );
  XNOR U8253 ( .A(n7813), .B(n7812), .Z(n7815) );
  XOR U8254 ( .A(n7883), .B(n7882), .Z(n7789) );
  XNOR U8255 ( .A(n7790), .B(n7789), .Z(n7791) );
  XNOR U8256 ( .A(n7792), .B(n7791), .Z(n7904) );
  XNOR U8257 ( .A(n7905), .B(n7904), .Z(n7907) );
  OR U8258 ( .A(n7760), .B(n7759), .Z(n7764) );
  NANDN U8259 ( .A(n7762), .B(n7761), .Z(n7763) );
  AND U8260 ( .A(n7764), .B(n7763), .Z(n7906) );
  XOR U8261 ( .A(n7907), .B(n7906), .Z(n7912) );
  XNOR U8262 ( .A(n7913), .B(n7912), .Z(n7923) );
  XOR U8263 ( .A(n7922), .B(n7923), .Z(n7925) );
  NANDN U8264 ( .A(n7766), .B(n7765), .Z(n7770) );
  OR U8265 ( .A(n7768), .B(n7767), .Z(n7769) );
  NAND U8266 ( .A(n7770), .B(n7769), .Z(n7784) );
  OR U8267 ( .A(n7772), .B(n7771), .Z(n7776) );
  NANDN U8268 ( .A(n7774), .B(n7773), .Z(n7775) );
  AND U8269 ( .A(n7776), .B(n7775), .Z(n7783) );
  XOR U8270 ( .A(n7784), .B(n7783), .Z(n7785) );
  NANDN U8271 ( .A(n7778), .B(n7777), .Z(n7782) );
  OR U8272 ( .A(n7780), .B(n7779), .Z(n7781) );
  NAND U8273 ( .A(n7782), .B(n7781), .Z(n7786) );
  XNOR U8274 ( .A(n7925), .B(n7924), .Z(n7919) );
  XOR U8275 ( .A(n7918), .B(n7919), .Z(N185) );
  OR U8276 ( .A(n7784), .B(n7783), .Z(n7788) );
  NANDN U8277 ( .A(n7786), .B(n7785), .Z(n7787) );
  AND U8278 ( .A(n7788), .B(n7787), .Z(n7936) );
  OR U8279 ( .A(n7790), .B(n7789), .Z(n7794) );
  OR U8280 ( .A(n7792), .B(n7791), .Z(n7793) );
  NAND U8281 ( .A(n7794), .B(n7793), .Z(n8061) );
  OR U8282 ( .A(n7796), .B(n7795), .Z(n7800) );
  OR U8283 ( .A(n7798), .B(n7797), .Z(n7799) );
  NAND U8284 ( .A(n7800), .B(n7799), .Z(n7975) );
  AND U8285 ( .A(y[720]), .B(x[139]), .Z(n8330) );
  NAND U8286 ( .A(n7801), .B(n8330), .Z(n7805) );
  NANDN U8287 ( .A(n7803), .B(n7802), .Z(n7804) );
  AND U8288 ( .A(n7805), .B(n7804), .Z(n8027) );
  NAND U8289 ( .A(y[718]), .B(x[139]), .Z(n8001) );
  AND U8290 ( .A(x[140]), .B(y[717]), .Z(n7998) );
  AND U8291 ( .A(x[135]), .B(y[722]), .Z(n7999) );
  XNOR U8292 ( .A(n7998), .B(n7999), .Z(n8000) );
  XOR U8293 ( .A(n8001), .B(n8000), .Z(n8024) );
  NAND U8294 ( .A(x[141]), .B(y[716]), .Z(n8019) );
  AND U8295 ( .A(y[728]), .B(x[129]), .Z(n8018) );
  XNOR U8296 ( .A(n8019), .B(n8018), .Z(n8020) );
  ANDN U8297 ( .B(y[705]), .A(n175), .Z(n7997) );
  XNOR U8298 ( .A(o[89]), .B(n7997), .Z(n8021) );
  XNOR U8299 ( .A(n8027), .B(n8026), .Z(n7974) );
  XNOR U8300 ( .A(n7975), .B(n7974), .Z(n7977) );
  NAND U8301 ( .A(n7807), .B(n7806), .Z(n7811) );
  NANDN U8302 ( .A(n7809), .B(n7808), .Z(n7810) );
  AND U8303 ( .A(n7811), .B(n7810), .Z(n7949) );
  NANDN U8304 ( .A(n7813), .B(n7812), .Z(n7817) );
  NAND U8305 ( .A(n7815), .B(n7814), .Z(n7816) );
  AND U8306 ( .A(n7817), .B(n7816), .Z(n7946) );
  AND U8307 ( .A(y[711]), .B(x[146]), .Z(n7986) );
  NAND U8308 ( .A(n7986), .B(n7818), .Z(n7822) );
  NANDN U8309 ( .A(n7820), .B(n7819), .Z(n7821) );
  AND U8310 ( .A(n7822), .B(n7821), .Z(n7954) );
  NAND U8311 ( .A(y[721]), .B(x[136]), .Z(n7965) );
  XOR U8312 ( .A(n7965), .B(n7964), .Z(n7952) );
  AND U8313 ( .A(n7823), .B(o[88]), .Z(n7961) );
  AND U8314 ( .A(y[704]), .B(x[153]), .Z(n7958) );
  AND U8315 ( .A(y[729]), .B(x[128]), .Z(n7959) );
  XNOR U8316 ( .A(n7958), .B(n7959), .Z(n7960) );
  XOR U8317 ( .A(n7961), .B(n7960), .Z(n7953) );
  XNOR U8318 ( .A(n7952), .B(n7953), .Z(n7955) );
  XNOR U8319 ( .A(n7954), .B(n7955), .Z(n7947) );
  XNOR U8320 ( .A(n7946), .B(n7947), .Z(n7948) );
  XNOR U8321 ( .A(n7949), .B(n7948), .Z(n7976) );
  XNOR U8322 ( .A(n7977), .B(n7976), .Z(n8056) );
  NANDN U8323 ( .A(n7825), .B(n7824), .Z(n7829) );
  NANDN U8324 ( .A(n7827), .B(n7826), .Z(n7828) );
  AND U8325 ( .A(n7829), .B(n7828), .Z(n8032) );
  NANDN U8326 ( .A(n7831), .B(n7830), .Z(n7835) );
  NANDN U8327 ( .A(n7833), .B(n7832), .Z(n7834) );
  AND U8328 ( .A(n7835), .B(n7834), .Z(n8030) );
  AND U8329 ( .A(y[726]), .B(x[131]), .Z(n8012) );
  XOR U8330 ( .A(n8013), .B(n8012), .Z(n8015) );
  AND U8331 ( .A(y[727]), .B(x[130]), .Z(n8014) );
  XNOR U8332 ( .A(n8015), .B(n8014), .Z(n8031) );
  XNOR U8333 ( .A(n8030), .B(n8031), .Z(n8033) );
  XNOR U8334 ( .A(n8032), .B(n8033), .Z(n8054) );
  OR U8335 ( .A(n7837), .B(n7836), .Z(n7841) );
  NANDN U8336 ( .A(n7839), .B(n7838), .Z(n7840) );
  NAND U8337 ( .A(n7841), .B(n7840), .Z(n8055) );
  XOR U8338 ( .A(n8054), .B(n8055), .Z(n8057) );
  XNOR U8339 ( .A(n8056), .B(n8057), .Z(n8060) );
  XOR U8340 ( .A(n8061), .B(n8060), .Z(n8063) );
  NANDN U8341 ( .A(n7843), .B(n7842), .Z(n7847) );
  OR U8342 ( .A(n7845), .B(n7844), .Z(n7846) );
  AND U8343 ( .A(n7847), .B(n7846), .Z(n8062) );
  XOR U8344 ( .A(n8063), .B(n8062), .Z(n7941) );
  OR U8345 ( .A(n7849), .B(n7848), .Z(n7853) );
  NANDN U8346 ( .A(n7851), .B(n7850), .Z(n7852) );
  NAND U8347 ( .A(n7853), .B(n7852), .Z(n8067) );
  NANDN U8348 ( .A(n7855), .B(n7854), .Z(n7859) );
  NANDN U8349 ( .A(n7857), .B(n7856), .Z(n7858) );
  AND U8350 ( .A(n7859), .B(n7858), .Z(n8044) );
  NAND U8351 ( .A(y[707]), .B(x[150]), .Z(n8004) );
  AND U8352 ( .A(x[133]), .B(y[724]), .Z(n8002) );
  AND U8353 ( .A(x[145]), .B(y[712]), .Z(n8003) );
  XOR U8354 ( .A(n8002), .B(n8003), .Z(n8005) );
  XNOR U8355 ( .A(n8004), .B(n8005), .Z(n8042) );
  AND U8356 ( .A(x[147]), .B(y[710]), .Z(n7861) );
  NAND U8357 ( .A(x[149]), .B(y[708]), .Z(n7860) );
  XOR U8358 ( .A(n7861), .B(n7860), .Z(n7994) );
  AND U8359 ( .A(y[709]), .B(x[148]), .Z(n7993) );
  XOR U8360 ( .A(n7994), .B(n7993), .Z(n8043) );
  XOR U8361 ( .A(n8042), .B(n8043), .Z(n8045) );
  XOR U8362 ( .A(n8044), .B(n8045), .Z(n7968) );
  NAND U8363 ( .A(x[151]), .B(y[706]), .Z(n8011) );
  AND U8364 ( .A(y[725]), .B(x[132]), .Z(n8008) );
  AND U8365 ( .A(x[144]), .B(y[713]), .Z(n8009) );
  XNOR U8366 ( .A(n8008), .B(n8009), .Z(n8010) );
  XOR U8367 ( .A(n8011), .B(n8010), .Z(n8038) );
  NAND U8368 ( .A(y[714]), .B(x[143]), .Z(n7989) );
  AND U8369 ( .A(y[723]), .B(x[134]), .Z(n7987) );
  XOR U8370 ( .A(n7989), .B(n7988), .Z(n8036) );
  NANDN U8371 ( .A(n7863), .B(n7862), .Z(n7867) );
  NANDN U8372 ( .A(n7865), .B(n7864), .Z(n7866) );
  AND U8373 ( .A(n7867), .B(n7866), .Z(n8037) );
  XOR U8374 ( .A(n8036), .B(n8037), .Z(n8039) );
  XOR U8375 ( .A(n8038), .B(n8039), .Z(n7969) );
  XNOR U8376 ( .A(n7968), .B(n7969), .Z(n7971) );
  NANDN U8377 ( .A(n7869), .B(n7868), .Z(n7873) );
  OR U8378 ( .A(n7871), .B(n7870), .Z(n7872) );
  NAND U8379 ( .A(n7873), .B(n7872), .Z(n7970) );
  XOR U8380 ( .A(n7971), .B(n7970), .Z(n7983) );
  NANDN U8381 ( .A(n7875), .B(n7874), .Z(n7879) );
  OR U8382 ( .A(n7877), .B(n7876), .Z(n7878) );
  AND U8383 ( .A(n7879), .B(n7878), .Z(n7980) );
  NANDN U8384 ( .A(n7881), .B(n7880), .Z(n7885) );
  NANDN U8385 ( .A(n7883), .B(n7882), .Z(n7884) );
  AND U8386 ( .A(n7885), .B(n7884), .Z(n7981) );
  XOR U8387 ( .A(n7980), .B(n7981), .Z(n7982) );
  OR U8388 ( .A(n7887), .B(n7886), .Z(n7891) );
  NANDN U8389 ( .A(n7889), .B(n7888), .Z(n7890) );
  NAND U8390 ( .A(n7891), .B(n7890), .Z(n8049) );
  NANDN U8391 ( .A(n7893), .B(n7892), .Z(n7897) );
  OR U8392 ( .A(n7895), .B(n7894), .Z(n7896) );
  NAND U8393 ( .A(n7897), .B(n7896), .Z(n8048) );
  XOR U8394 ( .A(n8049), .B(n8048), .Z(n8050) );
  XOR U8395 ( .A(n8067), .B(n8066), .Z(n8069) );
  OR U8396 ( .A(n7899), .B(n7898), .Z(n7903) );
  NANDN U8397 ( .A(n7901), .B(n7900), .Z(n7902) );
  AND U8398 ( .A(n7903), .B(n7902), .Z(n8068) );
  XOR U8399 ( .A(n8069), .B(n8068), .Z(n7940) );
  XOR U8400 ( .A(n7941), .B(n7940), .Z(n7943) );
  OR U8401 ( .A(n7905), .B(n7904), .Z(n7909) );
  OR U8402 ( .A(n7907), .B(n7906), .Z(n7908) );
  AND U8403 ( .A(n7909), .B(n7908), .Z(n7942) );
  XOR U8404 ( .A(n7943), .B(n7942), .Z(n7934) );
  OR U8405 ( .A(n7911), .B(n7910), .Z(n7915) );
  OR U8406 ( .A(n7913), .B(n7912), .Z(n7914) );
  AND U8407 ( .A(n7915), .B(n7914), .Z(n7935) );
  XNOR U8408 ( .A(n7934), .B(n7935), .Z(n7937) );
  XOR U8409 ( .A(n7936), .B(n7937), .Z(n7930) );
  NANDN U8410 ( .A(n7917), .B(n7916), .Z(n7921) );
  NANDN U8411 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U8412 ( .A(n7921), .B(n7920), .Z(n7928) );
  OR U8413 ( .A(n7923), .B(n7922), .Z(n7927) );
  NAND U8414 ( .A(n7925), .B(n7924), .Z(n7926) );
  AND U8415 ( .A(n7927), .B(n7926), .Z(n7929) );
  XNOR U8416 ( .A(n7928), .B(n7929), .Z(n7931) );
  XNOR U8417 ( .A(n7930), .B(n7931), .Z(N186) );
  NANDN U8418 ( .A(n7929), .B(n7928), .Z(n7933) );
  NAND U8419 ( .A(n7931), .B(n7930), .Z(n7932) );
  NAND U8420 ( .A(n7933), .B(n7932), .Z(n8072) );
  OR U8421 ( .A(n7935), .B(n7934), .Z(n7939) );
  OR U8422 ( .A(n7937), .B(n7936), .Z(n7938) );
  AND U8423 ( .A(n7939), .B(n7938), .Z(n8073) );
  XNOR U8424 ( .A(n8072), .B(n8073), .Z(n8074) );
  NANDN U8425 ( .A(n7941), .B(n7940), .Z(n7945) );
  OR U8426 ( .A(n7943), .B(n7942), .Z(n7944) );
  NAND U8427 ( .A(n7945), .B(n7944), .Z(n8079) );
  OR U8428 ( .A(n7947), .B(n7946), .Z(n7951) );
  OR U8429 ( .A(n7949), .B(n7948), .Z(n7950) );
  AND U8430 ( .A(n7951), .B(n7950), .Z(n8186) );
  OR U8431 ( .A(n7953), .B(n7952), .Z(n7957) );
  OR U8432 ( .A(n7955), .B(n7954), .Z(n7956) );
  AND U8433 ( .A(n7957), .B(n7956), .Z(n8184) );
  NAND U8434 ( .A(x[130]), .B(y[728]), .Z(n8133) );
  XOR U8435 ( .A(n8133), .B(n8132), .Z(n8135) );
  ANDN U8436 ( .B(y[706]), .A(n175), .Z(n8134) );
  XNOR U8437 ( .A(n8135), .B(n8134), .Z(n8096) );
  XOR U8438 ( .A(n8096), .B(n8097), .Z(n8099) );
  OR U8439 ( .A(n7963), .B(n7962), .Z(n7967) );
  NAND U8440 ( .A(n7965), .B(n7964), .Z(n7966) );
  NAND U8441 ( .A(n7967), .B(n7966), .Z(n8098) );
  XNOR U8442 ( .A(n8099), .B(n8098), .Z(n8185) );
  XNOR U8443 ( .A(n8184), .B(n8185), .Z(n8187) );
  XNOR U8444 ( .A(n8186), .B(n8187), .Z(n8174) );
  OR U8445 ( .A(n7969), .B(n7968), .Z(n7973) );
  OR U8446 ( .A(n7971), .B(n7970), .Z(n7972) );
  AND U8447 ( .A(n7973), .B(n7972), .Z(n8172) );
  OR U8448 ( .A(n7975), .B(n7974), .Z(n7979) );
  OR U8449 ( .A(n7977), .B(n7976), .Z(n7978) );
  NAND U8450 ( .A(n7979), .B(n7978), .Z(n8173) );
  XOR U8451 ( .A(n8172), .B(n8173), .Z(n8175) );
  XNOR U8452 ( .A(n8174), .B(n8175), .Z(n8087) );
  OR U8453 ( .A(n7981), .B(n7980), .Z(n7985) );
  NANDN U8454 ( .A(n7983), .B(n7982), .Z(n7984) );
  AND U8455 ( .A(n7985), .B(n7984), .Z(n8168) );
  ANDN U8456 ( .B(y[726]), .A(n155), .Z(n8139) );
  XNOR U8457 ( .A(n8138), .B(n8139), .Z(n8141) );
  XOR U8458 ( .A(n8140), .B(n8141), .Z(n8144) );
  OR U8459 ( .A(n7987), .B(n7986), .Z(n7991) );
  NAND U8460 ( .A(n7989), .B(n7988), .Z(n7990) );
  NAND U8461 ( .A(n7991), .B(n7990), .Z(n8145) );
  XNOR U8462 ( .A(n8144), .B(n8145), .Z(n8147) );
  NAND U8463 ( .A(x[147]), .B(y[711]), .Z(n8197) );
  AND U8464 ( .A(x[139]), .B(y[719]), .Z(n8196) );
  XNOR U8465 ( .A(n8197), .B(n8196), .Z(n8199) );
  AND U8466 ( .A(y[727]), .B(x[131]), .Z(n8198) );
  XOR U8467 ( .A(n8147), .B(n8146), .Z(n8120) );
  NOR U8468 ( .A(n172), .B(n148), .Z(n8269) );
  NAND U8469 ( .A(n8269), .B(n7992), .Z(n7996) );
  NANDN U8470 ( .A(n7994), .B(n7993), .Z(n7995) );
  NAND U8471 ( .A(n7996), .B(n7995), .Z(n8155) );
  NAND U8472 ( .A(x[150]), .B(y[708]), .Z(n8129) );
  NAND U8473 ( .A(y[707]), .B(x[151]), .Z(n8126) );
  XNOR U8474 ( .A(n8127), .B(n8126), .Z(n8128) );
  XNOR U8475 ( .A(n8129), .B(n8128), .Z(n8154) );
  XNOR U8476 ( .A(n8155), .B(n8154), .Z(n8157) );
  NAND U8477 ( .A(y[710]), .B(x[148]), .Z(n8211) );
  NAND U8478 ( .A(x[149]), .B(y[709]), .Z(n8208) );
  XNOR U8479 ( .A(n8209), .B(n8208), .Z(n8210) );
  XNOR U8480 ( .A(n8211), .B(n8210), .Z(n8156) );
  XNOR U8481 ( .A(n8157), .B(n8156), .Z(n8121) );
  XOR U8482 ( .A(n8120), .B(n8121), .Z(n8122) );
  AND U8483 ( .A(n7997), .B(o[89]), .Z(n8204) );
  ANDN U8484 ( .B(y[716]), .A(n165), .Z(n8202) );
  ANDN U8485 ( .B(y[729]), .A(n152), .Z(n8203) );
  XNOR U8486 ( .A(n8202), .B(n8203), .Z(n8205) );
  XNOR U8487 ( .A(n8204), .B(n8205), .Z(n8102) );
  NAND U8488 ( .A(x[128]), .B(y[730]), .Z(n8115) );
  AND U8489 ( .A(y[704]), .B(x[154]), .Z(n8114) );
  XNOR U8490 ( .A(n8115), .B(n8114), .Z(n8117) );
  NAND U8491 ( .A(x[153]), .B(y[705]), .Z(n8214) );
  XNOR U8492 ( .A(n8214), .B(o[90]), .Z(n8116) );
  XNOR U8493 ( .A(n8117), .B(n8116), .Z(n8103) );
  XOR U8494 ( .A(n8102), .B(n8103), .Z(n8105) );
  XOR U8495 ( .A(n8105), .B(n8104), .Z(n8153) );
  OR U8496 ( .A(n8003), .B(n8002), .Z(n8007) );
  NAND U8497 ( .A(n8005), .B(n8004), .Z(n8006) );
  AND U8498 ( .A(n8007), .B(n8006), .Z(n8150) );
  XOR U8499 ( .A(n8150), .B(n8151), .Z(n8152) );
  XOR U8500 ( .A(n8153), .B(n8152), .Z(n8123) );
  NAND U8501 ( .A(n8013), .B(n8012), .Z(n8017) );
  NAND U8502 ( .A(n8015), .B(n8014), .Z(n8016) );
  NAND U8503 ( .A(n8017), .B(n8016), .Z(n8161) );
  NANDN U8504 ( .A(n8019), .B(n8018), .Z(n8023) );
  NANDN U8505 ( .A(n8021), .B(n8020), .Z(n8022) );
  NAND U8506 ( .A(n8023), .B(n8022), .Z(n8160) );
  XOR U8507 ( .A(n8161), .B(n8160), .Z(n8162) );
  IV U8508 ( .A(y[721]), .Z(n8482) );
  NANDN U8509 ( .A(n8482), .B(x[137]), .Z(n8217) );
  IV U8510 ( .A(y[724]), .Z(n8445) );
  NANDN U8511 ( .A(n8445), .B(x[134]), .Z(n8215) );
  XNOR U8512 ( .A(n8215), .B(n8216), .Z(n8218) );
  XOR U8513 ( .A(n8217), .B(n8218), .Z(n8193) );
  NAND U8514 ( .A(x[135]), .B(y[723]), .Z(n8190) );
  NAND U8515 ( .A(x[138]), .B(y[720]), .Z(n8111) );
  AND U8516 ( .A(x[140]), .B(y[718]), .Z(n8108) );
  AND U8517 ( .A(y[725]), .B(x[133]), .Z(n8109) );
  XOR U8518 ( .A(n8108), .B(n8109), .Z(n8110) );
  XNOR U8519 ( .A(n8111), .B(n8110), .Z(n8191) );
  XNOR U8520 ( .A(n8190), .B(n8191), .Z(n8192) );
  XOR U8521 ( .A(n8193), .B(n8192), .Z(n8163) );
  NANDN U8522 ( .A(n8025), .B(n8024), .Z(n8029) );
  OR U8523 ( .A(n8027), .B(n8026), .Z(n8028) );
  AND U8524 ( .A(n8029), .B(n8028), .Z(n8091) );
  XOR U8525 ( .A(n8090), .B(n8091), .Z(n8092) );
  OR U8526 ( .A(n8031), .B(n8030), .Z(n8035) );
  OR U8527 ( .A(n8033), .B(n8032), .Z(n8034) );
  NAND U8528 ( .A(n8035), .B(n8034), .Z(n8181) );
  OR U8529 ( .A(n8037), .B(n8036), .Z(n8041) );
  NAND U8530 ( .A(n8039), .B(n8038), .Z(n8040) );
  NAND U8531 ( .A(n8041), .B(n8040), .Z(n8179) );
  NANDN U8532 ( .A(n8043), .B(n8042), .Z(n8047) );
  OR U8533 ( .A(n8045), .B(n8044), .Z(n8046) );
  NAND U8534 ( .A(n8047), .B(n8046), .Z(n8178) );
  XNOR U8535 ( .A(n8179), .B(n8178), .Z(n8180) );
  XOR U8536 ( .A(n8181), .B(n8180), .Z(n8166) );
  XNOR U8537 ( .A(n8167), .B(n8166), .Z(n8169) );
  XOR U8538 ( .A(n8168), .B(n8169), .Z(n8085) );
  OR U8539 ( .A(n8049), .B(n8048), .Z(n8053) );
  NANDN U8540 ( .A(n8051), .B(n8050), .Z(n8052) );
  AND U8541 ( .A(n8053), .B(n8052), .Z(n8084) );
  XNOR U8542 ( .A(n8085), .B(n8084), .Z(n8086) );
  XNOR U8543 ( .A(n8087), .B(n8086), .Z(n8224) );
  NANDN U8544 ( .A(n8055), .B(n8054), .Z(n8059) );
  NANDN U8545 ( .A(n8057), .B(n8056), .Z(n8058) );
  AND U8546 ( .A(n8059), .B(n8058), .Z(n8221) );
  NANDN U8547 ( .A(n8061), .B(n8060), .Z(n8065) );
  OR U8548 ( .A(n8063), .B(n8062), .Z(n8064) );
  AND U8549 ( .A(n8065), .B(n8064), .Z(n8222) );
  XOR U8550 ( .A(n8221), .B(n8222), .Z(n8223) );
  XOR U8551 ( .A(n8079), .B(n8078), .Z(n8081) );
  NANDN U8552 ( .A(n8067), .B(n8066), .Z(n8071) );
  OR U8553 ( .A(n8069), .B(n8068), .Z(n8070) );
  NAND U8554 ( .A(n8071), .B(n8070), .Z(n8080) );
  XOR U8555 ( .A(n8081), .B(n8080), .Z(n8075) );
  XNOR U8556 ( .A(n8074), .B(n8075), .Z(N187) );
  NANDN U8557 ( .A(n8073), .B(n8072), .Z(n8077) );
  NAND U8558 ( .A(n8075), .B(n8074), .Z(n8076) );
  NAND U8559 ( .A(n8077), .B(n8076), .Z(n8227) );
  NANDN U8560 ( .A(n8079), .B(n8078), .Z(n8083) );
  OR U8561 ( .A(n8081), .B(n8080), .Z(n8082) );
  AND U8562 ( .A(n8083), .B(n8082), .Z(n8228) );
  XNOR U8563 ( .A(n8227), .B(n8228), .Z(n8229) );
  OR U8564 ( .A(n8085), .B(n8084), .Z(n8089) );
  OR U8565 ( .A(n8087), .B(n8086), .Z(n8088) );
  AND U8566 ( .A(n8089), .B(n8088), .Z(n8233) );
  OR U8567 ( .A(n8091), .B(n8090), .Z(n8095) );
  NANDN U8568 ( .A(n8093), .B(n8092), .Z(n8094) );
  AND U8569 ( .A(n8095), .B(n8094), .Z(n8248) );
  NANDN U8570 ( .A(n8097), .B(n8096), .Z(n8101) );
  OR U8571 ( .A(n8099), .B(n8098), .Z(n8100) );
  NAND U8572 ( .A(n8101), .B(n8100), .Z(n8360) );
  NANDN U8573 ( .A(n8103), .B(n8102), .Z(n8107) );
  OR U8574 ( .A(n8105), .B(n8104), .Z(n8106) );
  NAND U8575 ( .A(n8107), .B(n8106), .Z(n8358) );
  ANDN U8576 ( .B(y[719]), .A(n163), .Z(n8345) );
  ANDN U8577 ( .B(y[718]), .A(n164), .Z(n8346) );
  XNOR U8578 ( .A(n8345), .B(n8346), .Z(n8348) );
  NAND U8579 ( .A(x[144]), .B(y[715]), .Z(n8327) );
  XOR U8580 ( .A(n8328), .B(n8327), .Z(n8329) );
  XOR U8581 ( .A(n8330), .B(n8329), .Z(n8347) );
  XNOR U8582 ( .A(n8348), .B(n8347), .Z(n8295) );
  ANDN U8583 ( .B(y[728]), .A(n154), .Z(n8353) );
  ANDN U8584 ( .B(y[729]), .A(n153), .Z(n8351) );
  ANDN U8585 ( .B(y[716]), .A(n166), .Z(n8352) );
  XNOR U8586 ( .A(n8351), .B(n8352), .Z(n8354) );
  XOR U8587 ( .A(n8353), .B(n8354), .Z(n8293) );
  NAND U8588 ( .A(x[134]), .B(y[725]), .Z(n8285) );
  ANDN U8589 ( .B(y[706]), .A(n14372), .Z(n8284) );
  NAND U8590 ( .A(y[712]), .B(x[147]), .Z(n8283) );
  XOR U8591 ( .A(n8284), .B(n8283), .Z(n8286) );
  XNOR U8592 ( .A(n8285), .B(n8286), .Z(n8294) );
  XNOR U8593 ( .A(n8293), .B(n8294), .Z(n8296) );
  XNOR U8594 ( .A(n8295), .B(n8296), .Z(n8323) );
  OR U8595 ( .A(n8109), .B(n8108), .Z(n8113) );
  NAND U8596 ( .A(n8111), .B(n8110), .Z(n8112) );
  AND U8597 ( .A(n8113), .B(n8112), .Z(n8321) );
  NANDN U8598 ( .A(n8115), .B(n8114), .Z(n8119) );
  NAND U8599 ( .A(n8117), .B(n8116), .Z(n8118) );
  NAND U8600 ( .A(n8119), .B(n8118), .Z(n8322) );
  XNOR U8601 ( .A(n8321), .B(n8322), .Z(n8324) );
  XOR U8602 ( .A(n8323), .B(n8324), .Z(n8357) );
  XNOR U8603 ( .A(n8358), .B(n8357), .Z(n8359) );
  XOR U8604 ( .A(n8360), .B(n8359), .Z(n8245) );
  OR U8605 ( .A(n8121), .B(n8120), .Z(n8125) );
  NANDN U8606 ( .A(n8123), .B(n8122), .Z(n8124) );
  NAND U8607 ( .A(n8125), .B(n8124), .Z(n8246) );
  XOR U8608 ( .A(n8245), .B(n8246), .Z(n8247) );
  XOR U8609 ( .A(n8248), .B(n8247), .Z(n8382) );
  NANDN U8610 ( .A(n8127), .B(n8126), .Z(n8131) );
  NAND U8611 ( .A(n8129), .B(n8128), .Z(n8130) );
  AND U8612 ( .A(n8131), .B(n8130), .Z(n8315) );
  NANDN U8613 ( .A(n8133), .B(n8132), .Z(n8137) );
  NANDN U8614 ( .A(n8135), .B(n8134), .Z(n8136) );
  NAND U8615 ( .A(n8137), .B(n8136), .Z(n8316) );
  XOR U8616 ( .A(n8315), .B(n8316), .Z(n8317) );
  OR U8617 ( .A(n8139), .B(n8138), .Z(n8143) );
  OR U8618 ( .A(n8141), .B(n8140), .Z(n8142) );
  AND U8619 ( .A(n8143), .B(n8142), .Z(n8309) );
  ANDN U8620 ( .B(y[722]), .A(n160), .Z(n8272) );
  ANDN U8621 ( .B(y[713]), .A(n169), .Z(n8271) );
  XNOR U8622 ( .A(n8269), .B(n8271), .Z(n8273) );
  XNOR U8623 ( .A(n8272), .B(n8273), .Z(n8310) );
  XOR U8624 ( .A(n8309), .B(n8310), .Z(n8311) );
  ANDN U8625 ( .B(y[731]), .A(n151), .Z(n8259) );
  ANDN U8626 ( .B(y[705]), .A(n176), .Z(n8276) );
  XOR U8627 ( .A(o[91]), .B(n8276), .Z(n8257) );
  ANDN U8628 ( .B(y[704]), .A(n177), .Z(n8258) );
  XNOR U8629 ( .A(n8257), .B(n8258), .Z(n8260) );
  XNOR U8630 ( .A(n8259), .B(n8260), .Z(n8312) );
  XOR U8631 ( .A(n8317), .B(n8318), .Z(n8363) );
  OR U8632 ( .A(n8145), .B(n8144), .Z(n8149) );
  OR U8633 ( .A(n8147), .B(n8146), .Z(n8148) );
  AND U8634 ( .A(n8149), .B(n8148), .Z(n8364) );
  XOR U8635 ( .A(n8363), .B(n8364), .Z(n8366) );
  XOR U8636 ( .A(n8366), .B(n8365), .Z(n8251) );
  OR U8637 ( .A(n8155), .B(n8154), .Z(n8159) );
  OR U8638 ( .A(n8157), .B(n8156), .Z(n8158) );
  NAND U8639 ( .A(n8159), .B(n8158), .Z(n8252) );
  XOR U8640 ( .A(n8251), .B(n8252), .Z(n8254) );
  OR U8641 ( .A(n8161), .B(n8160), .Z(n8165) );
  NANDN U8642 ( .A(n8163), .B(n8162), .Z(n8164) );
  NAND U8643 ( .A(n8165), .B(n8164), .Z(n8253) );
  XNOR U8644 ( .A(n8254), .B(n8253), .Z(n8380) );
  OR U8645 ( .A(n8167), .B(n8166), .Z(n8171) );
  OR U8646 ( .A(n8169), .B(n8168), .Z(n8170) );
  AND U8647 ( .A(n8171), .B(n8170), .Z(n8379) );
  XNOR U8648 ( .A(n8380), .B(n8379), .Z(n8381) );
  XNOR U8649 ( .A(n8382), .B(n8381), .Z(n8375) );
  OR U8650 ( .A(n8173), .B(n8172), .Z(n8177) );
  NAND U8651 ( .A(n8175), .B(n8174), .Z(n8176) );
  AND U8652 ( .A(n8177), .B(n8176), .Z(n8373) );
  OR U8653 ( .A(n8179), .B(n8178), .Z(n8183) );
  OR U8654 ( .A(n8181), .B(n8180), .Z(n8182) );
  NAND U8655 ( .A(n8183), .B(n8182), .Z(n8370) );
  OR U8656 ( .A(n8185), .B(n8184), .Z(n8189) );
  OR U8657 ( .A(n8187), .B(n8186), .Z(n8188) );
  AND U8658 ( .A(n8189), .B(n8188), .Z(n8367) );
  NANDN U8659 ( .A(n8191), .B(n8190), .Z(n8195) );
  NANDN U8660 ( .A(n8193), .B(n8192), .Z(n8194) );
  NAND U8661 ( .A(n8195), .B(n8194), .Z(n8241) );
  NANDN U8662 ( .A(n8197), .B(n8196), .Z(n8201) );
  NAND U8663 ( .A(n8199), .B(n8198), .Z(n8200) );
  AND U8664 ( .A(n8201), .B(n8200), .Z(n8301) );
  ANDN U8665 ( .B(y[709]), .A(n173), .Z(n8335) );
  ANDN U8666 ( .B(y[708]), .A(n174), .Z(n8333) );
  ANDN U8667 ( .B(y[723]), .A(n159), .Z(n8334) );
  XNOR U8668 ( .A(n8333), .B(n8334), .Z(n8336) );
  XOR U8669 ( .A(n8335), .B(n8336), .Z(n8299) );
  AND U8670 ( .A(x[135]), .B(y[724]), .Z(n8279) );
  NANDN U8671 ( .A(n147), .B(x[152]), .Z(n8277) );
  XOR U8672 ( .A(n8278), .B(n8277), .Z(n8280) );
  XOR U8673 ( .A(n8279), .B(n8280), .Z(n8300) );
  XOR U8674 ( .A(n8299), .B(n8300), .Z(n8302) );
  XOR U8675 ( .A(n8301), .B(n8302), .Z(n8239) );
  OR U8676 ( .A(n8203), .B(n8202), .Z(n8207) );
  OR U8677 ( .A(n8205), .B(n8204), .Z(n8206) );
  NAND U8678 ( .A(n8207), .B(n8206), .Z(n8290) );
  NANDN U8679 ( .A(n8209), .B(n8208), .Z(n8213) );
  NAND U8680 ( .A(n8211), .B(n8210), .Z(n8212) );
  NAND U8681 ( .A(n8213), .B(n8212), .Z(n8289) );
  XOR U8682 ( .A(n8290), .B(n8289), .Z(n8292) );
  ANDN U8683 ( .B(y[717]), .A(n165), .Z(n8341) );
  ANDN U8684 ( .B(o[90]), .A(n8214), .Z(n8339) );
  ANDN U8685 ( .B(y[730]), .A(n152), .Z(n8340) );
  XNOR U8686 ( .A(n8339), .B(n8340), .Z(n8342) );
  XOR U8687 ( .A(n8341), .B(n8342), .Z(n8304) );
  NAND U8688 ( .A(x[145]), .B(y[714]), .Z(n8264) );
  ANDN U8689 ( .B(y[727]), .A(n155), .Z(n8263) );
  XNOR U8690 ( .A(n8264), .B(n8263), .Z(n8266) );
  ANDN U8691 ( .B(y[726]), .A(n156), .Z(n8265) );
  XOR U8692 ( .A(n8266), .B(n8265), .Z(n8303) );
  XOR U8693 ( .A(n8304), .B(n8303), .Z(n8306) );
  NAND U8694 ( .A(n8216), .B(n8215), .Z(n8220) );
  NANDN U8695 ( .A(n8218), .B(n8217), .Z(n8219) );
  NAND U8696 ( .A(n8220), .B(n8219), .Z(n8305) );
  XOR U8697 ( .A(n8306), .B(n8305), .Z(n8291) );
  XOR U8698 ( .A(n8292), .B(n8291), .Z(n8240) );
  XNOR U8699 ( .A(n8367), .B(n8368), .Z(n8369) );
  XOR U8700 ( .A(n8370), .B(n8369), .Z(n8374) );
  XOR U8701 ( .A(n8373), .B(n8374), .Z(n8376) );
  XNOR U8702 ( .A(n8375), .B(n8376), .Z(n8234) );
  XOR U8703 ( .A(n8233), .B(n8234), .Z(n8235) );
  OR U8704 ( .A(n8222), .B(n8221), .Z(n8226) );
  NANDN U8705 ( .A(n8224), .B(n8223), .Z(n8225) );
  AND U8706 ( .A(n8226), .B(n8225), .Z(n8236) );
  XOR U8707 ( .A(n8229), .B(n8230), .Z(N188) );
  NANDN U8708 ( .A(n8228), .B(n8227), .Z(n8232) );
  NANDN U8709 ( .A(n8230), .B(n8229), .Z(n8231) );
  NAND U8710 ( .A(n8232), .B(n8231), .Z(n8385) );
  OR U8711 ( .A(n8234), .B(n8233), .Z(n8238) );
  NANDN U8712 ( .A(n8236), .B(n8235), .Z(n8237) );
  AND U8713 ( .A(n8238), .B(n8237), .Z(n8386) );
  XNOR U8714 ( .A(n8385), .B(n8386), .Z(n8387) );
  NANDN U8715 ( .A(n8240), .B(n8239), .Z(n8244) );
  NAND U8716 ( .A(n8242), .B(n8241), .Z(n8243) );
  NAND U8717 ( .A(n8244), .B(n8243), .Z(n8549) );
  OR U8718 ( .A(n8246), .B(n8245), .Z(n8250) );
  NANDN U8719 ( .A(n8248), .B(n8247), .Z(n8249) );
  NAND U8720 ( .A(n8250), .B(n8249), .Z(n8548) );
  NANDN U8721 ( .A(n8252), .B(n8251), .Z(n8256) );
  OR U8722 ( .A(n8254), .B(n8253), .Z(n8255) );
  NAND U8723 ( .A(n8256), .B(n8255), .Z(n8547) );
  XNOR U8724 ( .A(n8548), .B(n8547), .Z(n8550) );
  XNOR U8725 ( .A(n8549), .B(n8550), .Z(n8544) );
  OR U8726 ( .A(n8258), .B(n8257), .Z(n8262) );
  OR U8727 ( .A(n8260), .B(n8259), .Z(n8261) );
  AND U8728 ( .A(n8262), .B(n8261), .Z(n8495) );
  NANDN U8729 ( .A(n8264), .B(n8263), .Z(n8268) );
  NAND U8730 ( .A(n8266), .B(n8265), .Z(n8267) );
  NAND U8731 ( .A(n8268), .B(n8267), .Z(n8496) );
  XOR U8732 ( .A(n8495), .B(n8496), .Z(n8498) );
  IV U8733 ( .A(n8269), .Z(n8270) );
  NANDN U8734 ( .A(n8271), .B(n8270), .Z(n8275) );
  OR U8735 ( .A(n8273), .B(n8272), .Z(n8274) );
  AND U8736 ( .A(n8275), .B(n8274), .Z(n8458) );
  ANDN U8737 ( .B(y[722]), .A(n161), .Z(n8478) );
  ANDN U8738 ( .B(y[723]), .A(n160), .Z(n8476) );
  ANDN U8739 ( .B(y[724]), .A(n159), .Z(n8477) );
  XNOR U8740 ( .A(n8476), .B(n8477), .Z(n8479) );
  XNOR U8741 ( .A(n8478), .B(n8479), .Z(n8459) );
  XOR U8742 ( .A(n8458), .B(n8459), .Z(n8460) );
  ANDN U8743 ( .B(y[732]), .A(n151), .Z(n8466) );
  AND U8744 ( .A(n8276), .B(o[91]), .Z(n8464) );
  ANDN U8745 ( .B(y[704]), .A(n14373), .Z(n8465) );
  XNOR U8746 ( .A(n8464), .B(n8465), .Z(n8467) );
  XNOR U8747 ( .A(n8466), .B(n8467), .Z(n8461) );
  XNOR U8748 ( .A(n8498), .B(n8497), .Z(n8486) );
  ANDN U8749 ( .B(y[731]), .A(n152), .Z(n8397) );
  ANDN U8750 ( .B(y[707]), .A(n14372), .Z(n8398) );
  XNOR U8751 ( .A(n8397), .B(n8398), .Z(n8400) );
  XNOR U8752 ( .A(n8399), .B(n8400), .Z(n8491) );
  ANDN U8753 ( .B(y[716]), .A(n167), .Z(n8405) );
  ANDN U8754 ( .B(y[730]), .A(n153), .Z(n8403) );
  ANDN U8755 ( .B(y[708]), .A(n175), .Z(n8404) );
  XNOR U8756 ( .A(n8403), .B(n8404), .Z(n8406) );
  XOR U8757 ( .A(n8405), .B(n8406), .Z(n8489) );
  NANDN U8758 ( .A(n8278), .B(n8277), .Z(n8282) );
  OR U8759 ( .A(n8280), .B(n8279), .Z(n8281) );
  NAND U8760 ( .A(n8282), .B(n8281), .Z(n8490) );
  XNOR U8761 ( .A(n8489), .B(n8490), .Z(n8492) );
  XNOR U8762 ( .A(n8491), .B(n8492), .Z(n8484) );
  ANDN U8763 ( .B(y[709]), .A(n174), .Z(n8433) );
  ANDN U8764 ( .B(y[729]), .A(n154), .Z(n8434) );
  XNOR U8765 ( .A(n8433), .B(n8434), .Z(n8436) );
  XOR U8766 ( .A(n8435), .B(n8436), .Z(n8503) );
  ANDN U8767 ( .B(y[727]), .A(n156), .Z(n8417) );
  ANDN U8768 ( .B(y[712]), .A(n171), .Z(n8415) );
  ANDN U8769 ( .B(y[711]), .A(n172), .Z(n8416) );
  XNOR U8770 ( .A(n8415), .B(n8416), .Z(n8418) );
  XOR U8771 ( .A(n8417), .B(n8418), .Z(n8501) );
  NANDN U8772 ( .A(n8284), .B(n8283), .Z(n8288) );
  NANDN U8773 ( .A(n8286), .B(n8285), .Z(n8287) );
  NAND U8774 ( .A(n8288), .B(n8287), .Z(n8502) );
  XNOR U8775 ( .A(n8501), .B(n8502), .Z(n8504) );
  XNOR U8776 ( .A(n8503), .B(n8504), .Z(n8483) );
  XOR U8777 ( .A(n8484), .B(n8483), .Z(n8485) );
  XNOR U8778 ( .A(n8486), .B(n8485), .Z(n8536) );
  OR U8779 ( .A(n8294), .B(n8293), .Z(n8298) );
  OR U8780 ( .A(n8296), .B(n8295), .Z(n8297) );
  NAND U8781 ( .A(n8298), .B(n8297), .Z(n8520) );
  XOR U8782 ( .A(n8520), .B(n8519), .Z(n8521) );
  XOR U8783 ( .A(n8536), .B(n8535), .Z(n8538) );
  NANDN U8784 ( .A(n8304), .B(n8303), .Z(n8308) );
  OR U8785 ( .A(n8306), .B(n8305), .Z(n8307) );
  AND U8786 ( .A(n8308), .B(n8307), .Z(n8507) );
  OR U8787 ( .A(n8310), .B(n8309), .Z(n8314) );
  NANDN U8788 ( .A(n8312), .B(n8311), .Z(n8313) );
  NAND U8789 ( .A(n8314), .B(n8313), .Z(n8508) );
  XOR U8790 ( .A(n8507), .B(n8508), .Z(n8509) );
  OR U8791 ( .A(n8316), .B(n8315), .Z(n8320) );
  NANDN U8792 ( .A(n8318), .B(n8317), .Z(n8319) );
  NAND U8793 ( .A(n8320), .B(n8319), .Z(n8510) );
  OR U8794 ( .A(n8322), .B(n8321), .Z(n8326) );
  NANDN U8795 ( .A(n8324), .B(n8323), .Z(n8325) );
  AND U8796 ( .A(n8326), .B(n8325), .Z(n8526) );
  ANDN U8797 ( .B(y[725]), .A(n158), .Z(n8411) );
  ANDN U8798 ( .B(y[721]), .A(n162), .Z(n8409) );
  ANDN U8799 ( .B(y[720]), .A(n163), .Z(n8410) );
  XNOR U8800 ( .A(n8409), .B(n8410), .Z(n8412) );
  XOR U8801 ( .A(n8411), .B(n8412), .Z(n8427) );
  NANDN U8802 ( .A(n8328), .B(n8327), .Z(n8332) );
  OR U8803 ( .A(n8330), .B(n8329), .Z(n8331) );
  NAND U8804 ( .A(n8332), .B(n8331), .Z(n8428) );
  XNOR U8805 ( .A(n8427), .B(n8428), .Z(n8430) );
  NAND U8806 ( .A(x[154]), .B(y[706]), .Z(n8440) );
  AND U8807 ( .A(x[143]), .B(y[717]), .Z(n8439) );
  XNOR U8808 ( .A(n8440), .B(n8439), .Z(n8441) );
  AND U8809 ( .A(y[705]), .B(x[155]), .Z(n8644) );
  XNOR U8810 ( .A(o[92]), .B(n8644), .Z(n8442) );
  XOR U8811 ( .A(n8430), .B(n8429), .Z(n8513) );
  OR U8812 ( .A(n8334), .B(n8333), .Z(n8338) );
  OR U8813 ( .A(n8336), .B(n8335), .Z(n8337) );
  AND U8814 ( .A(n8338), .B(n8337), .Z(n8446) );
  ANDN U8815 ( .B(y[726]), .A(n157), .Z(n8425) );
  ANDN U8816 ( .B(y[713]), .A(n170), .Z(n8424) );
  XNOR U8817 ( .A(n8423), .B(n8424), .Z(n8426) );
  XNOR U8818 ( .A(n8425), .B(n8426), .Z(n8447) );
  XOR U8819 ( .A(n8446), .B(n8447), .Z(n8449) );
  NAND U8820 ( .A(x[145]), .B(y[715]), .Z(n8472) );
  ANDN U8821 ( .B(y[728]), .A(n155), .Z(n8471) );
  NAND U8822 ( .A(y[710]), .B(x[150]), .Z(n8470) );
  XOR U8823 ( .A(n8471), .B(n8470), .Z(n8473) );
  XNOR U8824 ( .A(n8472), .B(n8473), .Z(n8448) );
  XNOR U8825 ( .A(n8449), .B(n8448), .Z(n8514) );
  XNOR U8826 ( .A(n8513), .B(n8514), .Z(n8516) );
  OR U8827 ( .A(n8340), .B(n8339), .Z(n8344) );
  OR U8828 ( .A(n8342), .B(n8341), .Z(n8343) );
  AND U8829 ( .A(n8344), .B(n8343), .Z(n8455) );
  OR U8830 ( .A(n8346), .B(n8345), .Z(n8350) );
  NANDN U8831 ( .A(n8348), .B(n8347), .Z(n8349) );
  AND U8832 ( .A(n8350), .B(n8349), .Z(n8452) );
  OR U8833 ( .A(n8352), .B(n8351), .Z(n8356) );
  OR U8834 ( .A(n8354), .B(n8353), .Z(n8355) );
  AND U8835 ( .A(n8356), .B(n8355), .Z(n8453) );
  XOR U8836 ( .A(n8452), .B(n8453), .Z(n8454) );
  XOR U8837 ( .A(n8516), .B(n8515), .Z(n8525) );
  XOR U8838 ( .A(n8526), .B(n8525), .Z(n8528) );
  XOR U8839 ( .A(n8527), .B(n8528), .Z(n8537) );
  XNOR U8840 ( .A(n8538), .B(n8537), .Z(n8534) );
  OR U8841 ( .A(n8358), .B(n8357), .Z(n8362) );
  OR U8842 ( .A(n8360), .B(n8359), .Z(n8361) );
  AND U8843 ( .A(n8362), .B(n8361), .Z(n8531) );
  XOR U8844 ( .A(n8531), .B(n8532), .Z(n8533) );
  XNOR U8845 ( .A(n8534), .B(n8533), .Z(n8541) );
  OR U8846 ( .A(n8368), .B(n8367), .Z(n8372) );
  OR U8847 ( .A(n8370), .B(n8369), .Z(n8371) );
  AND U8848 ( .A(n8372), .B(n8371), .Z(n8542) );
  XOR U8849 ( .A(n8541), .B(n8542), .Z(n8543) );
  XNOR U8850 ( .A(n8544), .B(n8543), .Z(n8391) );
  OR U8851 ( .A(n8374), .B(n8373), .Z(n8378) );
  NAND U8852 ( .A(n8376), .B(n8375), .Z(n8377) );
  AND U8853 ( .A(n8378), .B(n8377), .Z(n8392) );
  XNOR U8854 ( .A(n8391), .B(n8392), .Z(n8394) );
  OR U8855 ( .A(n8380), .B(n8379), .Z(n8384) );
  OR U8856 ( .A(n8382), .B(n8381), .Z(n8383) );
  NAND U8857 ( .A(n8384), .B(n8383), .Z(n8393) );
  XOR U8858 ( .A(n8394), .B(n8393), .Z(n8388) );
  XNOR U8859 ( .A(n8387), .B(n8388), .Z(N189) );
  NANDN U8860 ( .A(n8386), .B(n8385), .Z(n8390) );
  NAND U8861 ( .A(n8388), .B(n8387), .Z(n8389) );
  NAND U8862 ( .A(n8390), .B(n8389), .Z(n8553) );
  OR U8863 ( .A(n8392), .B(n8391), .Z(n8396) );
  OR U8864 ( .A(n8394), .B(n8393), .Z(n8395) );
  AND U8865 ( .A(n8396), .B(n8395), .Z(n8554) );
  XNOR U8866 ( .A(n8553), .B(n8554), .Z(n8555) );
  OR U8867 ( .A(n8398), .B(n8397), .Z(n8402) );
  OR U8868 ( .A(n8400), .B(n8399), .Z(n8401) );
  AND U8869 ( .A(n8402), .B(n8401), .Z(n8572) );
  OR U8870 ( .A(n8404), .B(n8403), .Z(n8408) );
  OR U8871 ( .A(n8406), .B(n8405), .Z(n8407) );
  AND U8872 ( .A(n8408), .B(n8407), .Z(n8569) );
  ANDN U8873 ( .B(y[710]), .A(n174), .Z(n8655) );
  ANDN U8874 ( .B(y[709]), .A(n175), .Z(n8902) );
  XNOR U8875 ( .A(n8655), .B(n8902), .Z(n8657) );
  ANDN U8876 ( .B(y[720]), .A(n164), .Z(n8656) );
  XNOR U8877 ( .A(n8657), .B(n8656), .Z(n8627) );
  OR U8878 ( .A(n8410), .B(n8409), .Z(n8414) );
  OR U8879 ( .A(n8412), .B(n8411), .Z(n8413) );
  AND U8880 ( .A(n8414), .B(n8413), .Z(n8625) );
  ANDN U8881 ( .B(y[722]), .A(n162), .Z(n8649) );
  ANDN U8882 ( .B(y[716]), .A(n168), .Z(n8650) );
  XNOR U8883 ( .A(n8649), .B(n8650), .Z(n8652) );
  ANDN U8884 ( .B(y[730]), .A(n154), .Z(n8651) );
  XOR U8885 ( .A(n8652), .B(n8651), .Z(n8624) );
  XOR U8886 ( .A(n8625), .B(n8624), .Z(n8626) );
  XNOR U8887 ( .A(n8627), .B(n8626), .Z(n8570) );
  XOR U8888 ( .A(n8569), .B(n8570), .Z(n8571) );
  ANDN U8889 ( .B(y[715]), .A(n169), .Z(n8636) );
  ANDN U8890 ( .B(y[714]), .A(n170), .Z(n8637) );
  XNOR U8891 ( .A(n8636), .B(n8637), .Z(n8639) );
  ANDN U8892 ( .B(y[731]), .A(n153), .Z(n8638) );
  XNOR U8893 ( .A(n8639), .B(n8638), .Z(n8671) );
  OR U8894 ( .A(n8416), .B(n8415), .Z(n8420) );
  OR U8895 ( .A(n8418), .B(n8417), .Z(n8419) );
  AND U8896 ( .A(n8420), .B(n8419), .Z(n8669) );
  NAND U8897 ( .A(y[705]), .B(o[92]), .Z(n8421) );
  XNOR U8898 ( .A(y[706]), .B(n8421), .Z(n8422) );
  NAND U8899 ( .A(x[155]), .B(n8422), .Z(n8643) );
  ANDN U8900 ( .B(y[717]), .A(n167), .Z(n8642) );
  XOR U8901 ( .A(n8643), .B(n8642), .Z(n8668) );
  XOR U8902 ( .A(n8669), .B(n8668), .Z(n8670) );
  XNOR U8903 ( .A(n8671), .B(n8670), .Z(n8704) );
  ANDN U8904 ( .B(y[705]), .A(n14373), .Z(n8690) );
  XOR U8905 ( .A(o[93]), .B(n8690), .Z(n8594) );
  ANDN U8906 ( .B(y[704]), .A(n11441), .Z(n8595) );
  XNOR U8907 ( .A(n8594), .B(n8595), .Z(n8597) );
  ANDN U8908 ( .B(y[733]), .A(n151), .Z(n8596) );
  XOR U8909 ( .A(n8597), .B(n8596), .Z(n8581) );
  ANDN U8910 ( .B(y[708]), .A(n14372), .Z(n8674) );
  ANDN U8911 ( .B(y[707]), .A(n176), .Z(n8675) );
  XNOR U8912 ( .A(n8674), .B(n8675), .Z(n8677) );
  ANDN U8913 ( .B(y[719]), .A(n165), .Z(n8676) );
  XOR U8914 ( .A(n8677), .B(n8676), .Z(n8582) );
  XNOR U8915 ( .A(n8581), .B(n8582), .Z(n8584) );
  XOR U8916 ( .A(n8584), .B(n8583), .Z(n8703) );
  XNOR U8917 ( .A(n8704), .B(n8703), .Z(n8705) );
  XOR U8918 ( .A(n8706), .B(n8705), .Z(n8691) );
  OR U8919 ( .A(n8428), .B(n8427), .Z(n8432) );
  OR U8920 ( .A(n8430), .B(n8429), .Z(n8431) );
  AND U8921 ( .A(n8432), .B(n8431), .Z(n8692) );
  XNOR U8922 ( .A(n8691), .B(n8692), .Z(n8694) );
  OR U8923 ( .A(n8434), .B(n8433), .Z(n8438) );
  OR U8924 ( .A(n8436), .B(n8435), .Z(n8437) );
  AND U8925 ( .A(n8438), .B(n8437), .Z(n8618) );
  NANDN U8926 ( .A(n8440), .B(n8439), .Z(n8444) );
  NANDN U8927 ( .A(n8442), .B(n8441), .Z(n8443) );
  NAND U8928 ( .A(n8444), .B(n8443), .Z(n8619) );
  XOR U8929 ( .A(n8618), .B(n8619), .Z(n8620) );
  NOR U8930 ( .A(n160), .B(n8445), .Z(n8813) );
  ANDN U8931 ( .B(y[728]), .A(n156), .Z(n8630) );
  ANDN U8932 ( .B(y[723]), .A(n161), .Z(n8631) );
  XNOR U8933 ( .A(n8630), .B(n8631), .Z(n8633) );
  ANDN U8934 ( .B(y[729]), .A(n155), .Z(n8632) );
  XNOR U8935 ( .A(n8633), .B(n8632), .Z(n8587) );
  XNOR U8936 ( .A(n8813), .B(n8587), .Z(n8589) );
  ANDN U8937 ( .B(y[725]), .A(n159), .Z(n8660) );
  ANDN U8938 ( .B(y[726]), .A(n158), .Z(n8661) );
  XNOR U8939 ( .A(n8660), .B(n8661), .Z(n8663) );
  ANDN U8940 ( .B(y[727]), .A(n157), .Z(n8662) );
  XNOR U8941 ( .A(n8663), .B(n8662), .Z(n8588) );
  XNOR U8942 ( .A(n8589), .B(n8588), .Z(n8621) );
  XOR U8943 ( .A(n8694), .B(n8693), .Z(n8614) );
  OR U8944 ( .A(n8447), .B(n8446), .Z(n8451) );
  NAND U8945 ( .A(n8449), .B(n8448), .Z(n8450) );
  AND U8946 ( .A(n8451), .B(n8450), .Z(n8612) );
  OR U8947 ( .A(n8453), .B(n8452), .Z(n8457) );
  NANDN U8948 ( .A(n8455), .B(n8454), .Z(n8456) );
  AND U8949 ( .A(n8457), .B(n8456), .Z(n8608) );
  OR U8950 ( .A(n8459), .B(n8458), .Z(n8463) );
  NANDN U8951 ( .A(n8461), .B(n8460), .Z(n8462) );
  AND U8952 ( .A(n8463), .B(n8462), .Z(n8606) );
  OR U8953 ( .A(n8465), .B(n8464), .Z(n8469) );
  OR U8954 ( .A(n8467), .B(n8466), .Z(n8468) );
  AND U8955 ( .A(n8469), .B(n8468), .Z(n8603) );
  NANDN U8956 ( .A(n8471), .B(n8470), .Z(n8475) );
  NANDN U8957 ( .A(n8473), .B(n8472), .Z(n8474) );
  AND U8958 ( .A(n8475), .B(n8474), .Z(n8600) );
  OR U8959 ( .A(n8477), .B(n8476), .Z(n8481) );
  OR U8960 ( .A(n8479), .B(n8478), .Z(n8480) );
  AND U8961 ( .A(n8481), .B(n8480), .Z(n8575) );
  ANDN U8962 ( .B(y[713]), .A(n171), .Z(n8683) );
  ANDN U8963 ( .B(y[712]), .A(n172), .Z(n8824) );
  XNOR U8964 ( .A(n8683), .B(n8824), .Z(n8685) );
  ANDN U8965 ( .B(y[718]), .A(n166), .Z(n8684) );
  XNOR U8966 ( .A(n8685), .B(n8684), .Z(n8576) );
  XOR U8967 ( .A(n8575), .B(n8576), .Z(n8578) );
  ANDN U8968 ( .B(y[711]), .A(n173), .Z(n8680) );
  ANDN U8969 ( .B(y[732]), .A(n152), .Z(n8681) );
  XNOR U8970 ( .A(n8680), .B(n8681), .Z(n8682) );
  NOR U8971 ( .A(n163), .B(n8482), .Z(n8946) );
  XOR U8972 ( .A(n8682), .B(n8946), .Z(n8577) );
  XNOR U8973 ( .A(n8578), .B(n8577), .Z(n8601) );
  XOR U8974 ( .A(n8600), .B(n8601), .Z(n8602) );
  XNOR U8975 ( .A(n8606), .B(n8607), .Z(n8609) );
  XNOR U8976 ( .A(n8608), .B(n8609), .Z(n8613) );
  XNOR U8977 ( .A(n8612), .B(n8613), .Z(n8615) );
  XOR U8978 ( .A(n8614), .B(n8615), .Z(n8723) );
  NANDN U8979 ( .A(n8484), .B(n8483), .Z(n8488) );
  OR U8980 ( .A(n8486), .B(n8485), .Z(n8487) );
  AND U8981 ( .A(n8488), .B(n8487), .Z(n8717) );
  OR U8982 ( .A(n8490), .B(n8489), .Z(n8494) );
  NANDN U8983 ( .A(n8492), .B(n8491), .Z(n8493) );
  NAND U8984 ( .A(n8494), .B(n8493), .Z(n8700) );
  OR U8985 ( .A(n8496), .B(n8495), .Z(n8500) );
  NAND U8986 ( .A(n8498), .B(n8497), .Z(n8499) );
  AND U8987 ( .A(n8500), .B(n8499), .Z(n8697) );
  OR U8988 ( .A(n8502), .B(n8501), .Z(n8506) );
  OR U8989 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U8990 ( .A(n8506), .B(n8505), .Z(n8698) );
  XNOR U8991 ( .A(n8697), .B(n8698), .Z(n8699) );
  XOR U8992 ( .A(n8700), .B(n8699), .Z(n8712) );
  OR U8993 ( .A(n8508), .B(n8507), .Z(n8512) );
  NANDN U8994 ( .A(n8510), .B(n8509), .Z(n8511) );
  AND U8995 ( .A(n8512), .B(n8511), .Z(n8709) );
  OR U8996 ( .A(n8514), .B(n8513), .Z(n8518) );
  OR U8997 ( .A(n8516), .B(n8515), .Z(n8517) );
  NAND U8998 ( .A(n8518), .B(n8517), .Z(n8710) );
  XOR U8999 ( .A(n8709), .B(n8710), .Z(n8711) );
  OR U9000 ( .A(n8520), .B(n8519), .Z(n8524) );
  NANDN U9001 ( .A(n8522), .B(n8521), .Z(n8523) );
  AND U9002 ( .A(n8524), .B(n8523), .Z(n8716) );
  XNOR U9003 ( .A(n8715), .B(n8716), .Z(n8718) );
  XOR U9004 ( .A(n8717), .B(n8718), .Z(n8721) );
  NANDN U9005 ( .A(n8526), .B(n8525), .Z(n8530) );
  NANDN U9006 ( .A(n8528), .B(n8527), .Z(n8529) );
  NAND U9007 ( .A(n8530), .B(n8529), .Z(n8722) );
  XNOR U9008 ( .A(n8721), .B(n8722), .Z(n8724) );
  XOR U9009 ( .A(n8723), .B(n8724), .Z(n8568) );
  NANDN U9010 ( .A(n8536), .B(n8535), .Z(n8540) );
  OR U9011 ( .A(n8538), .B(n8537), .Z(n8539) );
  NAND U9012 ( .A(n8540), .B(n8539), .Z(n8566) );
  XOR U9013 ( .A(n8565), .B(n8566), .Z(n8567) );
  XOR U9014 ( .A(n8568), .B(n8567), .Z(n8561) );
  OR U9015 ( .A(n8542), .B(n8541), .Z(n8546) );
  NANDN U9016 ( .A(n8544), .B(n8543), .Z(n8545) );
  AND U9017 ( .A(n8546), .B(n8545), .Z(n8559) );
  OR U9018 ( .A(n8548), .B(n8547), .Z(n8552) );
  NANDN U9019 ( .A(n8550), .B(n8549), .Z(n8551) );
  NAND U9020 ( .A(n8552), .B(n8551), .Z(n8560) );
  XNOR U9021 ( .A(n8559), .B(n8560), .Z(n8562) );
  XOR U9022 ( .A(n8561), .B(n8562), .Z(n8556) );
  XOR U9023 ( .A(n8555), .B(n8556), .Z(N190) );
  NANDN U9024 ( .A(n8554), .B(n8553), .Z(n8558) );
  NANDN U9025 ( .A(n8556), .B(n8555), .Z(n8557) );
  AND U9026 ( .A(n8558), .B(n8557), .Z(n8729) );
  OR U9027 ( .A(n8560), .B(n8559), .Z(n8564) );
  OR U9028 ( .A(n8562), .B(n8561), .Z(n8563) );
  NAND U9029 ( .A(n8564), .B(n8563), .Z(n8730) );
  XNOR U9030 ( .A(n8729), .B(n8730), .Z(n8728) );
  OR U9031 ( .A(n8570), .B(n8569), .Z(n8574) );
  NANDN U9032 ( .A(n8572), .B(n8571), .Z(n8573) );
  AND U9033 ( .A(n8574), .B(n8573), .Z(n8747) );
  OR U9034 ( .A(n8576), .B(n8575), .Z(n8580) );
  NAND U9035 ( .A(n8578), .B(n8577), .Z(n8579) );
  AND U9036 ( .A(n8580), .B(n8579), .Z(n8748) );
  XOR U9037 ( .A(n8747), .B(n8748), .Z(n8745) );
  OR U9038 ( .A(n8582), .B(n8581), .Z(n8586) );
  OR U9039 ( .A(n8584), .B(n8583), .Z(n8585) );
  NAND U9040 ( .A(n8586), .B(n8585), .Z(n8746) );
  XNOR U9041 ( .A(n8745), .B(n8746), .Z(n9001) );
  NAND U9042 ( .A(x[155]), .B(y[707]), .Z(n8952) );
  NAND U9043 ( .A(x[129]), .B(y[733]), .Z(n8951) );
  XNOR U9044 ( .A(n8952), .B(n8951), .Z(n8950) );
  XNOR U9045 ( .A(n8949), .B(n8950), .Z(n8799) );
  AND U9046 ( .A(x[140]), .B(y[722]), .Z(n8591) );
  XNOR U9047 ( .A(n8591), .B(n8590), .Z(n8944) );
  XOR U9048 ( .A(n8943), .B(n8944), .Z(n8812) );
  AND U9049 ( .A(x[138]), .B(y[724]), .Z(n8593) );
  AND U9050 ( .A(y[725]), .B(x[137]), .Z(n8592) );
  XNOR U9051 ( .A(n8593), .B(n8592), .Z(n8811) );
  XOR U9052 ( .A(n8812), .B(n8811), .Z(n8801) );
  OR U9053 ( .A(n8595), .B(n8594), .Z(n8599) );
  OR U9054 ( .A(n8597), .B(n8596), .Z(n8598) );
  AND U9055 ( .A(n8599), .B(n8598), .Z(n8802) );
  XNOR U9056 ( .A(n8801), .B(n8802), .Z(n8800) );
  XOR U9057 ( .A(n8799), .B(n8800), .Z(n8755) );
  XNOR U9058 ( .A(n8756), .B(n8755), .Z(n8754) );
  OR U9059 ( .A(n8601), .B(n8600), .Z(n8605) );
  NANDN U9060 ( .A(n8603), .B(n8602), .Z(n8604) );
  NAND U9061 ( .A(n8605), .B(n8604), .Z(n8753) );
  XOR U9062 ( .A(n8754), .B(n8753), .Z(n9002) );
  XOR U9063 ( .A(n9001), .B(n9002), .Z(n9003) );
  OR U9064 ( .A(n8607), .B(n8606), .Z(n8611) );
  OR U9065 ( .A(n8609), .B(n8608), .Z(n8610) );
  NAND U9066 ( .A(n8611), .B(n8610), .Z(n9004) );
  XOR U9067 ( .A(n9003), .B(n9004), .Z(n8735) );
  OR U9068 ( .A(n8613), .B(n8612), .Z(n8617) );
  OR U9069 ( .A(n8615), .B(n8614), .Z(n8616) );
  NAND U9070 ( .A(n8617), .B(n8616), .Z(n8736) );
  OR U9071 ( .A(n8619), .B(n8618), .Z(n8623) );
  NANDN U9072 ( .A(n8621), .B(n8620), .Z(n8622) );
  AND U9073 ( .A(n8623), .B(n8622), .Z(n8979) );
  NANDN U9074 ( .A(n8625), .B(n8624), .Z(n8629) );
  OR U9075 ( .A(n8627), .B(n8626), .Z(n8628) );
  AND U9076 ( .A(n8629), .B(n8628), .Z(n8981) );
  OR U9077 ( .A(n8631), .B(n8630), .Z(n8635) );
  OR U9078 ( .A(n8633), .B(n8632), .Z(n8634) );
  AND U9079 ( .A(n8635), .B(n8634), .Z(n8772) );
  NAND U9080 ( .A(x[134]), .B(y[728]), .Z(n8906) );
  NAND U9081 ( .A(x[133]), .B(y[729]), .Z(n8908) );
  NAND U9082 ( .A(x[147]), .B(y[715]), .Z(n8907) );
  XNOR U9083 ( .A(n8908), .B(n8907), .Z(n8905) );
  XNOR U9084 ( .A(n8906), .B(n8905), .Z(n8791) );
  OR U9085 ( .A(n8637), .B(n8636), .Z(n8641) );
  OR U9086 ( .A(n8639), .B(n8638), .Z(n8640) );
  AND U9087 ( .A(n8641), .B(n8640), .Z(n8793) );
  NAND U9088 ( .A(x[132]), .B(y[730]), .Z(n8832) );
  NAND U9089 ( .A(x[131]), .B(y[731]), .Z(n8830) );
  AND U9090 ( .A(y[716]), .B(x[146]), .Z(n8829) );
  XNOR U9091 ( .A(n8830), .B(n8829), .Z(n8831) );
  XNOR U9092 ( .A(n8832), .B(n8831), .Z(n8794) );
  XOR U9093 ( .A(n8793), .B(n8794), .Z(n8792) );
  XNOR U9094 ( .A(n8791), .B(n8792), .Z(n8771) );
  XOR U9095 ( .A(n8772), .B(n8771), .Z(n8774) );
  OR U9096 ( .A(n8643), .B(n8642), .Z(n8648) );
  NAND U9097 ( .A(n8644), .B(o[92]), .Z(n8646) );
  NAND U9098 ( .A(x[155]), .B(y[706]), .Z(n8645) );
  AND U9099 ( .A(n8646), .B(n8645), .Z(n8647) );
  ANDN U9100 ( .B(n8648), .A(n8647), .Z(n8773) );
  XNOR U9101 ( .A(n8981), .B(n8982), .Z(n8980) );
  XNOR U9102 ( .A(n8979), .B(n8980), .Z(n8976) );
  OR U9103 ( .A(n8650), .B(n8649), .Z(n8654) );
  OR U9104 ( .A(n8652), .B(n8651), .Z(n8653) );
  NAND U9105 ( .A(n8654), .B(n8653), .Z(n8780) );
  NAND U9106 ( .A(x[148]), .B(y[714]), .Z(n8938) );
  AND U9107 ( .A(y[720]), .B(x[142]), .Z(n8937) );
  XOR U9108 ( .A(n8938), .B(n8937), .Z(n8936) );
  AND U9109 ( .A(y[726]), .B(x[136]), .Z(n8935) );
  XOR U9110 ( .A(n8936), .B(n8935), .Z(n8782) );
  NAND U9111 ( .A(y[704]), .B(x[158]), .Z(n8808) );
  NAND U9112 ( .A(x[157]), .B(y[705]), .Z(n8861) );
  XNOR U9113 ( .A(o[94]), .B(n8861), .Z(n8807) );
  XOR U9114 ( .A(n8808), .B(n8807), .Z(n8806) );
  AND U9115 ( .A(y[734]), .B(x[128]), .Z(n8805) );
  XNOR U9116 ( .A(n8806), .B(n8805), .Z(n8781) );
  XOR U9117 ( .A(n8780), .B(n8779), .Z(n8761) );
  OR U9118 ( .A(n8902), .B(n8655), .Z(n8659) );
  OR U9119 ( .A(n8657), .B(n8656), .Z(n8658) );
  AND U9120 ( .A(n8659), .B(n8658), .Z(n8762) );
  XNOR U9121 ( .A(n8761), .B(n8762), .Z(n8760) );
  OR U9122 ( .A(n8661), .B(n8660), .Z(n8665) );
  OR U9123 ( .A(n8663), .B(n8662), .Z(n8664) );
  AND U9124 ( .A(n8665), .B(n8664), .Z(n8856) );
  NAND U9125 ( .A(x[145]), .B(y[717]), .Z(n8930) );
  NAND U9126 ( .A(x[130]), .B(y[732]), .Z(n8932) );
  NAND U9127 ( .A(x[154]), .B(y[708]), .Z(n8931) );
  XNOR U9128 ( .A(n8932), .B(n8931), .Z(n8929) );
  XNOR U9129 ( .A(n8930), .B(n8929), .Z(n8858) );
  NAND U9130 ( .A(x[135]), .B(y[727]), .Z(n8825) );
  AND U9131 ( .A(x[150]), .B(y[712]), .Z(n8667) );
  AND U9132 ( .A(x[149]), .B(y[713]), .Z(n8666) );
  XNOR U9133 ( .A(n8667), .B(n8666), .Z(n8826) );
  XOR U9134 ( .A(n8825), .B(n8826), .Z(n8857) );
  XNOR U9135 ( .A(n8858), .B(n8857), .Z(n8855) );
  XOR U9136 ( .A(n8856), .B(n8855), .Z(n8759) );
  XNOR U9137 ( .A(n8760), .B(n8759), .Z(n8739) );
  NANDN U9138 ( .A(n8669), .B(n8668), .Z(n8673) );
  OR U9139 ( .A(n8671), .B(n8670), .Z(n8672) );
  NAND U9140 ( .A(n8673), .B(n8672), .Z(n8742) );
  OR U9141 ( .A(n8675), .B(n8674), .Z(n8679) );
  OR U9142 ( .A(n8677), .B(n8676), .Z(n8678) );
  AND U9143 ( .A(n8679), .B(n8678), .Z(n8765) );
  OR U9144 ( .A(n8824), .B(n8683), .Z(n8687) );
  OR U9145 ( .A(n8685), .B(n8684), .Z(n8686) );
  AND U9146 ( .A(n8687), .B(n8686), .Z(n8785) );
  NAND U9147 ( .A(x[151]), .B(y[711]), .Z(n8901) );
  AND U9148 ( .A(y[709]), .B(x[153]), .Z(n8689) );
  AND U9149 ( .A(x[152]), .B(y[710]), .Z(n8688) );
  XNOR U9150 ( .A(n8689), .B(n8688), .Z(n8900) );
  XOR U9151 ( .A(n8901), .B(n8900), .Z(n8787) );
  NAND U9152 ( .A(n8690), .B(o[93]), .Z(n8820) );
  NAND U9153 ( .A(x[156]), .B(y[706]), .Z(n8818) );
  AND U9154 ( .A(x[144]), .B(y[718]), .Z(n8819) );
  XNOR U9155 ( .A(n8818), .B(n8819), .Z(n8821) );
  XNOR U9156 ( .A(n8820), .B(n8821), .Z(n8788) );
  XNOR U9157 ( .A(n8787), .B(n8788), .Z(n8786) );
  XOR U9158 ( .A(n8785), .B(n8786), .Z(n8767) );
  XOR U9159 ( .A(n8765), .B(n8766), .Z(n8741) );
  XNOR U9160 ( .A(n8742), .B(n8741), .Z(n8740) );
  XNOR U9161 ( .A(n8739), .B(n8740), .Z(n8975) );
  XNOR U9162 ( .A(n8976), .B(n8975), .Z(n8974) );
  OR U9163 ( .A(n8692), .B(n8691), .Z(n8696) );
  OR U9164 ( .A(n8694), .B(n8693), .Z(n8695) );
  NAND U9165 ( .A(n8696), .B(n8695), .Z(n8973) );
  XNOR U9166 ( .A(n8974), .B(n8973), .Z(n8995) );
  OR U9167 ( .A(n8698), .B(n8697), .Z(n8702) );
  OR U9168 ( .A(n8700), .B(n8699), .Z(n8701) );
  NAND U9169 ( .A(n8702), .B(n8701), .Z(n8998) );
  OR U9170 ( .A(n8704), .B(n8703), .Z(n8708) );
  OR U9171 ( .A(n8706), .B(n8705), .Z(n8707) );
  NAND U9172 ( .A(n8708), .B(n8707), .Z(n8997) );
  XNOR U9173 ( .A(n8998), .B(n8997), .Z(n8996) );
  XOR U9174 ( .A(n8995), .B(n8996), .Z(n8733) );
  XNOR U9175 ( .A(n8734), .B(n8733), .Z(n9015) );
  OR U9176 ( .A(n8710), .B(n8709), .Z(n8714) );
  NANDN U9177 ( .A(n8712), .B(n8711), .Z(n8713) );
  NAND U9178 ( .A(n8714), .B(n8713), .Z(n9020) );
  OR U9179 ( .A(n8716), .B(n8715), .Z(n8720) );
  OR U9180 ( .A(n8718), .B(n8717), .Z(n8719) );
  AND U9181 ( .A(n8720), .B(n8719), .Z(n9021) );
  OR U9182 ( .A(n8722), .B(n8721), .Z(n8726) );
  OR U9183 ( .A(n8724), .B(n8723), .Z(n8725) );
  NAND U9184 ( .A(n8726), .B(n8725), .Z(n9022) );
  XNOR U9185 ( .A(n9021), .B(n9022), .Z(n9019) );
  XOR U9186 ( .A(n9020), .B(n9019), .Z(n9016) );
  XNOR U9187 ( .A(n9015), .B(n9016), .Z(n9014) );
  XOR U9188 ( .A(n9013), .B(n9014), .Z(n8727) );
  XOR U9189 ( .A(n8728), .B(n8727), .Z(N191) );
  NANDN U9190 ( .A(n8728), .B(n8727), .Z(n8732) );
  OR U9191 ( .A(n8730), .B(n8729), .Z(n8731) );
  AND U9192 ( .A(n8732), .B(n8731), .Z(n9012) );
  OR U9193 ( .A(n8734), .B(n8733), .Z(n8738) );
  NANDN U9194 ( .A(n8736), .B(n8735), .Z(n8737) );
  AND U9195 ( .A(n8738), .B(n8737), .Z(n8994) );
  NANDN U9196 ( .A(n8740), .B(n8739), .Z(n8744) );
  OR U9197 ( .A(n8742), .B(n8741), .Z(n8743) );
  AND U9198 ( .A(n8744), .B(n8743), .Z(n8752) );
  NANDN U9199 ( .A(n8746), .B(n8745), .Z(n8750) );
  OR U9200 ( .A(n8748), .B(n8747), .Z(n8749) );
  NAND U9201 ( .A(n8750), .B(n8749), .Z(n8751) );
  XNOR U9202 ( .A(n8752), .B(n8751), .Z(n8992) );
  OR U9203 ( .A(n8754), .B(n8753), .Z(n8758) );
  OR U9204 ( .A(n8756), .B(n8755), .Z(n8757) );
  AND U9205 ( .A(n8758), .B(n8757), .Z(n8990) );
  OR U9206 ( .A(n8760), .B(n8759), .Z(n8764) );
  OR U9207 ( .A(n8762), .B(n8761), .Z(n8763) );
  AND U9208 ( .A(n8764), .B(n8763), .Z(n8972) );
  OR U9209 ( .A(n8766), .B(n8765), .Z(n8770) );
  NANDN U9210 ( .A(n8768), .B(n8767), .Z(n8769) );
  AND U9211 ( .A(n8770), .B(n8769), .Z(n8778) );
  NOR U9212 ( .A(n8772), .B(n8771), .Z(n8776) );
  ANDN U9213 ( .B(n8774), .A(n8773), .Z(n8775) );
  OR U9214 ( .A(n8776), .B(n8775), .Z(n8777) );
  XNOR U9215 ( .A(n8778), .B(n8777), .Z(n8970) );
  OR U9216 ( .A(n8780), .B(n8779), .Z(n8784) );
  NANDN U9217 ( .A(n8782), .B(n8781), .Z(n8783) );
  AND U9218 ( .A(n8784), .B(n8783), .Z(n8968) );
  OR U9219 ( .A(n8786), .B(n8785), .Z(n8790) );
  OR U9220 ( .A(n8788), .B(n8787), .Z(n8789) );
  AND U9221 ( .A(n8790), .B(n8789), .Z(n8798) );
  NAND U9222 ( .A(n8792), .B(n8791), .Z(n8796) );
  OR U9223 ( .A(n8794), .B(n8793), .Z(n8795) );
  NAND U9224 ( .A(n8796), .B(n8795), .Z(n8797) );
  XNOR U9225 ( .A(n8798), .B(n8797), .Z(n8966) );
  OR U9226 ( .A(n8800), .B(n8799), .Z(n8804) );
  OR U9227 ( .A(n8802), .B(n8801), .Z(n8803) );
  AND U9228 ( .A(n8804), .B(n8803), .Z(n8964) );
  NANDN U9229 ( .A(n8806), .B(n8805), .Z(n8810) );
  NANDN U9230 ( .A(n8808), .B(n8807), .Z(n8809) );
  AND U9231 ( .A(n8810), .B(n8809), .Z(n8817) );
  OR U9232 ( .A(n8812), .B(n8811), .Z(n8815) );
  NAND U9233 ( .A(x[138]), .B(y[725]), .Z(n8863) );
  NANDN U9234 ( .A(n8863), .B(n8813), .Z(n8814) );
  NAND U9235 ( .A(n8815), .B(n8814), .Z(n8816) );
  XNOR U9236 ( .A(n8817), .B(n8816), .Z(n8962) );
  ANDN U9237 ( .B(n8819), .A(n8818), .Z(n8823) );
  ANDN U9238 ( .B(n8821), .A(n8820), .Z(n8822) );
  NOR U9239 ( .A(n8823), .B(n8822), .Z(n8854) );
  NAND U9240 ( .A(x[150]), .B(y[713]), .Z(n8862) );
  ANDN U9241 ( .B(n8824), .A(n8862), .Z(n8828) );
  NOR U9242 ( .A(n8826), .B(n8825), .Z(n8827) );
  NOR U9243 ( .A(n8828), .B(n8827), .Z(n8836) );
  NANDN U9244 ( .A(n8830), .B(n8829), .Z(n8834) );
  NANDN U9245 ( .A(n8832), .B(n8831), .Z(n8833) );
  AND U9246 ( .A(n8834), .B(n8833), .Z(n8835) );
  XNOR U9247 ( .A(n8836), .B(n8835), .Z(n8852) );
  AND U9248 ( .A(y[732]), .B(x[131]), .Z(n8838) );
  NAND U9249 ( .A(x[129]), .B(y[734]), .Z(n8837) );
  XNOR U9250 ( .A(n8838), .B(n8837), .Z(n8842) );
  AND U9251 ( .A(x[159]), .B(y[704]), .Z(n8840) );
  NAND U9252 ( .A(x[146]), .B(y[717]), .Z(n8839) );
  XNOR U9253 ( .A(n8840), .B(n8839), .Z(n8841) );
  XOR U9254 ( .A(n8842), .B(n8841), .Z(n8850) );
  AND U9255 ( .A(y[706]), .B(x[157]), .Z(n8844) );
  NAND U9256 ( .A(x[128]), .B(y[735]), .Z(n8843) );
  XNOR U9257 ( .A(n8844), .B(n8843), .Z(n8848) );
  AND U9258 ( .A(y[720]), .B(x[143]), .Z(n8846) );
  NAND U9259 ( .A(x[156]), .B(y[707]), .Z(n8845) );
  XNOR U9260 ( .A(n8846), .B(n8845), .Z(n8847) );
  XNOR U9261 ( .A(n8848), .B(n8847), .Z(n8849) );
  XNOR U9262 ( .A(n8850), .B(n8849), .Z(n8851) );
  XOR U9263 ( .A(n8852), .B(n8851), .Z(n8853) );
  XNOR U9264 ( .A(n8854), .B(n8853), .Z(n8928) );
  NANDN U9265 ( .A(n8856), .B(n8855), .Z(n8860) );
  ANDN U9266 ( .B(n8858), .A(n8857), .Z(n8859) );
  ANDN U9267 ( .B(n8860), .A(n8859), .Z(n8926) );
  AND U9268 ( .A(y[727]), .B(x[136]), .Z(n8869) );
  ANDN U9269 ( .B(o[94]), .A(n8861), .Z(n8867) );
  XNOR U9270 ( .A(n8862), .B(o[95]), .Z(n8865) );
  XOR U9271 ( .A(n8945), .B(n8863), .Z(n8864) );
  XNOR U9272 ( .A(n8865), .B(n8864), .Z(n8866) );
  XNOR U9273 ( .A(n8867), .B(n8866), .Z(n8868) );
  XNOR U9274 ( .A(n8869), .B(n8868), .Z(n8877) );
  AND U9275 ( .A(y[729]), .B(x[134]), .Z(n8871) );
  NAND U9276 ( .A(x[152]), .B(y[711]), .Z(n8870) );
  XNOR U9277 ( .A(n8871), .B(n8870), .Z(n8875) );
  AND U9278 ( .A(y[716]), .B(x[147]), .Z(n8873) );
  NAND U9279 ( .A(x[149]), .B(y[714]), .Z(n8872) );
  XNOR U9280 ( .A(n8873), .B(n8872), .Z(n8874) );
  XNOR U9281 ( .A(n8875), .B(n8874), .Z(n8876) );
  XNOR U9282 ( .A(n8877), .B(n8876), .Z(n8924) );
  AND U9283 ( .A(y[726]), .B(x[137]), .Z(n8879) );
  NAND U9284 ( .A(x[132]), .B(y[731]), .Z(n8878) );
  XNOR U9285 ( .A(n8879), .B(n8878), .Z(n8883) );
  AND U9286 ( .A(y[709]), .B(x[154]), .Z(n8881) );
  NAND U9287 ( .A(x[142]), .B(y[721]), .Z(n8880) );
  XNOR U9288 ( .A(n8881), .B(n8880), .Z(n8882) );
  XOR U9289 ( .A(n8883), .B(n8882), .Z(n8891) );
  AND U9290 ( .A(y[723]), .B(x[140]), .Z(n8885) );
  NAND U9291 ( .A(x[139]), .B(y[724]), .Z(n8884) );
  XNOR U9292 ( .A(n8885), .B(n8884), .Z(n8889) );
  AND U9293 ( .A(y[715]), .B(x[148]), .Z(n8887) );
  NAND U9294 ( .A(x[144]), .B(y[719]), .Z(n8886) );
  XNOR U9295 ( .A(n8887), .B(n8886), .Z(n8888) );
  XNOR U9296 ( .A(n8889), .B(n8888), .Z(n8890) );
  XNOR U9297 ( .A(n8891), .B(n8890), .Z(n8899) );
  AND U9298 ( .A(x[158]), .B(y[705]), .Z(n8893) );
  NAND U9299 ( .A(x[155]), .B(y[708]), .Z(n8892) );
  XNOR U9300 ( .A(n8893), .B(n8892), .Z(n8897) );
  AND U9301 ( .A(x[151]), .B(y[712]), .Z(n8895) );
  NAND U9302 ( .A(x[145]), .B(y[718]), .Z(n8894) );
  XNOR U9303 ( .A(n8895), .B(n8894), .Z(n8896) );
  XNOR U9304 ( .A(n8897), .B(n8896), .Z(n8898) );
  XNOR U9305 ( .A(n8899), .B(n8898), .Z(n8914) );
  OR U9306 ( .A(n8901), .B(n8900), .Z(n8904) );
  NAND U9307 ( .A(x[153]), .B(y[710]), .Z(n8920) );
  NANDN U9308 ( .A(n8920), .B(n8902), .Z(n8903) );
  AND U9309 ( .A(n8904), .B(n8903), .Z(n8912) );
  OR U9310 ( .A(n8906), .B(n8905), .Z(n8910) );
  OR U9311 ( .A(n8908), .B(n8907), .Z(n8909) );
  NAND U9312 ( .A(n8910), .B(n8909), .Z(n8911) );
  XNOR U9313 ( .A(n8912), .B(n8911), .Z(n8913) );
  XOR U9314 ( .A(n8914), .B(n8913), .Z(n8922) );
  AND U9315 ( .A(y[730]), .B(x[133]), .Z(n8916) );
  NAND U9316 ( .A(x[130]), .B(y[733]), .Z(n8915) );
  XNOR U9317 ( .A(n8916), .B(n8915), .Z(n8918) );
  NAND U9318 ( .A(x[135]), .B(y[728]), .Z(n8917) );
  XNOR U9319 ( .A(n8918), .B(n8917), .Z(n8919) );
  XOR U9320 ( .A(n8920), .B(n8919), .Z(n8921) );
  XNOR U9321 ( .A(n8922), .B(n8921), .Z(n8923) );
  XNOR U9322 ( .A(n8924), .B(n8923), .Z(n8925) );
  XNOR U9323 ( .A(n8926), .B(n8925), .Z(n8927) );
  XOR U9324 ( .A(n8928), .B(n8927), .Z(n8960) );
  OR U9325 ( .A(n8930), .B(n8929), .Z(n8934) );
  OR U9326 ( .A(n8932), .B(n8931), .Z(n8933) );
  AND U9327 ( .A(n8934), .B(n8933), .Z(n8942) );
  NANDN U9328 ( .A(n8936), .B(n8935), .Z(n8940) );
  NANDN U9329 ( .A(n8938), .B(n8937), .Z(n8939) );
  NAND U9330 ( .A(n8940), .B(n8939), .Z(n8941) );
  XNOR U9331 ( .A(n8942), .B(n8941), .Z(n8958) );
  NANDN U9332 ( .A(n8944), .B(n8943), .Z(n8948) );
  NAND U9333 ( .A(n8946), .B(n8945), .Z(n8947) );
  AND U9334 ( .A(n8948), .B(n8947), .Z(n8956) );
  NANDN U9335 ( .A(n8950), .B(n8949), .Z(n8954) );
  OR U9336 ( .A(n8952), .B(n8951), .Z(n8953) );
  NAND U9337 ( .A(n8954), .B(n8953), .Z(n8955) );
  XNOR U9338 ( .A(n8956), .B(n8955), .Z(n8957) );
  XNOR U9339 ( .A(n8958), .B(n8957), .Z(n8959) );
  XNOR U9340 ( .A(n8960), .B(n8959), .Z(n8961) );
  XNOR U9341 ( .A(n8962), .B(n8961), .Z(n8963) );
  XNOR U9342 ( .A(n8964), .B(n8963), .Z(n8965) );
  XNOR U9343 ( .A(n8966), .B(n8965), .Z(n8967) );
  XNOR U9344 ( .A(n8968), .B(n8967), .Z(n8969) );
  XNOR U9345 ( .A(n8970), .B(n8969), .Z(n8971) );
  XNOR U9346 ( .A(n8972), .B(n8971), .Z(n8988) );
  OR U9347 ( .A(n8974), .B(n8973), .Z(n8978) );
  OR U9348 ( .A(n8976), .B(n8975), .Z(n8977) );
  AND U9349 ( .A(n8978), .B(n8977), .Z(n8986) );
  OR U9350 ( .A(n8980), .B(n8979), .Z(n8984) );
  OR U9351 ( .A(n8982), .B(n8981), .Z(n8983) );
  NAND U9352 ( .A(n8984), .B(n8983), .Z(n8985) );
  XNOR U9353 ( .A(n8986), .B(n8985), .Z(n8987) );
  XNOR U9354 ( .A(n8988), .B(n8987), .Z(n8989) );
  XNOR U9355 ( .A(n8990), .B(n8989), .Z(n8991) );
  XNOR U9356 ( .A(n8992), .B(n8991), .Z(n8993) );
  XNOR U9357 ( .A(n8994), .B(n8993), .Z(n9010) );
  NANDN U9358 ( .A(n8996), .B(n8995), .Z(n9000) );
  OR U9359 ( .A(n8998), .B(n8997), .Z(n8999) );
  AND U9360 ( .A(n9000), .B(n8999), .Z(n9008) );
  ANDN U9361 ( .B(n9002), .A(n9001), .Z(n9006) );
  NOR U9362 ( .A(n9004), .B(n9003), .Z(n9005) );
  OR U9363 ( .A(n9006), .B(n9005), .Z(n9007) );
  XNOR U9364 ( .A(n9008), .B(n9007), .Z(n9009) );
  XNOR U9365 ( .A(n9010), .B(n9009), .Z(n9011) );
  XNOR U9366 ( .A(n9012), .B(n9011), .Z(n9028) );
  OR U9367 ( .A(n9014), .B(n9013), .Z(n9018) );
  NAND U9368 ( .A(n9016), .B(n9015), .Z(n9017) );
  AND U9369 ( .A(n9018), .B(n9017), .Z(n9026) );
  OR U9370 ( .A(n9020), .B(n9019), .Z(n9024) );
  OR U9371 ( .A(n9022), .B(n9021), .Z(n9023) );
  NAND U9372 ( .A(n9024), .B(n9023), .Z(n9025) );
  XNOR U9373 ( .A(n9026), .B(n9025), .Z(n9027) );
  XNOR U9374 ( .A(n9028), .B(n9027), .Z(N192) );
  AND U9375 ( .A(y[736]), .B(x[128]), .Z(n9710) );
  XOR U9376 ( .A(n9710), .B(o[96]), .Z(N225) );
  AND U9377 ( .A(y[736]), .B(x[129]), .Z(n9029) );
  NAND U9378 ( .A(x[128]), .B(y[737]), .Z(n9035) );
  XNOR U9379 ( .A(n9035), .B(o[97]), .Z(n9030) );
  XOR U9380 ( .A(n9029), .B(n9030), .Z(n9031) );
  AND U9381 ( .A(o[96]), .B(n9710), .Z(n9032) );
  XOR U9382 ( .A(n9031), .B(n9032), .Z(N226) );
  OR U9383 ( .A(n9030), .B(n9029), .Z(n9034) );
  NANDN U9384 ( .A(n9032), .B(n9031), .Z(n9033) );
  NAND U9385 ( .A(n9034), .B(n9033), .Z(n9037) );
  NAND U9386 ( .A(x[128]), .B(y[738]), .Z(n9048) );
  XOR U9387 ( .A(n9048), .B(o[98]), .Z(n9036) );
  XNOR U9388 ( .A(n9037), .B(n9036), .Z(n9039) );
  ANDN U9389 ( .B(o[97]), .A(n9035), .Z(n9042) );
  ANDN U9390 ( .B(y[736]), .A(n153), .Z(n9043) );
  XNOR U9391 ( .A(n9042), .B(n9043), .Z(n9045) );
  ANDN U9392 ( .B(y[737]), .A(n152), .Z(n9044) );
  XNOR U9393 ( .A(n9045), .B(n9044), .Z(n9038) );
  XNOR U9394 ( .A(n9039), .B(n9038), .Z(N227) );
  NAND U9395 ( .A(n9037), .B(n9036), .Z(n9041) );
  OR U9396 ( .A(n9039), .B(n9038), .Z(n9040) );
  NAND U9397 ( .A(n9041), .B(n9040), .Z(n9052) );
  OR U9398 ( .A(n9043), .B(n9042), .Z(n9047) );
  OR U9399 ( .A(n9045), .B(n9044), .Z(n9046) );
  AND U9400 ( .A(n9047), .B(n9046), .Z(n9053) );
  XNOR U9401 ( .A(n9052), .B(n9053), .Z(n9054) );
  NAND U9402 ( .A(x[130]), .B(y[737]), .Z(n9060) );
  XNOR U9403 ( .A(n9060), .B(o[99]), .Z(n9058) );
  NANDN U9404 ( .A(n9048), .B(o[98]), .Z(n9064) );
  AND U9405 ( .A(y[736]), .B(x[131]), .Z(n9050) );
  NAND U9406 ( .A(x[128]), .B(y[739]), .Z(n9049) );
  XOR U9407 ( .A(n9050), .B(n9049), .Z(n9063) );
  XNOR U9408 ( .A(n9064), .B(n9063), .Z(n9059) );
  ANDN U9409 ( .B(y[738]), .A(n152), .Z(n9088) );
  XOR U9410 ( .A(n9059), .B(n9088), .Z(n9051) );
  XOR U9411 ( .A(n9058), .B(n9051), .Z(n9055) );
  XNOR U9412 ( .A(n9054), .B(n9055), .Z(N228) );
  NANDN U9413 ( .A(n9053), .B(n9052), .Z(n9057) );
  NAND U9414 ( .A(n9055), .B(n9054), .Z(n9056) );
  NAND U9415 ( .A(n9057), .B(n9056), .Z(n9069) );
  XNOR U9416 ( .A(n9069), .B(n9070), .Z(n9071) );
  NANDN U9417 ( .A(n9060), .B(o[99]), .Z(n9085) );
  AND U9418 ( .A(y[736]), .B(x[132]), .Z(n9062) );
  AND U9419 ( .A(y[740]), .B(x[128]), .Z(n9061) );
  XNOR U9420 ( .A(n9062), .B(n9061), .Z(n9084) );
  XOR U9421 ( .A(n9085), .B(n9084), .Z(n9077) );
  ANDN U9422 ( .B(y[739]), .A(n154), .Z(n9136) );
  NAND U9423 ( .A(n9710), .B(n9136), .Z(n9066) );
  OR U9424 ( .A(n9064), .B(n9063), .Z(n9065) );
  NAND U9425 ( .A(n9066), .B(n9065), .Z(n9075) );
  AND U9426 ( .A(x[129]), .B(y[739]), .Z(n9068) );
  NAND U9427 ( .A(x[130]), .B(y[738]), .Z(n9067) );
  XOR U9428 ( .A(n9068), .B(n9067), .Z(n9090) );
  NAND U9429 ( .A(x[131]), .B(y[737]), .Z(n9081) );
  XNOR U9430 ( .A(n9081), .B(o[100]), .Z(n9089) );
  XOR U9431 ( .A(n9090), .B(n9089), .Z(n9076) );
  XOR U9432 ( .A(n9077), .B(n9078), .Z(n9072) );
  XOR U9433 ( .A(n9071), .B(n9072), .Z(N229) );
  NANDN U9434 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U9435 ( .A(n9072), .B(n9071), .Z(n9073) );
  NAND U9436 ( .A(n9074), .B(n9073), .Z(n9093) );
  NANDN U9437 ( .A(n9076), .B(n9075), .Z(n9080) );
  NAND U9438 ( .A(n9078), .B(n9077), .Z(n9079) );
  NAND U9439 ( .A(n9080), .B(n9079), .Z(n9094) );
  XNOR U9440 ( .A(n9093), .B(n9094), .Z(n9095) );
  NANDN U9441 ( .A(n9081), .B(o[100]), .Z(n9112) );
  AND U9442 ( .A(y[736]), .B(x[133]), .Z(n9083) );
  AND U9443 ( .A(y[741]), .B(x[128]), .Z(n9082) );
  XNOR U9444 ( .A(n9083), .B(n9082), .Z(n9111) );
  XOR U9445 ( .A(n9112), .B(n9111), .Z(n9107) );
  ANDN U9446 ( .B(y[739]), .A(n153), .Z(n9105) );
  ANDN U9447 ( .B(y[740]), .A(n152), .Z(n9120) );
  ANDN U9448 ( .B(y[737]), .A(n155), .Z(n9115) );
  XOR U9449 ( .A(o[101]), .B(n9115), .Z(n9118) );
  ANDN U9450 ( .B(y[738]), .A(n154), .Z(n9119) );
  XNOR U9451 ( .A(n9118), .B(n9119), .Z(n9121) );
  XNOR U9452 ( .A(n9120), .B(n9121), .Z(n9106) );
  XNOR U9453 ( .A(n9105), .B(n9106), .Z(n9108) );
  XNOR U9454 ( .A(n9107), .B(n9108), .Z(n9102) );
  ANDN U9455 ( .B(y[740]), .A(n155), .Z(n9198) );
  NAND U9456 ( .A(n9710), .B(n9198), .Z(n9087) );
  OR U9457 ( .A(n9085), .B(n9084), .Z(n9086) );
  NAND U9458 ( .A(n9087), .B(n9086), .Z(n9100) );
  NAND U9459 ( .A(n9088), .B(n9105), .Z(n9092) );
  NANDN U9460 ( .A(n9090), .B(n9089), .Z(n9091) );
  NAND U9461 ( .A(n9092), .B(n9091), .Z(n9099) );
  XNOR U9462 ( .A(n9100), .B(n9099), .Z(n9101) );
  XNOR U9463 ( .A(n9102), .B(n9101), .Z(n9096) );
  XOR U9464 ( .A(n9095), .B(n9096), .Z(N230) );
  NANDN U9465 ( .A(n9094), .B(n9093), .Z(n9098) );
  NANDN U9466 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U9467 ( .A(n9098), .B(n9097), .Z(n9124) );
  OR U9468 ( .A(n9100), .B(n9099), .Z(n9104) );
  OR U9469 ( .A(n9102), .B(n9101), .Z(n9103) );
  AND U9470 ( .A(n9104), .B(n9103), .Z(n9125) );
  XNOR U9471 ( .A(n9124), .B(n9125), .Z(n9126) );
  OR U9472 ( .A(n9106), .B(n9105), .Z(n9110) );
  OR U9473 ( .A(n9108), .B(n9107), .Z(n9109) );
  AND U9474 ( .A(n9110), .B(n9109), .Z(n9130) );
  NAND U9475 ( .A(x[133]), .B(y[741]), .Z(n9462) );
  NANDN U9476 ( .A(n9462), .B(n9710), .Z(n9114) );
  OR U9477 ( .A(n9112), .B(n9111), .Z(n9113) );
  NAND U9478 ( .A(n9114), .B(n9113), .Z(n9152) );
  NAND U9479 ( .A(n9115), .B(o[101]), .Z(n9142) );
  AND U9480 ( .A(y[736]), .B(x[134]), .Z(n9117) );
  AND U9481 ( .A(x[128]), .B(y[742]), .Z(n9116) );
  XNOR U9482 ( .A(n9117), .B(n9116), .Z(n9141) );
  XOR U9483 ( .A(n9142), .B(n9141), .Z(n9151) );
  XNOR U9484 ( .A(n9152), .B(n9151), .Z(n9154) );
  AND U9485 ( .A(y[741]), .B(x[129]), .Z(n9422) );
  NAND U9486 ( .A(x[133]), .B(y[737]), .Z(n9145) );
  XNOR U9487 ( .A(n9145), .B(o[102]), .Z(n9146) );
  XNOR U9488 ( .A(n9422), .B(n9146), .Z(n9148) );
  AND U9489 ( .A(y[738]), .B(x[132]), .Z(n9147) );
  XOR U9490 ( .A(n9148), .B(n9147), .Z(n9137) );
  AND U9491 ( .A(y[740]), .B(x[130]), .Z(n9451) );
  XNOR U9492 ( .A(n9136), .B(n9451), .Z(n9138) );
  XOR U9493 ( .A(n9137), .B(n9138), .Z(n9153) );
  XNOR U9494 ( .A(n9154), .B(n9153), .Z(n9131) );
  XOR U9495 ( .A(n9130), .B(n9131), .Z(n9132) );
  OR U9496 ( .A(n9119), .B(n9118), .Z(n9123) );
  OR U9497 ( .A(n9121), .B(n9120), .Z(n9122) );
  AND U9498 ( .A(n9123), .B(n9122), .Z(n9133) );
  XOR U9499 ( .A(n9126), .B(n9127), .Z(N231) );
  NANDN U9500 ( .A(n9125), .B(n9124), .Z(n9129) );
  NANDN U9501 ( .A(n9127), .B(n9126), .Z(n9128) );
  NAND U9502 ( .A(n9129), .B(n9128), .Z(n9186) );
  OR U9503 ( .A(n9131), .B(n9130), .Z(n9135) );
  NANDN U9504 ( .A(n9133), .B(n9132), .Z(n9134) );
  AND U9505 ( .A(n9135), .B(n9134), .Z(n9187) );
  XNOR U9506 ( .A(n9186), .B(n9187), .Z(n9188) );
  OR U9507 ( .A(n9136), .B(n9451), .Z(n9140) );
  NANDN U9508 ( .A(n9138), .B(n9137), .Z(n9139) );
  NAND U9509 ( .A(n9140), .B(n9139), .Z(n9183) );
  AND U9510 ( .A(y[742]), .B(x[134]), .Z(n9410) );
  NAND U9511 ( .A(n9710), .B(n9410), .Z(n9144) );
  OR U9512 ( .A(n9142), .B(n9141), .Z(n9143) );
  AND U9513 ( .A(n9144), .B(n9143), .Z(n9181) );
  ANDN U9514 ( .B(y[738]), .A(n156), .Z(n9319) );
  AND U9515 ( .A(y[742]), .B(x[129]), .Z(n9538) );
  NAND U9516 ( .A(x[134]), .B(y[737]), .Z(n9175) );
  XNOR U9517 ( .A(o[103]), .B(n9175), .Z(n9176) );
  XNOR U9518 ( .A(n9538), .B(n9176), .Z(n9177) );
  XNOR U9519 ( .A(n9319), .B(n9177), .Z(n9180) );
  XOR U9520 ( .A(n9181), .B(n9180), .Z(n9182) );
  XNOR U9521 ( .A(n9183), .B(n9182), .Z(n9192) );
  ANDN U9522 ( .B(y[741]), .A(n153), .Z(n9600) );
  ANDN U9523 ( .B(y[739]), .A(n155), .Z(n9341) );
  ANDN U9524 ( .B(y[740]), .A(n154), .Z(n9165) );
  XNOR U9525 ( .A(n9341), .B(n9165), .Z(n9166) );
  XOR U9526 ( .A(n9600), .B(n9166), .Z(n9169) );
  NAND U9527 ( .A(x[128]), .B(y[743]), .Z(n9161) );
  ANDN U9528 ( .B(o[102]), .A(n9145), .Z(n9160) );
  NAND U9529 ( .A(x[135]), .B(y[736]), .Z(n9159) );
  XOR U9530 ( .A(n9160), .B(n9159), .Z(n9162) );
  XNOR U9531 ( .A(n9161), .B(n9162), .Z(n9170) );
  XNOR U9532 ( .A(n9169), .B(n9170), .Z(n9172) );
  NAND U9533 ( .A(n9422), .B(n9146), .Z(n9150) );
  NANDN U9534 ( .A(n9148), .B(n9147), .Z(n9149) );
  AND U9535 ( .A(n9150), .B(n9149), .Z(n9171) );
  XOR U9536 ( .A(n9172), .B(n9171), .Z(n9193) );
  XOR U9537 ( .A(n9192), .B(n9193), .Z(n9195) );
  OR U9538 ( .A(n9152), .B(n9151), .Z(n9156) );
  OR U9539 ( .A(n9154), .B(n9153), .Z(n9155) );
  AND U9540 ( .A(n9156), .B(n9155), .Z(n9194) );
  XOR U9541 ( .A(n9195), .B(n9194), .Z(n9189) );
  XNOR U9542 ( .A(n9188), .B(n9189), .Z(N232) );
  AND U9543 ( .A(y[736]), .B(x[136]), .Z(n9158) );
  NAND U9544 ( .A(x[128]), .B(y[744]), .Z(n9157) );
  XOR U9545 ( .A(n9158), .B(n9157), .Z(n9207) );
  NAND U9546 ( .A(x[135]), .B(y[737]), .Z(n9210) );
  XNOR U9547 ( .A(n9210), .B(o[104]), .Z(n9206) );
  XOR U9548 ( .A(n9207), .B(n9206), .Z(n9227) );
  NANDN U9549 ( .A(n9160), .B(n9159), .Z(n9164) );
  NANDN U9550 ( .A(n9162), .B(n9161), .Z(n9163) );
  NAND U9551 ( .A(n9164), .B(n9163), .Z(n9226) );
  XOR U9552 ( .A(n9227), .B(n9226), .Z(n9228) );
  OR U9553 ( .A(n9165), .B(n9341), .Z(n9168) );
  OR U9554 ( .A(n9166), .B(n9600), .Z(n9167) );
  NAND U9555 ( .A(n9168), .B(n9167), .Z(n9229) );
  XNOR U9556 ( .A(n9228), .B(n9229), .Z(n9240) );
  OR U9557 ( .A(n9170), .B(n9169), .Z(n9174) );
  OR U9558 ( .A(n9172), .B(n9171), .Z(n9173) );
  AND U9559 ( .A(n9174), .B(n9173), .Z(n9222) );
  ANDN U9560 ( .B(y[738]), .A(n157), .Z(n9199) );
  XNOR U9561 ( .A(n9198), .B(n9199), .Z(n9200) );
  XNOR U9562 ( .A(n9200), .B(n9726), .Z(n9201) );
  ANDN U9563 ( .B(y[741]), .A(n154), .Z(n10021) );
  XNOR U9564 ( .A(n9201), .B(n10021), .Z(n9203) );
  NANDN U9565 ( .A(n9175), .B(o[103]), .Z(n9217) );
  AND U9566 ( .A(x[133]), .B(y[739]), .Z(n9845) );
  AND U9567 ( .A(y[743]), .B(x[129]), .Z(n9705) );
  XNOR U9568 ( .A(n9845), .B(n9705), .Z(n9216) );
  XOR U9569 ( .A(n9217), .B(n9216), .Z(n9202) );
  XNOR U9570 ( .A(n9203), .B(n9202), .Z(n9220) );
  NAND U9571 ( .A(n9538), .B(n9176), .Z(n9179) );
  NANDN U9572 ( .A(n9177), .B(n9319), .Z(n9178) );
  AND U9573 ( .A(n9179), .B(n9178), .Z(n9221) );
  XOR U9574 ( .A(n9220), .B(n9221), .Z(n9223) );
  XOR U9575 ( .A(n9222), .B(n9223), .Z(n9238) );
  NANDN U9576 ( .A(n9181), .B(n9180), .Z(n9185) );
  OR U9577 ( .A(n9183), .B(n9182), .Z(n9184) );
  NAND U9578 ( .A(n9185), .B(n9184), .Z(n9239) );
  XNOR U9579 ( .A(n9238), .B(n9239), .Z(n9241) );
  XNOR U9580 ( .A(n9240), .B(n9241), .Z(n9235) );
  NANDN U9581 ( .A(n9187), .B(n9186), .Z(n9191) );
  NAND U9582 ( .A(n9189), .B(n9188), .Z(n9190) );
  NAND U9583 ( .A(n9191), .B(n9190), .Z(n9232) );
  NANDN U9584 ( .A(n9193), .B(n9192), .Z(n9197) );
  OR U9585 ( .A(n9195), .B(n9194), .Z(n9196) );
  AND U9586 ( .A(n9197), .B(n9196), .Z(n9233) );
  XNOR U9587 ( .A(n9232), .B(n9233), .Z(n9234) );
  XOR U9588 ( .A(n9235), .B(n9234), .Z(N233) );
  OR U9589 ( .A(n9201), .B(n10021), .Z(n9205) );
  OR U9590 ( .A(n9203), .B(n9202), .Z(n9204) );
  NAND U9591 ( .A(n9205), .B(n9204), .Z(n9272) );
  XOR U9592 ( .A(n9273), .B(n9272), .Z(n9274) );
  AND U9593 ( .A(y[744]), .B(x[136]), .Z(n9723) );
  NAND U9594 ( .A(n9710), .B(n9723), .Z(n9209) );
  NANDN U9595 ( .A(n9207), .B(n9206), .Z(n9208) );
  NAND U9596 ( .A(n9209), .B(n9208), .Z(n9259) );
  NANDN U9597 ( .A(n9210), .B(o[104]), .Z(n9290) );
  AND U9598 ( .A(y[740]), .B(x[133]), .Z(n9211) );
  AND U9599 ( .A(y[738]), .B(x[135]), .Z(n9604) );
  XNOR U9600 ( .A(n9211), .B(n9604), .Z(n9289) );
  XOR U9601 ( .A(n9290), .B(n9289), .Z(n9257) );
  AND U9602 ( .A(y[736]), .B(x[137]), .Z(n9213) );
  NAND U9603 ( .A(x[128]), .B(y[745]), .Z(n9212) );
  XOR U9604 ( .A(n9213), .B(n9212), .Z(n9284) );
  NAND U9605 ( .A(x[136]), .B(y[737]), .Z(n9278) );
  XOR U9606 ( .A(n9278), .B(o[105]), .Z(n9283) );
  XNOR U9607 ( .A(n9284), .B(n9283), .Z(n9256) );
  XOR U9608 ( .A(n9257), .B(n9256), .Z(n9258) );
  XNOR U9609 ( .A(n9259), .B(n9258), .Z(n9268) );
  AND U9610 ( .A(y[741]), .B(x[132]), .Z(n9717) );
  AND U9611 ( .A(x[134]), .B(y[739]), .Z(n9215) );
  NAND U9612 ( .A(x[129]), .B(y[744]), .Z(n9214) );
  XNOR U9613 ( .A(n9215), .B(n9214), .Z(n9280) );
  XOR U9614 ( .A(n9717), .B(n9280), .Z(n9262) );
  ANDN U9615 ( .B(y[743]), .A(n153), .Z(n9917) );
  NAND U9616 ( .A(y[742]), .B(x[131]), .Z(n9631) );
  XOR U9617 ( .A(n9917), .B(n9631), .Z(n9263) );
  XNOR U9618 ( .A(n9262), .B(n9263), .Z(n9266) );
  NAND U9619 ( .A(x[129]), .B(y[739]), .Z(n9279) );
  AND U9620 ( .A(y[743]), .B(x[133]), .Z(n9412) );
  NANDN U9621 ( .A(n9279), .B(n9412), .Z(n9219) );
  OR U9622 ( .A(n9217), .B(n9216), .Z(n9218) );
  AND U9623 ( .A(n9219), .B(n9218), .Z(n9267) );
  XOR U9624 ( .A(n9266), .B(n9267), .Z(n9269) );
  XOR U9625 ( .A(n9268), .B(n9269), .Z(n9275) );
  NANDN U9626 ( .A(n9221), .B(n9220), .Z(n9225) );
  OR U9627 ( .A(n9223), .B(n9222), .Z(n9224) );
  NAND U9628 ( .A(n9225), .B(n9224), .Z(n9251) );
  OR U9629 ( .A(n9227), .B(n9226), .Z(n9231) );
  NANDN U9630 ( .A(n9229), .B(n9228), .Z(n9230) );
  NAND U9631 ( .A(n9231), .B(n9230), .Z(n9250) );
  XOR U9632 ( .A(n9251), .B(n9250), .Z(n9253) );
  XNOR U9633 ( .A(n9252), .B(n9253), .Z(n9247) );
  NANDN U9634 ( .A(n9233), .B(n9232), .Z(n9237) );
  NANDN U9635 ( .A(n9235), .B(n9234), .Z(n9236) );
  NAND U9636 ( .A(n9237), .B(n9236), .Z(n9244) );
  OR U9637 ( .A(n9239), .B(n9238), .Z(n9243) );
  OR U9638 ( .A(n9241), .B(n9240), .Z(n9242) );
  AND U9639 ( .A(n9243), .B(n9242), .Z(n9245) );
  XNOR U9640 ( .A(n9244), .B(n9245), .Z(n9246) );
  XOR U9641 ( .A(n9247), .B(n9246), .Z(N234) );
  NANDN U9642 ( .A(n9245), .B(n9244), .Z(n9249) );
  NANDN U9643 ( .A(n9247), .B(n9246), .Z(n9248) );
  NAND U9644 ( .A(n9249), .B(n9248), .Z(n9293) );
  OR U9645 ( .A(n9251), .B(n9250), .Z(n9255) );
  NAND U9646 ( .A(n9253), .B(n9252), .Z(n9254) );
  AND U9647 ( .A(n9255), .B(n9254), .Z(n9294) );
  XNOR U9648 ( .A(n9293), .B(n9294), .Z(n9295) );
  NANDN U9649 ( .A(n9257), .B(n9256), .Z(n9261) );
  OR U9650 ( .A(n9259), .B(n9258), .Z(n9260) );
  NAND U9651 ( .A(n9261), .B(n9260), .Z(n9353) );
  NANDN U9652 ( .A(n9917), .B(n9631), .Z(n9265) );
  OR U9653 ( .A(n9263), .B(n9262), .Z(n9264) );
  NAND U9654 ( .A(n9265), .B(n9264), .Z(n9352) );
  XOR U9655 ( .A(n9353), .B(n9352), .Z(n9354) );
  NANDN U9656 ( .A(n9267), .B(n9266), .Z(n9271) );
  NANDN U9657 ( .A(n9269), .B(n9268), .Z(n9270) );
  AND U9658 ( .A(n9271), .B(n9270), .Z(n9355) );
  XNOR U9659 ( .A(n9354), .B(n9355), .Z(n9301) );
  OR U9660 ( .A(n9273), .B(n9272), .Z(n9277) );
  NANDN U9661 ( .A(n9275), .B(n9274), .Z(n9276) );
  NAND U9662 ( .A(n9277), .B(n9276), .Z(n9300) );
  ANDN U9663 ( .B(y[746]), .A(n151), .Z(n9338) );
  NANDN U9664 ( .A(n9278), .B(o[105]), .Z(n9335) );
  ANDN U9665 ( .B(y[736]), .A(n161), .Z(n9336) );
  XNOR U9666 ( .A(n9338), .B(n9337), .Z(n9327) );
  ANDN U9667 ( .B(y[745]), .A(n152), .Z(n10230) );
  ANDN U9668 ( .B(y[743]), .A(n154), .Z(n10260) );
  IV U9669 ( .A(y[744]), .Z(n11414) );
  NANDN U9670 ( .A(n11414), .B(x[130]), .Z(n9315) );
  XNOR U9671 ( .A(n10260), .B(n9315), .Z(n9316) );
  XNOR U9672 ( .A(n10230), .B(n9316), .Z(n9325) );
  ANDN U9673 ( .B(y[744]), .A(n157), .Z(n9616) );
  NANDN U9674 ( .A(n9279), .B(n9616), .Z(n9282) );
  NAND U9675 ( .A(n9280), .B(n9717), .Z(n9281) );
  AND U9676 ( .A(n9282), .B(n9281), .Z(n9324) );
  XOR U9677 ( .A(n9325), .B(n9324), .Z(n9326) );
  XOR U9678 ( .A(n9327), .B(n9326), .Z(n9346) );
  ANDN U9679 ( .B(y[745]), .A(n160), .Z(n9984) );
  NAND U9680 ( .A(n9710), .B(n9984), .Z(n9286) );
  OR U9681 ( .A(n9284), .B(n9283), .Z(n9285) );
  NAND U9682 ( .A(n9286), .B(n9285), .Z(n9347) );
  XNOR U9683 ( .A(n9346), .B(n9347), .Z(n9349) );
  AND U9684 ( .A(y[738]), .B(x[136]), .Z(n9403) );
  XOR U9685 ( .A(n9403), .B(n9462), .Z(n9321) );
  NAND U9686 ( .A(x[137]), .B(y[737]), .Z(n9330) );
  XOR U9687 ( .A(o[106]), .B(n9330), .Z(n9320) );
  XOR U9688 ( .A(n9321), .B(n9320), .Z(n9305) );
  AND U9689 ( .A(y[740]), .B(x[134]), .Z(n9555) );
  AND U9690 ( .A(x[132]), .B(y[742]), .Z(n9288) );
  NAND U9691 ( .A(x[135]), .B(y[739]), .Z(n9287) );
  XOR U9692 ( .A(n9288), .B(n9287), .Z(n9343) );
  XNOR U9693 ( .A(n9555), .B(n9343), .Z(n9306) );
  XNOR U9694 ( .A(n9305), .B(n9306), .Z(n9308) );
  ANDN U9695 ( .B(y[740]), .A(n158), .Z(n9404) );
  NAND U9696 ( .A(n9319), .B(n9404), .Z(n9292) );
  OR U9697 ( .A(n9290), .B(n9289), .Z(n9291) );
  NAND U9698 ( .A(n9292), .B(n9291), .Z(n9307) );
  XOR U9699 ( .A(n9308), .B(n9307), .Z(n9348) );
  XOR U9700 ( .A(n9300), .B(n9299), .Z(n9302) );
  XNOR U9701 ( .A(n9301), .B(n9302), .Z(n9296) );
  XOR U9702 ( .A(n9295), .B(n9296), .Z(N235) );
  NANDN U9703 ( .A(n9294), .B(n9293), .Z(n9298) );
  NANDN U9704 ( .A(n9296), .B(n9295), .Z(n9297) );
  NAND U9705 ( .A(n9298), .B(n9297), .Z(n9358) );
  NANDN U9706 ( .A(n9300), .B(n9299), .Z(n9304) );
  OR U9707 ( .A(n9302), .B(n9301), .Z(n9303) );
  AND U9708 ( .A(n9304), .B(n9303), .Z(n9359) );
  XNOR U9709 ( .A(n9358), .B(n9359), .Z(n9360) );
  OR U9710 ( .A(n9306), .B(n9305), .Z(n9310) );
  OR U9711 ( .A(n9308), .B(n9307), .Z(n9309) );
  NAND U9712 ( .A(n9310), .B(n9309), .Z(n9373) );
  AND U9713 ( .A(y[744]), .B(x[131]), .Z(n10419) );
  AND U9714 ( .A(x[133]), .B(y[742]), .Z(n9312) );
  NAND U9715 ( .A(x[130]), .B(y[745]), .Z(n9311) );
  XOR U9716 ( .A(n9312), .B(n9311), .Z(n9419) );
  NAND U9717 ( .A(x[132]), .B(y[743]), .Z(n9418) );
  XNOR U9718 ( .A(n9419), .B(n9418), .Z(n9388) );
  XOR U9719 ( .A(n10419), .B(n9388), .Z(n9390) );
  AND U9720 ( .A(x[136]), .B(y[739]), .Z(n9314) );
  NAND U9721 ( .A(x[137]), .B(y[738]), .Z(n9313) );
  XNOR U9722 ( .A(n9314), .B(n9313), .Z(n9405) );
  XNOR U9723 ( .A(n9404), .B(n9405), .Z(n9389) );
  XOR U9724 ( .A(n9390), .B(n9389), .Z(n9396) );
  NANDN U9725 ( .A(n10260), .B(n9315), .Z(n9318) );
  NANDN U9726 ( .A(n10230), .B(n9316), .Z(n9317) );
  NAND U9727 ( .A(n9318), .B(n9317), .Z(n9393) );
  ANDN U9728 ( .B(y[741]), .A(n159), .Z(n10161) );
  NAND U9729 ( .A(n10161), .B(n9319), .Z(n9323) );
  OR U9730 ( .A(n9321), .B(n9320), .Z(n9322) );
  NAND U9731 ( .A(n9323), .B(n9322), .Z(n9394) );
  XNOR U9732 ( .A(n9396), .B(n9395), .Z(n9371) );
  OR U9733 ( .A(n9325), .B(n9324), .Z(n9329) );
  NAND U9734 ( .A(n9327), .B(n9326), .Z(n9328) );
  NAND U9735 ( .A(n9329), .B(n9328), .Z(n9379) );
  NANDN U9736 ( .A(n9330), .B(o[106]), .Z(n9400) );
  AND U9737 ( .A(y[736]), .B(x[139]), .Z(n9332) );
  NAND U9738 ( .A(x[128]), .B(y[747]), .Z(n9331) );
  XNOR U9739 ( .A(n9332), .B(n9331), .Z(n9399) );
  AND U9740 ( .A(y[741]), .B(x[134]), .Z(n9334) );
  NAND U9741 ( .A(x[129]), .B(y[746]), .Z(n9333) );
  XOR U9742 ( .A(n9334), .B(n9333), .Z(n9424) );
  NAND U9743 ( .A(x[138]), .B(y[737]), .Z(n9408) );
  XOR U9744 ( .A(o[107]), .B(n9408), .Z(n9423) );
  XOR U9745 ( .A(n9424), .B(n9423), .Z(n9382) );
  NANDN U9746 ( .A(n9336), .B(n9335), .Z(n9340) );
  OR U9747 ( .A(n9338), .B(n9337), .Z(n9339) );
  NAND U9748 ( .A(n9340), .B(n9339), .Z(n9385) );
  XOR U9749 ( .A(n9384), .B(n9385), .Z(n9376) );
  AND U9750 ( .A(y[742]), .B(x[135]), .Z(n9342) );
  NAND U9751 ( .A(n9342), .B(n9341), .Z(n9345) );
  NANDN U9752 ( .A(n9343), .B(n9555), .Z(n9344) );
  NAND U9753 ( .A(n9345), .B(n9344), .Z(n9377) );
  XOR U9754 ( .A(n9379), .B(n9378), .Z(n9370) );
  XOR U9755 ( .A(n9371), .B(n9370), .Z(n9372) );
  XOR U9756 ( .A(n9373), .B(n9372), .Z(n9364) );
  OR U9757 ( .A(n9347), .B(n9346), .Z(n9351) );
  NANDN U9758 ( .A(n9349), .B(n9348), .Z(n9350) );
  AND U9759 ( .A(n9351), .B(n9350), .Z(n9365) );
  XNOR U9760 ( .A(n9364), .B(n9365), .Z(n9367) );
  OR U9761 ( .A(n9353), .B(n9352), .Z(n9357) );
  NANDN U9762 ( .A(n9355), .B(n9354), .Z(n9356) );
  NAND U9763 ( .A(n9357), .B(n9356), .Z(n9366) );
  XOR U9764 ( .A(n9367), .B(n9366), .Z(n9361) );
  XNOR U9765 ( .A(n9360), .B(n9361), .Z(N236) );
  NANDN U9766 ( .A(n9359), .B(n9358), .Z(n9363) );
  NAND U9767 ( .A(n9361), .B(n9360), .Z(n9362) );
  NAND U9768 ( .A(n9363), .B(n9362), .Z(n9427) );
  OR U9769 ( .A(n9365), .B(n9364), .Z(n9369) );
  OR U9770 ( .A(n9367), .B(n9366), .Z(n9368) );
  AND U9771 ( .A(n9369), .B(n9368), .Z(n9428) );
  XNOR U9772 ( .A(n9427), .B(n9428), .Z(n9429) );
  NANDN U9773 ( .A(n9371), .B(n9370), .Z(n9375) );
  OR U9774 ( .A(n9373), .B(n9372), .Z(n9374) );
  NAND U9775 ( .A(n9375), .B(n9374), .Z(n9434) );
  NANDN U9776 ( .A(n9377), .B(n9376), .Z(n9381) );
  NANDN U9777 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND U9778 ( .A(n9381), .B(n9380), .Z(n9442) );
  NAND U9779 ( .A(n9383), .B(n9382), .Z(n9387) );
  NANDN U9780 ( .A(n9385), .B(n9384), .Z(n9386) );
  NAND U9781 ( .A(n9387), .B(n9386), .Z(n9440) );
  NANDN U9782 ( .A(n9388), .B(n10419), .Z(n9392) );
  OR U9783 ( .A(n9390), .B(n9389), .Z(n9391) );
  AND U9784 ( .A(n9392), .B(n9391), .Z(n9439) );
  XNOR U9785 ( .A(n9442), .B(n9441), .Z(n9433) );
  XNOR U9786 ( .A(n9434), .B(n9433), .Z(n9436) );
  NANDN U9787 ( .A(n9394), .B(n9393), .Z(n9398) );
  NANDN U9788 ( .A(n9396), .B(n9395), .Z(n9397) );
  NAND U9789 ( .A(n9398), .B(n9397), .Z(n9501) );
  ANDN U9790 ( .B(y[747]), .A(n162), .Z(n10560) );
  NAND U9791 ( .A(n9710), .B(n10560), .Z(n9402) );
  NANDN U9792 ( .A(n9400), .B(n9399), .Z(n9401) );
  NAND U9793 ( .A(n9402), .B(n9401), .Z(n9475) );
  NAND U9794 ( .A(x[137]), .B(y[739]), .Z(n10110) );
  NANDN U9795 ( .A(n10110), .B(n9403), .Z(n9407) );
  NAND U9796 ( .A(n9405), .B(n9404), .Z(n9406) );
  NAND U9797 ( .A(n9407), .B(n9406), .Z(n9473) );
  NANDN U9798 ( .A(n9408), .B(o[107]), .Z(n9480) );
  NAND U9799 ( .A(x[129]), .B(y[747]), .Z(n9409) );
  XNOR U9800 ( .A(n9410), .B(n9409), .Z(n9479) );
  XOR U9801 ( .A(n9473), .B(n9474), .Z(n9476) );
  NAND U9802 ( .A(x[135]), .B(y[741]), .Z(n9411) );
  XOR U9803 ( .A(n9412), .B(n9411), .Z(n9464) );
  AND U9804 ( .A(y[738]), .B(x[138]), .Z(n9413) );
  XOR U9805 ( .A(n9413), .B(n10110), .Z(n9492) );
  NAND U9806 ( .A(x[132]), .B(y[744]), .Z(n9491) );
  XNOR U9807 ( .A(n9492), .B(n9491), .Z(n9463) );
  XOR U9808 ( .A(n9464), .B(n9463), .Z(n9469) );
  AND U9809 ( .A(y[736]), .B(x[140]), .Z(n9415) );
  NAND U9810 ( .A(x[128]), .B(y[748]), .Z(n9414) );
  XOR U9811 ( .A(n9415), .B(n9414), .Z(n9484) );
  NAND U9812 ( .A(x[139]), .B(y[737]), .Z(n9458) );
  XOR U9813 ( .A(o[108]), .B(n9458), .Z(n9483) );
  XOR U9814 ( .A(n9484), .B(n9483), .Z(n9467) );
  AND U9815 ( .A(y[740]), .B(x[136]), .Z(n9417) );
  NAND U9816 ( .A(x[130]), .B(y[746]), .Z(n9416) );
  XOR U9817 ( .A(n9417), .B(n9416), .Z(n9453) );
  NAND U9818 ( .A(x[131]), .B(y[745]), .Z(n9452) );
  XNOR U9819 ( .A(n9453), .B(n9452), .Z(n9468) );
  XOR U9820 ( .A(n9467), .B(n9468), .Z(n9470) );
  ANDN U9821 ( .B(y[745]), .A(n156), .Z(n9632) );
  NAND U9822 ( .A(n9726), .B(n9632), .Z(n9421) );
  OR U9823 ( .A(n9419), .B(n9418), .Z(n9420) );
  NAND U9824 ( .A(n9421), .B(n9420), .Z(n9446) );
  AND U9825 ( .A(y[746]), .B(x[134]), .Z(n9716) );
  NAND U9826 ( .A(n9716), .B(n9422), .Z(n9426) );
  OR U9827 ( .A(n9424), .B(n9423), .Z(n9425) );
  NAND U9828 ( .A(n9426), .B(n9425), .Z(n9445) );
  XOR U9829 ( .A(n9446), .B(n9445), .Z(n9448) );
  XNOR U9830 ( .A(n9447), .B(n9448), .Z(n9500) );
  XOR U9831 ( .A(n9499), .B(n9500), .Z(n9502) );
  XOR U9832 ( .A(n9501), .B(n9502), .Z(n9435) );
  XNOR U9833 ( .A(n9436), .B(n9435), .Z(n9430) );
  XOR U9834 ( .A(n9429), .B(n9430), .Z(N237) );
  NANDN U9835 ( .A(n9428), .B(n9427), .Z(n9432) );
  NANDN U9836 ( .A(n9430), .B(n9429), .Z(n9431) );
  NAND U9837 ( .A(n9432), .B(n9431), .Z(n9570) );
  OR U9838 ( .A(n9434), .B(n9433), .Z(n9438) );
  OR U9839 ( .A(n9436), .B(n9435), .Z(n9437) );
  AND U9840 ( .A(n9438), .B(n9437), .Z(n9571) );
  XNOR U9841 ( .A(n9570), .B(n9571), .Z(n9572) );
  NANDN U9842 ( .A(n9440), .B(n9439), .Z(n9444) );
  NAND U9843 ( .A(n9442), .B(n9441), .Z(n9443) );
  NAND U9844 ( .A(n9444), .B(n9443), .Z(n9579) );
  OR U9845 ( .A(n9446), .B(n9445), .Z(n9450) );
  NAND U9846 ( .A(n9448), .B(n9447), .Z(n9449) );
  AND U9847 ( .A(n9450), .B(n9449), .Z(n9511) );
  AND U9848 ( .A(y[746]), .B(x[136]), .Z(n9906) );
  NAND U9849 ( .A(n9906), .B(n9451), .Z(n9455) );
  OR U9850 ( .A(n9453), .B(n9452), .Z(n9454) );
  NAND U9851 ( .A(n9455), .B(n9454), .Z(n9532) );
  AND U9852 ( .A(y[743]), .B(x[134]), .Z(n9457) );
  NAND U9853 ( .A(x[137]), .B(y[740]), .Z(n9456) );
  XOR U9854 ( .A(n9457), .B(n9456), .Z(n9557) );
  NAND U9855 ( .A(x[130]), .B(y[747]), .Z(n9556) );
  XOR U9856 ( .A(n9557), .B(n9556), .Z(n9530) );
  NANDN U9857 ( .A(n9458), .B(o[108]), .Z(n9541) );
  AND U9858 ( .A(y[748]), .B(x[129]), .Z(n9460) );
  NAND U9859 ( .A(x[135]), .B(y[742]), .Z(n9459) );
  XNOR U9860 ( .A(n9460), .B(n9459), .Z(n9540) );
  XNOR U9861 ( .A(n9532), .B(n9531), .Z(n9506) );
  AND U9862 ( .A(y[743]), .B(x[135]), .Z(n9461) );
  NANDN U9863 ( .A(n9462), .B(n9461), .Z(n9466) );
  OR U9864 ( .A(n9464), .B(n9463), .Z(n9465) );
  AND U9865 ( .A(n9466), .B(n9465), .Z(n9505) );
  XOR U9866 ( .A(n9506), .B(n9505), .Z(n9507) );
  NANDN U9867 ( .A(n9468), .B(n9467), .Z(n9472) );
  NANDN U9868 ( .A(n9470), .B(n9469), .Z(n9471) );
  AND U9869 ( .A(n9472), .B(n9471), .Z(n9508) );
  XNOR U9870 ( .A(n9507), .B(n9508), .Z(n9512) );
  XOR U9871 ( .A(n9511), .B(n9512), .Z(n9513) );
  NANDN U9872 ( .A(n9474), .B(n9473), .Z(n9478) );
  NANDN U9873 ( .A(n9476), .B(n9475), .Z(n9477) );
  NAND U9874 ( .A(n9478), .B(n9477), .Z(n9520) );
  ANDN U9875 ( .B(y[747]), .A(n157), .Z(n9924) );
  NAND U9876 ( .A(n9538), .B(n9924), .Z(n9482) );
  NANDN U9877 ( .A(n9480), .B(n9479), .Z(n9481) );
  NAND U9878 ( .A(n9482), .B(n9481), .Z(n9525) );
  ANDN U9879 ( .B(y[748]), .A(n163), .Z(n10754) );
  NAND U9880 ( .A(n9710), .B(n10754), .Z(n9486) );
  OR U9881 ( .A(n9484), .B(n9483), .Z(n9485) );
  NAND U9882 ( .A(n9486), .B(n9485), .Z(n9523) );
  AND U9883 ( .A(y[738]), .B(x[139]), .Z(n9488) );
  NAND U9884 ( .A(x[138]), .B(y[739]), .Z(n9487) );
  XNOR U9885 ( .A(n9488), .B(n9487), .Z(n9544) );
  XNOR U9886 ( .A(n10161), .B(n9544), .Z(n9524) );
  XOR U9887 ( .A(n9525), .B(n9526), .Z(n9517) );
  AND U9888 ( .A(y[738]), .B(x[137]), .Z(n9490) );
  AND U9889 ( .A(y[739]), .B(x[138]), .Z(n9489) );
  NAND U9890 ( .A(n9490), .B(n9489), .Z(n9494) );
  OR U9891 ( .A(n9492), .B(n9491), .Z(n9493) );
  NAND U9892 ( .A(n9494), .B(n9493), .Z(n9567) );
  AND U9893 ( .A(y[736]), .B(x[141]), .Z(n9496) );
  NAND U9894 ( .A(x[128]), .B(y[749]), .Z(n9495) );
  XOR U9895 ( .A(n9496), .B(n9495), .Z(n9552) );
  NAND U9896 ( .A(x[140]), .B(y[737]), .Z(n9561) );
  XOR U9897 ( .A(o[109]), .B(n9561), .Z(n9551) );
  XOR U9898 ( .A(n9552), .B(n9551), .Z(n9565) );
  AND U9899 ( .A(x[131]), .B(y[746]), .Z(n9498) );
  NAND U9900 ( .A(x[133]), .B(y[744]), .Z(n9497) );
  XOR U9901 ( .A(n9498), .B(n9497), .Z(n9548) );
  NAND U9902 ( .A(x[132]), .B(y[745]), .Z(n9547) );
  XOR U9903 ( .A(n9548), .B(n9547), .Z(n9564) );
  XOR U9904 ( .A(n9567), .B(n9566), .Z(n9518) );
  XNOR U9905 ( .A(n9517), .B(n9518), .Z(n9519) );
  XOR U9906 ( .A(n9520), .B(n9519), .Z(n9514) );
  XNOR U9907 ( .A(n9513), .B(n9514), .Z(n9576) );
  NANDN U9908 ( .A(n9500), .B(n9499), .Z(n9504) );
  NANDN U9909 ( .A(n9502), .B(n9501), .Z(n9503) );
  NAND U9910 ( .A(n9504), .B(n9503), .Z(n9577) );
  XOR U9911 ( .A(n9576), .B(n9577), .Z(n9578) );
  XNOR U9912 ( .A(n9579), .B(n9578), .Z(n9573) );
  XOR U9913 ( .A(n9572), .B(n9573), .Z(N238) );
  OR U9914 ( .A(n9506), .B(n9505), .Z(n9510) );
  NANDN U9915 ( .A(n9508), .B(n9507), .Z(n9509) );
  NAND U9916 ( .A(n9510), .B(n9509), .Z(n9591) );
  OR U9917 ( .A(n9512), .B(n9511), .Z(n9516) );
  NANDN U9918 ( .A(n9514), .B(n9513), .Z(n9515) );
  AND U9919 ( .A(n9516), .B(n9515), .Z(n9588) );
  NANDN U9920 ( .A(n9518), .B(n9517), .Z(n9522) );
  NANDN U9921 ( .A(n9520), .B(n9519), .Z(n9521) );
  AND U9922 ( .A(n9522), .B(n9521), .Z(n9667) );
  NANDN U9923 ( .A(n9524), .B(n9523), .Z(n9528) );
  NANDN U9924 ( .A(n9526), .B(n9525), .Z(n9527) );
  NAND U9925 ( .A(n9528), .B(n9527), .Z(n9596) );
  NAND U9926 ( .A(n9530), .B(n9529), .Z(n9534) );
  NAND U9927 ( .A(n9532), .B(n9531), .Z(n9533) );
  NAND U9928 ( .A(n9534), .B(n9533), .Z(n9594) );
  ANDN U9929 ( .B(y[746]), .A(n155), .Z(n9647) );
  AND U9930 ( .A(y[740]), .B(x[138]), .Z(n10266) );
  AND U9931 ( .A(y[741]), .B(x[137]), .Z(n10224) );
  NAND U9932 ( .A(x[130]), .B(y[748]), .Z(n9535) );
  XOR U9933 ( .A(n10224), .B(n9535), .Z(n9601) );
  XNOR U9934 ( .A(n10266), .B(n9601), .Z(n9646) );
  XOR U9935 ( .A(n9647), .B(n9646), .Z(n9649) );
  AND U9936 ( .A(y[747]), .B(x[131]), .Z(n9537) );
  NAND U9937 ( .A(x[136]), .B(y[742]), .Z(n9536) );
  XOR U9938 ( .A(n9537), .B(n9536), .Z(n9633) );
  XOR U9939 ( .A(n9632), .B(n9633), .Z(n9648) );
  AND U9940 ( .A(y[748]), .B(x[135]), .Z(n9539) );
  NAND U9941 ( .A(n9539), .B(n9538), .Z(n9543) );
  NANDN U9942 ( .A(n9541), .B(n9540), .Z(n9542) );
  NAND U9943 ( .A(n9543), .B(n9542), .Z(n9652) );
  NAND U9944 ( .A(x[138]), .B(y[738]), .Z(n10166) );
  ANDN U9945 ( .B(y[739]), .A(n162), .Z(n9749) );
  NANDN U9946 ( .A(n10166), .B(n9749), .Z(n9546) );
  NAND U9947 ( .A(n9544), .B(n10161), .Z(n9545) );
  AND U9948 ( .A(n9546), .B(n9545), .Z(n9653) );
  XOR U9949 ( .A(n9655), .B(n9654), .Z(n9595) );
  XOR U9950 ( .A(n9596), .B(n9597), .Z(n9664) );
  ANDN U9951 ( .B(y[746]), .A(n156), .Z(n9700) );
  NAND U9952 ( .A(n9700), .B(n10419), .Z(n9550) );
  OR U9953 ( .A(n9548), .B(n9547), .Z(n9549) );
  NAND U9954 ( .A(n9550), .B(n9549), .Z(n9627) );
  XOR U9955 ( .A(n9749), .B(n9614), .Z(n9615) );
  XOR U9956 ( .A(n9616), .B(n9615), .Z(n9626) );
  AND U9957 ( .A(x[141]), .B(y[749]), .Z(n11149) );
  NAND U9958 ( .A(n9710), .B(n11149), .Z(n9554) );
  OR U9959 ( .A(n9552), .B(n9551), .Z(n9553) );
  AND U9960 ( .A(n9554), .B(n9553), .Z(n9625) );
  XNOR U9961 ( .A(n9626), .B(n9625), .Z(n9628) );
  XOR U9962 ( .A(n9627), .B(n9628), .Z(n9660) );
  AND U9963 ( .A(y[743]), .B(x[137]), .Z(n9755) );
  NAND U9964 ( .A(n9755), .B(n9555), .Z(n9559) );
  OR U9965 ( .A(n9557), .B(n9556), .Z(n9558) );
  AND U9966 ( .A(n9559), .B(n9558), .Z(n9622) );
  NAND U9967 ( .A(x[141]), .B(y[737]), .Z(n9611) );
  XOR U9968 ( .A(o[110]), .B(n9611), .Z(n9606) );
  AND U9969 ( .A(y[738]), .B(x[140]), .Z(n10219) );
  NAND U9970 ( .A(x[135]), .B(y[743]), .Z(n9560) );
  XNOR U9971 ( .A(n10219), .B(n9560), .Z(n9605) );
  NANDN U9972 ( .A(n9561), .B(o[109]), .Z(n9637) );
  AND U9973 ( .A(y[750]), .B(x[128]), .Z(n9563) );
  AND U9974 ( .A(y[736]), .B(x[142]), .Z(n9562) );
  XNOR U9975 ( .A(n9563), .B(n9562), .Z(n9636) );
  XOR U9976 ( .A(n9637), .B(n9636), .Z(n9619) );
  XOR U9977 ( .A(n9622), .B(n9621), .Z(n9658) );
  NAND U9978 ( .A(n9565), .B(n9564), .Z(n9569) );
  NAND U9979 ( .A(n9567), .B(n9566), .Z(n9568) );
  NAND U9980 ( .A(n9569), .B(n9568), .Z(n9659) );
  XOR U9981 ( .A(n9658), .B(n9659), .Z(n9661) );
  XNOR U9982 ( .A(n9660), .B(n9661), .Z(n9665) );
  XOR U9983 ( .A(n9667), .B(n9666), .Z(n9589) );
  XNOR U9984 ( .A(n9588), .B(n9589), .Z(n9590) );
  XNOR U9985 ( .A(n9591), .B(n9590), .Z(n9585) );
  NANDN U9986 ( .A(n9571), .B(n9570), .Z(n9575) );
  NANDN U9987 ( .A(n9573), .B(n9572), .Z(n9574) );
  NAND U9988 ( .A(n9575), .B(n9574), .Z(n9582) );
  OR U9989 ( .A(n9577), .B(n9576), .Z(n9581) );
  NANDN U9990 ( .A(n9579), .B(n9578), .Z(n9580) );
  NAND U9991 ( .A(n9581), .B(n9580), .Z(n9583) );
  XNOR U9992 ( .A(n9582), .B(n9583), .Z(n9584) );
  XOR U9993 ( .A(n9585), .B(n9584), .Z(N239) );
  NANDN U9994 ( .A(n9583), .B(n9582), .Z(n9587) );
  NANDN U9995 ( .A(n9585), .B(n9584), .Z(n9586) );
  NAND U9996 ( .A(n9587), .B(n9586), .Z(n9670) );
  OR U9997 ( .A(n9589), .B(n9588), .Z(n9593) );
  OR U9998 ( .A(n9591), .B(n9590), .Z(n9592) );
  AND U9999 ( .A(n9593), .B(n9592), .Z(n9671) );
  XNOR U10000 ( .A(n9670), .B(n9671), .Z(n9672) );
  NANDN U10001 ( .A(n9595), .B(n9594), .Z(n9599) );
  NANDN U10002 ( .A(n9597), .B(n9596), .Z(n9598) );
  NAND U10003 ( .A(n9599), .B(n9598), .Z(n9761) );
  ANDN U10004 ( .B(y[748]), .A(n160), .Z(n10362) );
  NAND U10005 ( .A(n9600), .B(n10362), .Z(n9603) );
  NANDN U10006 ( .A(n9601), .B(n10266), .Z(n9602) );
  AND U10007 ( .A(n9603), .B(n9602), .Z(n9688) );
  AND U10008 ( .A(y[743]), .B(x[140]), .Z(n9989) );
  NAND U10009 ( .A(n9604), .B(n9989), .Z(n9608) );
  NANDN U10010 ( .A(n9606), .B(n9605), .Z(n9607) );
  NAND U10011 ( .A(n9608), .B(n9607), .Z(n9740) );
  AND U10012 ( .A(x[140]), .B(y[739]), .Z(n9610) );
  NAND U10013 ( .A(x[139]), .B(y[740]), .Z(n9609) );
  XOR U10014 ( .A(n9610), .B(n9609), .Z(n9751) );
  NAND U10015 ( .A(x[141]), .B(y[738]), .Z(n9750) );
  XOR U10016 ( .A(n9751), .B(n9750), .Z(n9737) );
  NANDN U10017 ( .A(n9611), .B(o[110]), .Z(n9712) );
  AND U10018 ( .A(y[736]), .B(x[143]), .Z(n9613) );
  NAND U10019 ( .A(x[128]), .B(y[751]), .Z(n9612) );
  XOR U10020 ( .A(n9613), .B(n9612), .Z(n9711) );
  XOR U10021 ( .A(n9712), .B(n9711), .Z(n9738) );
  XNOR U10022 ( .A(n9737), .B(n9738), .Z(n9739) );
  XOR U10023 ( .A(n9740), .B(n9739), .Z(n9689) );
  XOR U10024 ( .A(n9688), .B(n9689), .Z(n9690) );
  NANDN U10025 ( .A(n9749), .B(n9614), .Z(n9618) );
  OR U10026 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U10027 ( .A(n9618), .B(n9617), .Z(n9691) );
  NAND U10028 ( .A(n9620), .B(n9619), .Z(n9624) );
  NANDN U10029 ( .A(n9622), .B(n9621), .Z(n9623) );
  AND U10030 ( .A(n9624), .B(n9623), .Z(n9682) );
  XNOR U10031 ( .A(n9683), .B(n9682), .Z(n9685) );
  OR U10032 ( .A(n9626), .B(n9625), .Z(n9630) );
  NANDN U10033 ( .A(n9628), .B(n9627), .Z(n9629) );
  AND U10034 ( .A(n9630), .B(n9629), .Z(n9684) );
  XOR U10035 ( .A(n9685), .B(n9684), .Z(n9759) );
  NAND U10036 ( .A(x[136]), .B(y[747]), .Z(n10030) );
  OR U10037 ( .A(n10030), .B(n9631), .Z(n9635) );
  NANDN U10038 ( .A(n9633), .B(n9632), .Z(n9634) );
  NAND U10039 ( .A(n9635), .B(n9634), .Z(n9732) );
  AND U10040 ( .A(y[750]), .B(x[142]), .Z(n11417) );
  NAND U10041 ( .A(n9710), .B(n11417), .Z(n9639) );
  OR U10042 ( .A(n9637), .B(n9636), .Z(n9638) );
  NAND U10043 ( .A(n9639), .B(n9638), .Z(n9731) );
  XOR U10044 ( .A(n9732), .B(n9731), .Z(n9733) );
  NAND U10045 ( .A(x[135]), .B(y[744]), .Z(n10125) );
  AND U10046 ( .A(y[741]), .B(x[138]), .Z(n9641) );
  NAND U10047 ( .A(x[132]), .B(y[747]), .Z(n9640) );
  XNOR U10048 ( .A(n9641), .B(n9640), .Z(n9718) );
  XNOR U10049 ( .A(n10125), .B(n9718), .Z(n9701) );
  NAND U10050 ( .A(x[134]), .B(y[745]), .Z(n9828) );
  XOR U10051 ( .A(n9700), .B(n9828), .Z(n9702) );
  XNOR U10052 ( .A(n9701), .B(n9702), .Z(n9746) );
  AND U10053 ( .A(y[737]), .B(x[142]), .Z(n9721) );
  XNOR U10054 ( .A(o[111]), .B(n9721), .Z(n9707) );
  AND U10055 ( .A(y[743]), .B(x[136]), .Z(n9643) );
  NAND U10056 ( .A(x[129]), .B(y[750]), .Z(n9642) );
  XNOR U10057 ( .A(n9643), .B(n9642), .Z(n9706) );
  XNOR U10058 ( .A(n9707), .B(n9706), .Z(n9743) );
  NAND U10059 ( .A(x[131]), .B(y[748]), .Z(n9728) );
  AND U10060 ( .A(x[137]), .B(y[742]), .Z(n9645) );
  NAND U10061 ( .A(x[130]), .B(y[749]), .Z(n9644) );
  XOR U10062 ( .A(n9645), .B(n9644), .Z(n9727) );
  XOR U10063 ( .A(n9728), .B(n9727), .Z(n9744) );
  XNOR U10064 ( .A(n9743), .B(n9744), .Z(n9745) );
  XNOR U10065 ( .A(n9746), .B(n9745), .Z(n9734) );
  OR U10066 ( .A(n9647), .B(n9646), .Z(n9651) );
  NAND U10067 ( .A(n9649), .B(n9648), .Z(n9650) );
  NAND U10068 ( .A(n9651), .B(n9650), .Z(n9695) );
  XNOR U10069 ( .A(n9694), .B(n9695), .Z(n9697) );
  NANDN U10070 ( .A(n9653), .B(n9652), .Z(n9657) );
  NANDN U10071 ( .A(n9655), .B(n9654), .Z(n9656) );
  AND U10072 ( .A(n9657), .B(n9656), .Z(n9696) );
  XOR U10073 ( .A(n9697), .B(n9696), .Z(n9758) );
  XOR U10074 ( .A(n9759), .B(n9758), .Z(n9760) );
  XOR U10075 ( .A(n9761), .B(n9760), .Z(n9676) );
  NANDN U10076 ( .A(n9659), .B(n9658), .Z(n9663) );
  NANDN U10077 ( .A(n9661), .B(n9660), .Z(n9662) );
  NAND U10078 ( .A(n9663), .B(n9662), .Z(n9677) );
  NAND U10079 ( .A(n9665), .B(n9664), .Z(n9669) );
  NANDN U10080 ( .A(n9667), .B(n9666), .Z(n9668) );
  NAND U10081 ( .A(n9669), .B(n9668), .Z(n9679) );
  XNOR U10082 ( .A(n9678), .B(n9679), .Z(n9673) );
  XOR U10083 ( .A(n9672), .B(n9673), .Z(N240) );
  NANDN U10084 ( .A(n9671), .B(n9670), .Z(n9675) );
  NANDN U10085 ( .A(n9673), .B(n9672), .Z(n9674) );
  NAND U10086 ( .A(n9675), .B(n9674), .Z(n9764) );
  NANDN U10087 ( .A(n9677), .B(n9676), .Z(n9681) );
  NANDN U10088 ( .A(n9679), .B(n9678), .Z(n9680) );
  NAND U10089 ( .A(n9681), .B(n9680), .Z(n9765) );
  XNOR U10090 ( .A(n9764), .B(n9765), .Z(n9766) );
  OR U10091 ( .A(n9683), .B(n9682), .Z(n9687) );
  OR U10092 ( .A(n9685), .B(n9684), .Z(n9686) );
  NAND U10093 ( .A(n9687), .B(n9686), .Z(n9855) );
  OR U10094 ( .A(n9689), .B(n9688), .Z(n9693) );
  NANDN U10095 ( .A(n9691), .B(n9690), .Z(n9692) );
  NAND U10096 ( .A(n9693), .B(n9692), .Z(n9853) );
  OR U10097 ( .A(n9695), .B(n9694), .Z(n9699) );
  OR U10098 ( .A(n9697), .B(n9696), .Z(n9698) );
  NAND U10099 ( .A(n9699), .B(n9698), .Z(n9852) );
  XOR U10100 ( .A(n9853), .B(n9852), .Z(n9854) );
  XNOR U10101 ( .A(n9855), .B(n9854), .Z(n9773) );
  NANDN U10102 ( .A(n9700), .B(n9828), .Z(n9704) );
  OR U10103 ( .A(n9702), .B(n9701), .Z(n9703) );
  AND U10104 ( .A(n9704), .B(n9703), .Z(n9810) );
  NAND U10105 ( .A(x[136]), .B(y[750]), .Z(n10706) );
  NANDN U10106 ( .A(n10706), .B(n9705), .Z(n9709) );
  NANDN U10107 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U10108 ( .A(n9709), .B(n9708), .Z(n9776) );
  NAND U10109 ( .A(y[751]), .B(x[143]), .Z(n11759) );
  NANDN U10110 ( .A(n11759), .B(n9710), .Z(n9714) );
  OR U10111 ( .A(n9712), .B(n9711), .Z(n9713) );
  AND U10112 ( .A(n9714), .B(n9713), .Z(n9777) );
  NAND U10113 ( .A(x[128]), .B(y[752]), .Z(n9840) );
  AND U10114 ( .A(y[736]), .B(x[144]), .Z(n9839) );
  XNOR U10115 ( .A(n9840), .B(n9839), .Z(n9842) );
  NAND U10116 ( .A(x[143]), .B(y[737]), .Z(n9849) );
  XNOR U10117 ( .A(n9849), .B(o[112]), .Z(n9841) );
  XNOR U10118 ( .A(n9842), .B(n9841), .Z(n9823) );
  NAND U10119 ( .A(x[135]), .B(y[745]), .Z(n9715) );
  XOR U10120 ( .A(n9716), .B(n9715), .Z(n9830) );
  NAND U10121 ( .A(x[138]), .B(y[742]), .Z(n9829) );
  XNOR U10122 ( .A(n9830), .B(n9829), .Z(n9822) );
  XNOR U10123 ( .A(n9823), .B(n9822), .Z(n9825) );
  ANDN U10124 ( .B(y[747]), .A(n161), .Z(n10408) );
  NAND U10125 ( .A(n9717), .B(n10408), .Z(n9720) );
  NANDN U10126 ( .A(n10125), .B(n9718), .Z(n9719) );
  AND U10127 ( .A(n9720), .B(n9719), .Z(n9824) );
  XOR U10128 ( .A(n9825), .B(n9824), .Z(n9779) );
  XOR U10129 ( .A(n9778), .B(n9779), .Z(n9811) );
  XOR U10130 ( .A(n9810), .B(n9811), .Z(n9812) );
  NAND U10131 ( .A(n9721), .B(o[111]), .Z(n9834) );
  NAND U10132 ( .A(x[129]), .B(y[751]), .Z(n9722) );
  XOR U10133 ( .A(n9723), .B(n9722), .Z(n9833) );
  XNOR U10134 ( .A(n9834), .B(n9833), .Z(n9818) );
  AND U10135 ( .A(y[741]), .B(x[139]), .Z(n9725) );
  NAND U10136 ( .A(x[142]), .B(y[738]), .Z(n9724) );
  XOR U10137 ( .A(n9725), .B(n9724), .Z(n9789) );
  NAND U10138 ( .A(x[132]), .B(y[748]), .Z(n9788) );
  XOR U10139 ( .A(n9789), .B(n9788), .Z(n9817) );
  ANDN U10140 ( .B(y[749]), .A(n160), .Z(n10519) );
  NAND U10141 ( .A(n9726), .B(n10519), .Z(n9730) );
  OR U10142 ( .A(n9728), .B(n9727), .Z(n9729) );
  NAND U10143 ( .A(n9730), .B(n9729), .Z(n9816) );
  XNOR U10144 ( .A(n9817), .B(n9816), .Z(n9819) );
  XOR U10145 ( .A(n9818), .B(n9819), .Z(n9813) );
  XOR U10146 ( .A(n9812), .B(n9813), .Z(n9805) );
  OR U10147 ( .A(n9732), .B(n9731), .Z(n9736) );
  NANDN U10148 ( .A(n9734), .B(n9733), .Z(n9735) );
  AND U10149 ( .A(n9736), .B(n9735), .Z(n9804) );
  XOR U10150 ( .A(n9805), .B(n9804), .Z(n9806) );
  OR U10151 ( .A(n9738), .B(n9737), .Z(n9742) );
  OR U10152 ( .A(n9740), .B(n9739), .Z(n9741) );
  AND U10153 ( .A(n9742), .B(n9741), .Z(n9801) );
  OR U10154 ( .A(n9744), .B(n9743), .Z(n9748) );
  OR U10155 ( .A(n9746), .B(n9745), .Z(n9747) );
  AND U10156 ( .A(n9748), .B(n9747), .Z(n9798) );
  NAND U10157 ( .A(x[140]), .B(y[740]), .Z(n10523) );
  NANDN U10158 ( .A(n10523), .B(n9749), .Z(n9753) );
  OR U10159 ( .A(n9751), .B(n9750), .Z(n9752) );
  NAND U10160 ( .A(n9753), .B(n9752), .Z(n9795) );
  NAND U10161 ( .A(x[130]), .B(y[750]), .Z(n9754) );
  XOR U10162 ( .A(n9755), .B(n9754), .Z(n9784) );
  NAND U10163 ( .A(y[749]), .B(x[131]), .Z(n9783) );
  XOR U10164 ( .A(n9784), .B(n9783), .Z(n9793) );
  AND U10165 ( .A(x[141]), .B(y[739]), .Z(n9757) );
  AND U10166 ( .A(y[747]), .B(x[133]), .Z(n9756) );
  XNOR U10167 ( .A(n9757), .B(n9756), .Z(n9846) );
  XOR U10168 ( .A(n10523), .B(n9846), .Z(n9792) );
  XOR U10169 ( .A(n9795), .B(n9794), .Z(n9799) );
  XOR U10170 ( .A(n9798), .B(n9799), .Z(n9800) );
  XNOR U10171 ( .A(n9806), .B(n9807), .Z(n9770) );
  OR U10172 ( .A(n9759), .B(n9758), .Z(n9763) );
  NANDN U10173 ( .A(n9761), .B(n9760), .Z(n9762) );
  NAND U10174 ( .A(n9763), .B(n9762), .Z(n9771) );
  XOR U10175 ( .A(n9770), .B(n9771), .Z(n9772) );
  XNOR U10176 ( .A(n9773), .B(n9772), .Z(n9767) );
  XOR U10177 ( .A(n9766), .B(n9767), .Z(N241) );
  NANDN U10178 ( .A(n9765), .B(n9764), .Z(n9769) );
  NANDN U10179 ( .A(n9767), .B(n9766), .Z(n9768) );
  NAND U10180 ( .A(n9769), .B(n9768), .Z(n9858) );
  OR U10181 ( .A(n9771), .B(n9770), .Z(n9775) );
  NANDN U10182 ( .A(n9773), .B(n9772), .Z(n9774) );
  NAND U10183 ( .A(n9775), .B(n9774), .Z(n9859) );
  XNOR U10184 ( .A(n9858), .B(n9859), .Z(n9860) );
  NANDN U10185 ( .A(n9777), .B(n9776), .Z(n9781) );
  NAND U10186 ( .A(n9779), .B(n9778), .Z(n9780) );
  NAND U10187 ( .A(n9781), .B(n9780), .Z(n9949) );
  ANDN U10188 ( .B(y[746]), .A(n158), .Z(n10029) );
  ANDN U10189 ( .B(y[745]), .A(n159), .Z(n9925) );
  XNOR U10190 ( .A(n9924), .B(n9925), .Z(n9927) );
  ANDN U10191 ( .B(y[748]), .A(n156), .Z(n9926) );
  XOR U10192 ( .A(n9927), .B(n9926), .Z(n9913) );
  ANDN U10193 ( .B(y[749]), .A(n155), .Z(n9890) );
  ANDN U10194 ( .B(y[742]), .A(n162), .Z(n9888) );
  ANDN U10195 ( .B(y[740]), .A(n164), .Z(n9889) );
  XNOR U10196 ( .A(n9888), .B(n9889), .Z(n9891) );
  XNOR U10197 ( .A(n9890), .B(n9891), .Z(n9912) );
  XOR U10198 ( .A(n9913), .B(n9912), .Z(n9914) );
  XOR U10199 ( .A(n10029), .B(n9914), .Z(n9936) );
  AND U10200 ( .A(y[750]), .B(x[137]), .Z(n9782) );
  NAND U10201 ( .A(n9782), .B(n9917), .Z(n9786) );
  OR U10202 ( .A(n9784), .B(n9783), .Z(n9785) );
  NAND U10203 ( .A(n9786), .B(n9785), .Z(n9935) );
  NAND U10204 ( .A(x[139]), .B(y[738]), .Z(n9991) );
  AND U10205 ( .A(y[741]), .B(x[142]), .Z(n9787) );
  NANDN U10206 ( .A(n9991), .B(n9787), .Z(n9791) );
  OR U10207 ( .A(n9789), .B(n9788), .Z(n9790) );
  NAND U10208 ( .A(n9791), .B(n9790), .Z(n9934) );
  XNOR U10209 ( .A(n9935), .B(n9934), .Z(n9937) );
  XNOR U10210 ( .A(n9936), .B(n9937), .Z(n9947) );
  NAND U10211 ( .A(n9793), .B(n9792), .Z(n9797) );
  NAND U10212 ( .A(n9795), .B(n9794), .Z(n9796) );
  AND U10213 ( .A(n9797), .B(n9796), .Z(n9946) );
  XOR U10214 ( .A(n9947), .B(n9946), .Z(n9948) );
  XNOR U10215 ( .A(n9949), .B(n9948), .Z(n9953) );
  OR U10216 ( .A(n9799), .B(n9798), .Z(n9803) );
  NANDN U10217 ( .A(n9801), .B(n9800), .Z(n9802) );
  NAND U10218 ( .A(n9803), .B(n9802), .Z(n9952) );
  XOR U10219 ( .A(n9953), .B(n9952), .Z(n9954) );
  OR U10220 ( .A(n9805), .B(n9804), .Z(n9809) );
  NANDN U10221 ( .A(n9807), .B(n9806), .Z(n9808) );
  NAND U10222 ( .A(n9809), .B(n9808), .Z(n9955) );
  XNOR U10223 ( .A(n9954), .B(n9955), .Z(n9864) );
  OR U10224 ( .A(n9811), .B(n9810), .Z(n9815) );
  NANDN U10225 ( .A(n9813), .B(n9812), .Z(n9814) );
  NAND U10226 ( .A(n9815), .B(n9814), .Z(n9961) );
  OR U10227 ( .A(n9817), .B(n9816), .Z(n9821) );
  NANDN U10228 ( .A(n9819), .B(n9818), .Z(n9820) );
  NAND U10229 ( .A(n9821), .B(n9820), .Z(n9959) );
  OR U10230 ( .A(n9823), .B(n9822), .Z(n9827) );
  OR U10231 ( .A(n9825), .B(n9824), .Z(n9826) );
  NAND U10232 ( .A(n9827), .B(n9826), .Z(n9942) );
  NANDN U10233 ( .A(n9828), .B(n10029), .Z(n9832) );
  OR U10234 ( .A(n9830), .B(n9829), .Z(n9831) );
  AND U10235 ( .A(n9832), .B(n9831), .Z(n9882) );
  NAND U10236 ( .A(x[136]), .B(y[751]), .Z(n10518) );
  ANDN U10237 ( .B(y[744]), .A(n152), .Z(n10008) );
  NANDN U10238 ( .A(n10518), .B(n10008), .Z(n9836) );
  OR U10239 ( .A(n9834), .B(n9833), .Z(n9835) );
  AND U10240 ( .A(n9836), .B(n9835), .Z(n9883) );
  XOR U10241 ( .A(n9882), .B(n9883), .Z(n9884) );
  NAND U10242 ( .A(x[144]), .B(y[737]), .Z(n9896) );
  XOR U10243 ( .A(o[113]), .B(n9896), .Z(n9900) );
  AND U10244 ( .A(y[736]), .B(x[145]), .Z(n9899) );
  XOR U10245 ( .A(n9900), .B(n9899), .Z(n9902) );
  AND U10246 ( .A(x[128]), .B(y[753]), .Z(n9901) );
  XOR U10247 ( .A(n9902), .B(n9901), .Z(n9879) );
  AND U10248 ( .A(y[743]), .B(x[138]), .Z(n9838) );
  NAND U10249 ( .A(x[130]), .B(y[751]), .Z(n9837) );
  XOR U10250 ( .A(n9838), .B(n9837), .Z(n9919) );
  AND U10251 ( .A(y[750]), .B(x[131]), .Z(n9918) );
  XNOR U10252 ( .A(n9919), .B(n9918), .Z(n9876) );
  NANDN U10253 ( .A(n9840), .B(n9839), .Z(n9844) );
  NAND U10254 ( .A(n9842), .B(n9841), .Z(n9843) );
  AND U10255 ( .A(n9844), .B(n9843), .Z(n9877) );
  XOR U10256 ( .A(n9879), .B(n9878), .Z(n9885) );
  XNOR U10257 ( .A(n9884), .B(n9885), .Z(n9941) );
  ANDN U10258 ( .B(y[747]), .A(n164), .Z(n10746) );
  NAND U10259 ( .A(n9845), .B(n10746), .Z(n9848) );
  OR U10260 ( .A(n9846), .B(n10523), .Z(n9847) );
  AND U10261 ( .A(n9848), .B(n9847), .Z(n9873) );
  ANDN U10262 ( .B(y[741]), .A(n163), .Z(n9910) );
  NOR U10263 ( .A(n165), .B(n149), .Z(n9983) );
  ANDN U10264 ( .B(y[738]), .A(n166), .Z(n9909) );
  XNOR U10265 ( .A(n9983), .B(n9909), .Z(n9911) );
  XOR U10266 ( .A(n9910), .B(n9911), .Z(n9871) );
  NANDN U10267 ( .A(n9849), .B(o[112]), .Z(n9931) );
  AND U10268 ( .A(x[137]), .B(y[744]), .Z(n9851) );
  NAND U10269 ( .A(x[129]), .B(y[752]), .Z(n9850) );
  XOR U10270 ( .A(n9851), .B(n9850), .Z(n9930) );
  XNOR U10271 ( .A(n9931), .B(n9930), .Z(n9870) );
  XOR U10272 ( .A(n9871), .B(n9870), .Z(n9872) );
  XOR U10273 ( .A(n9873), .B(n9872), .Z(n9940) );
  XOR U10274 ( .A(n9941), .B(n9940), .Z(n9943) );
  XOR U10275 ( .A(n9942), .B(n9943), .Z(n9958) );
  XNOR U10276 ( .A(n9959), .B(n9958), .Z(n9960) );
  XOR U10277 ( .A(n9961), .B(n9960), .Z(n9865) );
  XNOR U10278 ( .A(n9864), .B(n9865), .Z(n9867) );
  OR U10279 ( .A(n9853), .B(n9852), .Z(n9857) );
  NANDN U10280 ( .A(n9855), .B(n9854), .Z(n9856) );
  AND U10281 ( .A(n9857), .B(n9856), .Z(n9866) );
  XOR U10282 ( .A(n9867), .B(n9866), .Z(n9861) );
  XNOR U10283 ( .A(n9860), .B(n9861), .Z(N242) );
  NANDN U10284 ( .A(n9859), .B(n9858), .Z(n9863) );
  NAND U10285 ( .A(n9861), .B(n9860), .Z(n9862) );
  NAND U10286 ( .A(n9863), .B(n9862), .Z(n9964) );
  OR U10287 ( .A(n9865), .B(n9864), .Z(n9869) );
  OR U10288 ( .A(n9867), .B(n9866), .Z(n9868) );
  AND U10289 ( .A(n9869), .B(n9868), .Z(n9965) );
  XNOR U10290 ( .A(n9964), .B(n9965), .Z(n9966) );
  OR U10291 ( .A(n9871), .B(n9870), .Z(n9875) );
  NANDN U10292 ( .A(n9873), .B(n9872), .Z(n9874) );
  AND U10293 ( .A(n9875), .B(n9874), .Z(n10044) );
  NANDN U10294 ( .A(n9877), .B(n9876), .Z(n9881) );
  NANDN U10295 ( .A(n9879), .B(n9878), .Z(n9880) );
  AND U10296 ( .A(n9881), .B(n9880), .Z(n10045) );
  XOR U10297 ( .A(n10044), .B(n10045), .Z(n10046) );
  OR U10298 ( .A(n9883), .B(n9882), .Z(n9887) );
  NANDN U10299 ( .A(n9885), .B(n9884), .Z(n9886) );
  AND U10300 ( .A(n9887), .B(n9886), .Z(n10047) );
  XNOR U10301 ( .A(n10046), .B(n10047), .Z(n10076) );
  OR U10302 ( .A(n9889), .B(n9888), .Z(n9893) );
  OR U10303 ( .A(n9891), .B(n9890), .Z(n9892) );
  NAND U10304 ( .A(n9893), .B(n9892), .Z(n9999) );
  AND U10305 ( .A(x[143]), .B(y[739]), .Z(n9895) );
  NAND U10306 ( .A(x[142]), .B(y[740]), .Z(n9894) );
  XNOR U10307 ( .A(n9895), .B(n9894), .Z(n9985) );
  XNOR U10308 ( .A(n9984), .B(n9985), .Z(n9997) );
  NANDN U10309 ( .A(n9896), .B(o[113]), .Z(n10010) );
  AND U10310 ( .A(x[138]), .B(y[744]), .Z(n9898) );
  NAND U10311 ( .A(x[129]), .B(y[753]), .Z(n9897) );
  XNOR U10312 ( .A(n9898), .B(n9897), .Z(n10009) );
  XOR U10313 ( .A(n9999), .B(n9998), .Z(n10063) );
  NANDN U10314 ( .A(n9900), .B(n9899), .Z(n9904) );
  NANDN U10315 ( .A(n9902), .B(n9901), .Z(n9903) );
  NAND U10316 ( .A(n9904), .B(n9903), .Z(n10051) );
  NAND U10317 ( .A(x[135]), .B(y[747]), .Z(n9905) );
  XOR U10318 ( .A(n9906), .B(n9905), .Z(n10032) );
  NAND U10319 ( .A(x[132]), .B(y[750]), .Z(n10031) );
  XNOR U10320 ( .A(n10032), .B(n10031), .Z(n9977) );
  AND U10321 ( .A(x[133]), .B(y[749]), .Z(n10151) );
  NAND U10322 ( .A(x[134]), .B(y[748]), .Z(n9976) );
  XNOR U10323 ( .A(n10151), .B(n9976), .Z(n9978) );
  XOR U10324 ( .A(n10051), .B(n10050), .Z(n10053) );
  NAND U10325 ( .A(x[130]), .B(y[752]), .Z(n9993) );
  AND U10326 ( .A(y[743]), .B(x[139]), .Z(n9908) );
  AND U10327 ( .A(y[738]), .B(x[144]), .Z(n9907) );
  XNOR U10328 ( .A(n9908), .B(n9907), .Z(n9992) );
  XOR U10329 ( .A(n9993), .B(n9992), .Z(n10052) );
  XNOR U10330 ( .A(n10053), .B(n10052), .Z(n10062) );
  XOR U10331 ( .A(n10063), .B(n10062), .Z(n10065) );
  XOR U10332 ( .A(n10065), .B(n10064), .Z(n10075) );
  NANDN U10333 ( .A(n9913), .B(n9912), .Z(n9916) );
  NANDN U10334 ( .A(n9914), .B(n10029), .Z(n9915) );
  NAND U10335 ( .A(n9916), .B(n9915), .Z(n10039) );
  IV U10336 ( .A(y[751]), .Z(n10692) );
  NOR U10337 ( .A(n161), .B(n10692), .Z(n10903) );
  NAND U10338 ( .A(n10903), .B(n9917), .Z(n9921) );
  NANDN U10339 ( .A(n9919), .B(n9918), .Z(n9920) );
  AND U10340 ( .A(n9921), .B(n9920), .Z(n10004) );
  NAND U10341 ( .A(x[128]), .B(y[754]), .Z(n10014) );
  NAND U10342 ( .A(x[146]), .B(y[736]), .Z(n10013) );
  XOR U10343 ( .A(n10014), .B(n10013), .Z(n10015) );
  NAND U10344 ( .A(x[145]), .B(y[737]), .Z(n10037) );
  XOR U10345 ( .A(o[114]), .B(n10037), .Z(n10016) );
  XOR U10346 ( .A(n10015), .B(n10016), .Z(n10003) );
  ANDN U10347 ( .B(y[742]), .A(n163), .Z(n10115) );
  AND U10348 ( .A(x[131]), .B(y[751]), .Z(n9923) );
  NAND U10349 ( .A(x[141]), .B(y[741]), .Z(n9922) );
  XOR U10350 ( .A(n9923), .B(n9922), .Z(n10022) );
  XOR U10351 ( .A(n10115), .B(n10022), .Z(n10002) );
  XNOR U10352 ( .A(n10003), .B(n10002), .Z(n10005) );
  XOR U10353 ( .A(n10004), .B(n10005), .Z(n10056) );
  OR U10354 ( .A(n9925), .B(n9924), .Z(n9929) );
  OR U10355 ( .A(n9927), .B(n9926), .Z(n9928) );
  AND U10356 ( .A(n9929), .B(n9928), .Z(n10057) );
  XNOR U10357 ( .A(n10056), .B(n10057), .Z(n10059) );
  AND U10358 ( .A(y[752]), .B(x[137]), .Z(n10904) );
  NAND U10359 ( .A(n10008), .B(n10904), .Z(n9933) );
  OR U10360 ( .A(n9931), .B(n9930), .Z(n9932) );
  NAND U10361 ( .A(n9933), .B(n9932), .Z(n10058) );
  XNOR U10362 ( .A(n10059), .B(n10058), .Z(n10038) );
  XNOR U10363 ( .A(n10039), .B(n10038), .Z(n10041) );
  OR U10364 ( .A(n9935), .B(n9934), .Z(n9939) );
  NANDN U10365 ( .A(n9937), .B(n9936), .Z(n9938) );
  AND U10366 ( .A(n9939), .B(n9938), .Z(n10040) );
  XOR U10367 ( .A(n10041), .B(n10040), .Z(n10074) );
  XOR U10368 ( .A(n10075), .B(n10074), .Z(n10077) );
  XNOR U10369 ( .A(n10076), .B(n10077), .Z(n10071) );
  NANDN U10370 ( .A(n9941), .B(n9940), .Z(n9945) );
  OR U10371 ( .A(n9943), .B(n9942), .Z(n9944) );
  NAND U10372 ( .A(n9945), .B(n9944), .Z(n10068) );
  OR U10373 ( .A(n9947), .B(n9946), .Z(n9951) );
  NAND U10374 ( .A(n9949), .B(n9948), .Z(n9950) );
  NAND U10375 ( .A(n9951), .B(n9950), .Z(n10069) );
  XOR U10376 ( .A(n10071), .B(n10070), .Z(n9973) );
  OR U10377 ( .A(n9953), .B(n9952), .Z(n9957) );
  NANDN U10378 ( .A(n9955), .B(n9954), .Z(n9956) );
  NAND U10379 ( .A(n9957), .B(n9956), .Z(n9971) );
  OR U10380 ( .A(n9959), .B(n9958), .Z(n9963) );
  OR U10381 ( .A(n9961), .B(n9960), .Z(n9962) );
  NAND U10382 ( .A(n9963), .B(n9962), .Z(n9970) );
  XNOR U10383 ( .A(n9971), .B(n9970), .Z(n9972) );
  XNOR U10384 ( .A(n9973), .B(n9972), .Z(n9967) );
  XOR U10385 ( .A(n9966), .B(n9967), .Z(N243) );
  NANDN U10386 ( .A(n9965), .B(n9964), .Z(n9969) );
  NANDN U10387 ( .A(n9967), .B(n9966), .Z(n9968) );
  NAND U10388 ( .A(n9969), .B(n9968), .Z(n10189) );
  OR U10389 ( .A(n9971), .B(n9970), .Z(n9975) );
  OR U10390 ( .A(n9973), .B(n9972), .Z(n9974) );
  AND U10391 ( .A(n9975), .B(n9974), .Z(n10190) );
  XNOR U10392 ( .A(n10189), .B(n10190), .Z(n10191) );
  NANDN U10393 ( .A(n10151), .B(n9976), .Z(n9980) );
  NAND U10394 ( .A(n9978), .B(n9977), .Z(n9979) );
  AND U10395 ( .A(n9980), .B(n9979), .Z(n10185) );
  AND U10396 ( .A(y[747]), .B(x[136]), .Z(n9982) );
  NAND U10397 ( .A(x[142]), .B(y[741]), .Z(n9981) );
  XOR U10398 ( .A(n9982), .B(n9981), .Z(n10163) );
  NAND U10399 ( .A(y[754]), .B(x[129]), .Z(n10162) );
  XOR U10400 ( .A(n10163), .B(n10162), .Z(n10100) );
  ANDN U10401 ( .B(y[740]), .A(n166), .Z(n10111) );
  NAND U10402 ( .A(n9983), .B(n10111), .Z(n9987) );
  NAND U10403 ( .A(n9985), .B(n9984), .Z(n9986) );
  NAND U10404 ( .A(n9987), .B(n9986), .Z(n10098) );
  NAND U10405 ( .A(x[141]), .B(y[742]), .Z(n9988) );
  XOR U10406 ( .A(n9989), .B(n9988), .Z(n10118) );
  NAND U10407 ( .A(y[753]), .B(x[130]), .Z(n10117) );
  XNOR U10408 ( .A(n10118), .B(n10117), .Z(n10099) );
  XOR U10409 ( .A(n10098), .B(n10099), .Z(n10101) );
  XNOR U10410 ( .A(n10100), .B(n10101), .Z(n10183) );
  AND U10411 ( .A(y[743]), .B(x[144]), .Z(n9990) );
  NANDN U10412 ( .A(n9991), .B(n9990), .Z(n9995) );
  OR U10413 ( .A(n9993), .B(n9992), .Z(n9994) );
  NAND U10414 ( .A(n9995), .B(n9994), .Z(n10184) );
  XNOR U10415 ( .A(n10183), .B(n10184), .Z(n10186) );
  XOR U10416 ( .A(n10185), .B(n10186), .Z(n10092) );
  NANDN U10417 ( .A(n9997), .B(n9996), .Z(n10001) );
  NANDN U10418 ( .A(n9999), .B(n9998), .Z(n10000) );
  NAND U10419 ( .A(n10001), .B(n10000), .Z(n10178) );
  OR U10420 ( .A(n10003), .B(n10002), .Z(n10007) );
  OR U10421 ( .A(n10005), .B(n10004), .Z(n10006) );
  NAND U10422 ( .A(n10007), .B(n10006), .Z(n10177) );
  XOR U10423 ( .A(n10178), .B(n10177), .Z(n10179) );
  AND U10424 ( .A(x[138]), .B(y[753]), .Z(n11285) );
  NAND U10425 ( .A(n10008), .B(n11285), .Z(n10012) );
  NANDN U10426 ( .A(n10010), .B(n10009), .Z(n10011) );
  NAND U10427 ( .A(n10012), .B(n10011), .Z(n10142) );
  OR U10428 ( .A(n10014), .B(n10013), .Z(n10018) );
  NANDN U10429 ( .A(n10016), .B(n10015), .Z(n10017) );
  NAND U10430 ( .A(n10018), .B(n10017), .Z(n10139) );
  AND U10431 ( .A(x[137]), .B(y[746]), .Z(n10020) );
  NAND U10432 ( .A(x[144]), .B(y[739]), .Z(n10019) );
  XNOR U10433 ( .A(n10020), .B(n10019), .Z(n10112) );
  XNOR U10434 ( .A(n10111), .B(n10112), .Z(n10140) );
  XOR U10435 ( .A(n10142), .B(n10141), .Z(n10173) );
  NOR U10436 ( .A(n164), .B(n10692), .Z(n11450) );
  NAND U10437 ( .A(n11450), .B(n10021), .Z(n10024) );
  NANDN U10438 ( .A(n10022), .B(n10115), .Z(n10023) );
  NAND U10439 ( .A(n10024), .B(n10023), .Z(n10136) );
  AND U10440 ( .A(x[139]), .B(y[744]), .Z(n10026) );
  NAND U10441 ( .A(x[135]), .B(y[748]), .Z(n10025) );
  XOR U10442 ( .A(n10026), .B(n10025), .Z(n10127) );
  NAND U10443 ( .A(x[131]), .B(y[752]), .Z(n10126) );
  XOR U10444 ( .A(n10127), .B(n10126), .Z(n10134) );
  NAND U10445 ( .A(x[146]), .B(y[737]), .Z(n10132) );
  XOR U10446 ( .A(o[115]), .B(n10132), .Z(n10168) );
  AND U10447 ( .A(y[745]), .B(x[138]), .Z(n10028) );
  NAND U10448 ( .A(x[145]), .B(y[738]), .Z(n10027) );
  XNOR U10449 ( .A(n10028), .B(n10027), .Z(n10167) );
  XOR U10450 ( .A(n10136), .B(n10135), .Z(n10171) );
  NANDN U10451 ( .A(n10030), .B(n10029), .Z(n10034) );
  OR U10452 ( .A(n10032), .B(n10031), .Z(n10033) );
  NAND U10453 ( .A(n10034), .B(n10033), .Z(n10105) );
  NAND U10454 ( .A(x[132]), .B(y[751]), .Z(n10249) );
  AND U10455 ( .A(x[134]), .B(y[749]), .Z(n10036) );
  NAND U10456 ( .A(x[133]), .B(y[750]), .Z(n10035) );
  XNOR U10457 ( .A(n10036), .B(n10035), .Z(n10152) );
  XNOR U10458 ( .A(n10105), .B(n10104), .Z(n10106) );
  NANDN U10459 ( .A(n10037), .B(o[114]), .Z(n10148) );
  NAND U10460 ( .A(x[128]), .B(y[755]), .Z(n10146) );
  NAND U10461 ( .A(x[147]), .B(y[736]), .Z(n10145) );
  XOR U10462 ( .A(n10146), .B(n10145), .Z(n10147) );
  XOR U10463 ( .A(n10148), .B(n10147), .Z(n10107) );
  XOR U10464 ( .A(n10106), .B(n10107), .Z(n10172) );
  XNOR U10465 ( .A(n10171), .B(n10172), .Z(n10174) );
  XNOR U10466 ( .A(n10173), .B(n10174), .Z(n10180) );
  XNOR U10467 ( .A(n10179), .B(n10180), .Z(n10093) );
  XNOR U10468 ( .A(n10092), .B(n10093), .Z(n10095) );
  OR U10469 ( .A(n10039), .B(n10038), .Z(n10043) );
  OR U10470 ( .A(n10041), .B(n10040), .Z(n10042) );
  NAND U10471 ( .A(n10043), .B(n10042), .Z(n10094) );
  XOR U10472 ( .A(n10095), .B(n10094), .Z(n10089) );
  OR U10473 ( .A(n10045), .B(n10044), .Z(n10049) );
  NANDN U10474 ( .A(n10047), .B(n10046), .Z(n10048) );
  NAND U10475 ( .A(n10049), .B(n10048), .Z(n10087) );
  NANDN U10476 ( .A(n10051), .B(n10050), .Z(n10055) );
  OR U10477 ( .A(n10053), .B(n10052), .Z(n10054) );
  AND U10478 ( .A(n10055), .B(n10054), .Z(n10083) );
  OR U10479 ( .A(n10057), .B(n10056), .Z(n10061) );
  OR U10480 ( .A(n10059), .B(n10058), .Z(n10060) );
  AND U10481 ( .A(n10061), .B(n10060), .Z(n10080) );
  NANDN U10482 ( .A(n10063), .B(n10062), .Z(n10067) );
  OR U10483 ( .A(n10065), .B(n10064), .Z(n10066) );
  NAND U10484 ( .A(n10067), .B(n10066), .Z(n10081) );
  XOR U10485 ( .A(n10080), .B(n10081), .Z(n10082) );
  XOR U10486 ( .A(n10087), .B(n10086), .Z(n10088) );
  XNOR U10487 ( .A(n10089), .B(n10088), .Z(n10198) );
  NANDN U10488 ( .A(n10069), .B(n10068), .Z(n10073) );
  NANDN U10489 ( .A(n10071), .B(n10070), .Z(n10072) );
  NAND U10490 ( .A(n10073), .B(n10072), .Z(n10196) );
  NANDN U10491 ( .A(n10075), .B(n10074), .Z(n10079) );
  OR U10492 ( .A(n10077), .B(n10076), .Z(n10078) );
  AND U10493 ( .A(n10079), .B(n10078), .Z(n10195) );
  XNOR U10494 ( .A(n10198), .B(n10197), .Z(n10192) );
  XOR U10495 ( .A(n10191), .B(n10192), .Z(N244) );
  OR U10496 ( .A(n10081), .B(n10080), .Z(n10085) );
  NANDN U10497 ( .A(n10083), .B(n10082), .Z(n10084) );
  AND U10498 ( .A(n10085), .B(n10084), .Z(n10315) );
  OR U10499 ( .A(n10087), .B(n10086), .Z(n10091) );
  NANDN U10500 ( .A(n10089), .B(n10088), .Z(n10090) );
  AND U10501 ( .A(n10091), .B(n10090), .Z(n10314) );
  OR U10502 ( .A(n10093), .B(n10092), .Z(n10097) );
  OR U10503 ( .A(n10095), .B(n10094), .Z(n10096) );
  AND U10504 ( .A(n10097), .B(n10096), .Z(n10298) );
  NANDN U10505 ( .A(n10099), .B(n10098), .Z(n10103) );
  NANDN U10506 ( .A(n10101), .B(n10100), .Z(n10102) );
  NAND U10507 ( .A(n10103), .B(n10102), .Z(n10201) );
  NAND U10508 ( .A(n10105), .B(n10104), .Z(n10109) );
  OR U10509 ( .A(n10107), .B(n10106), .Z(n10108) );
  AND U10510 ( .A(n10109), .B(n10108), .Z(n10202) );
  AND U10511 ( .A(x[144]), .B(y[746]), .Z(n11040) );
  NANDN U10512 ( .A(n10110), .B(n11040), .Z(n10114) );
  NAND U10513 ( .A(n10112), .B(n10111), .Z(n10113) );
  NAND U10514 ( .A(n10114), .B(n10113), .Z(n10241) );
  AND U10515 ( .A(y[743]), .B(x[141]), .Z(n10116) );
  NAND U10516 ( .A(n10116), .B(n10115), .Z(n10120) );
  OR U10517 ( .A(n10118), .B(n10117), .Z(n10119) );
  NAND U10518 ( .A(n10120), .B(n10119), .Z(n10280) );
  AND U10519 ( .A(x[138]), .B(y[746]), .Z(n10122) );
  NAND U10520 ( .A(x[144]), .B(y[740]), .Z(n10121) );
  XOR U10521 ( .A(n10122), .B(n10121), .Z(n10268) );
  NAND U10522 ( .A(y[754]), .B(x[130]), .Z(n10267) );
  XOR U10523 ( .A(n10268), .B(n10267), .Z(n10278) );
  AND U10524 ( .A(y[741]), .B(x[143]), .Z(n10124) );
  NAND U10525 ( .A(x[137]), .B(y[747]), .Z(n10123) );
  XOR U10526 ( .A(n10124), .B(n10123), .Z(n10226) );
  AND U10527 ( .A(x[142]), .B(y[742]), .Z(n10225) );
  XNOR U10528 ( .A(n10226), .B(n10225), .Z(n10277) );
  XNOR U10529 ( .A(n10280), .B(n10279), .Z(n10242) );
  ANDN U10530 ( .B(y[748]), .A(n162), .Z(n10713) );
  NANDN U10531 ( .A(n10125), .B(n10713), .Z(n10129) );
  OR U10532 ( .A(n10127), .B(n10126), .Z(n10128) );
  AND U10533 ( .A(n10129), .B(n10128), .Z(n10285) );
  AND U10534 ( .A(y[745]), .B(x[139]), .Z(n10131) );
  NAND U10535 ( .A(x[129]), .B(y[755]), .Z(n10130) );
  XOR U10536 ( .A(n10131), .B(n10130), .Z(n10232) );
  NAND U10537 ( .A(x[147]), .B(y[737]), .Z(n10229) );
  XNOR U10538 ( .A(n10229), .B(o[116]), .Z(n10231) );
  XOR U10539 ( .A(n10232), .B(n10231), .Z(n10284) );
  NANDN U10540 ( .A(n10132), .B(o[115]), .Z(n10257) );
  NAND U10541 ( .A(x[128]), .B(y[756]), .Z(n10255) );
  NAND U10542 ( .A(x[148]), .B(y[736]), .Z(n10254) );
  XOR U10543 ( .A(n10255), .B(n10254), .Z(n10256) );
  XNOR U10544 ( .A(n10257), .B(n10256), .Z(n10283) );
  XOR U10545 ( .A(n10284), .B(n10283), .Z(n10286) );
  XOR U10546 ( .A(n10285), .B(n10286), .Z(n10243) );
  NAND U10547 ( .A(n10134), .B(n10133), .Z(n10138) );
  NAND U10548 ( .A(n10136), .B(n10135), .Z(n10137) );
  NAND U10549 ( .A(n10138), .B(n10137), .Z(n10290) );
  NANDN U10550 ( .A(n10140), .B(n10139), .Z(n10144) );
  NAND U10551 ( .A(n10142), .B(n10141), .Z(n10143) );
  NAND U10552 ( .A(n10144), .B(n10143), .Z(n10238) );
  OR U10553 ( .A(n10146), .B(n10145), .Z(n10150) );
  NANDN U10554 ( .A(n10148), .B(n10147), .Z(n10149) );
  NAND U10555 ( .A(n10150), .B(n10149), .Z(n10209) );
  ANDN U10556 ( .B(y[750]), .A(n157), .Z(n10213) );
  NAND U10557 ( .A(n10213), .B(n10151), .Z(n10154) );
  NANDN U10558 ( .A(n10249), .B(n10152), .Z(n10153) );
  NAND U10559 ( .A(n10154), .B(n10153), .Z(n10207) );
  AND U10560 ( .A(x[140]), .B(y[744]), .Z(n10156) );
  NAND U10561 ( .A(x[146]), .B(y[738]), .Z(n10155) );
  XOR U10562 ( .A(n10156), .B(n10155), .Z(n10221) );
  NAND U10563 ( .A(y[739]), .B(x[145]), .Z(n10220) );
  XNOR U10564 ( .A(n10221), .B(n10220), .Z(n10208) );
  XOR U10565 ( .A(n10207), .B(n10208), .Z(n10210) );
  AND U10566 ( .A(x[131]), .B(y[753]), .Z(n10158) );
  NAND U10567 ( .A(x[141]), .B(y[743]), .Z(n10157) );
  XOR U10568 ( .A(n10158), .B(n10157), .Z(n10263) );
  NAND U10569 ( .A(x[136]), .B(y[748]), .Z(n10262) );
  XOR U10570 ( .A(n10263), .B(n10262), .Z(n10215) );
  AND U10571 ( .A(x[133]), .B(y[751]), .Z(n10160) );
  NAND U10572 ( .A(x[132]), .B(y[752]), .Z(n10159) );
  XOR U10573 ( .A(n10160), .B(n10159), .Z(n10251) );
  NAND U10574 ( .A(x[135]), .B(y[749]), .Z(n10250) );
  XNOR U10575 ( .A(n10251), .B(n10250), .Z(n10214) );
  XNOR U10576 ( .A(n10215), .B(n10216), .Z(n10274) );
  ANDN U10577 ( .B(y[747]), .A(n165), .Z(n10957) );
  NAND U10578 ( .A(n10957), .B(n10161), .Z(n10165) );
  OR U10579 ( .A(n10163), .B(n10162), .Z(n10164) );
  NAND U10580 ( .A(n10165), .B(n10164), .Z(n10272) );
  AND U10581 ( .A(y[745]), .B(x[145]), .Z(n11054) );
  NANDN U10582 ( .A(n10166), .B(n11054), .Z(n10170) );
  NANDN U10583 ( .A(n10168), .B(n10167), .Z(n10169) );
  AND U10584 ( .A(n10170), .B(n10169), .Z(n10271) );
  XOR U10585 ( .A(n10274), .B(n10273), .Z(n10236) );
  XNOR U10586 ( .A(n10235), .B(n10236), .Z(n10237) );
  XNOR U10587 ( .A(n10238), .B(n10237), .Z(n10289) );
  XOR U10588 ( .A(n10290), .B(n10289), .Z(n10291) );
  XNOR U10589 ( .A(n10292), .B(n10291), .Z(n10296) );
  OR U10590 ( .A(n10172), .B(n10171), .Z(n10176) );
  OR U10591 ( .A(n10174), .B(n10173), .Z(n10175) );
  NAND U10592 ( .A(n10176), .B(n10175), .Z(n10302) );
  OR U10593 ( .A(n10178), .B(n10177), .Z(n10182) );
  NANDN U10594 ( .A(n10180), .B(n10179), .Z(n10181) );
  NAND U10595 ( .A(n10182), .B(n10181), .Z(n10301) );
  XOR U10596 ( .A(n10302), .B(n10301), .Z(n10303) );
  OR U10597 ( .A(n10184), .B(n10183), .Z(n10188) );
  OR U10598 ( .A(n10186), .B(n10185), .Z(n10187) );
  NAND U10599 ( .A(n10188), .B(n10187), .Z(n10304) );
  XOR U10600 ( .A(n10296), .B(n10295), .Z(n10297) );
  XOR U10601 ( .A(n10298), .B(n10297), .Z(n10313) );
  XOR U10602 ( .A(n10315), .B(n10316), .Z(n10309) );
  NANDN U10603 ( .A(n10190), .B(n10189), .Z(n10194) );
  NANDN U10604 ( .A(n10192), .B(n10191), .Z(n10193) );
  NAND U10605 ( .A(n10194), .B(n10193), .Z(n10307) );
  NANDN U10606 ( .A(n10196), .B(n10195), .Z(n10200) );
  NANDN U10607 ( .A(n10198), .B(n10197), .Z(n10199) );
  NAND U10608 ( .A(n10200), .B(n10199), .Z(n10308) );
  XNOR U10609 ( .A(n10307), .B(n10308), .Z(n10310) );
  XNOR U10610 ( .A(n10309), .B(n10310), .Z(N245) );
  NANDN U10611 ( .A(n10202), .B(n10201), .Z(n10206) );
  NAND U10612 ( .A(n10204), .B(n10203), .Z(n10205) );
  NAND U10613 ( .A(n10206), .B(n10205), .Z(n10339) );
  NANDN U10614 ( .A(n10208), .B(n10207), .Z(n10212) );
  NANDN U10615 ( .A(n10210), .B(n10209), .Z(n10211) );
  NAND U10616 ( .A(n10212), .B(n10211), .Z(n10426) );
  NANDN U10617 ( .A(n10214), .B(n10213), .Z(n10218) );
  NANDN U10618 ( .A(n10216), .B(n10215), .Z(n10217) );
  NAND U10619 ( .A(n10218), .B(n10217), .Z(n10425) );
  NOR U10620 ( .A(n169), .B(n11414), .Z(n11051) );
  NAND U10621 ( .A(n11051), .B(n10219), .Z(n10223) );
  OR U10622 ( .A(n10221), .B(n10220), .Z(n10222) );
  AND U10623 ( .A(n10223), .B(n10222), .Z(n10432) );
  AND U10624 ( .A(y[752]), .B(x[133]), .Z(n10412) );
  NAND U10625 ( .A(x[144]), .B(y[741]), .Z(n10413) );
  XOR U10626 ( .A(n10412), .B(n10413), .Z(n10415) );
  NAND U10627 ( .A(x[143]), .B(y[742]), .Z(n10414) );
  XNOR U10628 ( .A(n10415), .B(n10414), .Z(n10381) );
  ANDN U10629 ( .B(y[747]), .A(n166), .Z(n11045) );
  NAND U10630 ( .A(n10224), .B(n11045), .Z(n10228) );
  NANDN U10631 ( .A(n10226), .B(n10225), .Z(n10227) );
  NAND U10632 ( .A(n10228), .B(n10227), .Z(n10382) );
  ANDN U10633 ( .B(y[757]), .A(n151), .Z(n10402) );
  ANDN U10634 ( .B(o[116]), .A(n10229), .Z(n10400) );
  ANDN U10635 ( .B(y[736]), .A(n172), .Z(n10401) );
  XNOR U10636 ( .A(n10400), .B(n10401), .Z(n10403) );
  XOR U10637 ( .A(n10402), .B(n10403), .Z(n10384) );
  XOR U10638 ( .A(n10383), .B(n10384), .Z(n10430) );
  NAND U10639 ( .A(x[139]), .B(y[755]), .Z(n11883) );
  NANDN U10640 ( .A(n11883), .B(n10230), .Z(n10234) );
  NANDN U10641 ( .A(n10232), .B(n10231), .Z(n10233) );
  AND U10642 ( .A(n10234), .B(n10233), .Z(n10431) );
  XNOR U10643 ( .A(n10430), .B(n10431), .Z(n10433) );
  XOR U10644 ( .A(n10432), .B(n10433), .Z(n10424) );
  XNOR U10645 ( .A(n10425), .B(n10424), .Z(n10427) );
  NANDN U10646 ( .A(n10236), .B(n10235), .Z(n10240) );
  NANDN U10647 ( .A(n10238), .B(n10237), .Z(n10239) );
  AND U10648 ( .A(n10240), .B(n10239), .Z(n10338) );
  XNOR U10649 ( .A(n10337), .B(n10338), .Z(n10340) );
  NANDN U10650 ( .A(n10242), .B(n10241), .Z(n10246) );
  NAND U10651 ( .A(n10244), .B(n10243), .Z(n10245) );
  NAND U10652 ( .A(n10246), .B(n10245), .Z(n10346) );
  ANDN U10653 ( .B(y[751]), .A(n157), .Z(n10394) );
  ANDN U10654 ( .B(y[750]), .A(n158), .Z(n10517) );
  ANDN U10655 ( .B(y[743]), .A(n165), .Z(n10393) );
  XNOR U10656 ( .A(n10517), .B(n10393), .Z(n10395) );
  XNOR U10657 ( .A(n10394), .B(n10395), .Z(n10364) );
  NAND U10658 ( .A(y[749]), .B(x[136]), .Z(n10361) );
  XNOR U10659 ( .A(n10362), .B(n10361), .Z(n10363) );
  XNOR U10660 ( .A(n10364), .B(n10363), .Z(n10389) );
  NAND U10661 ( .A(x[132]), .B(y[753]), .Z(n10421) );
  AND U10662 ( .A(x[131]), .B(y[754]), .Z(n10248) );
  AND U10663 ( .A(x[141]), .B(y[744]), .Z(n10247) );
  XNOR U10664 ( .A(n10248), .B(n10247), .Z(n10420) );
  XOR U10665 ( .A(n10421), .B(n10420), .Z(n10387) );
  ANDN U10666 ( .B(y[745]), .A(n163), .Z(n10369) );
  ANDN U10667 ( .B(y[755]), .A(n153), .Z(n10367) );
  ANDN U10668 ( .B(y[740]), .A(n168), .Z(n10368) );
  XNOR U10669 ( .A(n10367), .B(n10368), .Z(n10370) );
  XOR U10670 ( .A(n10369), .B(n10370), .Z(n10388) );
  XOR U10671 ( .A(n10387), .B(n10388), .Z(n10390) );
  XNOR U10672 ( .A(n10389), .B(n10390), .Z(n10439) );
  NANDN U10673 ( .A(n10249), .B(n10412), .Z(n10253) );
  OR U10674 ( .A(n10251), .B(n10250), .Z(n10252) );
  AND U10675 ( .A(n10253), .B(n10252), .Z(n10437) );
  OR U10676 ( .A(n10255), .B(n10254), .Z(n10259) );
  NANDN U10677 ( .A(n10257), .B(n10256), .Z(n10258) );
  AND U10678 ( .A(n10259), .B(n10258), .Z(n10436) );
  XNOR U10679 ( .A(n10437), .B(n10436), .Z(n10438) );
  XOR U10680 ( .A(n10439), .B(n10438), .Z(n10358) );
  AND U10681 ( .A(y[753]), .B(x[141]), .Z(n10261) );
  NAND U10682 ( .A(n10261), .B(n10260), .Z(n10265) );
  OR U10683 ( .A(n10263), .B(n10262), .Z(n10264) );
  AND U10684 ( .A(n10265), .B(n10264), .Z(n10444) );
  ANDN U10685 ( .B(y[756]), .A(n152), .Z(n10406) );
  ANDN U10686 ( .B(y[739]), .A(n169), .Z(n10407) );
  XNOR U10687 ( .A(n10406), .B(n10407), .Z(n10409) );
  XNOR U10688 ( .A(n10408), .B(n10409), .Z(n10442) );
  NAND U10689 ( .A(x[139]), .B(y[746]), .Z(n10378) );
  NAND U10690 ( .A(x[148]), .B(y[737]), .Z(n10418) );
  XOR U10691 ( .A(o[117]), .B(n10418), .Z(n10376) );
  NAND U10692 ( .A(x[147]), .B(y[738]), .Z(n10375) );
  XNOR U10693 ( .A(n10376), .B(n10375), .Z(n10377) );
  XNOR U10694 ( .A(n10378), .B(n10377), .Z(n10443) );
  XOR U10695 ( .A(n10442), .B(n10443), .Z(n10445) );
  XOR U10696 ( .A(n10444), .B(n10445), .Z(n10356) );
  NAND U10697 ( .A(n10266), .B(n11040), .Z(n10270) );
  OR U10698 ( .A(n10268), .B(n10267), .Z(n10269) );
  NAND U10699 ( .A(n10270), .B(n10269), .Z(n10355) );
  XNOR U10700 ( .A(n10356), .B(n10355), .Z(n10357) );
  XOR U10701 ( .A(n10358), .B(n10357), .Z(n10344) );
  NANDN U10702 ( .A(n10272), .B(n10271), .Z(n10276) );
  NANDN U10703 ( .A(n10274), .B(n10273), .Z(n10275) );
  AND U10704 ( .A(n10276), .B(n10275), .Z(n10349) );
  NAND U10705 ( .A(n10278), .B(n10277), .Z(n10282) );
  NAND U10706 ( .A(n10280), .B(n10279), .Z(n10281) );
  NAND U10707 ( .A(n10282), .B(n10281), .Z(n10350) );
  XOR U10708 ( .A(n10349), .B(n10350), .Z(n10351) );
  NANDN U10709 ( .A(n10284), .B(n10283), .Z(n10288) );
  OR U10710 ( .A(n10286), .B(n10285), .Z(n10287) );
  NAND U10711 ( .A(n10288), .B(n10287), .Z(n10352) );
  XNOR U10712 ( .A(n10351), .B(n10352), .Z(n10343) );
  XOR U10713 ( .A(n10344), .B(n10343), .Z(n10345) );
  XNOR U10714 ( .A(n10346), .B(n10345), .Z(n10332) );
  NANDN U10715 ( .A(n10290), .B(n10289), .Z(n10294) );
  OR U10716 ( .A(n10292), .B(n10291), .Z(n10293) );
  AND U10717 ( .A(n10294), .B(n10293), .Z(n10331) );
  XOR U10718 ( .A(n10333), .B(n10334), .Z(n10328) );
  NAND U10719 ( .A(n10296), .B(n10295), .Z(n10300) );
  NANDN U10720 ( .A(n10298), .B(n10297), .Z(n10299) );
  NAND U10721 ( .A(n10300), .B(n10299), .Z(n10326) );
  OR U10722 ( .A(n10302), .B(n10301), .Z(n10306) );
  NANDN U10723 ( .A(n10304), .B(n10303), .Z(n10305) );
  NAND U10724 ( .A(n10306), .B(n10305), .Z(n10325) );
  XOR U10725 ( .A(n10326), .B(n10325), .Z(n10327) );
  XOR U10726 ( .A(n10328), .B(n10327), .Z(n10322) );
  NANDN U10727 ( .A(n10308), .B(n10307), .Z(n10312) );
  NAND U10728 ( .A(n10310), .B(n10309), .Z(n10311) );
  NAND U10729 ( .A(n10312), .B(n10311), .Z(n10319) );
  NANDN U10730 ( .A(n10314), .B(n10313), .Z(n10318) );
  OR U10731 ( .A(n10316), .B(n10315), .Z(n10317) );
  AND U10732 ( .A(n10318), .B(n10317), .Z(n10320) );
  XNOR U10733 ( .A(n10319), .B(n10320), .Z(n10321) );
  XOR U10734 ( .A(n10322), .B(n10321), .Z(N246) );
  NANDN U10735 ( .A(n10320), .B(n10319), .Z(n10324) );
  NANDN U10736 ( .A(n10322), .B(n10321), .Z(n10323) );
  NAND U10737 ( .A(n10324), .B(n10323), .Z(n10448) );
  OR U10738 ( .A(n10326), .B(n10325), .Z(n10330) );
  NANDN U10739 ( .A(n10328), .B(n10327), .Z(n10329) );
  AND U10740 ( .A(n10330), .B(n10329), .Z(n10449) );
  XNOR U10741 ( .A(n10448), .B(n10449), .Z(n10450) );
  NANDN U10742 ( .A(n10332), .B(n10331), .Z(n10336) );
  NAND U10743 ( .A(n10334), .B(n10333), .Z(n10335) );
  NAND U10744 ( .A(n10336), .B(n10335), .Z(n10457) );
  NAND U10745 ( .A(n10338), .B(n10337), .Z(n10342) );
  NANDN U10746 ( .A(n10340), .B(n10339), .Z(n10341) );
  NAND U10747 ( .A(n10342), .B(n10341), .Z(n10454) );
  OR U10748 ( .A(n10344), .B(n10343), .Z(n10348) );
  NAND U10749 ( .A(n10346), .B(n10345), .Z(n10347) );
  AND U10750 ( .A(n10348), .B(n10347), .Z(n10578) );
  OR U10751 ( .A(n10350), .B(n10349), .Z(n10354) );
  NANDN U10752 ( .A(n10352), .B(n10351), .Z(n10353) );
  NAND U10753 ( .A(n10354), .B(n10353), .Z(n10579) );
  XOR U10754 ( .A(n10578), .B(n10579), .Z(n10581) );
  OR U10755 ( .A(n10356), .B(n10355), .Z(n10360) );
  OR U10756 ( .A(n10358), .B(n10357), .Z(n10359) );
  NAND U10757 ( .A(n10360), .B(n10359), .Z(n10469) );
  NANDN U10758 ( .A(n10362), .B(n10361), .Z(n10366) );
  NANDN U10759 ( .A(n10364), .B(n10363), .Z(n10365) );
  AND U10760 ( .A(n10366), .B(n10365), .Z(n10486) );
  OR U10761 ( .A(n10368), .B(n10367), .Z(n10372) );
  OR U10762 ( .A(n10370), .B(n10369), .Z(n10371) );
  NAND U10763 ( .A(n10372), .B(n10371), .Z(n10555) );
  AND U10764 ( .A(x[140]), .B(y[746]), .Z(n10374) );
  NAND U10765 ( .A(x[146]), .B(y[740]), .Z(n10373) );
  XOR U10766 ( .A(n10374), .B(n10373), .Z(n10525) );
  NAND U10767 ( .A(y[754]), .B(x[132]), .Z(n10524) );
  XOR U10768 ( .A(n10525), .B(n10524), .Z(n10552) );
  NAND U10769 ( .A(x[133]), .B(y[753]), .Z(n10491) );
  NAND U10770 ( .A(x[145]), .B(y[741]), .Z(n10490) );
  XOR U10771 ( .A(n10491), .B(n10490), .Z(n10492) );
  NAND U10772 ( .A(y[742]), .B(x[144]), .Z(n10493) );
  XOR U10773 ( .A(n10492), .B(n10493), .Z(n10553) );
  XOR U10774 ( .A(n10555), .B(n10554), .Z(n10484) );
  OR U10775 ( .A(n10376), .B(n10375), .Z(n10380) );
  OR U10776 ( .A(n10378), .B(n10377), .Z(n10379) );
  NAND U10777 ( .A(n10380), .B(n10379), .Z(n10485) );
  XNOR U10778 ( .A(n10484), .B(n10485), .Z(n10487) );
  XNOR U10779 ( .A(n10486), .B(n10487), .Z(n10466) );
  NANDN U10780 ( .A(n10382), .B(n10381), .Z(n10386) );
  NAND U10781 ( .A(n10384), .B(n10383), .Z(n10385) );
  NAND U10782 ( .A(n10386), .B(n10385), .Z(n10475) );
  NANDN U10783 ( .A(n10388), .B(n10387), .Z(n10392) );
  OR U10784 ( .A(n10390), .B(n10389), .Z(n10391) );
  AND U10785 ( .A(n10392), .B(n10391), .Z(n10472) );
  OR U10786 ( .A(n10393), .B(n10517), .Z(n10397) );
  OR U10787 ( .A(n10395), .B(n10394), .Z(n10396) );
  NAND U10788 ( .A(n10397), .B(n10396), .Z(n10543) );
  AND U10789 ( .A(y[750]), .B(x[136]), .Z(n10399) );
  NAND U10790 ( .A(x[135]), .B(y[751]), .Z(n10398) );
  XNOR U10791 ( .A(n10399), .B(n10398), .Z(n10520) );
  XNOR U10792 ( .A(n10519), .B(n10520), .Z(n10541) );
  NAND U10793 ( .A(x[128]), .B(y[758]), .Z(n10529) );
  NAND U10794 ( .A(x[150]), .B(y[736]), .Z(n10528) );
  XOR U10795 ( .A(n10529), .B(n10528), .Z(n10530) );
  NAND U10796 ( .A(x[149]), .B(y[737]), .Z(n10496) );
  XOR U10797 ( .A(o[118]), .B(n10496), .Z(n10531) );
  XOR U10798 ( .A(n10530), .B(n10531), .Z(n10540) );
  XOR U10799 ( .A(n10541), .B(n10540), .Z(n10542) );
  XNOR U10800 ( .A(n10543), .B(n10542), .Z(n10549) );
  OR U10801 ( .A(n10401), .B(n10400), .Z(n10405) );
  OR U10802 ( .A(n10403), .B(n10402), .Z(n10404) );
  AND U10803 ( .A(n10405), .B(n10404), .Z(n10546) );
  OR U10804 ( .A(n10407), .B(n10406), .Z(n10411) );
  OR U10805 ( .A(n10409), .B(n10408), .Z(n10410) );
  AND U10806 ( .A(n10411), .B(n10410), .Z(n10547) );
  XOR U10807 ( .A(n10546), .B(n10547), .Z(n10548) );
  XOR U10808 ( .A(n10549), .B(n10548), .Z(n10481) );
  NAND U10809 ( .A(x[130]), .B(y[756]), .Z(n10504) );
  NAND U10810 ( .A(x[148]), .B(y[738]), .Z(n10503) );
  XOR U10811 ( .A(n10504), .B(n10503), .Z(n10505) );
  NAND U10812 ( .A(x[141]), .B(y[745]), .Z(n10506) );
  XOR U10813 ( .A(n10505), .B(n10506), .Z(n10511) );
  NANDN U10814 ( .A(n10413), .B(n10412), .Z(n10417) );
  OR U10815 ( .A(n10415), .B(n10414), .Z(n10416) );
  NAND U10816 ( .A(n10417), .B(n10416), .Z(n10509) );
  NAND U10817 ( .A(x[134]), .B(y[752]), .Z(n10498) );
  NAND U10818 ( .A(x[138]), .B(y[748]), .Z(n10497) );
  XOR U10819 ( .A(n10498), .B(n10497), .Z(n10499) );
  NAND U10820 ( .A(x[143]), .B(y[743]), .Z(n10500) );
  XOR U10821 ( .A(n10499), .B(n10500), .Z(n10510) );
  XOR U10822 ( .A(n10511), .B(n10512), .Z(n10478) );
  NANDN U10823 ( .A(n10418), .B(o[117]), .Z(n10563) );
  NAND U10824 ( .A(x[129]), .B(y[757]), .Z(n10561) );
  XOR U10825 ( .A(n10560), .B(n10561), .Z(n10562) );
  XOR U10826 ( .A(n10563), .B(n10562), .Z(n10536) );
  ANDN U10827 ( .B(y[754]), .A(n164), .Z(n11886) );
  NAND U10828 ( .A(n10419), .B(n11886), .Z(n10423) );
  OR U10829 ( .A(n10421), .B(n10420), .Z(n10422) );
  AND U10830 ( .A(n10423), .B(n10422), .Z(n10534) );
  NAND U10831 ( .A(x[142]), .B(y[744]), .Z(n10567) );
  NAND U10832 ( .A(x[131]), .B(y[755]), .Z(n10566) );
  XOR U10833 ( .A(n10567), .B(n10566), .Z(n10568) );
  NAND U10834 ( .A(y[739]), .B(x[147]), .Z(n10569) );
  XOR U10835 ( .A(n10568), .B(n10569), .Z(n10535) );
  XNOR U10836 ( .A(n10534), .B(n10535), .Z(n10537) );
  XNOR U10837 ( .A(n10536), .B(n10537), .Z(n10479) );
  XNOR U10838 ( .A(n10478), .B(n10479), .Z(n10480) );
  XOR U10839 ( .A(n10481), .B(n10480), .Z(n10473) );
  XOR U10840 ( .A(n10472), .B(n10473), .Z(n10474) );
  XNOR U10841 ( .A(n10469), .B(n10468), .Z(n10462) );
  NAND U10842 ( .A(n10425), .B(n10424), .Z(n10429) );
  NANDN U10843 ( .A(n10427), .B(n10426), .Z(n10428) );
  NAND U10844 ( .A(n10429), .B(n10428), .Z(n10461) );
  OR U10845 ( .A(n10431), .B(n10430), .Z(n10435) );
  OR U10846 ( .A(n10433), .B(n10432), .Z(n10434) );
  NAND U10847 ( .A(n10435), .B(n10434), .Z(n10575) );
  OR U10848 ( .A(n10437), .B(n10436), .Z(n10441) );
  OR U10849 ( .A(n10439), .B(n10438), .Z(n10440) );
  NAND U10850 ( .A(n10441), .B(n10440), .Z(n10573) );
  NANDN U10851 ( .A(n10443), .B(n10442), .Z(n10447) );
  OR U10852 ( .A(n10445), .B(n10444), .Z(n10446) );
  NAND U10853 ( .A(n10447), .B(n10446), .Z(n10572) );
  XOR U10854 ( .A(n10573), .B(n10572), .Z(n10574) );
  XOR U10855 ( .A(n10461), .B(n10460), .Z(n10463) );
  XNOR U10856 ( .A(n10462), .B(n10463), .Z(n10580) );
  XNOR U10857 ( .A(n10581), .B(n10580), .Z(n10455) );
  XOR U10858 ( .A(n10457), .B(n10456), .Z(n10451) );
  XOR U10859 ( .A(n10450), .B(n10451), .Z(N247) );
  NANDN U10860 ( .A(n10449), .B(n10448), .Z(n10453) );
  NANDN U10861 ( .A(n10451), .B(n10450), .Z(n10452) );
  NAND U10862 ( .A(n10453), .B(n10452), .Z(n10584) );
  NANDN U10863 ( .A(n10455), .B(n10454), .Z(n10459) );
  NAND U10864 ( .A(n10457), .B(n10456), .Z(n10458) );
  NAND U10865 ( .A(n10459), .B(n10458), .Z(n10585) );
  XNOR U10866 ( .A(n10584), .B(n10585), .Z(n10586) );
  NANDN U10867 ( .A(n10461), .B(n10460), .Z(n10465) );
  OR U10868 ( .A(n10463), .B(n10462), .Z(n10464) );
  AND U10869 ( .A(n10465), .B(n10464), .Z(n10590) );
  NAND U10870 ( .A(n10467), .B(n10466), .Z(n10471) );
  NANDN U10871 ( .A(n10469), .B(n10468), .Z(n10470) );
  NAND U10872 ( .A(n10471), .B(n10470), .Z(n10615) );
  OR U10873 ( .A(n10473), .B(n10472), .Z(n10477) );
  NANDN U10874 ( .A(n10475), .B(n10474), .Z(n10476) );
  NAND U10875 ( .A(n10477), .B(n10476), .Z(n10611) );
  OR U10876 ( .A(n10479), .B(n10478), .Z(n10483) );
  OR U10877 ( .A(n10481), .B(n10480), .Z(n10482) );
  AND U10878 ( .A(n10483), .B(n10482), .Z(n10608) );
  OR U10879 ( .A(n10485), .B(n10484), .Z(n10489) );
  OR U10880 ( .A(n10487), .B(n10486), .Z(n10488) );
  AND U10881 ( .A(n10489), .B(n10488), .Z(n10609) );
  XOR U10882 ( .A(n10608), .B(n10609), .Z(n10610) );
  XOR U10883 ( .A(n10615), .B(n10614), .Z(n10617) );
  NAND U10884 ( .A(x[141]), .B(y[746]), .Z(n10645) );
  NAND U10885 ( .A(x[130]), .B(y[757]), .Z(n10644) );
  XOR U10886 ( .A(n10645), .B(n10644), .Z(n10646) );
  NAND U10887 ( .A(x[149]), .B(y[738]), .Z(n10647) );
  XNOR U10888 ( .A(n10646), .B(n10647), .Z(n10676) );
  OR U10889 ( .A(n10491), .B(n10490), .Z(n10495) );
  NANDN U10890 ( .A(n10493), .B(n10492), .Z(n10494) );
  NAND U10891 ( .A(n10495), .B(n10494), .Z(n10674) );
  NANDN U10892 ( .A(n10496), .B(o[118]), .Z(n10702) );
  NAND U10893 ( .A(x[140]), .B(y[747]), .Z(n10700) );
  NAND U10894 ( .A(x[129]), .B(y[758]), .Z(n10699) );
  XOR U10895 ( .A(n10700), .B(n10699), .Z(n10701) );
  XOR U10896 ( .A(n10702), .B(n10701), .Z(n10675) );
  XOR U10897 ( .A(n10674), .B(n10675), .Z(n10677) );
  XOR U10898 ( .A(n10676), .B(n10677), .Z(n10688) );
  NAND U10899 ( .A(x[142]), .B(y[745]), .Z(n10639) );
  NAND U10900 ( .A(y[756]), .B(x[131]), .Z(n10638) );
  XOR U10901 ( .A(n10639), .B(n10638), .Z(n10640) );
  NAND U10902 ( .A(x[132]), .B(y[755]), .Z(n10641) );
  XNOR U10903 ( .A(n10640), .B(n10641), .Z(n10658) );
  OR U10904 ( .A(n10498), .B(n10497), .Z(n10502) );
  NANDN U10905 ( .A(n10500), .B(n10499), .Z(n10501) );
  NAND U10906 ( .A(n10502), .B(n10501), .Z(n10656) );
  NAND U10907 ( .A(x[133]), .B(y[754]), .Z(n10633) );
  NAND U10908 ( .A(x[146]), .B(y[741]), .Z(n10632) );
  XOR U10909 ( .A(n10633), .B(n10632), .Z(n10634) );
  NAND U10910 ( .A(y[742]), .B(x[145]), .Z(n10635) );
  XOR U10911 ( .A(n10634), .B(n10635), .Z(n10657) );
  XOR U10912 ( .A(n10656), .B(n10657), .Z(n10659) );
  XOR U10913 ( .A(n10658), .B(n10659), .Z(n10686) );
  OR U10914 ( .A(n10504), .B(n10503), .Z(n10508) );
  NANDN U10915 ( .A(n10506), .B(n10505), .Z(n10507) );
  NAND U10916 ( .A(n10508), .B(n10507), .Z(n10687) );
  XOR U10917 ( .A(n10688), .B(n10689), .Z(n10680) );
  NANDN U10918 ( .A(n10510), .B(n10509), .Z(n10514) );
  OR U10919 ( .A(n10512), .B(n10511), .Z(n10513) );
  AND U10920 ( .A(n10514), .B(n10513), .Z(n10681) );
  XOR U10921 ( .A(n10680), .B(n10681), .Z(n10683) );
  NAND U10922 ( .A(x[128]), .B(y[759]), .Z(n10694) );
  NAND U10923 ( .A(x[151]), .B(y[736]), .Z(n10693) );
  XOR U10924 ( .A(n10694), .B(n10693), .Z(n10695) );
  NAND U10925 ( .A(x[150]), .B(y[737]), .Z(n10721) );
  XOR U10926 ( .A(o[119]), .B(n10721), .Z(n10696) );
  XOR U10927 ( .A(n10695), .B(n10696), .Z(n10664) );
  ANDN U10928 ( .B(y[740]), .A(n170), .Z(n10952) );
  AND U10929 ( .A(x[148]), .B(y[739]), .Z(n10516) );
  NAND U10930 ( .A(x[144]), .B(y[743]), .Z(n10515) );
  XOR U10931 ( .A(n10516), .B(n10515), .Z(n10718) );
  XOR U10932 ( .A(n10952), .B(n10718), .Z(n10662) );
  NANDN U10933 ( .A(n10518), .B(n10517), .Z(n10522) );
  NAND U10934 ( .A(n10520), .B(n10519), .Z(n10521) );
  NAND U10935 ( .A(n10522), .B(n10521), .Z(n10663) );
  XOR U10936 ( .A(n10664), .B(n10665), .Z(n10670) );
  NANDN U10937 ( .A(n10523), .B(n11442), .Z(n10527) );
  OR U10938 ( .A(n10525), .B(n10524), .Z(n10526) );
  NAND U10939 ( .A(n10527), .B(n10526), .Z(n10668) );
  OR U10940 ( .A(n10529), .B(n10528), .Z(n10533) );
  NANDN U10941 ( .A(n10531), .B(n10530), .Z(n10532) );
  AND U10942 ( .A(n10533), .B(n10532), .Z(n10669) );
  XNOR U10943 ( .A(n10683), .B(n10682), .Z(n10596) );
  OR U10944 ( .A(n10535), .B(n10534), .Z(n10539) );
  NANDN U10945 ( .A(n10537), .B(n10536), .Z(n10538) );
  AND U10946 ( .A(n10539), .B(n10538), .Z(n10620) );
  OR U10947 ( .A(n10541), .B(n10540), .Z(n10545) );
  NANDN U10948 ( .A(n10543), .B(n10542), .Z(n10544) );
  AND U10949 ( .A(n10545), .B(n10544), .Z(n10621) );
  XOR U10950 ( .A(n10620), .B(n10621), .Z(n10622) );
  OR U10951 ( .A(n10547), .B(n10546), .Z(n10551) );
  NANDN U10952 ( .A(n10549), .B(n10548), .Z(n10550) );
  NAND U10953 ( .A(n10551), .B(n10550), .Z(n10623) );
  NANDN U10954 ( .A(n10553), .B(n10552), .Z(n10557) );
  OR U10955 ( .A(n10555), .B(n10554), .Z(n10556) );
  AND U10956 ( .A(n10557), .B(n10556), .Z(n10602) );
  AND U10957 ( .A(x[136]), .B(y[751]), .Z(n10559) );
  NAND U10958 ( .A(x[137]), .B(y[750]), .Z(n10558) );
  XOR U10959 ( .A(n10559), .B(n10558), .Z(n10708) );
  NAND U10960 ( .A(x[135]), .B(y[752]), .Z(n10707) );
  XOR U10961 ( .A(n10708), .B(n10707), .Z(n10650) );
  NAND U10962 ( .A(y[749]), .B(x[138]), .Z(n10651) );
  XNOR U10963 ( .A(n10650), .B(n10651), .Z(n10652) );
  NAND U10964 ( .A(x[134]), .B(y[753]), .Z(n10712) );
  NAND U10965 ( .A(y[744]), .B(x[143]), .Z(n10711) );
  XOR U10966 ( .A(n10712), .B(n10711), .Z(n10714) );
  XNOR U10967 ( .A(n10713), .B(n10714), .Z(n10653) );
  XOR U10968 ( .A(n10652), .B(n10653), .Z(n10629) );
  NANDN U10969 ( .A(n10561), .B(n10560), .Z(n10565) );
  OR U10970 ( .A(n10563), .B(n10562), .Z(n10564) );
  NAND U10971 ( .A(n10565), .B(n10564), .Z(n10627) );
  OR U10972 ( .A(n10567), .B(n10566), .Z(n10571) );
  NANDN U10973 ( .A(n10569), .B(n10568), .Z(n10570) );
  AND U10974 ( .A(n10571), .B(n10570), .Z(n10626) );
  XOR U10975 ( .A(n10629), .B(n10628), .Z(n10603) );
  XOR U10976 ( .A(n10602), .B(n10603), .Z(n10604) );
  XNOR U10977 ( .A(n10605), .B(n10604), .Z(n10597) );
  XNOR U10978 ( .A(n10596), .B(n10597), .Z(n10599) );
  OR U10979 ( .A(n10573), .B(n10572), .Z(n10577) );
  NANDN U10980 ( .A(n10575), .B(n10574), .Z(n10576) );
  AND U10981 ( .A(n10577), .B(n10576), .Z(n10598) );
  XNOR U10982 ( .A(n10599), .B(n10598), .Z(n10616) );
  XNOR U10983 ( .A(n10617), .B(n10616), .Z(n10591) );
  XOR U10984 ( .A(n10590), .B(n10591), .Z(n10592) );
  OR U10985 ( .A(n10579), .B(n10578), .Z(n10583) );
  NAND U10986 ( .A(n10581), .B(n10580), .Z(n10582) );
  NAND U10987 ( .A(n10583), .B(n10582), .Z(n10593) );
  XOR U10988 ( .A(n10586), .B(n10587), .Z(N248) );
  NANDN U10989 ( .A(n10585), .B(n10584), .Z(n10589) );
  NANDN U10990 ( .A(n10587), .B(n10586), .Z(n10588) );
  NAND U10991 ( .A(n10589), .B(n10588), .Z(n10722) );
  OR U10992 ( .A(n10591), .B(n10590), .Z(n10595) );
  NANDN U10993 ( .A(n10593), .B(n10592), .Z(n10594) );
  AND U10994 ( .A(n10595), .B(n10594), .Z(n10723) );
  XNOR U10995 ( .A(n10722), .B(n10723), .Z(n10724) );
  OR U10996 ( .A(n10597), .B(n10596), .Z(n10601) );
  OR U10997 ( .A(n10599), .B(n10598), .Z(n10600) );
  AND U10998 ( .A(n10601), .B(n10600), .Z(n10860) );
  OR U10999 ( .A(n10603), .B(n10602), .Z(n10607) );
  NANDN U11000 ( .A(n10605), .B(n10604), .Z(n10606) );
  NAND U11001 ( .A(n10607), .B(n10606), .Z(n10858) );
  OR U11002 ( .A(n10609), .B(n10608), .Z(n10613) );
  NANDN U11003 ( .A(n10611), .B(n10610), .Z(n10612) );
  AND U11004 ( .A(n10613), .B(n10612), .Z(n10857) );
  XOR U11005 ( .A(n10858), .B(n10857), .Z(n10859) );
  NANDN U11006 ( .A(n10615), .B(n10614), .Z(n10619) );
  OR U11007 ( .A(n10617), .B(n10616), .Z(n10618) );
  AND U11008 ( .A(n10619), .B(n10618), .Z(n10729) );
  OR U11009 ( .A(n10621), .B(n10620), .Z(n10625) );
  NANDN U11010 ( .A(n10623), .B(n10622), .Z(n10624) );
  NAND U11011 ( .A(n10625), .B(n10624), .Z(n10864) );
  NANDN U11012 ( .A(n10627), .B(n10626), .Z(n10631) );
  NAND U11013 ( .A(n10629), .B(n10628), .Z(n10630) );
  NAND U11014 ( .A(n10631), .B(n10630), .Z(n10742) );
  OR U11015 ( .A(n10633), .B(n10632), .Z(n10637) );
  NANDN U11016 ( .A(n10635), .B(n10634), .Z(n10636) );
  NAND U11017 ( .A(n10637), .B(n10636), .Z(n10828) );
  NAND U11018 ( .A(x[128]), .B(y[760]), .Z(n10784) );
  AND U11019 ( .A(y[736]), .B(x[152]), .Z(n10783) );
  XNOR U11020 ( .A(n10784), .B(n10783), .Z(n10785) );
  NAND U11021 ( .A(x[151]), .B(y[737]), .Z(n10764) );
  XOR U11022 ( .A(o[120]), .B(n10764), .Z(n10786) );
  NAND U11023 ( .A(x[135]), .B(y[753]), .Z(n10759) );
  NAND U11024 ( .A(x[145]), .B(y[743]), .Z(n10758) );
  XOR U11025 ( .A(n10759), .B(n10758), .Z(n10760) );
  NAND U11026 ( .A(y[742]), .B(x[146]), .Z(n10761) );
  XNOR U11027 ( .A(n10760), .B(n10761), .Z(n10825) );
  XNOR U11028 ( .A(n10826), .B(n10825), .Z(n10827) );
  XNOR U11029 ( .A(n10828), .B(n10827), .Z(n10854) );
  OR U11030 ( .A(n10639), .B(n10638), .Z(n10643) );
  NANDN U11031 ( .A(n10641), .B(n10640), .Z(n10642) );
  NAND U11032 ( .A(n10643), .B(n10642), .Z(n10851) );
  OR U11033 ( .A(n10645), .B(n10644), .Z(n10649) );
  NANDN U11034 ( .A(n10647), .B(n10646), .Z(n10648) );
  AND U11035 ( .A(n10649), .B(n10648), .Z(n10852) );
  XOR U11036 ( .A(n10854), .B(n10853), .Z(n10740) );
  NANDN U11037 ( .A(n10651), .B(n10650), .Z(n10655) );
  NANDN U11038 ( .A(n10653), .B(n10652), .Z(n10654) );
  NAND U11039 ( .A(n10655), .B(n10654), .Z(n10741) );
  XOR U11040 ( .A(n10742), .B(n10743), .Z(n10804) );
  NANDN U11041 ( .A(n10657), .B(n10656), .Z(n10661) );
  NANDN U11042 ( .A(n10659), .B(n10658), .Z(n10660) );
  NAND U11043 ( .A(n10661), .B(n10660), .Z(n10810) );
  NANDN U11044 ( .A(n10663), .B(n10662), .Z(n10667) );
  NANDN U11045 ( .A(n10665), .B(n10664), .Z(n10666) );
  AND U11046 ( .A(n10667), .B(n10666), .Z(n10807) );
  NANDN U11047 ( .A(n10669), .B(n10668), .Z(n10673) );
  NAND U11048 ( .A(n10671), .B(n10670), .Z(n10672) );
  NAND U11049 ( .A(n10673), .B(n10672), .Z(n10808) );
  XOR U11050 ( .A(n10807), .B(n10808), .Z(n10809) );
  XNOR U11051 ( .A(n10810), .B(n10809), .Z(n10802) );
  NANDN U11052 ( .A(n10675), .B(n10674), .Z(n10679) );
  NANDN U11053 ( .A(n10677), .B(n10676), .Z(n10678) );
  AND U11054 ( .A(n10679), .B(n10678), .Z(n10801) );
  XOR U11055 ( .A(n10802), .B(n10801), .Z(n10803) );
  XOR U11056 ( .A(n10804), .B(n10803), .Z(n10863) );
  XNOR U11057 ( .A(n10864), .B(n10863), .Z(n10866) );
  NANDN U11058 ( .A(n10681), .B(n10680), .Z(n10685) );
  NANDN U11059 ( .A(n10683), .B(n10682), .Z(n10684) );
  NAND U11060 ( .A(n10685), .B(n10684), .Z(n10737) );
  NANDN U11061 ( .A(n10687), .B(n10686), .Z(n10691) );
  NANDN U11062 ( .A(n10689), .B(n10688), .Z(n10690) );
  NAND U11063 ( .A(n10691), .B(n10690), .Z(n10734) );
  NAND U11064 ( .A(x[136]), .B(y[752]), .Z(n10772) );
  AND U11065 ( .A(x[139]), .B(y[749]), .Z(n10771) );
  XNOR U11066 ( .A(n10772), .B(n10771), .Z(n10773) );
  NAND U11067 ( .A(x[142]), .B(y[746]), .Z(n10774) );
  XNOR U11068 ( .A(n10773), .B(n10774), .Z(n10768) );
  NOR U11069 ( .A(n160), .B(n10692), .Z(n10705) );
  IV U11070 ( .A(n10705), .Z(n10765) );
  ANDN U11071 ( .B(y[750]), .A(n161), .Z(n10766) );
  XNOR U11072 ( .A(n10765), .B(n10766), .Z(n10767) );
  XNOR U11073 ( .A(n10768), .B(n10767), .Z(n10790) );
  OR U11074 ( .A(n10694), .B(n10693), .Z(n10698) );
  NANDN U11075 ( .A(n10696), .B(n10695), .Z(n10697) );
  AND U11076 ( .A(n10698), .B(n10697), .Z(n10789) );
  XOR U11077 ( .A(n10790), .B(n10789), .Z(n10792) );
  NAND U11078 ( .A(x[143]), .B(y[745]), .Z(n10778) );
  NAND U11079 ( .A(x[131]), .B(y[757]), .Z(n10777) );
  XOR U11080 ( .A(n10778), .B(n10777), .Z(n10779) );
  NAND U11081 ( .A(y[756]), .B(x[132]), .Z(n10780) );
  XNOR U11082 ( .A(n10779), .B(n10780), .Z(n10791) );
  OR U11083 ( .A(n10700), .B(n10699), .Z(n10704) );
  NANDN U11084 ( .A(n10702), .B(n10701), .Z(n10703) );
  NAND U11085 ( .A(n10704), .B(n10703), .Z(n10847) );
  NANDN U11086 ( .A(n10706), .B(n10705), .Z(n10710) );
  OR U11087 ( .A(n10708), .B(n10707), .Z(n10709) );
  NAND U11088 ( .A(n10710), .B(n10709), .Z(n10845) );
  NAND U11089 ( .A(x[149]), .B(y[739]), .Z(n10832) );
  NAND U11090 ( .A(x[133]), .B(y[755]), .Z(n10831) );
  XOR U11091 ( .A(n10832), .B(n10831), .Z(n10833) );
  NAND U11092 ( .A(y[744]), .B(x[144]), .Z(n10834) );
  XOR U11093 ( .A(n10833), .B(n10834), .Z(n10822) );
  OR U11094 ( .A(n10712), .B(n10711), .Z(n10716) );
  NAND U11095 ( .A(n10714), .B(n10713), .Z(n10715) );
  AND U11096 ( .A(n10716), .B(n10715), .Z(n10819) );
  NAND U11097 ( .A(x[134]), .B(y[754]), .Z(n10840) );
  NAND U11098 ( .A(x[147]), .B(y[741]), .Z(n10839) );
  XOR U11099 ( .A(n10840), .B(n10839), .Z(n10841) );
  NAND U11100 ( .A(x[148]), .B(y[740]), .Z(n10842) );
  XOR U11101 ( .A(n10841), .B(n10842), .Z(n10820) );
  XNOR U11102 ( .A(n10819), .B(n10820), .Z(n10821) );
  XNOR U11103 ( .A(n10822), .B(n10821), .Z(n10846) );
  NAND U11104 ( .A(x[150]), .B(y[738]), .Z(n10753) );
  NAND U11105 ( .A(x[130]), .B(y[758]), .Z(n10752) );
  XOR U11106 ( .A(n10753), .B(n10752), .Z(n10755) );
  XNOR U11107 ( .A(n10754), .B(n10755), .Z(n10816) );
  AND U11108 ( .A(y[739]), .B(x[144]), .Z(n10717) );
  AND U11109 ( .A(y[743]), .B(x[148]), .Z(n11223) );
  NAND U11110 ( .A(n10717), .B(n11223), .Z(n10720) );
  NANDN U11111 ( .A(n10718), .B(n10952), .Z(n10719) );
  NAND U11112 ( .A(n10720), .B(n10719), .Z(n10814) );
  NANDN U11113 ( .A(n10721), .B(o[119]), .Z(n10749) );
  NAND U11114 ( .A(x[129]), .B(y[759]), .Z(n10747) );
  XOR U11115 ( .A(n10746), .B(n10747), .Z(n10748) );
  XOR U11116 ( .A(n10749), .B(n10748), .Z(n10813) );
  XNOR U11117 ( .A(n10814), .B(n10813), .Z(n10815) );
  XOR U11118 ( .A(n10816), .B(n10815), .Z(n10796) );
  XOR U11119 ( .A(n10795), .B(n10796), .Z(n10797) );
  XNOR U11120 ( .A(n10798), .B(n10797), .Z(n10735) );
  XOR U11121 ( .A(n10737), .B(n10736), .Z(n10865) );
  XOR U11122 ( .A(n10866), .B(n10865), .Z(n10728) );
  XOR U11123 ( .A(n10729), .B(n10728), .Z(n10730) );
  XNOR U11124 ( .A(n10731), .B(n10730), .Z(n10725) );
  XOR U11125 ( .A(n10724), .B(n10725), .Z(N249) );
  NANDN U11126 ( .A(n10723), .B(n10722), .Z(n10727) );
  NANDN U11127 ( .A(n10725), .B(n10724), .Z(n10726) );
  NAND U11128 ( .A(n10727), .B(n10726), .Z(n10869) );
  NANDN U11129 ( .A(n10729), .B(n10728), .Z(n10733) );
  OR U11130 ( .A(n10731), .B(n10730), .Z(n10732) );
  AND U11131 ( .A(n10733), .B(n10732), .Z(n10870) );
  XNOR U11132 ( .A(n10869), .B(n10870), .Z(n10871) );
  NANDN U11133 ( .A(n10735), .B(n10734), .Z(n10739) );
  NANDN U11134 ( .A(n10737), .B(n10736), .Z(n10738) );
  NAND U11135 ( .A(n10739), .B(n10738), .Z(n11007) );
  NANDN U11136 ( .A(n10741), .B(n10740), .Z(n10745) );
  NANDN U11137 ( .A(n10743), .B(n10742), .Z(n10744) );
  NAND U11138 ( .A(n10745), .B(n10744), .Z(n11001) );
  NANDN U11139 ( .A(n10747), .B(n10746), .Z(n10751) );
  OR U11140 ( .A(n10749), .B(n10748), .Z(n10750) );
  NAND U11141 ( .A(n10751), .B(n10750), .Z(n10889) );
  OR U11142 ( .A(n10753), .B(n10752), .Z(n10757) );
  NAND U11143 ( .A(n10755), .B(n10754), .Z(n10756) );
  NAND U11144 ( .A(n10757), .B(n10756), .Z(n10887) );
  OR U11145 ( .A(n10759), .B(n10758), .Z(n10763) );
  NANDN U11146 ( .A(n10761), .B(n10760), .Z(n10762) );
  AND U11147 ( .A(n10763), .B(n10762), .Z(n10895) );
  NAND U11148 ( .A(y[753]), .B(x[136]), .Z(n10906) );
  XOR U11149 ( .A(n10906), .B(n10905), .Z(n10894) );
  NANDN U11150 ( .A(n10764), .B(o[120]), .Z(n10902) );
  AND U11151 ( .A(y[736]), .B(x[153]), .Z(n10899) );
  AND U11152 ( .A(y[761]), .B(x[128]), .Z(n10900) );
  XNOR U11153 ( .A(n10899), .B(n10900), .Z(n10901) );
  XOR U11154 ( .A(n10902), .B(n10901), .Z(n10893) );
  XNOR U11155 ( .A(n10895), .B(n10896), .Z(n10888) );
  XOR U11156 ( .A(n10889), .B(n10890), .Z(n10912) );
  NANDN U11157 ( .A(n10766), .B(n10765), .Z(n10770) );
  NANDN U11158 ( .A(n10768), .B(n10767), .Z(n10769) );
  NAND U11159 ( .A(n10770), .B(n10769), .Z(n10909) );
  NAND U11160 ( .A(x[139]), .B(y[750]), .Z(n10937) );
  AND U11161 ( .A(x[140]), .B(y[749]), .Z(n10934) );
  AND U11162 ( .A(x[135]), .B(y[754]), .Z(n10935) );
  XNOR U11163 ( .A(n10934), .B(n10935), .Z(n10936) );
  XOR U11164 ( .A(n10937), .B(n10936), .Z(n10969) );
  NANDN U11165 ( .A(n10772), .B(n10771), .Z(n10776) );
  NANDN U11166 ( .A(n10774), .B(n10773), .Z(n10775) );
  AND U11167 ( .A(n10776), .B(n10775), .Z(n10970) );
  NAND U11168 ( .A(x[141]), .B(y[748]), .Z(n10964) );
  AND U11169 ( .A(y[760]), .B(x[129]), .Z(n10963) );
  XNOR U11170 ( .A(n10964), .B(n10963), .Z(n10965) );
  ANDN U11171 ( .B(y[737]), .A(n175), .Z(n10933) );
  XNOR U11172 ( .A(o[121]), .B(n10933), .Z(n10966) );
  XNOR U11173 ( .A(n10971), .B(n10972), .Z(n10910) );
  XOR U11174 ( .A(n10912), .B(n10911), .Z(n10995) );
  OR U11175 ( .A(n10778), .B(n10777), .Z(n10782) );
  NANDN U11176 ( .A(n10780), .B(n10779), .Z(n10781) );
  NAND U11177 ( .A(n10782), .B(n10781), .Z(n10977) );
  NANDN U11178 ( .A(n10784), .B(n10783), .Z(n10788) );
  NANDN U11179 ( .A(n10786), .B(n10785), .Z(n10787) );
  NAND U11180 ( .A(n10788), .B(n10787), .Z(n10976) );
  NAND U11181 ( .A(x[130]), .B(y[759]), .Z(n10958) );
  XOR U11182 ( .A(n10957), .B(n10958), .Z(n10960) );
  NAND U11183 ( .A(x[131]), .B(y[758]), .Z(n10959) );
  XOR U11184 ( .A(n10960), .B(n10959), .Z(n10975) );
  XNOR U11185 ( .A(n10976), .B(n10975), .Z(n10978) );
  XNOR U11186 ( .A(n10977), .B(n10978), .Z(n10993) );
  OR U11187 ( .A(n10790), .B(n10789), .Z(n10794) );
  NAND U11188 ( .A(n10792), .B(n10791), .Z(n10793) );
  AND U11189 ( .A(n10794), .B(n10793), .Z(n10994) );
  XOR U11190 ( .A(n10993), .B(n10994), .Z(n10996) );
  XOR U11191 ( .A(n10995), .B(n10996), .Z(n11000) );
  NANDN U11192 ( .A(n10796), .B(n10795), .Z(n10800) );
  OR U11193 ( .A(n10798), .B(n10797), .Z(n10799) );
  AND U11194 ( .A(n10800), .B(n10799), .Z(n10999) );
  XNOR U11195 ( .A(n11000), .B(n10999), .Z(n11002) );
  XOR U11196 ( .A(n11001), .B(n11002), .Z(n11005) );
  OR U11197 ( .A(n10802), .B(n10801), .Z(n10806) );
  NAND U11198 ( .A(n10804), .B(n10803), .Z(n10805) );
  NAND U11199 ( .A(n10806), .B(n10805), .Z(n10884) );
  OR U11200 ( .A(n10808), .B(n10807), .Z(n10812) );
  NANDN U11201 ( .A(n10810), .B(n10809), .Z(n10811) );
  AND U11202 ( .A(n10812), .B(n10811), .Z(n10882) );
  NAND U11203 ( .A(n10814), .B(n10813), .Z(n10818) );
  OR U11204 ( .A(n10816), .B(n10815), .Z(n10817) );
  AND U11205 ( .A(n10818), .B(n10817), .Z(n10930) );
  OR U11206 ( .A(n10820), .B(n10819), .Z(n10824) );
  OR U11207 ( .A(n10822), .B(n10821), .Z(n10823) );
  AND U11208 ( .A(n10824), .B(n10823), .Z(n10928) );
  NANDN U11209 ( .A(n10826), .B(n10825), .Z(n10830) );
  NAND U11210 ( .A(n10828), .B(n10827), .Z(n10829) );
  AND U11211 ( .A(n10830), .B(n10829), .Z(n10917) );
  OR U11212 ( .A(n10832), .B(n10831), .Z(n10836) );
  NANDN U11213 ( .A(n10834), .B(n10833), .Z(n10835) );
  AND U11214 ( .A(n10836), .B(n10835), .Z(n10983) );
  NAND U11215 ( .A(y[739]), .B(x[150]), .Z(n10940) );
  AND U11216 ( .A(x[133]), .B(y[756]), .Z(n10938) );
  AND U11217 ( .A(x[145]), .B(y[744]), .Z(n10939) );
  XOR U11218 ( .A(n10938), .B(n10939), .Z(n10941) );
  XNOR U11219 ( .A(n10940), .B(n10941), .Z(n10981) );
  AND U11220 ( .A(x[147]), .B(y[742]), .Z(n10838) );
  NAND U11221 ( .A(x[149]), .B(y[740]), .Z(n10837) );
  XOR U11222 ( .A(n10838), .B(n10837), .Z(n10954) );
  AND U11223 ( .A(y[741]), .B(x[148]), .Z(n10953) );
  XOR U11224 ( .A(n10954), .B(n10953), .Z(n10982) );
  XOR U11225 ( .A(n10981), .B(n10982), .Z(n10984) );
  XNOR U11226 ( .A(n10983), .B(n10984), .Z(n10916) );
  NAND U11227 ( .A(x[151]), .B(y[738]), .Z(n10947) );
  AND U11228 ( .A(y[757]), .B(x[132]), .Z(n10944) );
  AND U11229 ( .A(y[745]), .B(x[144]), .Z(n10945) );
  XNOR U11230 ( .A(n10944), .B(n10945), .Z(n10946) );
  XNOR U11231 ( .A(n10947), .B(n10946), .Z(n10989) );
  NAND U11232 ( .A(y[746]), .B(x[143]), .Z(n10951) );
  AND U11233 ( .A(y[743]), .B(x[146]), .Z(n10948) );
  AND U11234 ( .A(y[755]), .B(x[134]), .Z(n10949) );
  XNOR U11235 ( .A(n10948), .B(n10949), .Z(n10950) );
  XOR U11236 ( .A(n10951), .B(n10950), .Z(n10987) );
  OR U11237 ( .A(n10840), .B(n10839), .Z(n10844) );
  NANDN U11238 ( .A(n10842), .B(n10841), .Z(n10843) );
  AND U11239 ( .A(n10844), .B(n10843), .Z(n10988) );
  XOR U11240 ( .A(n10989), .B(n10990), .Z(n10915) );
  XOR U11241 ( .A(n10916), .B(n10915), .Z(n10918) );
  XOR U11242 ( .A(n10917), .B(n10918), .Z(n10927) );
  XNOR U11243 ( .A(n10928), .B(n10927), .Z(n10929) );
  XOR U11244 ( .A(n10930), .B(n10929), .Z(n10923) );
  NANDN U11245 ( .A(n10846), .B(n10845), .Z(n10850) );
  NANDN U11246 ( .A(n10848), .B(n10847), .Z(n10849) );
  NAND U11247 ( .A(n10850), .B(n10849), .Z(n10922) );
  NANDN U11248 ( .A(n10852), .B(n10851), .Z(n10856) );
  NANDN U11249 ( .A(n10854), .B(n10853), .Z(n10855) );
  AND U11250 ( .A(n10856), .B(n10855), .Z(n10921) );
  XOR U11251 ( .A(n10882), .B(n10881), .Z(n10883) );
  XOR U11252 ( .A(n10884), .B(n10883), .Z(n11006) );
  XOR U11253 ( .A(n11005), .B(n11006), .Z(n11008) );
  XOR U11254 ( .A(n11007), .B(n11008), .Z(n10878) );
  OR U11255 ( .A(n10858), .B(n10857), .Z(n10862) );
  NANDN U11256 ( .A(n10860), .B(n10859), .Z(n10861) );
  AND U11257 ( .A(n10862), .B(n10861), .Z(n10875) );
  OR U11258 ( .A(n10864), .B(n10863), .Z(n10868) );
  OR U11259 ( .A(n10866), .B(n10865), .Z(n10867) );
  AND U11260 ( .A(n10868), .B(n10867), .Z(n10876) );
  XOR U11261 ( .A(n10875), .B(n10876), .Z(n10877) );
  XOR U11262 ( .A(n10878), .B(n10877), .Z(n10872) );
  XOR U11263 ( .A(n10871), .B(n10872), .Z(N250) );
  NANDN U11264 ( .A(n10870), .B(n10869), .Z(n10874) );
  NANDN U11265 ( .A(n10872), .B(n10871), .Z(n10873) );
  NAND U11266 ( .A(n10874), .B(n10873), .Z(n11011) );
  OR U11267 ( .A(n10876), .B(n10875), .Z(n10880) );
  NANDN U11268 ( .A(n10878), .B(n10877), .Z(n10879) );
  AND U11269 ( .A(n10880), .B(n10879), .Z(n11012) );
  XNOR U11270 ( .A(n11011), .B(n11012), .Z(n11013) );
  NANDN U11271 ( .A(n10882), .B(n10881), .Z(n10886) );
  OR U11272 ( .A(n10884), .B(n10883), .Z(n10885) );
  NAND U11273 ( .A(n10886), .B(n10885), .Z(n11020) );
  NANDN U11274 ( .A(n10888), .B(n10887), .Z(n10892) );
  NANDN U11275 ( .A(n10890), .B(n10889), .Z(n10891) );
  AND U11276 ( .A(n10892), .B(n10891), .Z(n11126) );
  NANDN U11277 ( .A(n10894), .B(n10893), .Z(n10898) );
  OR U11278 ( .A(n10896), .B(n10895), .Z(n10897) );
  AND U11279 ( .A(n10898), .B(n10897), .Z(n11124) );
  NAND U11280 ( .A(x[130]), .B(y[760]), .Z(n11046) );
  XNOR U11281 ( .A(n11046), .B(n11045), .Z(n11048) );
  ANDN U11282 ( .B(y[738]), .A(n175), .Z(n11047) );
  XOR U11283 ( .A(n11048), .B(n11047), .Z(n11082) );
  XOR U11284 ( .A(n11082), .B(n11083), .Z(n11085) );
  OR U11285 ( .A(n10904), .B(n10903), .Z(n10908) );
  NAND U11286 ( .A(n10906), .B(n10905), .Z(n10907) );
  NAND U11287 ( .A(n10908), .B(n10907), .Z(n11084) );
  XNOR U11288 ( .A(n11085), .B(n11084), .Z(n11125) );
  XNOR U11289 ( .A(n11124), .B(n11125), .Z(n11127) );
  XNOR U11290 ( .A(n11126), .B(n11127), .Z(n11114) );
  NANDN U11291 ( .A(n10910), .B(n10909), .Z(n10914) );
  NAND U11292 ( .A(n10912), .B(n10911), .Z(n10913) );
  AND U11293 ( .A(n10914), .B(n10913), .Z(n11112) );
  NANDN U11294 ( .A(n10916), .B(n10915), .Z(n10920) );
  OR U11295 ( .A(n10918), .B(n10917), .Z(n10919) );
  NAND U11296 ( .A(n10920), .B(n10919), .Z(n11113) );
  XOR U11297 ( .A(n11112), .B(n11113), .Z(n11115) );
  XNOR U11298 ( .A(n11114), .B(n11115), .Z(n11026) );
  NANDN U11299 ( .A(n10922), .B(n10921), .Z(n10926) );
  NAND U11300 ( .A(n10924), .B(n10923), .Z(n10925) );
  AND U11301 ( .A(n10926), .B(n10925), .Z(n11023) );
  NANDN U11302 ( .A(n10928), .B(n10927), .Z(n10932) );
  NANDN U11303 ( .A(n10930), .B(n10929), .Z(n10931) );
  NAND U11304 ( .A(n10932), .B(n10931), .Z(n11073) );
  AND U11305 ( .A(n10933), .B(o[121]), .Z(n11144) );
  ANDN U11306 ( .B(y[748]), .A(n165), .Z(n11142) );
  ANDN U11307 ( .B(y[761]), .A(n152), .Z(n11143) );
  XNOR U11308 ( .A(n11142), .B(n11143), .Z(n11145) );
  XNOR U11309 ( .A(n11144), .B(n11145), .Z(n11088) );
  NAND U11310 ( .A(x[128]), .B(y[762]), .Z(n11101) );
  AND U11311 ( .A(y[736]), .B(x[154]), .Z(n11100) );
  XNOR U11312 ( .A(n11101), .B(n11100), .Z(n11103) );
  NAND U11313 ( .A(x[153]), .B(y[737]), .Z(n11160) );
  XNOR U11314 ( .A(n11160), .B(o[122]), .Z(n11102) );
  XNOR U11315 ( .A(n11103), .B(n11102), .Z(n11089) );
  XOR U11316 ( .A(n11088), .B(n11089), .Z(n11091) );
  XOR U11317 ( .A(n11091), .B(n11090), .Z(n11032) );
  OR U11318 ( .A(n10939), .B(n10938), .Z(n10943) );
  NAND U11319 ( .A(n10941), .B(n10940), .Z(n10942) );
  AND U11320 ( .A(n10943), .B(n10942), .Z(n11029) );
  XOR U11321 ( .A(n11029), .B(n11030), .Z(n11031) );
  XOR U11322 ( .A(n11032), .B(n11031), .Z(n11109) );
  ANDN U11323 ( .B(y[758]), .A(n155), .Z(n11053) );
  XNOR U11324 ( .A(n11051), .B(n11053), .Z(n11055) );
  XNOR U11325 ( .A(n11054), .B(n11055), .Z(n11033) );
  XOR U11326 ( .A(n11033), .B(n11034), .Z(n11036) );
  NAND U11327 ( .A(x[147]), .B(y[743]), .Z(n11137) );
  AND U11328 ( .A(x[139]), .B(y[751]), .Z(n11136) );
  XNOR U11329 ( .A(n11137), .B(n11136), .Z(n11139) );
  AND U11330 ( .A(y[759]), .B(x[131]), .Z(n11138) );
  XOR U11331 ( .A(n11036), .B(n11035), .Z(n11106) );
  ANDN U11332 ( .B(y[742]), .A(n172), .Z(n11209) );
  NAND U11333 ( .A(n11209), .B(n10952), .Z(n10956) );
  NANDN U11334 ( .A(n10954), .B(n10953), .Z(n10955) );
  NAND U11335 ( .A(n10956), .B(n10955), .Z(n11059) );
  NAND U11336 ( .A(x[150]), .B(y[740]), .Z(n11042) );
  NAND U11337 ( .A(y[739]), .B(x[151]), .Z(n11039) );
  XNOR U11338 ( .A(n11040), .B(n11039), .Z(n11041) );
  XNOR U11339 ( .A(n11042), .B(n11041), .Z(n11058) );
  XNOR U11340 ( .A(n11059), .B(n11058), .Z(n11061) );
  NAND U11341 ( .A(y[742]), .B(x[148]), .Z(n11151) );
  NAND U11342 ( .A(x[149]), .B(y[741]), .Z(n11148) );
  XNOR U11343 ( .A(n11149), .B(n11148), .Z(n11150) );
  XNOR U11344 ( .A(n11151), .B(n11150), .Z(n11060) );
  XNOR U11345 ( .A(n11061), .B(n11060), .Z(n11107) );
  XOR U11346 ( .A(n11106), .B(n11107), .Z(n11108) );
  NANDN U11347 ( .A(n10958), .B(n10957), .Z(n10962) );
  OR U11348 ( .A(n10960), .B(n10959), .Z(n10961) );
  NAND U11349 ( .A(n10962), .B(n10961), .Z(n11065) );
  NANDN U11350 ( .A(n10964), .B(n10963), .Z(n10968) );
  NANDN U11351 ( .A(n10966), .B(n10965), .Z(n10967) );
  NAND U11352 ( .A(n10968), .B(n10967), .Z(n11064) );
  XOR U11353 ( .A(n11065), .B(n11064), .Z(n11066) );
  IV U11354 ( .A(y[756]), .Z(n11458) );
  NANDN U11355 ( .A(n11458), .B(x[134]), .Z(n11154) );
  XNOR U11356 ( .A(n11154), .B(n11155), .Z(n11157) );
  XOR U11357 ( .A(n11156), .B(n11157), .Z(n11133) );
  NAND U11358 ( .A(x[135]), .B(y[755]), .Z(n11130) );
  NAND U11359 ( .A(x[138]), .B(y[752]), .Z(n11097) );
  AND U11360 ( .A(y[750]), .B(x[140]), .Z(n11094) );
  AND U11361 ( .A(y[757]), .B(x[133]), .Z(n11095) );
  XOR U11362 ( .A(n11094), .B(n11095), .Z(n11096) );
  XNOR U11363 ( .A(n11097), .B(n11096), .Z(n11131) );
  XNOR U11364 ( .A(n11130), .B(n11131), .Z(n11132) );
  XOR U11365 ( .A(n11133), .B(n11132), .Z(n11067) );
  NANDN U11366 ( .A(n10970), .B(n10969), .Z(n10974) );
  NANDN U11367 ( .A(n10972), .B(n10971), .Z(n10973) );
  AND U11368 ( .A(n10974), .B(n10973), .Z(n11077) );
  XOR U11369 ( .A(n11076), .B(n11077), .Z(n11078) );
  XNOR U11370 ( .A(n11079), .B(n11078), .Z(n11071) );
  NAND U11371 ( .A(n10976), .B(n10975), .Z(n10980) );
  NANDN U11372 ( .A(n10978), .B(n10977), .Z(n10979) );
  NAND U11373 ( .A(n10980), .B(n10979), .Z(n11121) );
  NANDN U11374 ( .A(n10982), .B(n10981), .Z(n10986) );
  OR U11375 ( .A(n10984), .B(n10983), .Z(n10985) );
  NAND U11376 ( .A(n10986), .B(n10985), .Z(n11119) );
  NANDN U11377 ( .A(n10988), .B(n10987), .Z(n10992) );
  OR U11378 ( .A(n10990), .B(n10989), .Z(n10991) );
  NAND U11379 ( .A(n10992), .B(n10991), .Z(n11118) );
  XNOR U11380 ( .A(n11119), .B(n11118), .Z(n11120) );
  XOR U11381 ( .A(n11121), .B(n11120), .Z(n11070) );
  XOR U11382 ( .A(n11071), .B(n11070), .Z(n11072) );
  XNOR U11383 ( .A(n11073), .B(n11072), .Z(n11024) );
  XNOR U11384 ( .A(n11023), .B(n11024), .Z(n11025) );
  XNOR U11385 ( .A(n11026), .B(n11025), .Z(n11164) );
  NANDN U11386 ( .A(n10994), .B(n10993), .Z(n10998) );
  OR U11387 ( .A(n10996), .B(n10995), .Z(n10997) );
  NAND U11388 ( .A(n10998), .B(n10997), .Z(n11162) );
  OR U11389 ( .A(n11000), .B(n10999), .Z(n11004) );
  NANDN U11390 ( .A(n11002), .B(n11001), .Z(n11003) );
  AND U11391 ( .A(n11004), .B(n11003), .Z(n11161) );
  XOR U11392 ( .A(n11162), .B(n11161), .Z(n11163) );
  XNOR U11393 ( .A(n11164), .B(n11163), .Z(n11018) );
  NANDN U11394 ( .A(n11006), .B(n11005), .Z(n11010) );
  OR U11395 ( .A(n11008), .B(n11007), .Z(n11009) );
  AND U11396 ( .A(n11010), .B(n11009), .Z(n11017) );
  XOR U11397 ( .A(n11018), .B(n11017), .Z(n11019) );
  XNOR U11398 ( .A(n11020), .B(n11019), .Z(n11014) );
  XOR U11399 ( .A(n11013), .B(n11014), .Z(N251) );
  NANDN U11400 ( .A(n11012), .B(n11011), .Z(n11016) );
  NANDN U11401 ( .A(n11014), .B(n11013), .Z(n11015) );
  NAND U11402 ( .A(n11016), .B(n11015), .Z(n11167) );
  OR U11403 ( .A(n11018), .B(n11017), .Z(n11022) );
  NANDN U11404 ( .A(n11020), .B(n11019), .Z(n11021) );
  NAND U11405 ( .A(n11022), .B(n11021), .Z(n11168) );
  XNOR U11406 ( .A(n11167), .B(n11168), .Z(n11169) );
  OR U11407 ( .A(n11024), .B(n11023), .Z(n11028) );
  OR U11408 ( .A(n11026), .B(n11025), .Z(n11027) );
  AND U11409 ( .A(n11028), .B(n11027), .Z(n11173) );
  NANDN U11410 ( .A(n11034), .B(n11033), .Z(n11038) );
  OR U11411 ( .A(n11036), .B(n11035), .Z(n11037) );
  NAND U11412 ( .A(n11038), .B(n11037), .Z(n11303) );
  NANDN U11413 ( .A(n11040), .B(n11039), .Z(n11044) );
  NAND U11414 ( .A(n11042), .B(n11041), .Z(n11043) );
  AND U11415 ( .A(n11044), .B(n11043), .Z(n11254) );
  NANDN U11416 ( .A(n11046), .B(n11045), .Z(n11050) );
  NAND U11417 ( .A(n11048), .B(n11047), .Z(n11049) );
  NAND U11418 ( .A(n11050), .B(n11049), .Z(n11255) );
  XOR U11419 ( .A(n11254), .B(n11255), .Z(n11257) );
  IV U11420 ( .A(n11051), .Z(n11052) );
  NANDN U11421 ( .A(n11053), .B(n11052), .Z(n11057) );
  OR U11422 ( .A(n11055), .B(n11054), .Z(n11056) );
  AND U11423 ( .A(n11057), .B(n11056), .Z(n11248) );
  ANDN U11424 ( .B(y[754]), .A(n160), .Z(n11211) );
  ANDN U11425 ( .B(y[745]), .A(n169), .Z(n11210) );
  XNOR U11426 ( .A(n11209), .B(n11210), .Z(n11212) );
  XNOR U11427 ( .A(n11211), .B(n11212), .Z(n11249) );
  XOR U11428 ( .A(n11248), .B(n11249), .Z(n11250) );
  ANDN U11429 ( .B(y[763]), .A(n151), .Z(n11199) );
  ANDN U11430 ( .B(y[737]), .A(n176), .Z(n11215) );
  XOR U11431 ( .A(o[123]), .B(n11215), .Z(n11197) );
  ANDN U11432 ( .B(y[736]), .A(n177), .Z(n11198) );
  XNOR U11433 ( .A(n11197), .B(n11198), .Z(n11200) );
  XNOR U11434 ( .A(n11199), .B(n11200), .Z(n11251) );
  XNOR U11435 ( .A(n11257), .B(n11256), .Z(n11302) );
  XNOR U11436 ( .A(n11303), .B(n11302), .Z(n11305) );
  XOR U11437 ( .A(n11304), .B(n11305), .Z(n11191) );
  OR U11438 ( .A(n11059), .B(n11058), .Z(n11063) );
  OR U11439 ( .A(n11061), .B(n11060), .Z(n11062) );
  NAND U11440 ( .A(n11063), .B(n11062), .Z(n11192) );
  XOR U11441 ( .A(n11191), .B(n11192), .Z(n11193) );
  OR U11442 ( .A(n11065), .B(n11064), .Z(n11069) );
  NANDN U11443 ( .A(n11067), .B(n11066), .Z(n11068) );
  NAND U11444 ( .A(n11069), .B(n11068), .Z(n11194) );
  XOR U11445 ( .A(n11193), .B(n11194), .Z(n11319) );
  NANDN U11446 ( .A(n11071), .B(n11070), .Z(n11075) );
  OR U11447 ( .A(n11073), .B(n11072), .Z(n11074) );
  NAND U11448 ( .A(n11075), .B(n11074), .Z(n11318) );
  XOR U11449 ( .A(n11319), .B(n11318), .Z(n11320) );
  OR U11450 ( .A(n11077), .B(n11076), .Z(n11081) );
  NANDN U11451 ( .A(n11079), .B(n11078), .Z(n11080) );
  AND U11452 ( .A(n11081), .B(n11080), .Z(n11188) );
  NANDN U11453 ( .A(n11083), .B(n11082), .Z(n11087) );
  OR U11454 ( .A(n11085), .B(n11084), .Z(n11086) );
  NAND U11455 ( .A(n11087), .B(n11086), .Z(n11299) );
  NANDN U11456 ( .A(n11089), .B(n11088), .Z(n11093) );
  OR U11457 ( .A(n11091), .B(n11090), .Z(n11092) );
  NAND U11458 ( .A(n11093), .B(n11092), .Z(n11297) );
  ANDN U11459 ( .B(y[751]), .A(n163), .Z(n11272) );
  ANDN U11460 ( .B(y[750]), .A(n164), .Z(n11273) );
  XNOR U11461 ( .A(n11272), .B(n11273), .Z(n11275) );
  NAND U11462 ( .A(x[139]), .B(y[752]), .Z(n11287) );
  NAND U11463 ( .A(x[144]), .B(y[747]), .Z(n11284) );
  XNOR U11464 ( .A(n11285), .B(n11284), .Z(n11286) );
  XNOR U11465 ( .A(n11287), .B(n11286), .Z(n11274) );
  XNOR U11466 ( .A(n11275), .B(n11274), .Z(n11234) );
  ANDN U11467 ( .B(y[760]), .A(n154), .Z(n11280) );
  ANDN U11468 ( .B(y[761]), .A(n153), .Z(n11278) );
  ANDN U11469 ( .B(y[748]), .A(n166), .Z(n11279) );
  XNOR U11470 ( .A(n11278), .B(n11279), .Z(n11281) );
  XOR U11471 ( .A(n11280), .B(n11281), .Z(n11232) );
  NAND U11472 ( .A(x[134]), .B(y[757]), .Z(n11218) );
  ANDN U11473 ( .B(y[738]), .A(n14372), .Z(n11217) );
  NAND U11474 ( .A(y[744]), .B(x[147]), .Z(n11216) );
  XOR U11475 ( .A(n11217), .B(n11216), .Z(n11219) );
  XNOR U11476 ( .A(n11218), .B(n11219), .Z(n11233) );
  XNOR U11477 ( .A(n11232), .B(n11233), .Z(n11235) );
  OR U11478 ( .A(n11095), .B(n11094), .Z(n11099) );
  NAND U11479 ( .A(n11097), .B(n11096), .Z(n11098) );
  AND U11480 ( .A(n11099), .B(n11098), .Z(n11260) );
  NANDN U11481 ( .A(n11101), .B(n11100), .Z(n11105) );
  NAND U11482 ( .A(n11103), .B(n11102), .Z(n11104) );
  NAND U11483 ( .A(n11105), .B(n11104), .Z(n11261) );
  XNOR U11484 ( .A(n11260), .B(n11261), .Z(n11262) );
  XNOR U11485 ( .A(n11263), .B(n11262), .Z(n11296) );
  XNOR U11486 ( .A(n11297), .B(n11296), .Z(n11298) );
  XOR U11487 ( .A(n11299), .B(n11298), .Z(n11185) );
  OR U11488 ( .A(n11107), .B(n11106), .Z(n11111) );
  NANDN U11489 ( .A(n11109), .B(n11108), .Z(n11110) );
  NAND U11490 ( .A(n11111), .B(n11110), .Z(n11186) );
  XOR U11491 ( .A(n11185), .B(n11186), .Z(n11187) );
  XOR U11492 ( .A(n11188), .B(n11187), .Z(n11321) );
  OR U11493 ( .A(n11113), .B(n11112), .Z(n11117) );
  NAND U11494 ( .A(n11115), .B(n11114), .Z(n11116) );
  AND U11495 ( .A(n11117), .B(n11116), .Z(n11312) );
  OR U11496 ( .A(n11119), .B(n11118), .Z(n11123) );
  OR U11497 ( .A(n11121), .B(n11120), .Z(n11122) );
  NAND U11498 ( .A(n11123), .B(n11122), .Z(n11309) );
  OR U11499 ( .A(n11125), .B(n11124), .Z(n11129) );
  OR U11500 ( .A(n11127), .B(n11126), .Z(n11128) );
  AND U11501 ( .A(n11129), .B(n11128), .Z(n11306) );
  NANDN U11502 ( .A(n11131), .B(n11130), .Z(n11135) );
  NANDN U11503 ( .A(n11133), .B(n11132), .Z(n11134) );
  NAND U11504 ( .A(n11135), .B(n11134), .Z(n11181) );
  NANDN U11505 ( .A(n11137), .B(n11136), .Z(n11141) );
  NAND U11506 ( .A(n11139), .B(n11138), .Z(n11140) );
  AND U11507 ( .A(n11141), .B(n11140), .Z(n11240) );
  ANDN U11508 ( .B(y[741]), .A(n173), .Z(n11292) );
  ANDN U11509 ( .B(y[740]), .A(n174), .Z(n11290) );
  ANDN U11510 ( .B(y[755]), .A(n159), .Z(n11291) );
  XNOR U11511 ( .A(n11290), .B(n11291), .Z(n11293) );
  XOR U11512 ( .A(n11292), .B(n11293), .Z(n11238) );
  AND U11513 ( .A(x[135]), .B(y[756]), .Z(n11224) );
  NANDN U11514 ( .A(n149), .B(x[152]), .Z(n11222) );
  XOR U11515 ( .A(n11223), .B(n11222), .Z(n11225) );
  XOR U11516 ( .A(n11224), .B(n11225), .Z(n11239) );
  XOR U11517 ( .A(n11238), .B(n11239), .Z(n11241) );
  XOR U11518 ( .A(n11240), .B(n11241), .Z(n11179) );
  OR U11519 ( .A(n11143), .B(n11142), .Z(n11147) );
  OR U11520 ( .A(n11145), .B(n11144), .Z(n11146) );
  NAND U11521 ( .A(n11147), .B(n11146), .Z(n11229) );
  NANDN U11522 ( .A(n11149), .B(n11148), .Z(n11153) );
  NAND U11523 ( .A(n11151), .B(n11150), .Z(n11152) );
  NAND U11524 ( .A(n11153), .B(n11152), .Z(n11228) );
  XOR U11525 ( .A(n11229), .B(n11228), .Z(n11230) );
  NAND U11526 ( .A(n11155), .B(n11154), .Z(n11159) );
  NANDN U11527 ( .A(n11157), .B(n11156), .Z(n11158) );
  NAND U11528 ( .A(n11159), .B(n11158), .Z(n11245) );
  NAND U11529 ( .A(x[145]), .B(y[746]), .Z(n11204) );
  ANDN U11530 ( .B(y[759]), .A(n155), .Z(n11203) );
  XNOR U11531 ( .A(n11204), .B(n11203), .Z(n11206) );
  ANDN U11532 ( .B(y[758]), .A(n156), .Z(n11205) );
  XOR U11533 ( .A(n11206), .B(n11205), .Z(n11242) );
  NAND U11534 ( .A(y[749]), .B(x[142]), .Z(n11268) );
  ANDN U11535 ( .B(o[122]), .A(n11160), .Z(n11267) );
  NAND U11536 ( .A(x[129]), .B(y[762]), .Z(n11266) );
  XOR U11537 ( .A(n11267), .B(n11266), .Z(n11269) );
  XNOR U11538 ( .A(n11268), .B(n11269), .Z(n11243) );
  XOR U11539 ( .A(n11245), .B(n11244), .Z(n11231) );
  XNOR U11540 ( .A(n11230), .B(n11231), .Z(n11180) );
  XNOR U11541 ( .A(n11306), .B(n11307), .Z(n11308) );
  XOR U11542 ( .A(n11309), .B(n11308), .Z(n11313) );
  XOR U11543 ( .A(n11312), .B(n11313), .Z(n11314) );
  XOR U11544 ( .A(n11315), .B(n11314), .Z(n11174) );
  XOR U11545 ( .A(n11173), .B(n11174), .Z(n11175) );
  OR U11546 ( .A(n11162), .B(n11161), .Z(n11166) );
  NANDN U11547 ( .A(n11164), .B(n11163), .Z(n11165) );
  AND U11548 ( .A(n11166), .B(n11165), .Z(n11176) );
  XOR U11549 ( .A(n11169), .B(n11170), .Z(N252) );
  NANDN U11550 ( .A(n11168), .B(n11167), .Z(n11172) );
  NANDN U11551 ( .A(n11170), .B(n11169), .Z(n11171) );
  NAND U11552 ( .A(n11172), .B(n11171), .Z(n11324) );
  OR U11553 ( .A(n11174), .B(n11173), .Z(n11178) );
  NANDN U11554 ( .A(n11176), .B(n11175), .Z(n11177) );
  AND U11555 ( .A(n11178), .B(n11177), .Z(n11325) );
  XNOR U11556 ( .A(n11324), .B(n11325), .Z(n11326) );
  NANDN U11557 ( .A(n11180), .B(n11179), .Z(n11184) );
  NAND U11558 ( .A(n11182), .B(n11181), .Z(n11183) );
  NAND U11559 ( .A(n11184), .B(n11183), .Z(n11489) );
  OR U11560 ( .A(n11186), .B(n11185), .Z(n11190) );
  NANDN U11561 ( .A(n11188), .B(n11187), .Z(n11189) );
  NAND U11562 ( .A(n11190), .B(n11189), .Z(n11488) );
  OR U11563 ( .A(n11192), .B(n11191), .Z(n11196) );
  NANDN U11564 ( .A(n11194), .B(n11193), .Z(n11195) );
  NAND U11565 ( .A(n11196), .B(n11195), .Z(n11487) );
  XNOR U11566 ( .A(n11488), .B(n11487), .Z(n11490) );
  XNOR U11567 ( .A(n11489), .B(n11490), .Z(n11484) );
  OR U11568 ( .A(n11198), .B(n11197), .Z(n11202) );
  OR U11569 ( .A(n11200), .B(n11199), .Z(n11201) );
  AND U11570 ( .A(n11202), .B(n11201), .Z(n11354) );
  NANDN U11571 ( .A(n11204), .B(n11203), .Z(n11208) );
  NAND U11572 ( .A(n11206), .B(n11205), .Z(n11207) );
  NAND U11573 ( .A(n11208), .B(n11207), .Z(n11355) );
  XOR U11574 ( .A(n11354), .B(n11355), .Z(n11357) );
  OR U11575 ( .A(n11210), .B(n11209), .Z(n11214) );
  OR U11576 ( .A(n11212), .B(n11211), .Z(n11213) );
  AND U11577 ( .A(n11214), .B(n11213), .Z(n11390) );
  ANDN U11578 ( .B(y[754]), .A(n161), .Z(n11410) );
  ANDN U11579 ( .B(y[755]), .A(n160), .Z(n11408) );
  ANDN U11580 ( .B(y[756]), .A(n159), .Z(n11409) );
  XNOR U11581 ( .A(n11408), .B(n11409), .Z(n11411) );
  XNOR U11582 ( .A(n11410), .B(n11411), .Z(n11391) );
  XOR U11583 ( .A(n11390), .B(n11391), .Z(n11392) );
  ANDN U11584 ( .B(y[764]), .A(n151), .Z(n11398) );
  AND U11585 ( .A(n11215), .B(o[123]), .Z(n11396) );
  ANDN U11586 ( .B(y[736]), .A(n14373), .Z(n11397) );
  XNOR U11587 ( .A(n11396), .B(n11397), .Z(n11399) );
  XNOR U11588 ( .A(n11398), .B(n11399), .Z(n11393) );
  XNOR U11589 ( .A(n11357), .B(n11356), .Z(n11339) );
  ANDN U11590 ( .B(y[759]), .A(n156), .Z(n11435) );
  ANDN U11591 ( .B(y[744]), .A(n171), .Z(n11433) );
  ANDN U11592 ( .B(y[743]), .A(n172), .Z(n11434) );
  XNOR U11593 ( .A(n11433), .B(n11434), .Z(n11436) );
  XOR U11594 ( .A(n11435), .B(n11436), .Z(n11360) );
  ANDN U11595 ( .B(y[741]), .A(n174), .Z(n11449) );
  NAND U11596 ( .A(x[131]), .B(y[761]), .Z(n11448) );
  XOR U11597 ( .A(n11449), .B(n11448), .Z(n11451) );
  XOR U11598 ( .A(n11450), .B(n11451), .Z(n11361) );
  XNOR U11599 ( .A(n11360), .B(n11361), .Z(n11363) );
  NANDN U11600 ( .A(n11217), .B(n11216), .Z(n11221) );
  NANDN U11601 ( .A(n11219), .B(n11218), .Z(n11220) );
  NAND U11602 ( .A(n11221), .B(n11220), .Z(n11362) );
  XOR U11603 ( .A(n11363), .B(n11362), .Z(n11337) );
  ANDN U11604 ( .B(y[763]), .A(n152), .Z(n11415) );
  ANDN U11605 ( .B(y[739]), .A(n14372), .Z(n11416) );
  XNOR U11606 ( .A(n11415), .B(n11416), .Z(n11418) );
  XOR U11607 ( .A(n11417), .B(n11418), .Z(n11368) );
  ANDN U11608 ( .B(y[748]), .A(n167), .Z(n11423) );
  ANDN U11609 ( .B(y[762]), .A(n153), .Z(n11421) );
  ANDN U11610 ( .B(y[740]), .A(n175), .Z(n11422) );
  XNOR U11611 ( .A(n11421), .B(n11422), .Z(n11424) );
  XOR U11612 ( .A(n11423), .B(n11424), .Z(n11366) );
  NANDN U11613 ( .A(n11223), .B(n11222), .Z(n11227) );
  OR U11614 ( .A(n11225), .B(n11224), .Z(n11226) );
  NAND U11615 ( .A(n11227), .B(n11226), .Z(n11367) );
  XNOR U11616 ( .A(n11366), .B(n11367), .Z(n11369) );
  XNOR U11617 ( .A(n11368), .B(n11369), .Z(n11336) );
  XOR U11618 ( .A(n11337), .B(n11336), .Z(n11338) );
  XNOR U11619 ( .A(n11339), .B(n11338), .Z(n11476) );
  OR U11620 ( .A(n11233), .B(n11232), .Z(n11237) );
  NANDN U11621 ( .A(n11235), .B(n11234), .Z(n11236) );
  NAND U11622 ( .A(n11237), .B(n11236), .Z(n11343) );
  XOR U11623 ( .A(n11343), .B(n11342), .Z(n11344) );
  XOR U11624 ( .A(n11476), .B(n11475), .Z(n11478) );
  NANDN U11625 ( .A(n11243), .B(n11242), .Z(n11247) );
  NANDN U11626 ( .A(n11245), .B(n11244), .Z(n11246) );
  AND U11627 ( .A(n11247), .B(n11246), .Z(n11372) );
  OR U11628 ( .A(n11249), .B(n11248), .Z(n11253) );
  NANDN U11629 ( .A(n11251), .B(n11250), .Z(n11252) );
  NAND U11630 ( .A(n11253), .B(n11252), .Z(n11373) );
  XOR U11631 ( .A(n11372), .B(n11373), .Z(n11374) );
  OR U11632 ( .A(n11255), .B(n11254), .Z(n11259) );
  NAND U11633 ( .A(n11257), .B(n11256), .Z(n11258) );
  NAND U11634 ( .A(n11259), .B(n11258), .Z(n11375) );
  OR U11635 ( .A(n11261), .B(n11260), .Z(n11265) );
  OR U11636 ( .A(n11263), .B(n11262), .Z(n11264) );
  AND U11637 ( .A(n11265), .B(n11264), .Z(n11379) );
  NANDN U11638 ( .A(n11267), .B(n11266), .Z(n11271) );
  NANDN U11639 ( .A(n11269), .B(n11268), .Z(n11270) );
  AND U11640 ( .A(n11271), .B(n11270), .Z(n11387) );
  OR U11641 ( .A(n11273), .B(n11272), .Z(n11277) );
  OR U11642 ( .A(n11275), .B(n11274), .Z(n11276) );
  AND U11643 ( .A(n11277), .B(n11276), .Z(n11384) );
  OR U11644 ( .A(n11279), .B(n11278), .Z(n11283) );
  OR U11645 ( .A(n11281), .B(n11280), .Z(n11282) );
  AND U11646 ( .A(n11283), .B(n11282), .Z(n11385) );
  XOR U11647 ( .A(n11384), .B(n11385), .Z(n11386) );
  ANDN U11648 ( .B(y[757]), .A(n158), .Z(n11429) );
  ANDN U11649 ( .B(y[753]), .A(n162), .Z(n11427) );
  ANDN U11650 ( .B(y[752]), .A(n163), .Z(n11428) );
  XNOR U11651 ( .A(n11427), .B(n11428), .Z(n11430) );
  XOR U11652 ( .A(n11429), .B(n11430), .Z(n11459) );
  NANDN U11653 ( .A(n11285), .B(n11284), .Z(n11289) );
  NAND U11654 ( .A(n11287), .B(n11286), .Z(n11288) );
  NAND U11655 ( .A(n11289), .B(n11288), .Z(n11460) );
  XNOR U11656 ( .A(n11459), .B(n11460), .Z(n11462) );
  NAND U11657 ( .A(x[143]), .B(y[749]), .Z(n11453) );
  AND U11658 ( .A(y[738]), .B(x[154]), .Z(n11452) );
  XNOR U11659 ( .A(n11453), .B(n11452), .Z(n11454) );
  AND U11660 ( .A(y[737]), .B(x[155]), .Z(n11583) );
  XNOR U11661 ( .A(o[124]), .B(n11583), .Z(n11455) );
  XOR U11662 ( .A(n11462), .B(n11461), .Z(n11348) );
  OR U11663 ( .A(n11291), .B(n11290), .Z(n11295) );
  OR U11664 ( .A(n11293), .B(n11292), .Z(n11294) );
  AND U11665 ( .A(n11295), .B(n11294), .Z(n11465) );
  ANDN U11666 ( .B(y[758]), .A(n157), .Z(n11444) );
  ANDN U11667 ( .B(y[745]), .A(n170), .Z(n11443) );
  XNOR U11668 ( .A(n11442), .B(n11443), .Z(n11445) );
  XNOR U11669 ( .A(n11444), .B(n11445), .Z(n11466) );
  XOR U11670 ( .A(n11465), .B(n11466), .Z(n11468) );
  NAND U11671 ( .A(x[145]), .B(y[747]), .Z(n11404) );
  ANDN U11672 ( .B(y[760]), .A(n155), .Z(n11403) );
  NAND U11673 ( .A(y[742]), .B(x[150]), .Z(n11402) );
  XOR U11674 ( .A(n11403), .B(n11402), .Z(n11405) );
  XNOR U11675 ( .A(n11404), .B(n11405), .Z(n11467) );
  XNOR U11676 ( .A(n11468), .B(n11467), .Z(n11349) );
  XNOR U11677 ( .A(n11348), .B(n11349), .Z(n11350) );
  XOR U11678 ( .A(n11351), .B(n11350), .Z(n11378) );
  XOR U11679 ( .A(n11379), .B(n11378), .Z(n11381) );
  XOR U11680 ( .A(n11380), .B(n11381), .Z(n11477) );
  XNOR U11681 ( .A(n11478), .B(n11477), .Z(n11474) );
  OR U11682 ( .A(n11297), .B(n11296), .Z(n11301) );
  OR U11683 ( .A(n11299), .B(n11298), .Z(n11300) );
  AND U11684 ( .A(n11301), .B(n11300), .Z(n11471) );
  XOR U11685 ( .A(n11471), .B(n11472), .Z(n11473) );
  XNOR U11686 ( .A(n11474), .B(n11473), .Z(n11481) );
  OR U11687 ( .A(n11307), .B(n11306), .Z(n11311) );
  OR U11688 ( .A(n11309), .B(n11308), .Z(n11310) );
  AND U11689 ( .A(n11311), .B(n11310), .Z(n11482) );
  XOR U11690 ( .A(n11481), .B(n11482), .Z(n11483) );
  XNOR U11691 ( .A(n11484), .B(n11483), .Z(n11330) );
  OR U11692 ( .A(n11313), .B(n11312), .Z(n11317) );
  NANDN U11693 ( .A(n11315), .B(n11314), .Z(n11316) );
  AND U11694 ( .A(n11317), .B(n11316), .Z(n11331) );
  XNOR U11695 ( .A(n11330), .B(n11331), .Z(n11333) );
  OR U11696 ( .A(n11319), .B(n11318), .Z(n11323) );
  NANDN U11697 ( .A(n11321), .B(n11320), .Z(n11322) );
  NAND U11698 ( .A(n11323), .B(n11322), .Z(n11332) );
  XOR U11699 ( .A(n11333), .B(n11332), .Z(n11327) );
  XNOR U11700 ( .A(n11326), .B(n11327), .Z(N253) );
  NANDN U11701 ( .A(n11325), .B(n11324), .Z(n11329) );
  NAND U11702 ( .A(n11327), .B(n11326), .Z(n11328) );
  NAND U11703 ( .A(n11329), .B(n11328), .Z(n11493) );
  OR U11704 ( .A(n11331), .B(n11330), .Z(n11335) );
  OR U11705 ( .A(n11333), .B(n11332), .Z(n11334) );
  AND U11706 ( .A(n11335), .B(n11334), .Z(n11494) );
  XNOR U11707 ( .A(n11493), .B(n11494), .Z(n11495) );
  NANDN U11708 ( .A(n11337), .B(n11336), .Z(n11341) );
  OR U11709 ( .A(n11339), .B(n11338), .Z(n11340) );
  AND U11710 ( .A(n11341), .B(n11340), .Z(n11651) );
  OR U11711 ( .A(n11343), .B(n11342), .Z(n11347) );
  NANDN U11712 ( .A(n11345), .B(n11344), .Z(n11346) );
  AND U11713 ( .A(n11347), .B(n11346), .Z(n11649) );
  OR U11714 ( .A(n11349), .B(n11348), .Z(n11353) );
  OR U11715 ( .A(n11351), .B(n11350), .Z(n11352) );
  AND U11716 ( .A(n11353), .B(n11352), .Z(n11661) );
  OR U11717 ( .A(n11355), .B(n11354), .Z(n11359) );
  NAND U11718 ( .A(n11357), .B(n11356), .Z(n11358) );
  NAND U11719 ( .A(n11359), .B(n11358), .Z(n11591) );
  OR U11720 ( .A(n11361), .B(n11360), .Z(n11365) );
  OR U11721 ( .A(n11363), .B(n11362), .Z(n11364) );
  AND U11722 ( .A(n11365), .B(n11364), .Z(n11588) );
  OR U11723 ( .A(n11367), .B(n11366), .Z(n11371) );
  OR U11724 ( .A(n11369), .B(n11368), .Z(n11370) );
  AND U11725 ( .A(n11371), .B(n11370), .Z(n11589) );
  XOR U11726 ( .A(n11588), .B(n11589), .Z(n11590) );
  XNOR U11727 ( .A(n11591), .B(n11590), .Z(n11662) );
  XOR U11728 ( .A(n11661), .B(n11662), .Z(n11663) );
  OR U11729 ( .A(n11373), .B(n11372), .Z(n11377) );
  NANDN U11730 ( .A(n11375), .B(n11374), .Z(n11376) );
  NAND U11731 ( .A(n11377), .B(n11376), .Z(n11664) );
  XNOR U11732 ( .A(n11649), .B(n11650), .Z(n11652) );
  XOR U11733 ( .A(n11651), .B(n11652), .Z(n11655) );
  NANDN U11734 ( .A(n11379), .B(n11378), .Z(n11383) );
  NANDN U11735 ( .A(n11381), .B(n11380), .Z(n11382) );
  NAND U11736 ( .A(n11383), .B(n11382), .Z(n11656) );
  XNOR U11737 ( .A(n11655), .B(n11656), .Z(n11658) );
  OR U11738 ( .A(n11385), .B(n11384), .Z(n11389) );
  NANDN U11739 ( .A(n11387), .B(n11386), .Z(n11388) );
  AND U11740 ( .A(n11389), .B(n11388), .Z(n11645) );
  OR U11741 ( .A(n11391), .B(n11390), .Z(n11395) );
  NANDN U11742 ( .A(n11393), .B(n11392), .Z(n11394) );
  AND U11743 ( .A(n11395), .B(n11394), .Z(n11643) );
  OR U11744 ( .A(n11397), .B(n11396), .Z(n11401) );
  OR U11745 ( .A(n11399), .B(n11398), .Z(n11400) );
  AND U11746 ( .A(n11401), .B(n11400), .Z(n11640) );
  NANDN U11747 ( .A(n11403), .B(n11402), .Z(n11407) );
  NANDN U11748 ( .A(n11405), .B(n11404), .Z(n11406) );
  AND U11749 ( .A(n11407), .B(n11406), .Z(n11637) );
  OR U11750 ( .A(n11409), .B(n11408), .Z(n11413) );
  OR U11751 ( .A(n11411), .B(n11410), .Z(n11412) );
  AND U11752 ( .A(n11413), .B(n11412), .Z(n11606) );
  ANDN U11753 ( .B(y[750]), .A(n166), .Z(n11540) );
  NOR U11754 ( .A(n172), .B(n11414), .Z(n11766) );
  ANDN U11755 ( .B(y[745]), .A(n171), .Z(n11539) );
  XNOR U11756 ( .A(n11766), .B(n11539), .Z(n11541) );
  XNOR U11757 ( .A(n11540), .B(n11541), .Z(n11607) );
  XOR U11758 ( .A(n11606), .B(n11607), .Z(n11608) );
  AND U11759 ( .A(x[140]), .B(y[753]), .Z(n11885) );
  ANDN U11760 ( .B(y[743]), .A(n173), .Z(n11535) );
  NAND U11761 ( .A(x[129]), .B(y[764]), .Z(n11534) );
  XOR U11762 ( .A(n11535), .B(n11534), .Z(n11536) );
  XNOR U11763 ( .A(n11885), .B(n11536), .Z(n11609) );
  XOR U11764 ( .A(n11608), .B(n11609), .Z(n11638) );
  XOR U11765 ( .A(n11637), .B(n11638), .Z(n11639) );
  XNOR U11766 ( .A(n11643), .B(n11644), .Z(n11646) );
  XNOR U11767 ( .A(n11645), .B(n11646), .Z(n11602) );
  OR U11768 ( .A(n11416), .B(n11415), .Z(n11420) );
  OR U11769 ( .A(n11418), .B(n11417), .Z(n11419) );
  AND U11770 ( .A(n11420), .B(n11419), .Z(n11615) );
  OR U11771 ( .A(n11422), .B(n11421), .Z(n11426) );
  OR U11772 ( .A(n11424), .B(n11423), .Z(n11425) );
  AND U11773 ( .A(n11426), .B(n11425), .Z(n11612) );
  ANDN U11774 ( .B(y[752]), .A(n164), .Z(n11522) );
  ANDN U11775 ( .B(y[742]), .A(n174), .Z(n11521) );
  AND U11776 ( .A(y[741]), .B(x[152]), .Z(n11877) );
  XNOR U11777 ( .A(n11521), .B(n11877), .Z(n11523) );
  XNOR U11778 ( .A(n11522), .B(n11523), .Z(n11566) );
  OR U11779 ( .A(n11428), .B(n11427), .Z(n11432) );
  OR U11780 ( .A(n11430), .B(n11429), .Z(n11431) );
  AND U11781 ( .A(n11432), .B(n11431), .Z(n11564) );
  NAND U11782 ( .A(x[131]), .B(y[762]), .Z(n11517) );
  ANDN U11783 ( .B(y[754]), .A(n162), .Z(n11516) );
  NAND U11784 ( .A(x[145]), .B(y[748]), .Z(n11515) );
  XOR U11785 ( .A(n11516), .B(n11515), .Z(n11518) );
  XNOR U11786 ( .A(n11517), .B(n11518), .Z(n11563) );
  XOR U11787 ( .A(n11564), .B(n11563), .Z(n11565) );
  XNOR U11788 ( .A(n11566), .B(n11565), .Z(n11613) );
  XOR U11789 ( .A(n11612), .B(n11613), .Z(n11614) );
  OR U11790 ( .A(n11434), .B(n11433), .Z(n11438) );
  OR U11791 ( .A(n11436), .B(n11435), .Z(n11437) );
  AND U11792 ( .A(n11438), .B(n11437), .Z(n11509) );
  NAND U11793 ( .A(y[737]), .B(o[124]), .Z(n11439) );
  XNOR U11794 ( .A(y[738]), .B(n11439), .Z(n11440) );
  NAND U11795 ( .A(x[155]), .B(n11440), .Z(n11582) );
  ANDN U11796 ( .B(y[749]), .A(n167), .Z(n11581) );
  XNOR U11797 ( .A(n11582), .B(n11581), .Z(n11510) );
  XOR U11798 ( .A(n11509), .B(n11510), .Z(n11512) );
  ANDN U11799 ( .B(y[747]), .A(n169), .Z(n11575) );
  ANDN U11800 ( .B(y[746]), .A(n170), .Z(n11576) );
  XNOR U11801 ( .A(n11575), .B(n11576), .Z(n11578) );
  ANDN U11802 ( .B(y[763]), .A(n153), .Z(n11577) );
  XOR U11803 ( .A(n11578), .B(n11577), .Z(n11511) );
  XNOR U11804 ( .A(n11512), .B(n11511), .Z(n11595) );
  ANDN U11805 ( .B(y[765]), .A(n151), .Z(n11633) );
  ANDN U11806 ( .B(y[737]), .A(n14373), .Z(n11544) );
  XOR U11807 ( .A(o[125]), .B(n11544), .Z(n11631) );
  ANDN U11808 ( .B(y[736]), .A(n11441), .Z(n11632) );
  XNOR U11809 ( .A(n11631), .B(n11632), .Z(n11634) );
  XOR U11810 ( .A(n11633), .B(n11634), .Z(n11618) );
  NAND U11811 ( .A(y[751]), .B(x[142]), .Z(n11547) );
  ANDN U11812 ( .B(y[740]), .A(n14372), .Z(n11546) );
  NAND U11813 ( .A(y[739]), .B(x[154]), .Z(n11545) );
  XOR U11814 ( .A(n11546), .B(n11545), .Z(n11548) );
  XNOR U11815 ( .A(n11547), .B(n11548), .Z(n11619) );
  XNOR U11816 ( .A(n11618), .B(n11619), .Z(n11621) );
  OR U11817 ( .A(n11443), .B(n11442), .Z(n11447) );
  OR U11818 ( .A(n11445), .B(n11444), .Z(n11446) );
  NAND U11819 ( .A(n11447), .B(n11446), .Z(n11620) );
  XOR U11820 ( .A(n11621), .B(n11620), .Z(n11594) );
  XNOR U11821 ( .A(n11595), .B(n11594), .Z(n11596) );
  XOR U11822 ( .A(n11597), .B(n11596), .Z(n11553) );
  NANDN U11823 ( .A(n11453), .B(n11452), .Z(n11457) );
  NANDN U11824 ( .A(n11455), .B(n11454), .Z(n11456) );
  NAND U11825 ( .A(n11457), .B(n11456), .Z(n11558) );
  XOR U11826 ( .A(n11557), .B(n11558), .Z(n11559) );
  NOR U11827 ( .A(n160), .B(n11458), .Z(n11747) );
  ANDN U11828 ( .B(y[760]), .A(n156), .Z(n11569) );
  ANDN U11829 ( .B(y[755]), .A(n161), .Z(n11570) );
  XNOR U11830 ( .A(n11569), .B(n11570), .Z(n11572) );
  ANDN U11831 ( .B(y[761]), .A(n155), .Z(n11571) );
  XNOR U11832 ( .A(n11572), .B(n11571), .Z(n11624) );
  XNOR U11833 ( .A(n11747), .B(n11624), .Z(n11626) );
  ANDN U11834 ( .B(y[759]), .A(n157), .Z(n11528) );
  ANDN U11835 ( .B(y[757]), .A(n159), .Z(n11526) );
  ANDN U11836 ( .B(y[758]), .A(n158), .Z(n11527) );
  XNOR U11837 ( .A(n11526), .B(n11527), .Z(n11529) );
  XNOR U11838 ( .A(n11528), .B(n11529), .Z(n11625) );
  XNOR U11839 ( .A(n11626), .B(n11625), .Z(n11560) );
  OR U11840 ( .A(n11460), .B(n11459), .Z(n11464) );
  OR U11841 ( .A(n11462), .B(n11461), .Z(n11463) );
  AND U11842 ( .A(n11464), .B(n11463), .Z(n11552) );
  XNOR U11843 ( .A(n11551), .B(n11552), .Z(n11554) );
  XNOR U11844 ( .A(n11553), .B(n11554), .Z(n11601) );
  OR U11845 ( .A(n11466), .B(n11465), .Z(n11470) );
  NAND U11846 ( .A(n11468), .B(n11467), .Z(n11469) );
  NAND U11847 ( .A(n11470), .B(n11469), .Z(n11600) );
  XNOR U11848 ( .A(n11601), .B(n11600), .Z(n11603) );
  XOR U11849 ( .A(n11602), .B(n11603), .Z(n11657) );
  XOR U11850 ( .A(n11658), .B(n11657), .Z(n11508) );
  NANDN U11851 ( .A(n11476), .B(n11475), .Z(n11480) );
  OR U11852 ( .A(n11478), .B(n11477), .Z(n11479) );
  NAND U11853 ( .A(n11480), .B(n11479), .Z(n11506) );
  XOR U11854 ( .A(n11505), .B(n11506), .Z(n11507) );
  XOR U11855 ( .A(n11508), .B(n11507), .Z(n11501) );
  OR U11856 ( .A(n11482), .B(n11481), .Z(n11486) );
  NANDN U11857 ( .A(n11484), .B(n11483), .Z(n11485) );
  AND U11858 ( .A(n11486), .B(n11485), .Z(n11499) );
  OR U11859 ( .A(n11488), .B(n11487), .Z(n11492) );
  NANDN U11860 ( .A(n11490), .B(n11489), .Z(n11491) );
  NAND U11861 ( .A(n11492), .B(n11491), .Z(n11500) );
  XNOR U11862 ( .A(n11499), .B(n11500), .Z(n11502) );
  XOR U11863 ( .A(n11501), .B(n11502), .Z(n11496) );
  XOR U11864 ( .A(n11495), .B(n11496), .Z(N254) );
  NANDN U11865 ( .A(n11494), .B(n11493), .Z(n11498) );
  NANDN U11866 ( .A(n11496), .B(n11495), .Z(n11497) );
  AND U11867 ( .A(n11498), .B(n11497), .Z(n11669) );
  OR U11868 ( .A(n11500), .B(n11499), .Z(n11504) );
  OR U11869 ( .A(n11502), .B(n11501), .Z(n11503) );
  NAND U11870 ( .A(n11504), .B(n11503), .Z(n11670) );
  XNOR U11871 ( .A(n11669), .B(n11670), .Z(n11668) );
  OR U11872 ( .A(n11510), .B(n11509), .Z(n11514) );
  NAND U11873 ( .A(n11512), .B(n11511), .Z(n11513) );
  NAND U11874 ( .A(n11514), .B(n11513), .Z(n11922) );
  NANDN U11875 ( .A(n11516), .B(n11515), .Z(n11520) );
  NANDN U11876 ( .A(n11518), .B(n11517), .Z(n11519) );
  NAND U11877 ( .A(n11520), .B(n11519), .Z(n11720) );
  NAND U11878 ( .A(x[148]), .B(y[746]), .Z(n11772) );
  AND U11879 ( .A(y[752]), .B(x[142]), .Z(n11771) );
  XOR U11880 ( .A(n11772), .B(n11771), .Z(n11770) );
  AND U11881 ( .A(y[758]), .B(x[136]), .Z(n11769) );
  XOR U11882 ( .A(n11770), .B(n11769), .Z(n11722) );
  NAND U11883 ( .A(y[736]), .B(x[158]), .Z(n11753) );
  NAND U11884 ( .A(x[157]), .B(y[737]), .Z(n11801) );
  XNOR U11885 ( .A(o[126]), .B(n11801), .Z(n11752) );
  XOR U11886 ( .A(n11753), .B(n11752), .Z(n11751) );
  AND U11887 ( .A(y[766]), .B(x[128]), .Z(n11750) );
  XNOR U11888 ( .A(n11751), .B(n11750), .Z(n11721) );
  XOR U11889 ( .A(n11720), .B(n11719), .Z(n11695) );
  OR U11890 ( .A(n11521), .B(n11877), .Z(n11525) );
  OR U11891 ( .A(n11523), .B(n11522), .Z(n11524) );
  AND U11892 ( .A(n11525), .B(n11524), .Z(n11696) );
  XNOR U11893 ( .A(n11695), .B(n11696), .Z(n11694) );
  OR U11894 ( .A(n11527), .B(n11526), .Z(n11531) );
  OR U11895 ( .A(n11529), .B(n11528), .Z(n11530) );
  AND U11896 ( .A(n11531), .B(n11530), .Z(n11733) );
  NAND U11897 ( .A(x[145]), .B(y[749]), .Z(n11846) );
  NAND U11898 ( .A(x[130]), .B(y[764]), .Z(n11848) );
  NAND U11899 ( .A(x[154]), .B(y[740]), .Z(n11847) );
  XNOR U11900 ( .A(n11848), .B(n11847), .Z(n11845) );
  XNOR U11901 ( .A(n11846), .B(n11845), .Z(n11732) );
  NAND U11902 ( .A(x[135]), .B(y[759]), .Z(n11765) );
  AND U11903 ( .A(y[744]), .B(x[150]), .Z(n11533) );
  AND U11904 ( .A(y[745]), .B(x[149]), .Z(n11532) );
  XNOR U11905 ( .A(n11533), .B(n11532), .Z(n11764) );
  XOR U11906 ( .A(n11765), .B(n11764), .Z(n11731) );
  XNOR U11907 ( .A(n11732), .B(n11731), .Z(n11734) );
  XOR U11908 ( .A(n11733), .B(n11734), .Z(n11693) );
  XNOR U11909 ( .A(n11694), .B(n11693), .Z(n11921) );
  XOR U11910 ( .A(n11922), .B(n11921), .Z(n11920) );
  NANDN U11911 ( .A(n11535), .B(n11534), .Z(n11538) );
  OR U11912 ( .A(n11536), .B(n11885), .Z(n11537) );
  AND U11913 ( .A(n11538), .B(n11537), .Z(n11714) );
  NAND U11914 ( .A(x[151]), .B(y[743]), .Z(n11876) );
  AND U11915 ( .A(y[741]), .B(x[153]), .Z(n11543) );
  AND U11916 ( .A(x[152]), .B(y[742]), .Z(n11542) );
  XNOR U11917 ( .A(n11543), .B(n11542), .Z(n11875) );
  XOR U11918 ( .A(n11876), .B(n11875), .Z(n11797) );
  NAND U11919 ( .A(n11544), .B(o[125]), .Z(n11840) );
  NAND U11920 ( .A(x[156]), .B(y[738]), .Z(n11842) );
  AND U11921 ( .A(y[750]), .B(x[144]), .Z(n11841) );
  XNOR U11922 ( .A(n11842), .B(n11841), .Z(n11839) );
  XNOR U11923 ( .A(n11840), .B(n11839), .Z(n11798) );
  XNOR U11924 ( .A(n11797), .B(n11798), .Z(n11796) );
  XOR U11925 ( .A(n11795), .B(n11796), .Z(n11713) );
  NANDN U11926 ( .A(n11546), .B(n11545), .Z(n11550) );
  NANDN U11927 ( .A(n11548), .B(n11547), .Z(n11549) );
  AND U11928 ( .A(n11550), .B(n11549), .Z(n11711) );
  XOR U11929 ( .A(n11712), .B(n11711), .Z(n11919) );
  XNOR U11930 ( .A(n11920), .B(n11919), .Z(n11676) );
  OR U11931 ( .A(n11552), .B(n11551), .Z(n11556) );
  OR U11932 ( .A(n11554), .B(n11553), .Z(n11555) );
  AND U11933 ( .A(n11556), .B(n11555), .Z(n11675) );
  XOR U11934 ( .A(n11676), .B(n11675), .Z(n11673) );
  OR U11935 ( .A(n11558), .B(n11557), .Z(n11562) );
  NANDN U11936 ( .A(n11560), .B(n11559), .Z(n11561) );
  AND U11937 ( .A(n11562), .B(n11561), .Z(n11685) );
  NANDN U11938 ( .A(n11564), .B(n11563), .Z(n11568) );
  OR U11939 ( .A(n11566), .B(n11565), .Z(n11567) );
  AND U11940 ( .A(n11568), .B(n11567), .Z(n11687) );
  OR U11941 ( .A(n11570), .B(n11569), .Z(n11574) );
  OR U11942 ( .A(n11572), .B(n11571), .Z(n11573) );
  AND U11943 ( .A(n11574), .B(n11573), .Z(n11707) );
  NAND U11944 ( .A(x[134]), .B(y[760]), .Z(n11870) );
  NAND U11945 ( .A(x[133]), .B(y[761]), .Z(n11872) );
  NAND U11946 ( .A(x[147]), .B(y[747]), .Z(n11871) );
  XNOR U11947 ( .A(n11872), .B(n11871), .Z(n11869) );
  XNOR U11948 ( .A(n11870), .B(n11869), .Z(n11725) );
  OR U11949 ( .A(n11576), .B(n11575), .Z(n11580) );
  OR U11950 ( .A(n11578), .B(n11577), .Z(n11579) );
  AND U11951 ( .A(n11580), .B(n11579), .Z(n11728) );
  NAND U11952 ( .A(x[132]), .B(y[762]), .Z(n11890) );
  NAND U11953 ( .A(x[131]), .B(y[763]), .Z(n11892) );
  AND U11954 ( .A(y[748]), .B(x[146]), .Z(n11891) );
  XNOR U11955 ( .A(n11892), .B(n11891), .Z(n11889) );
  XNOR U11956 ( .A(n11890), .B(n11889), .Z(n11727) );
  XOR U11957 ( .A(n11728), .B(n11727), .Z(n11726) );
  XNOR U11958 ( .A(n11725), .B(n11726), .Z(n11708) );
  XOR U11959 ( .A(n11707), .B(n11708), .Z(n11705) );
  OR U11960 ( .A(n11582), .B(n11581), .Z(n11587) );
  NAND U11961 ( .A(n11583), .B(o[124]), .Z(n11585) );
  NAND U11962 ( .A(x[155]), .B(y[738]), .Z(n11584) );
  AND U11963 ( .A(n11585), .B(n11584), .Z(n11586) );
  ANDN U11964 ( .B(n11587), .A(n11586), .Z(n11706) );
  XNOR U11965 ( .A(n11687), .B(n11688), .Z(n11686) );
  XOR U11966 ( .A(n11685), .B(n11686), .Z(n11674) );
  OR U11967 ( .A(n11589), .B(n11588), .Z(n11593) );
  NANDN U11968 ( .A(n11591), .B(n11590), .Z(n11592) );
  NAND U11969 ( .A(n11593), .B(n11592), .Z(n11944) );
  XNOR U11970 ( .A(n11943), .B(n11944), .Z(n11942) );
  OR U11971 ( .A(n11595), .B(n11594), .Z(n11599) );
  OR U11972 ( .A(n11597), .B(n11596), .Z(n11598) );
  AND U11973 ( .A(n11599), .B(n11598), .Z(n11941) );
  XOR U11974 ( .A(n11942), .B(n11941), .Z(n11935) );
  OR U11975 ( .A(n11601), .B(n11600), .Z(n11605) );
  NANDN U11976 ( .A(n11603), .B(n11602), .Z(n11604) );
  AND U11977 ( .A(n11605), .B(n11604), .Z(n11938) );
  OR U11978 ( .A(n11607), .B(n11606), .Z(n11611) );
  NANDN U11979 ( .A(n11609), .B(n11608), .Z(n11610) );
  AND U11980 ( .A(n11611), .B(n11610), .Z(n11681) );
  OR U11981 ( .A(n11613), .B(n11612), .Z(n11617) );
  NANDN U11982 ( .A(n11615), .B(n11614), .Z(n11616) );
  AND U11983 ( .A(n11617), .B(n11616), .Z(n11682) );
  XOR U11984 ( .A(n11681), .B(n11682), .Z(n11679) );
  OR U11985 ( .A(n11619), .B(n11618), .Z(n11623) );
  OR U11986 ( .A(n11621), .B(n11620), .Z(n11622) );
  NAND U11987 ( .A(n11623), .B(n11622), .Z(n11680) );
  XNOR U11988 ( .A(n11679), .B(n11680), .Z(n11916) );
  NAND U11989 ( .A(x[155]), .B(y[739]), .Z(n11761) );
  AND U11990 ( .A(y[765]), .B(x[129]), .Z(n11760) );
  XNOR U11991 ( .A(n11761), .B(n11760), .Z(n11758) );
  AND U11992 ( .A(x[140]), .B(y[754]), .Z(n11628) );
  NAND U11993 ( .A(x[141]), .B(y[753]), .Z(n11627) );
  XOR U11994 ( .A(n11628), .B(n11627), .Z(n11884) );
  XNOR U11995 ( .A(n11884), .B(n11883), .Z(n11746) );
  AND U11996 ( .A(x[138]), .B(y[756]), .Z(n11630) );
  AND U11997 ( .A(y[757]), .B(x[137]), .Z(n11629) );
  XNOR U11998 ( .A(n11630), .B(n11629), .Z(n11745) );
  XOR U11999 ( .A(n11746), .B(n11745), .Z(n11741) );
  OR U12000 ( .A(n11632), .B(n11631), .Z(n11636) );
  OR U12001 ( .A(n11634), .B(n11633), .Z(n11635) );
  AND U12002 ( .A(n11636), .B(n11635), .Z(n11742) );
  XNOR U12003 ( .A(n11741), .B(n11742), .Z(n11740) );
  XOR U12004 ( .A(n11739), .B(n11740), .Z(n11701) );
  XNOR U12005 ( .A(n11702), .B(n11701), .Z(n11700) );
  OR U12006 ( .A(n11638), .B(n11637), .Z(n11642) );
  NANDN U12007 ( .A(n11640), .B(n11639), .Z(n11641) );
  NAND U12008 ( .A(n11642), .B(n11641), .Z(n11699) );
  XOR U12009 ( .A(n11700), .B(n11699), .Z(n11915) );
  XOR U12010 ( .A(n11916), .B(n11915), .Z(n11914) );
  OR U12011 ( .A(n11644), .B(n11643), .Z(n11648) );
  OR U12012 ( .A(n11646), .B(n11645), .Z(n11647) );
  NAND U12013 ( .A(n11648), .B(n11647), .Z(n11913) );
  XOR U12014 ( .A(n11914), .B(n11913), .Z(n11937) );
  XOR U12015 ( .A(n11935), .B(n11936), .Z(n11955) );
  OR U12016 ( .A(n11650), .B(n11649), .Z(n11654) );
  OR U12017 ( .A(n11652), .B(n11651), .Z(n11653) );
  AND U12018 ( .A(n11654), .B(n11653), .Z(n11961) );
  OR U12019 ( .A(n11656), .B(n11655), .Z(n11660) );
  OR U12020 ( .A(n11658), .B(n11657), .Z(n11659) );
  NAND U12021 ( .A(n11660), .B(n11659), .Z(n11962) );
  XOR U12022 ( .A(n11961), .B(n11962), .Z(n11959) );
  OR U12023 ( .A(n11662), .B(n11661), .Z(n11666) );
  NANDN U12024 ( .A(n11664), .B(n11663), .Z(n11665) );
  AND U12025 ( .A(n11666), .B(n11665), .Z(n11960) );
  XNOR U12026 ( .A(n11955), .B(n11956), .Z(n11954) );
  XOR U12027 ( .A(n11953), .B(n11954), .Z(n11667) );
  XOR U12028 ( .A(n11668), .B(n11667), .Z(N255) );
  NANDN U12029 ( .A(n11668), .B(n11667), .Z(n11672) );
  OR U12030 ( .A(n11670), .B(n11669), .Z(n11671) );
  AND U12031 ( .A(n11672), .B(n11671), .Z(n11952) );
  NANDN U12032 ( .A(n11674), .B(n11673), .Z(n11678) );
  OR U12033 ( .A(n11676), .B(n11675), .Z(n11677) );
  AND U12034 ( .A(n11678), .B(n11677), .Z(n11934) );
  NANDN U12035 ( .A(n11680), .B(n11679), .Z(n11684) );
  OR U12036 ( .A(n11682), .B(n11681), .Z(n11683) );
  AND U12037 ( .A(n11684), .B(n11683), .Z(n11692) );
  OR U12038 ( .A(n11686), .B(n11685), .Z(n11690) );
  OR U12039 ( .A(n11688), .B(n11687), .Z(n11689) );
  NAND U12040 ( .A(n11690), .B(n11689), .Z(n11691) );
  XNOR U12041 ( .A(n11692), .B(n11691), .Z(n11932) );
  OR U12042 ( .A(n11694), .B(n11693), .Z(n11698) );
  OR U12043 ( .A(n11696), .B(n11695), .Z(n11697) );
  AND U12044 ( .A(n11698), .B(n11697), .Z(n11930) );
  OR U12045 ( .A(n11700), .B(n11699), .Z(n11704) );
  OR U12046 ( .A(n11702), .B(n11701), .Z(n11703) );
  AND U12047 ( .A(n11704), .B(n11703), .Z(n11912) );
  NANDN U12048 ( .A(n11706), .B(n11705), .Z(n11710) );
  OR U12049 ( .A(n11708), .B(n11707), .Z(n11709) );
  AND U12050 ( .A(n11710), .B(n11709), .Z(n11718) );
  OR U12051 ( .A(n11712), .B(n11711), .Z(n11716) );
  NANDN U12052 ( .A(n11714), .B(n11713), .Z(n11715) );
  NAND U12053 ( .A(n11716), .B(n11715), .Z(n11717) );
  XNOR U12054 ( .A(n11718), .B(n11717), .Z(n11910) );
  OR U12055 ( .A(n11720), .B(n11719), .Z(n11724) );
  NANDN U12056 ( .A(n11722), .B(n11721), .Z(n11723) );
  AND U12057 ( .A(n11724), .B(n11723), .Z(n11908) );
  NAND U12058 ( .A(n11726), .B(n11725), .Z(n11730) );
  NOR U12059 ( .A(n11728), .B(n11727), .Z(n11729) );
  ANDN U12060 ( .B(n11730), .A(n11729), .Z(n11738) );
  ANDN U12061 ( .B(n11732), .A(n11731), .Z(n11736) );
  ANDN U12062 ( .B(n11734), .A(n11733), .Z(n11735) );
  OR U12063 ( .A(n11736), .B(n11735), .Z(n11737) );
  XNOR U12064 ( .A(n11738), .B(n11737), .Z(n11906) );
  OR U12065 ( .A(n11740), .B(n11739), .Z(n11744) );
  OR U12066 ( .A(n11742), .B(n11741), .Z(n11743) );
  AND U12067 ( .A(n11744), .B(n11743), .Z(n11904) );
  OR U12068 ( .A(n11746), .B(n11745), .Z(n11749) );
  NAND U12069 ( .A(x[138]), .B(y[757]), .Z(n11860) );
  NANDN U12070 ( .A(n11860), .B(n11747), .Z(n11748) );
  AND U12071 ( .A(n11749), .B(n11748), .Z(n11757) );
  NANDN U12072 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U12073 ( .A(n11753), .B(n11752), .Z(n11754) );
  NAND U12074 ( .A(n11755), .B(n11754), .Z(n11756) );
  XNOR U12075 ( .A(n11757), .B(n11756), .Z(n11902) );
  NANDN U12076 ( .A(n11759), .B(n11758), .Z(n11763) );
  NANDN U12077 ( .A(n11761), .B(n11760), .Z(n11762) );
  AND U12078 ( .A(n11763), .B(n11762), .Z(n11794) );
  OR U12079 ( .A(n11765), .B(n11764), .Z(n11768) );
  NAND U12080 ( .A(x[150]), .B(y[745]), .Z(n11802) );
  NANDN U12081 ( .A(n11802), .B(n11766), .Z(n11767) );
  AND U12082 ( .A(n11768), .B(n11767), .Z(n11776) );
  NANDN U12083 ( .A(n11770), .B(n11769), .Z(n11774) );
  NANDN U12084 ( .A(n11772), .B(n11771), .Z(n11773) );
  NAND U12085 ( .A(n11774), .B(n11773), .Z(n11775) );
  XNOR U12086 ( .A(n11776), .B(n11775), .Z(n11792) );
  AND U12087 ( .A(x[151]), .B(y[744]), .Z(n11778) );
  NAND U12088 ( .A(x[133]), .B(y[762]), .Z(n11777) );
  XNOR U12089 ( .A(n11778), .B(n11777), .Z(n11782) );
  AND U12090 ( .A(y[759]), .B(x[136]), .Z(n11780) );
  NAND U12091 ( .A(x[135]), .B(y[760]), .Z(n11779) );
  XNOR U12092 ( .A(n11780), .B(n11779), .Z(n11781) );
  XOR U12093 ( .A(n11782), .B(n11781), .Z(n11790) );
  AND U12094 ( .A(y[740]), .B(x[155]), .Z(n11784) );
  NAND U12095 ( .A(x[130]), .B(y[765]), .Z(n11783) );
  XNOR U12096 ( .A(n11784), .B(n11783), .Z(n11788) );
  AND U12097 ( .A(x[146]), .B(y[749]), .Z(n11786) );
  NAND U12098 ( .A(x[145]), .B(y[750]), .Z(n11785) );
  XNOR U12099 ( .A(n11786), .B(n11785), .Z(n11787) );
  XNOR U12100 ( .A(n11788), .B(n11787), .Z(n11789) );
  XNOR U12101 ( .A(n11790), .B(n11789), .Z(n11791) );
  XNOR U12102 ( .A(n11792), .B(n11791), .Z(n11793) );
  XNOR U12103 ( .A(n11794), .B(n11793), .Z(n11868) );
  OR U12104 ( .A(n11796), .B(n11795), .Z(n11800) );
  OR U12105 ( .A(n11798), .B(n11797), .Z(n11799) );
  AND U12106 ( .A(n11800), .B(n11799), .Z(n11866) );
  AND U12107 ( .A(x[159]), .B(y[736]), .Z(n11808) );
  ANDN U12108 ( .B(o[126]), .A(n11801), .Z(n11806) );
  XOR U12109 ( .A(n11886), .B(o[127]), .Z(n11804) );
  NAND U12110 ( .A(x[153]), .B(y[742]), .Z(n11878) );
  XNOR U12111 ( .A(n11802), .B(n11878), .Z(n11803) );
  XNOR U12112 ( .A(n11804), .B(n11803), .Z(n11805) );
  XNOR U12113 ( .A(n11806), .B(n11805), .Z(n11807) );
  XNOR U12114 ( .A(n11808), .B(n11807), .Z(n11816) );
  AND U12115 ( .A(y[764]), .B(x[131]), .Z(n11810) );
  NAND U12116 ( .A(x[152]), .B(y[743]), .Z(n11809) );
  XNOR U12117 ( .A(n11810), .B(n11809), .Z(n11814) );
  AND U12118 ( .A(y[761]), .B(x[134]), .Z(n11812) );
  NAND U12119 ( .A(x[132]), .B(y[763]), .Z(n11811) );
  XNOR U12120 ( .A(n11812), .B(n11811), .Z(n11813) );
  XNOR U12121 ( .A(n11814), .B(n11813), .Z(n11815) );
  XNOR U12122 ( .A(n11816), .B(n11815), .Z(n11864) );
  AND U12123 ( .A(y[747]), .B(x[148]), .Z(n11818) );
  NAND U12124 ( .A(x[144]), .B(y[751]), .Z(n11817) );
  XNOR U12125 ( .A(n11818), .B(n11817), .Z(n11822) );
  AND U12126 ( .A(x[158]), .B(y[737]), .Z(n11820) );
  NAND U12127 ( .A(x[157]), .B(y[738]), .Z(n11819) );
  XNOR U12128 ( .A(n11820), .B(n11819), .Z(n11821) );
  XOR U12129 ( .A(n11822), .B(n11821), .Z(n11830) );
  AND U12130 ( .A(y[755]), .B(x[140]), .Z(n11824) );
  NAND U12131 ( .A(x[139]), .B(y[756]), .Z(n11823) );
  XNOR U12132 ( .A(n11824), .B(n11823), .Z(n11828) );
  AND U12133 ( .A(y[767]), .B(x[128]), .Z(n11826) );
  NAND U12134 ( .A(x[154]), .B(y[741]), .Z(n11825) );
  XNOR U12135 ( .A(n11826), .B(n11825), .Z(n11827) );
  XNOR U12136 ( .A(n11828), .B(n11827), .Z(n11829) );
  XNOR U12137 ( .A(n11830), .B(n11829), .Z(n11838) );
  AND U12138 ( .A(y[752]), .B(x[143]), .Z(n11832) );
  NAND U12139 ( .A(x[129]), .B(y[766]), .Z(n11831) );
  XNOR U12140 ( .A(n11832), .B(n11831), .Z(n11836) );
  AND U12141 ( .A(x[156]), .B(y[739]), .Z(n11834) );
  NAND U12142 ( .A(x[137]), .B(y[758]), .Z(n11833) );
  XNOR U12143 ( .A(n11834), .B(n11833), .Z(n11835) );
  XNOR U12144 ( .A(n11836), .B(n11835), .Z(n11837) );
  XNOR U12145 ( .A(n11838), .B(n11837), .Z(n11854) );
  NANDN U12146 ( .A(n11840), .B(n11839), .Z(n11844) );
  NANDN U12147 ( .A(n11842), .B(n11841), .Z(n11843) );
  AND U12148 ( .A(n11844), .B(n11843), .Z(n11852) );
  OR U12149 ( .A(n11846), .B(n11845), .Z(n11850) );
  OR U12150 ( .A(n11848), .B(n11847), .Z(n11849) );
  NAND U12151 ( .A(n11850), .B(n11849), .Z(n11851) );
  XNOR U12152 ( .A(n11852), .B(n11851), .Z(n11853) );
  XOR U12153 ( .A(n11854), .B(n11853), .Z(n11862) );
  AND U12154 ( .A(x[149]), .B(y[746]), .Z(n11856) );
  NAND U12155 ( .A(x[142]), .B(y[753]), .Z(n11855) );
  XNOR U12156 ( .A(n11856), .B(n11855), .Z(n11858) );
  NAND U12157 ( .A(x[147]), .B(y[748]), .Z(n11857) );
  XNOR U12158 ( .A(n11858), .B(n11857), .Z(n11859) );
  XOR U12159 ( .A(n11860), .B(n11859), .Z(n11861) );
  XNOR U12160 ( .A(n11862), .B(n11861), .Z(n11863) );
  XNOR U12161 ( .A(n11864), .B(n11863), .Z(n11865) );
  XNOR U12162 ( .A(n11866), .B(n11865), .Z(n11867) );
  XOR U12163 ( .A(n11868), .B(n11867), .Z(n11900) );
  OR U12164 ( .A(n11870), .B(n11869), .Z(n11874) );
  OR U12165 ( .A(n11872), .B(n11871), .Z(n11873) );
  AND U12166 ( .A(n11874), .B(n11873), .Z(n11882) );
  OR U12167 ( .A(n11876), .B(n11875), .Z(n11880) );
  NANDN U12168 ( .A(n11878), .B(n11877), .Z(n11879) );
  NAND U12169 ( .A(n11880), .B(n11879), .Z(n11881) );
  XNOR U12170 ( .A(n11882), .B(n11881), .Z(n11898) );
  OR U12171 ( .A(n11884), .B(n11883), .Z(n11888) );
  NAND U12172 ( .A(n11886), .B(n11885), .Z(n11887) );
  AND U12173 ( .A(n11888), .B(n11887), .Z(n11896) );
  NANDN U12174 ( .A(n11890), .B(n11889), .Z(n11894) );
  NANDN U12175 ( .A(n11892), .B(n11891), .Z(n11893) );
  NAND U12176 ( .A(n11894), .B(n11893), .Z(n11895) );
  XNOR U12177 ( .A(n11896), .B(n11895), .Z(n11897) );
  XNOR U12178 ( .A(n11898), .B(n11897), .Z(n11899) );
  XNOR U12179 ( .A(n11900), .B(n11899), .Z(n11901) );
  XNOR U12180 ( .A(n11902), .B(n11901), .Z(n11903) );
  XNOR U12181 ( .A(n11904), .B(n11903), .Z(n11905) );
  XNOR U12182 ( .A(n11906), .B(n11905), .Z(n11907) );
  XNOR U12183 ( .A(n11908), .B(n11907), .Z(n11909) );
  XNOR U12184 ( .A(n11910), .B(n11909), .Z(n11911) );
  XNOR U12185 ( .A(n11912), .B(n11911), .Z(n11928) );
  OR U12186 ( .A(n11914), .B(n11913), .Z(n11918) );
  NANDN U12187 ( .A(n11916), .B(n11915), .Z(n11917) );
  AND U12188 ( .A(n11918), .B(n11917), .Z(n11926) );
  OR U12189 ( .A(n11920), .B(n11919), .Z(n11924) );
  NANDN U12190 ( .A(n11922), .B(n11921), .Z(n11923) );
  NAND U12191 ( .A(n11924), .B(n11923), .Z(n11925) );
  XNOR U12192 ( .A(n11926), .B(n11925), .Z(n11927) );
  XNOR U12193 ( .A(n11928), .B(n11927), .Z(n11929) );
  XNOR U12194 ( .A(n11930), .B(n11929), .Z(n11931) );
  XNOR U12195 ( .A(n11932), .B(n11931), .Z(n11933) );
  XNOR U12196 ( .A(n11934), .B(n11933), .Z(n11950) );
  OR U12197 ( .A(n11936), .B(n11935), .Z(n11940) );
  NANDN U12198 ( .A(n11938), .B(n11937), .Z(n11939) );
  AND U12199 ( .A(n11940), .B(n11939), .Z(n11948) );
  OR U12200 ( .A(n11942), .B(n11941), .Z(n11946) );
  OR U12201 ( .A(n11944), .B(n11943), .Z(n11945) );
  NAND U12202 ( .A(n11946), .B(n11945), .Z(n11947) );
  XNOR U12203 ( .A(n11948), .B(n11947), .Z(n11949) );
  XNOR U12204 ( .A(n11950), .B(n11949), .Z(n11951) );
  XNOR U12205 ( .A(n11952), .B(n11951), .Z(n11968) );
  OR U12206 ( .A(n11954), .B(n11953), .Z(n11958) );
  OR U12207 ( .A(n11956), .B(n11955), .Z(n11957) );
  AND U12208 ( .A(n11958), .B(n11957), .Z(n11966) );
  NANDN U12209 ( .A(n11960), .B(n11959), .Z(n11964) );
  OR U12210 ( .A(n11962), .B(n11961), .Z(n11963) );
  NAND U12211 ( .A(n11964), .B(n11963), .Z(n11965) );
  XNOR U12212 ( .A(n11966), .B(n11965), .Z(n11967) );
  XNOR U12213 ( .A(n11968), .B(n11967), .Z(N256) );
  AND U12214 ( .A(y[768]), .B(x[128]), .Z(n12655) );
  XOR U12215 ( .A(n12655), .B(o[128]), .Z(N289) );
  AND U12216 ( .A(y[768]), .B(x[129]), .Z(n11969) );
  NAND U12217 ( .A(x[128]), .B(y[769]), .Z(n11975) );
  XNOR U12218 ( .A(n11975), .B(o[129]), .Z(n11970) );
  XOR U12219 ( .A(n11969), .B(n11970), .Z(n11971) );
  AND U12220 ( .A(o[128]), .B(n12655), .Z(n11972) );
  XOR U12221 ( .A(n11971), .B(n11972), .Z(N290) );
  OR U12222 ( .A(n11970), .B(n11969), .Z(n11974) );
  NANDN U12223 ( .A(n11972), .B(n11971), .Z(n11973) );
  NAND U12224 ( .A(n11974), .B(n11973), .Z(n11977) );
  NAND U12225 ( .A(x[128]), .B(y[770]), .Z(n11988) );
  XOR U12226 ( .A(n11988), .B(o[130]), .Z(n11976) );
  XNOR U12227 ( .A(n11977), .B(n11976), .Z(n11979) );
  ANDN U12228 ( .B(o[129]), .A(n11975), .Z(n11982) );
  ANDN U12229 ( .B(y[768]), .A(n153), .Z(n11983) );
  XNOR U12230 ( .A(n11982), .B(n11983), .Z(n11985) );
  ANDN U12231 ( .B(y[769]), .A(n152), .Z(n11984) );
  XNOR U12232 ( .A(n11985), .B(n11984), .Z(n11978) );
  XNOR U12233 ( .A(n11979), .B(n11978), .Z(N291) );
  NAND U12234 ( .A(n11977), .B(n11976), .Z(n11981) );
  OR U12235 ( .A(n11979), .B(n11978), .Z(n11980) );
  NAND U12236 ( .A(n11981), .B(n11980), .Z(n11992) );
  OR U12237 ( .A(n11983), .B(n11982), .Z(n11987) );
  OR U12238 ( .A(n11985), .B(n11984), .Z(n11986) );
  AND U12239 ( .A(n11987), .B(n11986), .Z(n11993) );
  XNOR U12240 ( .A(n11992), .B(n11993), .Z(n11994) );
  NAND U12241 ( .A(x[130]), .B(y[769]), .Z(n12004) );
  XNOR U12242 ( .A(n12004), .B(o[131]), .Z(n11998) );
  NANDN U12243 ( .A(n11988), .B(o[130]), .Z(n12001) );
  AND U12244 ( .A(y[768]), .B(x[131]), .Z(n11990) );
  NAND U12245 ( .A(x[128]), .B(y[771]), .Z(n11989) );
  XOR U12246 ( .A(n11990), .B(n11989), .Z(n12000) );
  XNOR U12247 ( .A(n12001), .B(n12000), .Z(n11999) );
  ANDN U12248 ( .B(y[770]), .A(n152), .Z(n12028) );
  XOR U12249 ( .A(n11999), .B(n12028), .Z(n11991) );
  XOR U12250 ( .A(n11998), .B(n11991), .Z(n11995) );
  XNOR U12251 ( .A(n11994), .B(n11995), .Z(N292) );
  NANDN U12252 ( .A(n11993), .B(n11992), .Z(n11997) );
  NAND U12253 ( .A(n11995), .B(n11994), .Z(n11996) );
  NAND U12254 ( .A(n11997), .B(n11996), .Z(n12009) );
  XNOR U12255 ( .A(n12009), .B(n12010), .Z(n12011) );
  ANDN U12256 ( .B(y[771]), .A(n154), .Z(n12076) );
  NAND U12257 ( .A(n12655), .B(n12076), .Z(n12003) );
  OR U12258 ( .A(n12001), .B(n12000), .Z(n12002) );
  NAND U12259 ( .A(n12003), .B(n12002), .Z(n12018) );
  NANDN U12260 ( .A(n12004), .B(o[131]), .Z(n12025) );
  AND U12261 ( .A(y[768]), .B(x[132]), .Z(n12006) );
  AND U12262 ( .A(y[772]), .B(x[128]), .Z(n12005) );
  XNOR U12263 ( .A(n12006), .B(n12005), .Z(n12024) );
  XOR U12264 ( .A(n12025), .B(n12024), .Z(n12016) );
  AND U12265 ( .A(x[129]), .B(y[771]), .Z(n12008) );
  NAND U12266 ( .A(x[130]), .B(y[770]), .Z(n12007) );
  XOR U12267 ( .A(n12008), .B(n12007), .Z(n12030) );
  NAND U12268 ( .A(x[131]), .B(y[769]), .Z(n12021) );
  XNOR U12269 ( .A(n12021), .B(o[132]), .Z(n12029) );
  XOR U12270 ( .A(n12018), .B(n12017), .Z(n12012) );
  XOR U12271 ( .A(n12011), .B(n12012), .Z(N293) );
  NANDN U12272 ( .A(n12010), .B(n12009), .Z(n12014) );
  NANDN U12273 ( .A(n12012), .B(n12011), .Z(n12013) );
  NAND U12274 ( .A(n12014), .B(n12013), .Z(n12033) );
  NAND U12275 ( .A(n12016), .B(n12015), .Z(n12020) );
  NAND U12276 ( .A(n12018), .B(n12017), .Z(n12019) );
  NAND U12277 ( .A(n12020), .B(n12019), .Z(n12034) );
  XNOR U12278 ( .A(n12033), .B(n12034), .Z(n12035) );
  NANDN U12279 ( .A(n12021), .B(o[132]), .Z(n12052) );
  AND U12280 ( .A(y[768]), .B(x[133]), .Z(n12023) );
  AND U12281 ( .A(y[773]), .B(x[128]), .Z(n12022) );
  XNOR U12282 ( .A(n12023), .B(n12022), .Z(n12051) );
  XOR U12283 ( .A(n12052), .B(n12051), .Z(n12047) );
  ANDN U12284 ( .B(y[771]), .A(n153), .Z(n12045) );
  ANDN U12285 ( .B(y[772]), .A(n152), .Z(n12060) );
  ANDN U12286 ( .B(y[769]), .A(n155), .Z(n12055) );
  XOR U12287 ( .A(o[133]), .B(n12055), .Z(n12058) );
  ANDN U12288 ( .B(y[770]), .A(n154), .Z(n12059) );
  XNOR U12289 ( .A(n12058), .B(n12059), .Z(n12061) );
  XNOR U12290 ( .A(n12060), .B(n12061), .Z(n12046) );
  XNOR U12291 ( .A(n12045), .B(n12046), .Z(n12048) );
  XNOR U12292 ( .A(n12047), .B(n12048), .Z(n12042) );
  ANDN U12293 ( .B(y[772]), .A(n155), .Z(n12150) );
  NAND U12294 ( .A(n12655), .B(n12150), .Z(n12027) );
  OR U12295 ( .A(n12025), .B(n12024), .Z(n12026) );
  NAND U12296 ( .A(n12027), .B(n12026), .Z(n12040) );
  NAND U12297 ( .A(n12028), .B(n12045), .Z(n12032) );
  NANDN U12298 ( .A(n12030), .B(n12029), .Z(n12031) );
  NAND U12299 ( .A(n12032), .B(n12031), .Z(n12039) );
  XNOR U12300 ( .A(n12040), .B(n12039), .Z(n12041) );
  XNOR U12301 ( .A(n12042), .B(n12041), .Z(n12036) );
  XOR U12302 ( .A(n12035), .B(n12036), .Z(N294) );
  NANDN U12303 ( .A(n12034), .B(n12033), .Z(n12038) );
  NANDN U12304 ( .A(n12036), .B(n12035), .Z(n12037) );
  NAND U12305 ( .A(n12038), .B(n12037), .Z(n12064) );
  OR U12306 ( .A(n12040), .B(n12039), .Z(n12044) );
  OR U12307 ( .A(n12042), .B(n12041), .Z(n12043) );
  AND U12308 ( .A(n12044), .B(n12043), .Z(n12065) );
  XNOR U12309 ( .A(n12064), .B(n12065), .Z(n12066) );
  OR U12310 ( .A(n12046), .B(n12045), .Z(n12050) );
  OR U12311 ( .A(n12048), .B(n12047), .Z(n12049) );
  AND U12312 ( .A(n12050), .B(n12049), .Z(n12070) );
  NAND U12313 ( .A(x[133]), .B(y[773]), .Z(n12426) );
  NANDN U12314 ( .A(n12426), .B(n12655), .Z(n12054) );
  OR U12315 ( .A(n12052), .B(n12051), .Z(n12053) );
  NAND U12316 ( .A(n12054), .B(n12053), .Z(n12092) );
  NAND U12317 ( .A(n12055), .B(o[133]), .Z(n12082) );
  AND U12318 ( .A(y[768]), .B(x[134]), .Z(n12057) );
  AND U12319 ( .A(x[128]), .B(y[774]), .Z(n12056) );
  XNOR U12320 ( .A(n12057), .B(n12056), .Z(n12081) );
  XOR U12321 ( .A(n12082), .B(n12081), .Z(n12091) );
  XNOR U12322 ( .A(n12092), .B(n12091), .Z(n12094) );
  AND U12323 ( .A(y[773]), .B(x[129]), .Z(n12360) );
  NAND U12324 ( .A(x[133]), .B(y[769]), .Z(n12085) );
  XNOR U12325 ( .A(n12085), .B(o[134]), .Z(n12086) );
  XNOR U12326 ( .A(n12360), .B(n12086), .Z(n12088) );
  AND U12327 ( .A(y[770]), .B(x[132]), .Z(n12087) );
  XOR U12328 ( .A(n12088), .B(n12087), .Z(n12077) );
  AND U12329 ( .A(y[772]), .B(x[130]), .Z(n12415) );
  XNOR U12330 ( .A(n12076), .B(n12415), .Z(n12078) );
  XOR U12331 ( .A(n12077), .B(n12078), .Z(n12093) );
  XNOR U12332 ( .A(n12094), .B(n12093), .Z(n12071) );
  XOR U12333 ( .A(n12070), .B(n12071), .Z(n12072) );
  OR U12334 ( .A(n12059), .B(n12058), .Z(n12063) );
  OR U12335 ( .A(n12061), .B(n12060), .Z(n12062) );
  AND U12336 ( .A(n12063), .B(n12062), .Z(n12073) );
  XOR U12337 ( .A(n12066), .B(n12067), .Z(N295) );
  NANDN U12338 ( .A(n12065), .B(n12064), .Z(n12069) );
  NANDN U12339 ( .A(n12067), .B(n12066), .Z(n12068) );
  NAND U12340 ( .A(n12069), .B(n12068), .Z(n12126) );
  OR U12341 ( .A(n12071), .B(n12070), .Z(n12075) );
  NANDN U12342 ( .A(n12073), .B(n12072), .Z(n12074) );
  AND U12343 ( .A(n12075), .B(n12074), .Z(n12127) );
  XNOR U12344 ( .A(n12126), .B(n12127), .Z(n12128) );
  OR U12345 ( .A(n12076), .B(n12415), .Z(n12080) );
  NANDN U12346 ( .A(n12078), .B(n12077), .Z(n12079) );
  NAND U12347 ( .A(n12080), .B(n12079), .Z(n12123) );
  AND U12348 ( .A(y[774]), .B(x[134]), .Z(n12348) );
  NAND U12349 ( .A(n12655), .B(n12348), .Z(n12084) );
  OR U12350 ( .A(n12082), .B(n12081), .Z(n12083) );
  AND U12351 ( .A(n12084), .B(n12083), .Z(n12121) );
  ANDN U12352 ( .B(y[770]), .A(n156), .Z(n12257) );
  AND U12353 ( .A(y[774]), .B(x[129]), .Z(n12476) );
  NAND U12354 ( .A(x[134]), .B(y[769]), .Z(n12109) );
  XNOR U12355 ( .A(o[135]), .B(n12109), .Z(n12110) );
  XNOR U12356 ( .A(n12476), .B(n12110), .Z(n12111) );
  XNOR U12357 ( .A(n12257), .B(n12111), .Z(n12120) );
  XOR U12358 ( .A(n12121), .B(n12120), .Z(n12122) );
  XNOR U12359 ( .A(n12123), .B(n12122), .Z(n12132) );
  AND U12360 ( .A(y[773]), .B(x[130]), .Z(n12583) );
  ANDN U12361 ( .B(y[771]), .A(n155), .Z(n12279) );
  ANDN U12362 ( .B(y[772]), .A(n154), .Z(n12105) );
  XNOR U12363 ( .A(n12279), .B(n12105), .Z(n12106) );
  XNOR U12364 ( .A(n12583), .B(n12106), .Z(n12114) );
  NAND U12365 ( .A(x[128]), .B(y[775]), .Z(n12101) );
  ANDN U12366 ( .B(o[134]), .A(n12085), .Z(n12100) );
  NAND U12367 ( .A(x[135]), .B(y[768]), .Z(n12099) );
  XOR U12368 ( .A(n12100), .B(n12099), .Z(n12102) );
  XNOR U12369 ( .A(n12101), .B(n12102), .Z(n12115) );
  XOR U12370 ( .A(n12114), .B(n12115), .Z(n12117) );
  NAND U12371 ( .A(n12360), .B(n12086), .Z(n12090) );
  NANDN U12372 ( .A(n12088), .B(n12087), .Z(n12089) );
  AND U12373 ( .A(n12090), .B(n12089), .Z(n12116) );
  XOR U12374 ( .A(n12117), .B(n12116), .Z(n12133) );
  XOR U12375 ( .A(n12132), .B(n12133), .Z(n12135) );
  OR U12376 ( .A(n12092), .B(n12091), .Z(n12096) );
  OR U12377 ( .A(n12094), .B(n12093), .Z(n12095) );
  AND U12378 ( .A(n12096), .B(n12095), .Z(n12134) );
  XOR U12379 ( .A(n12135), .B(n12134), .Z(n12129) );
  XNOR U12380 ( .A(n12128), .B(n12129), .Z(N296) );
  AND U12381 ( .A(y[768]), .B(x[136]), .Z(n12098) );
  NAND U12382 ( .A(x[128]), .B(y[776]), .Z(n12097) );
  XOR U12383 ( .A(n12098), .B(n12097), .Z(n12159) );
  NAND U12384 ( .A(x[135]), .B(y[769]), .Z(n12162) );
  XNOR U12385 ( .A(n12162), .B(o[136]), .Z(n12158) );
  XOR U12386 ( .A(n12159), .B(n12158), .Z(n12179) );
  NANDN U12387 ( .A(n12100), .B(n12099), .Z(n12104) );
  NANDN U12388 ( .A(n12102), .B(n12101), .Z(n12103) );
  NAND U12389 ( .A(n12104), .B(n12103), .Z(n12178) );
  XOR U12390 ( .A(n12179), .B(n12178), .Z(n12180) );
  OR U12391 ( .A(n12105), .B(n12279), .Z(n12108) );
  OR U12392 ( .A(n12106), .B(n12583), .Z(n12107) );
  NAND U12393 ( .A(n12108), .B(n12107), .Z(n12181) );
  XNOR U12394 ( .A(n12180), .B(n12181), .Z(n12146) );
  ANDN U12395 ( .B(y[770]), .A(n157), .Z(n12151) );
  XNOR U12396 ( .A(n12150), .B(n12151), .Z(n12152) );
  NOR U12397 ( .A(n153), .B(n150), .Z(n12665) );
  XNOR U12398 ( .A(n12152), .B(n12665), .Z(n12153) );
  ANDN U12399 ( .B(y[773]), .A(n154), .Z(n12970) );
  XNOR U12400 ( .A(n12153), .B(n12970), .Z(n12155) );
  NANDN U12401 ( .A(n12109), .B(o[135]), .Z(n12169) );
  AND U12402 ( .A(x[133]), .B(y[771]), .Z(n12767) );
  AND U12403 ( .A(y[775]), .B(x[129]), .Z(n12650) );
  XNOR U12404 ( .A(n12767), .B(n12650), .Z(n12168) );
  XOR U12405 ( .A(n12169), .B(n12168), .Z(n12154) );
  XNOR U12406 ( .A(n12155), .B(n12154), .Z(n12172) );
  NAND U12407 ( .A(n12476), .B(n12110), .Z(n12113) );
  NANDN U12408 ( .A(n12111), .B(n12257), .Z(n12112) );
  AND U12409 ( .A(n12113), .B(n12112), .Z(n12173) );
  XOR U12410 ( .A(n12172), .B(n12173), .Z(n12175) );
  NANDN U12411 ( .A(n12115), .B(n12114), .Z(n12119) );
  OR U12412 ( .A(n12117), .B(n12116), .Z(n12118) );
  AND U12413 ( .A(n12119), .B(n12118), .Z(n12174) );
  XOR U12414 ( .A(n12175), .B(n12174), .Z(n12144) );
  NANDN U12415 ( .A(n12121), .B(n12120), .Z(n12125) );
  OR U12416 ( .A(n12123), .B(n12122), .Z(n12124) );
  NAND U12417 ( .A(n12125), .B(n12124), .Z(n12145) );
  XNOR U12418 ( .A(n12144), .B(n12145), .Z(n12147) );
  XNOR U12419 ( .A(n12146), .B(n12147), .Z(n12141) );
  NANDN U12420 ( .A(n12127), .B(n12126), .Z(n12131) );
  NAND U12421 ( .A(n12129), .B(n12128), .Z(n12130) );
  NAND U12422 ( .A(n12131), .B(n12130), .Z(n12138) );
  NANDN U12423 ( .A(n12133), .B(n12132), .Z(n12137) );
  OR U12424 ( .A(n12135), .B(n12134), .Z(n12136) );
  AND U12425 ( .A(n12137), .B(n12136), .Z(n12139) );
  XNOR U12426 ( .A(n12138), .B(n12139), .Z(n12140) );
  XOR U12427 ( .A(n12141), .B(n12140), .Z(N297) );
  NANDN U12428 ( .A(n12139), .B(n12138), .Z(n12143) );
  NANDN U12429 ( .A(n12141), .B(n12140), .Z(n12142) );
  NAND U12430 ( .A(n12143), .B(n12142), .Z(n12184) );
  OR U12431 ( .A(n12145), .B(n12144), .Z(n12149) );
  OR U12432 ( .A(n12147), .B(n12146), .Z(n12148) );
  AND U12433 ( .A(n12149), .B(n12148), .Z(n12185) );
  XNOR U12434 ( .A(n12184), .B(n12185), .Z(n12186) );
  OR U12435 ( .A(n12153), .B(n12970), .Z(n12157) );
  OR U12436 ( .A(n12155), .B(n12154), .Z(n12156) );
  NAND U12437 ( .A(n12157), .B(n12156), .Z(n12212) );
  XOR U12438 ( .A(n12213), .B(n12212), .Z(n12214) );
  AND U12439 ( .A(y[776]), .B(x[136]), .Z(n12662) );
  NAND U12440 ( .A(n12655), .B(n12662), .Z(n12161) );
  NANDN U12441 ( .A(n12159), .B(n12158), .Z(n12160) );
  NAND U12442 ( .A(n12161), .B(n12160), .Z(n12199) );
  NANDN U12443 ( .A(n12162), .B(o[136]), .Z(n12219) );
  AND U12444 ( .A(y[772]), .B(x[133]), .Z(n12163) );
  AND U12445 ( .A(y[770]), .B(x[135]), .Z(n12587) );
  XNOR U12446 ( .A(n12163), .B(n12587), .Z(n12218) );
  XOR U12447 ( .A(n12219), .B(n12218), .Z(n12197) );
  AND U12448 ( .A(y[768]), .B(x[137]), .Z(n12165) );
  NAND U12449 ( .A(x[128]), .B(y[777]), .Z(n12164) );
  XOR U12450 ( .A(n12165), .B(n12164), .Z(n12230) );
  NAND U12451 ( .A(x[136]), .B(y[769]), .Z(n12224) );
  XOR U12452 ( .A(n12224), .B(o[137]), .Z(n12229) );
  XNOR U12453 ( .A(n12230), .B(n12229), .Z(n12196) );
  XOR U12454 ( .A(n12197), .B(n12196), .Z(n12198) );
  XNOR U12455 ( .A(n12199), .B(n12198), .Z(n12208) );
  NAND U12456 ( .A(x[132]), .B(y[773]), .Z(n12646) );
  AND U12457 ( .A(x[134]), .B(y[771]), .Z(n12167) );
  NAND U12458 ( .A(x[129]), .B(y[776]), .Z(n12166) );
  XNOR U12459 ( .A(n12167), .B(n12166), .Z(n12226) );
  XNOR U12460 ( .A(n12646), .B(n12226), .Z(n12202) );
  ANDN U12461 ( .B(y[775]), .A(n153), .Z(n12880) );
  NAND U12462 ( .A(y[774]), .B(x[131]), .Z(n12556) );
  XOR U12463 ( .A(n12880), .B(n12556), .Z(n12203) );
  XNOR U12464 ( .A(n12202), .B(n12203), .Z(n12206) );
  NAND U12465 ( .A(x[129]), .B(y[771]), .Z(n12225) );
  AND U12466 ( .A(y[775]), .B(x[133]), .Z(n12350) );
  NANDN U12467 ( .A(n12225), .B(n12350), .Z(n12171) );
  OR U12468 ( .A(n12169), .B(n12168), .Z(n12170) );
  AND U12469 ( .A(n12171), .B(n12170), .Z(n12207) );
  XOR U12470 ( .A(n12206), .B(n12207), .Z(n12209) );
  XOR U12471 ( .A(n12208), .B(n12209), .Z(n12215) );
  NANDN U12472 ( .A(n12173), .B(n12172), .Z(n12177) );
  OR U12473 ( .A(n12175), .B(n12174), .Z(n12176) );
  NAND U12474 ( .A(n12177), .B(n12176), .Z(n12191) );
  OR U12475 ( .A(n12179), .B(n12178), .Z(n12183) );
  NANDN U12476 ( .A(n12181), .B(n12180), .Z(n12182) );
  NAND U12477 ( .A(n12183), .B(n12182), .Z(n12190) );
  XOR U12478 ( .A(n12191), .B(n12190), .Z(n12193) );
  XNOR U12479 ( .A(n12192), .B(n12193), .Z(n12187) );
  XOR U12480 ( .A(n12186), .B(n12187), .Z(N298) );
  NANDN U12481 ( .A(n12185), .B(n12184), .Z(n12189) );
  NANDN U12482 ( .A(n12187), .B(n12186), .Z(n12188) );
  NAND U12483 ( .A(n12189), .B(n12188), .Z(n12233) );
  OR U12484 ( .A(n12191), .B(n12190), .Z(n12195) );
  NAND U12485 ( .A(n12193), .B(n12192), .Z(n12194) );
  AND U12486 ( .A(n12195), .B(n12194), .Z(n12234) );
  XNOR U12487 ( .A(n12233), .B(n12234), .Z(n12235) );
  NANDN U12488 ( .A(n12197), .B(n12196), .Z(n12201) );
  OR U12489 ( .A(n12199), .B(n12198), .Z(n12200) );
  NAND U12490 ( .A(n12201), .B(n12200), .Z(n12291) );
  NANDN U12491 ( .A(n12880), .B(n12556), .Z(n12205) );
  OR U12492 ( .A(n12203), .B(n12202), .Z(n12204) );
  NAND U12493 ( .A(n12205), .B(n12204), .Z(n12290) );
  XOR U12494 ( .A(n12291), .B(n12290), .Z(n12292) );
  NANDN U12495 ( .A(n12207), .B(n12206), .Z(n12211) );
  NANDN U12496 ( .A(n12209), .B(n12208), .Z(n12210) );
  AND U12497 ( .A(n12211), .B(n12210), .Z(n12293) );
  XNOR U12498 ( .A(n12292), .B(n12293), .Z(n12241) );
  OR U12499 ( .A(n12213), .B(n12212), .Z(n12217) );
  NANDN U12500 ( .A(n12215), .B(n12214), .Z(n12216) );
  NAND U12501 ( .A(n12217), .B(n12216), .Z(n12240) );
  ANDN U12502 ( .B(y[772]), .A(n158), .Z(n12342) );
  NAND U12503 ( .A(n12257), .B(n12342), .Z(n12221) );
  OR U12504 ( .A(n12219), .B(n12218), .Z(n12220) );
  AND U12505 ( .A(n12221), .B(n12220), .Z(n12247) );
  AND U12506 ( .A(y[770]), .B(x[136]), .Z(n12341) );
  XOR U12507 ( .A(n12341), .B(n12426), .Z(n12259) );
  NAND U12508 ( .A(x[137]), .B(y[769]), .Z(n12268) );
  XOR U12509 ( .A(o[138]), .B(n12268), .Z(n12258) );
  XOR U12510 ( .A(n12259), .B(n12258), .Z(n12245) );
  ANDN U12511 ( .B(y[772]), .A(n157), .Z(n12485) );
  AND U12512 ( .A(x[132]), .B(y[774]), .Z(n12223) );
  NAND U12513 ( .A(x[135]), .B(y[771]), .Z(n12222) );
  XOR U12514 ( .A(n12223), .B(n12222), .Z(n12281) );
  XOR U12515 ( .A(n12485), .B(n12281), .Z(n12246) );
  XNOR U12516 ( .A(n12247), .B(n12248), .Z(n12286) );
  ANDN U12517 ( .B(y[778]), .A(n151), .Z(n12276) );
  NANDN U12518 ( .A(n12224), .B(o[137]), .Z(n12273) );
  ANDN U12519 ( .B(y[768]), .A(n161), .Z(n12274) );
  XNOR U12520 ( .A(n12276), .B(n12275), .Z(n12264) );
  AND U12521 ( .A(y[775]), .B(x[131]), .Z(n13155) );
  ANDN U12522 ( .B(y[776]), .A(n153), .Z(n12255) );
  XOR U12523 ( .A(n13155), .B(n12255), .Z(n12256) );
  XNOR U12524 ( .A(n13212), .B(n12256), .Z(n12263) );
  ANDN U12525 ( .B(y[776]), .A(n157), .Z(n12580) );
  NANDN U12526 ( .A(n12225), .B(n12580), .Z(n12228) );
  NANDN U12527 ( .A(n12646), .B(n12226), .Z(n12227) );
  AND U12528 ( .A(n12228), .B(n12227), .Z(n12262) );
  XOR U12529 ( .A(n12263), .B(n12262), .Z(n12265) );
  AND U12530 ( .A(y[777]), .B(x[137]), .Z(n12858) );
  NAND U12531 ( .A(n12655), .B(n12858), .Z(n12232) );
  OR U12532 ( .A(n12230), .B(n12229), .Z(n12231) );
  NAND U12533 ( .A(n12232), .B(n12231), .Z(n12284) );
  XNOR U12534 ( .A(n12285), .B(n12284), .Z(n12287) );
  XOR U12535 ( .A(n12286), .B(n12287), .Z(n12239) );
  XNOR U12536 ( .A(n12240), .B(n12239), .Z(n12242) );
  XNOR U12537 ( .A(n12241), .B(n12242), .Z(n12236) );
  XOR U12538 ( .A(n12235), .B(n12236), .Z(N299) );
  NANDN U12539 ( .A(n12234), .B(n12233), .Z(n12238) );
  NANDN U12540 ( .A(n12236), .B(n12235), .Z(n12237) );
  NAND U12541 ( .A(n12238), .B(n12237), .Z(n12296) );
  OR U12542 ( .A(n12240), .B(n12239), .Z(n12244) );
  OR U12543 ( .A(n12242), .B(n12241), .Z(n12243) );
  AND U12544 ( .A(n12244), .B(n12243), .Z(n12297) );
  XNOR U12545 ( .A(n12296), .B(n12297), .Z(n12298) );
  NANDN U12546 ( .A(n12246), .B(n12245), .Z(n12250) );
  OR U12547 ( .A(n12248), .B(n12247), .Z(n12249) );
  AND U12548 ( .A(n12250), .B(n12249), .Z(n12310) );
  AND U12549 ( .A(y[776]), .B(x[131]), .Z(n13360) );
  AND U12550 ( .A(x[133]), .B(y[774]), .Z(n12252) );
  NAND U12551 ( .A(x[130]), .B(y[777]), .Z(n12251) );
  XOR U12552 ( .A(n12252), .B(n12251), .Z(n12357) );
  NAND U12553 ( .A(x[132]), .B(y[775]), .Z(n12356) );
  XNOR U12554 ( .A(n12357), .B(n12356), .Z(n12326) );
  XOR U12555 ( .A(n13360), .B(n12326), .Z(n12328) );
  AND U12556 ( .A(x[136]), .B(y[771]), .Z(n12254) );
  NAND U12557 ( .A(x[137]), .B(y[770]), .Z(n12253) );
  XNOR U12558 ( .A(n12254), .B(n12253), .Z(n12343) );
  XNOR U12559 ( .A(n12342), .B(n12343), .Z(n12327) );
  XOR U12560 ( .A(n12328), .B(n12327), .Z(n12334) );
  ANDN U12561 ( .B(y[773]), .A(n159), .Z(n13090) );
  NAND U12562 ( .A(n13090), .B(n12257), .Z(n12261) );
  OR U12563 ( .A(n12259), .B(n12258), .Z(n12260) );
  NAND U12564 ( .A(n12261), .B(n12260), .Z(n12332) );
  XNOR U12565 ( .A(n12334), .B(n12333), .Z(n12308) );
  OR U12566 ( .A(n12263), .B(n12262), .Z(n12267) );
  NAND U12567 ( .A(n12265), .B(n12264), .Z(n12266) );
  NAND U12568 ( .A(n12267), .B(n12266), .Z(n12317) );
  NANDN U12569 ( .A(n12268), .B(o[138]), .Z(n12338) );
  AND U12570 ( .A(y[768]), .B(x[139]), .Z(n12270) );
  NAND U12571 ( .A(x[128]), .B(y[779]), .Z(n12269) );
  XNOR U12572 ( .A(n12270), .B(n12269), .Z(n12337) );
  AND U12573 ( .A(y[773]), .B(x[134]), .Z(n12272) );
  NAND U12574 ( .A(x[129]), .B(y[778]), .Z(n12271) );
  XOR U12575 ( .A(n12272), .B(n12271), .Z(n12362) );
  NAND U12576 ( .A(x[138]), .B(y[769]), .Z(n12346) );
  XOR U12577 ( .A(o[139]), .B(n12346), .Z(n12361) );
  XOR U12578 ( .A(n12362), .B(n12361), .Z(n12320) );
  NANDN U12579 ( .A(n12274), .B(n12273), .Z(n12278) );
  OR U12580 ( .A(n12276), .B(n12275), .Z(n12277) );
  NAND U12581 ( .A(n12278), .B(n12277), .Z(n12323) );
  XOR U12582 ( .A(n12322), .B(n12323), .Z(n12314) );
  AND U12583 ( .A(y[774]), .B(x[135]), .Z(n12280) );
  NAND U12584 ( .A(n12280), .B(n12279), .Z(n12283) );
  NANDN U12585 ( .A(n12281), .B(n12485), .Z(n12282) );
  NAND U12586 ( .A(n12283), .B(n12282), .Z(n12315) );
  XNOR U12587 ( .A(n12317), .B(n12316), .Z(n12309) );
  XNOR U12588 ( .A(n12308), .B(n12309), .Z(n12311) );
  XOR U12589 ( .A(n12310), .B(n12311), .Z(n12302) );
  OR U12590 ( .A(n12285), .B(n12284), .Z(n12289) );
  NANDN U12591 ( .A(n12287), .B(n12286), .Z(n12288) );
  AND U12592 ( .A(n12289), .B(n12288), .Z(n12303) );
  XNOR U12593 ( .A(n12302), .B(n12303), .Z(n12305) );
  OR U12594 ( .A(n12291), .B(n12290), .Z(n12295) );
  NANDN U12595 ( .A(n12293), .B(n12292), .Z(n12294) );
  NAND U12596 ( .A(n12295), .B(n12294), .Z(n12304) );
  XOR U12597 ( .A(n12305), .B(n12304), .Z(n12299) );
  XNOR U12598 ( .A(n12298), .B(n12299), .Z(N300) );
  NANDN U12599 ( .A(n12297), .B(n12296), .Z(n12301) );
  NAND U12600 ( .A(n12299), .B(n12298), .Z(n12300) );
  NAND U12601 ( .A(n12301), .B(n12300), .Z(n12365) );
  OR U12602 ( .A(n12303), .B(n12302), .Z(n12307) );
  OR U12603 ( .A(n12305), .B(n12304), .Z(n12306) );
  AND U12604 ( .A(n12307), .B(n12306), .Z(n12366) );
  XNOR U12605 ( .A(n12365), .B(n12366), .Z(n12367) );
  OR U12606 ( .A(n12309), .B(n12308), .Z(n12313) );
  OR U12607 ( .A(n12311), .B(n12310), .Z(n12312) );
  NAND U12608 ( .A(n12313), .B(n12312), .Z(n12372) );
  NANDN U12609 ( .A(n12315), .B(n12314), .Z(n12319) );
  NANDN U12610 ( .A(n12317), .B(n12316), .Z(n12318) );
  NAND U12611 ( .A(n12319), .B(n12318), .Z(n12380) );
  NAND U12612 ( .A(n12321), .B(n12320), .Z(n12325) );
  NANDN U12613 ( .A(n12323), .B(n12322), .Z(n12324) );
  NAND U12614 ( .A(n12325), .B(n12324), .Z(n12378) );
  NANDN U12615 ( .A(n12326), .B(n13360), .Z(n12330) );
  OR U12616 ( .A(n12328), .B(n12327), .Z(n12329) );
  AND U12617 ( .A(n12330), .B(n12329), .Z(n12377) );
  XNOR U12618 ( .A(n12380), .B(n12379), .Z(n12371) );
  XNOR U12619 ( .A(n12372), .B(n12371), .Z(n12374) );
  NANDN U12620 ( .A(n12332), .B(n12331), .Z(n12336) );
  NANDN U12621 ( .A(n12334), .B(n12333), .Z(n12335) );
  NAND U12622 ( .A(n12336), .B(n12335), .Z(n12440) );
  ANDN U12623 ( .B(y[779]), .A(n162), .Z(n13476) );
  NAND U12624 ( .A(n12655), .B(n13476), .Z(n12340) );
  NANDN U12625 ( .A(n12338), .B(n12337), .Z(n12339) );
  AND U12626 ( .A(n12340), .B(n12339), .Z(n12405) );
  NAND U12627 ( .A(x[137]), .B(y[771]), .Z(n13033) );
  NANDN U12628 ( .A(n13033), .B(n12341), .Z(n12345) );
  NAND U12629 ( .A(n12343), .B(n12342), .Z(n12344) );
  AND U12630 ( .A(n12345), .B(n12344), .Z(n12403) );
  NANDN U12631 ( .A(n12346), .B(o[139]), .Z(n12384) );
  NAND U12632 ( .A(x[129]), .B(y[779]), .Z(n12347) );
  XOR U12633 ( .A(n12348), .B(n12347), .Z(n12383) );
  XNOR U12634 ( .A(n12384), .B(n12383), .Z(n12404) );
  XNOR U12635 ( .A(n12403), .B(n12404), .Z(n12406) );
  XNOR U12636 ( .A(n12405), .B(n12406), .Z(n12437) );
  NAND U12637 ( .A(x[135]), .B(y[773]), .Z(n12349) );
  XOR U12638 ( .A(n12350), .B(n12349), .Z(n12428) );
  NAND U12639 ( .A(x[132]), .B(y[776]), .Z(n12400) );
  AND U12640 ( .A(y[770]), .B(x[138]), .Z(n12351) );
  XOR U12641 ( .A(n12351), .B(n13033), .Z(n12399) );
  XNOR U12642 ( .A(n12400), .B(n12399), .Z(n12427) );
  XNOR U12643 ( .A(n12428), .B(n12427), .Z(n12434) );
  AND U12644 ( .A(y[768]), .B(x[140]), .Z(n12353) );
  NAND U12645 ( .A(x[128]), .B(y[780]), .Z(n12352) );
  XOR U12646 ( .A(n12353), .B(n12352), .Z(n12388) );
  NAND U12647 ( .A(x[139]), .B(y[769]), .Z(n12422) );
  XOR U12648 ( .A(o[140]), .B(n12422), .Z(n12387) );
  XOR U12649 ( .A(n12388), .B(n12387), .Z(n12431) );
  AND U12650 ( .A(y[772]), .B(x[136]), .Z(n12355) );
  NAND U12651 ( .A(x[130]), .B(y[778]), .Z(n12354) );
  XOR U12652 ( .A(n12355), .B(n12354), .Z(n12417) );
  NAND U12653 ( .A(y[777]), .B(x[131]), .Z(n12416) );
  XNOR U12654 ( .A(n12417), .B(n12416), .Z(n12432) );
  XOR U12655 ( .A(n12431), .B(n12432), .Z(n12433) );
  XOR U12656 ( .A(n12434), .B(n12433), .Z(n12412) );
  ANDN U12657 ( .B(y[777]), .A(n156), .Z(n12557) );
  NAND U12658 ( .A(n12665), .B(n12557), .Z(n12359) );
  OR U12659 ( .A(n12357), .B(n12356), .Z(n12358) );
  NAND U12660 ( .A(n12359), .B(n12358), .Z(n12410) );
  AND U12661 ( .A(y[778]), .B(x[134]), .Z(n12645) );
  NAND U12662 ( .A(n12645), .B(n12360), .Z(n12364) );
  OR U12663 ( .A(n12362), .B(n12361), .Z(n12363) );
  NAND U12664 ( .A(n12364), .B(n12363), .Z(n12409) );
  XOR U12665 ( .A(n12410), .B(n12409), .Z(n12411) );
  XOR U12666 ( .A(n12412), .B(n12411), .Z(n12438) );
  XNOR U12667 ( .A(n12440), .B(n12439), .Z(n12373) );
  XNOR U12668 ( .A(n12374), .B(n12373), .Z(n12368) );
  XOR U12669 ( .A(n12367), .B(n12368), .Z(N301) );
  NANDN U12670 ( .A(n12366), .B(n12365), .Z(n12370) );
  NANDN U12671 ( .A(n12368), .B(n12367), .Z(n12369) );
  NAND U12672 ( .A(n12370), .B(n12369), .Z(n12508) );
  OR U12673 ( .A(n12372), .B(n12371), .Z(n12376) );
  OR U12674 ( .A(n12374), .B(n12373), .Z(n12375) );
  AND U12675 ( .A(n12376), .B(n12375), .Z(n12509) );
  XNOR U12676 ( .A(n12508), .B(n12509), .Z(n12510) );
  NANDN U12677 ( .A(n12378), .B(n12377), .Z(n12382) );
  NAND U12678 ( .A(n12380), .B(n12379), .Z(n12381) );
  NAND U12679 ( .A(n12382), .B(n12381), .Z(n12517) );
  ANDN U12680 ( .B(y[779]), .A(n157), .Z(n12888) );
  NAND U12681 ( .A(n12476), .B(n12888), .Z(n12386) );
  OR U12682 ( .A(n12384), .B(n12383), .Z(n12385) );
  NAND U12683 ( .A(n12386), .B(n12385), .Z(n12464) );
  ANDN U12684 ( .B(y[780]), .A(n163), .Z(n13697) );
  NAND U12685 ( .A(n12655), .B(n13697), .Z(n12390) );
  OR U12686 ( .A(n12388), .B(n12387), .Z(n12389) );
  NAND U12687 ( .A(n12390), .B(n12389), .Z(n12461) );
  AND U12688 ( .A(y[770]), .B(x[139]), .Z(n12392) );
  NAND U12689 ( .A(x[138]), .B(y[771]), .Z(n12391) );
  XNOR U12690 ( .A(n12392), .B(n12391), .Z(n12482) );
  XNOR U12691 ( .A(n13090), .B(n12482), .Z(n12462) );
  XOR U12692 ( .A(n12464), .B(n12463), .Z(n12455) );
  AND U12693 ( .A(y[778]), .B(x[131]), .Z(n12394) );
  NAND U12694 ( .A(x[133]), .B(y[776]), .Z(n12393) );
  XOR U12695 ( .A(n12394), .B(n12393), .Z(n12495) );
  NAND U12696 ( .A(y[777]), .B(x[132]), .Z(n12494) );
  XOR U12697 ( .A(n12495), .B(n12494), .Z(n12502) );
  AND U12698 ( .A(y[768]), .B(x[141]), .Z(n12396) );
  NAND U12699 ( .A(x[128]), .B(y[781]), .Z(n12395) );
  XOR U12700 ( .A(n12396), .B(n12395), .Z(n12499) );
  NAND U12701 ( .A(x[140]), .B(y[769]), .Z(n12491) );
  XOR U12702 ( .A(o[141]), .B(n12491), .Z(n12498) );
  XNOR U12703 ( .A(n12499), .B(n12498), .Z(n12503) );
  AND U12704 ( .A(y[770]), .B(x[137]), .Z(n12398) );
  AND U12705 ( .A(y[771]), .B(x[138]), .Z(n12397) );
  NAND U12706 ( .A(n12398), .B(n12397), .Z(n12402) );
  OR U12707 ( .A(n12400), .B(n12399), .Z(n12401) );
  AND U12708 ( .A(n12402), .B(n12401), .Z(n12504) );
  XOR U12709 ( .A(n12505), .B(n12504), .Z(n12456) );
  XNOR U12710 ( .A(n12455), .B(n12456), .Z(n12458) );
  OR U12711 ( .A(n12404), .B(n12403), .Z(n12408) );
  OR U12712 ( .A(n12406), .B(n12405), .Z(n12407) );
  NAND U12713 ( .A(n12408), .B(n12407), .Z(n12457) );
  XOR U12714 ( .A(n12458), .B(n12457), .Z(n12452) );
  OR U12715 ( .A(n12410), .B(n12409), .Z(n12414) );
  NANDN U12716 ( .A(n12412), .B(n12411), .Z(n12413) );
  AND U12717 ( .A(n12414), .B(n12413), .Z(n12449) );
  AND U12718 ( .A(y[778]), .B(x[136]), .Z(n12845) );
  NAND U12719 ( .A(n12845), .B(n12415), .Z(n12419) );
  OR U12720 ( .A(n12417), .B(n12416), .Z(n12418) );
  NAND U12721 ( .A(n12419), .B(n12418), .Z(n12470) );
  AND U12722 ( .A(y[775]), .B(x[134]), .Z(n12421) );
  NAND U12723 ( .A(x[137]), .B(y[772]), .Z(n12420) );
  XOR U12724 ( .A(n12421), .B(n12420), .Z(n12487) );
  NAND U12725 ( .A(x[130]), .B(y[779]), .Z(n12486) );
  XOR U12726 ( .A(n12487), .B(n12486), .Z(n12468) );
  NANDN U12727 ( .A(n12422), .B(o[140]), .Z(n12479) );
  AND U12728 ( .A(y[780]), .B(x[129]), .Z(n12424) );
  NAND U12729 ( .A(x[135]), .B(y[774]), .Z(n12423) );
  XNOR U12730 ( .A(n12424), .B(n12423), .Z(n12478) );
  XNOR U12731 ( .A(n12470), .B(n12469), .Z(n12444) );
  AND U12732 ( .A(y[775]), .B(x[135]), .Z(n12425) );
  NANDN U12733 ( .A(n12426), .B(n12425), .Z(n12430) );
  OR U12734 ( .A(n12428), .B(n12427), .Z(n12429) );
  AND U12735 ( .A(n12430), .B(n12429), .Z(n12443) );
  XOR U12736 ( .A(n12444), .B(n12443), .Z(n12445) );
  NANDN U12737 ( .A(n12432), .B(n12431), .Z(n12436) );
  OR U12738 ( .A(n12434), .B(n12433), .Z(n12435) );
  AND U12739 ( .A(n12436), .B(n12435), .Z(n12446) );
  XNOR U12740 ( .A(n12445), .B(n12446), .Z(n12450) );
  XOR U12741 ( .A(n12449), .B(n12450), .Z(n12451) );
  XOR U12742 ( .A(n12452), .B(n12451), .Z(n12514) );
  NANDN U12743 ( .A(n12438), .B(n12437), .Z(n12442) );
  NAND U12744 ( .A(n12440), .B(n12439), .Z(n12441) );
  NAND U12745 ( .A(n12442), .B(n12441), .Z(n12515) );
  XOR U12746 ( .A(n12514), .B(n12515), .Z(n12516) );
  XNOR U12747 ( .A(n12517), .B(n12516), .Z(n12511) );
  XOR U12748 ( .A(n12510), .B(n12511), .Z(N302) );
  OR U12749 ( .A(n12444), .B(n12443), .Z(n12448) );
  NANDN U12750 ( .A(n12446), .B(n12445), .Z(n12447) );
  NAND U12751 ( .A(n12448), .B(n12447), .Z(n12529) );
  OR U12752 ( .A(n12450), .B(n12449), .Z(n12454) );
  NAND U12753 ( .A(n12452), .B(n12451), .Z(n12453) );
  AND U12754 ( .A(n12454), .B(n12453), .Z(n12526) );
  OR U12755 ( .A(n12456), .B(n12455), .Z(n12460) );
  OR U12756 ( .A(n12458), .B(n12457), .Z(n12459) );
  AND U12757 ( .A(n12460), .B(n12459), .Z(n12535) );
  NANDN U12758 ( .A(n12462), .B(n12461), .Z(n12466) );
  NAND U12759 ( .A(n12464), .B(n12463), .Z(n12465) );
  NAND U12760 ( .A(n12466), .B(n12465), .Z(n12546) );
  NAND U12761 ( .A(n12468), .B(n12467), .Z(n12472) );
  NAND U12762 ( .A(n12470), .B(n12469), .Z(n12471) );
  NAND U12763 ( .A(n12472), .B(n12471), .Z(n12544) );
  AND U12764 ( .A(y[779]), .B(x[131]), .Z(n12474) );
  NAND U12765 ( .A(x[136]), .B(y[774]), .Z(n12473) );
  XOR U12766 ( .A(n12474), .B(n12473), .Z(n12558) );
  XOR U12767 ( .A(n12557), .B(n12558), .Z(n12567) );
  ANDN U12768 ( .B(y[778]), .A(n155), .Z(n12566) );
  ANDN U12769 ( .B(y[772]), .A(n161), .Z(n13160) );
  AND U12770 ( .A(y[773]), .B(x[137]), .Z(n13201) );
  NAND U12771 ( .A(x[130]), .B(y[780]), .Z(n12475) );
  XOR U12772 ( .A(n13201), .B(n12475), .Z(n12584) );
  XOR U12773 ( .A(n13160), .B(n12584), .Z(n12565) );
  XNOR U12774 ( .A(n12567), .B(n12568), .Z(n12574) );
  AND U12775 ( .A(y[780]), .B(x[135]), .Z(n12477) );
  NAND U12776 ( .A(n12477), .B(n12476), .Z(n12481) );
  NANDN U12777 ( .A(n12479), .B(n12478), .Z(n12480) );
  NAND U12778 ( .A(n12481), .B(n12480), .Z(n12571) );
  NAND U12779 ( .A(x[138]), .B(y[770]), .Z(n13095) );
  NANDN U12780 ( .A(n13095), .B(n12680), .Z(n12484) );
  NAND U12781 ( .A(n12482), .B(n13090), .Z(n12483) );
  AND U12782 ( .A(n12484), .B(n12483), .Z(n12572) );
  XOR U12783 ( .A(n12574), .B(n12573), .Z(n12545) );
  XOR U12784 ( .A(n12544), .B(n12545), .Z(n12547) );
  AND U12785 ( .A(y[775]), .B(x[137]), .Z(n12679) );
  NAND U12786 ( .A(n12679), .B(n12485), .Z(n12489) );
  OR U12787 ( .A(n12487), .B(n12486), .Z(n12488) );
  NAND U12788 ( .A(n12489), .B(n12488), .Z(n12600) );
  AND U12789 ( .A(y[770]), .B(x[140]), .Z(n13207) );
  NAND U12790 ( .A(x[135]), .B(y[775]), .Z(n12490) );
  XOR U12791 ( .A(n13207), .B(n12490), .Z(n12589) );
  NAND U12792 ( .A(x[141]), .B(y[769]), .Z(n12592) );
  XOR U12793 ( .A(o[142]), .B(n12592), .Z(n12588) );
  XOR U12794 ( .A(n12589), .B(n12588), .Z(n12598) );
  NANDN U12795 ( .A(n12491), .B(o[141]), .Z(n12562) );
  AND U12796 ( .A(y[782]), .B(x[128]), .Z(n12493) );
  NAND U12797 ( .A(x[142]), .B(y[768]), .Z(n12492) );
  XNOR U12798 ( .A(n12493), .B(n12492), .Z(n12561) );
  XOR U12799 ( .A(n12600), .B(n12599), .Z(n12538) );
  ANDN U12800 ( .B(y[778]), .A(n156), .Z(n12639) );
  NAND U12801 ( .A(n13360), .B(n12639), .Z(n12497) );
  OR U12802 ( .A(n12495), .B(n12494), .Z(n12496) );
  NAND U12803 ( .A(n12497), .B(n12496), .Z(n12606) );
  IV U12804 ( .A(n12680), .Z(n12578) );
  IV U12805 ( .A(y[781]), .Z(n13714) );
  NANDN U12806 ( .A(n13714), .B(x[129]), .Z(n12577) );
  XNOR U12807 ( .A(n12578), .B(n12577), .Z(n12579) );
  XOR U12808 ( .A(n12580), .B(n12579), .Z(n12604) );
  ANDN U12809 ( .B(x[141]), .A(n13714), .Z(n14069) );
  NAND U12810 ( .A(n12655), .B(n14069), .Z(n12501) );
  OR U12811 ( .A(n12499), .B(n12498), .Z(n12500) );
  AND U12812 ( .A(n12501), .B(n12500), .Z(n12603) );
  XOR U12813 ( .A(n12604), .B(n12603), .Z(n12605) );
  XOR U12814 ( .A(n12606), .B(n12605), .Z(n12539) );
  XNOR U12815 ( .A(n12538), .B(n12539), .Z(n12541) );
  NANDN U12816 ( .A(n12503), .B(n12502), .Z(n12507) );
  OR U12817 ( .A(n12505), .B(n12504), .Z(n12506) );
  NAND U12818 ( .A(n12507), .B(n12506), .Z(n12540) );
  XNOR U12819 ( .A(n12541), .B(n12540), .Z(n12532) );
  XOR U12820 ( .A(n12533), .B(n12532), .Z(n12534) );
  XOR U12821 ( .A(n12535), .B(n12534), .Z(n12527) );
  XNOR U12822 ( .A(n12526), .B(n12527), .Z(n12528) );
  XNOR U12823 ( .A(n12529), .B(n12528), .Z(n12523) );
  NANDN U12824 ( .A(n12509), .B(n12508), .Z(n12513) );
  NANDN U12825 ( .A(n12511), .B(n12510), .Z(n12512) );
  NAND U12826 ( .A(n12513), .B(n12512), .Z(n12520) );
  OR U12827 ( .A(n12515), .B(n12514), .Z(n12519) );
  NANDN U12828 ( .A(n12517), .B(n12516), .Z(n12518) );
  NAND U12829 ( .A(n12519), .B(n12518), .Z(n12521) );
  XNOR U12830 ( .A(n12520), .B(n12521), .Z(n12522) );
  XOR U12831 ( .A(n12523), .B(n12522), .Z(N303) );
  NANDN U12832 ( .A(n12521), .B(n12520), .Z(n12525) );
  NANDN U12833 ( .A(n12523), .B(n12522), .Z(n12524) );
  NAND U12834 ( .A(n12525), .B(n12524), .Z(n12609) );
  OR U12835 ( .A(n12527), .B(n12526), .Z(n12531) );
  OR U12836 ( .A(n12529), .B(n12528), .Z(n12530) );
  AND U12837 ( .A(n12531), .B(n12530), .Z(n12610) );
  XNOR U12838 ( .A(n12609), .B(n12610), .Z(n12611) );
  OR U12839 ( .A(n12533), .B(n12532), .Z(n12537) );
  NANDN U12840 ( .A(n12535), .B(n12534), .Z(n12536) );
  AND U12841 ( .A(n12537), .B(n12536), .Z(n12615) );
  OR U12842 ( .A(n12539), .B(n12538), .Z(n12543) );
  OR U12843 ( .A(n12541), .B(n12540), .Z(n12542) );
  AND U12844 ( .A(n12543), .B(n12542), .Z(n12616) );
  XOR U12845 ( .A(n12615), .B(n12616), .Z(n12617) );
  NANDN U12846 ( .A(n12545), .B(n12544), .Z(n12549) );
  NANDN U12847 ( .A(n12547), .B(n12546), .Z(n12548) );
  NAND U12848 ( .A(n12549), .B(n12548), .Z(n12699) );
  NAND U12849 ( .A(x[142]), .B(y[769]), .Z(n12660) );
  XOR U12850 ( .A(o[143]), .B(n12660), .Z(n12652) );
  AND U12851 ( .A(y[775]), .B(x[136]), .Z(n12551) );
  NAND U12852 ( .A(x[129]), .B(y[782]), .Z(n12550) );
  XNOR U12853 ( .A(n12551), .B(n12550), .Z(n12651) );
  XNOR U12854 ( .A(n12652), .B(n12651), .Z(n12685) );
  NAND U12855 ( .A(x[131]), .B(y[780]), .Z(n12667) );
  AND U12856 ( .A(x[137]), .B(y[774]), .Z(n12553) );
  NAND U12857 ( .A(x[130]), .B(y[781]), .Z(n12552) );
  XOR U12858 ( .A(n12553), .B(n12552), .Z(n12666) );
  XOR U12859 ( .A(n12667), .B(n12666), .Z(n12686) );
  XNOR U12860 ( .A(n12685), .B(n12686), .Z(n12688) );
  ANDN U12861 ( .B(y[776]), .A(n158), .Z(n13048) );
  AND U12862 ( .A(y[773]), .B(x[138]), .Z(n12555) );
  NAND U12863 ( .A(x[132]), .B(y[779]), .Z(n12554) );
  XOR U12864 ( .A(n12555), .B(n12554), .Z(n12647) );
  XNOR U12865 ( .A(n13048), .B(n12647), .Z(n12640) );
  AND U12866 ( .A(x[134]), .B(y[777]), .Z(n12774) );
  XNOR U12867 ( .A(n12639), .B(n12774), .Z(n12641) );
  XOR U12868 ( .A(n12640), .B(n12641), .Z(n12687) );
  XOR U12869 ( .A(n12688), .B(n12687), .Z(n12673) );
  NAND U12870 ( .A(x[136]), .B(y[779]), .Z(n12977) );
  OR U12871 ( .A(n12977), .B(n12556), .Z(n12560) );
  NANDN U12872 ( .A(n12558), .B(n12557), .Z(n12559) );
  NAND U12873 ( .A(n12560), .B(n12559), .Z(n12671) );
  AND U12874 ( .A(y[782]), .B(x[142]), .Z(n14356) );
  NAND U12875 ( .A(n12655), .B(n14356), .Z(n12564) );
  NANDN U12876 ( .A(n12562), .B(n12561), .Z(n12563) );
  AND U12877 ( .A(n12564), .B(n12563), .Z(n12670) );
  XOR U12878 ( .A(n12673), .B(n12672), .Z(n12628) );
  NANDN U12879 ( .A(n12566), .B(n12565), .Z(n12570) );
  NANDN U12880 ( .A(n12568), .B(n12567), .Z(n12569) );
  AND U12881 ( .A(n12570), .B(n12569), .Z(n12627) );
  XNOR U12882 ( .A(n12628), .B(n12627), .Z(n12630) );
  NANDN U12883 ( .A(n12572), .B(n12571), .Z(n12576) );
  NANDN U12884 ( .A(n12574), .B(n12573), .Z(n12575) );
  NAND U12885 ( .A(n12576), .B(n12575), .Z(n12629) );
  XOR U12886 ( .A(n12630), .B(n12629), .Z(n12698) );
  NAND U12887 ( .A(n12578), .B(n12577), .Z(n12582) );
  OR U12888 ( .A(n12580), .B(n12579), .Z(n12581) );
  AND U12889 ( .A(n12582), .B(n12581), .Z(n12636) );
  ANDN U12890 ( .B(y[780]), .A(n160), .Z(n13314) );
  NAND U12891 ( .A(n13314), .B(n12583), .Z(n12586) );
  NANDN U12892 ( .A(n12584), .B(n13160), .Z(n12585) );
  NAND U12893 ( .A(n12586), .B(n12585), .Z(n12634) );
  AND U12894 ( .A(y[775]), .B(x[140]), .Z(n12934) );
  NAND U12895 ( .A(n12587), .B(n12934), .Z(n12591) );
  OR U12896 ( .A(n12589), .B(n12588), .Z(n12590) );
  NAND U12897 ( .A(n12591), .B(n12590), .Z(n12694) );
  NANDN U12898 ( .A(n12592), .B(o[142]), .Z(n12657) );
  AND U12899 ( .A(y[768]), .B(x[143]), .Z(n12594) );
  NAND U12900 ( .A(x[128]), .B(y[783]), .Z(n12593) );
  XOR U12901 ( .A(n12594), .B(n12593), .Z(n12656) );
  XNOR U12902 ( .A(n12657), .B(n12656), .Z(n12691) );
  AND U12903 ( .A(x[140]), .B(y[771]), .Z(n12596) );
  NAND U12904 ( .A(x[139]), .B(y[772]), .Z(n12595) );
  XOR U12905 ( .A(n12596), .B(n12595), .Z(n12682) );
  NAND U12906 ( .A(x[141]), .B(y[770]), .Z(n12681) );
  XOR U12907 ( .A(n12682), .B(n12681), .Z(n12692) );
  XOR U12908 ( .A(n12694), .B(n12693), .Z(n12633) );
  XOR U12909 ( .A(n12634), .B(n12633), .Z(n12635) );
  XNOR U12910 ( .A(n12636), .B(n12635), .Z(n12621) );
  NAND U12911 ( .A(n12598), .B(n12597), .Z(n12602) );
  NAND U12912 ( .A(n12600), .B(n12599), .Z(n12601) );
  AND U12913 ( .A(n12602), .B(n12601), .Z(n12622) );
  XNOR U12914 ( .A(n12621), .B(n12622), .Z(n12624) );
  OR U12915 ( .A(n12604), .B(n12603), .Z(n12608) );
  NAND U12916 ( .A(n12606), .B(n12605), .Z(n12607) );
  AND U12917 ( .A(n12608), .B(n12607), .Z(n12623) );
  XOR U12918 ( .A(n12624), .B(n12623), .Z(n12697) );
  XOR U12919 ( .A(n12698), .B(n12697), .Z(n12700) );
  XNOR U12920 ( .A(n12699), .B(n12700), .Z(n12618) );
  XOR U12921 ( .A(n12617), .B(n12618), .Z(n12612) );
  XOR U12922 ( .A(n12611), .B(n12612), .Z(N304) );
  NANDN U12923 ( .A(n12610), .B(n12609), .Z(n12614) );
  NANDN U12924 ( .A(n12612), .B(n12611), .Z(n12613) );
  NAND U12925 ( .A(n12614), .B(n12613), .Z(n12703) );
  OR U12926 ( .A(n12616), .B(n12615), .Z(n12620) );
  NANDN U12927 ( .A(n12618), .B(n12617), .Z(n12619) );
  AND U12928 ( .A(n12620), .B(n12619), .Z(n12704) );
  XNOR U12929 ( .A(n12703), .B(n12704), .Z(n12705) );
  OR U12930 ( .A(n12622), .B(n12621), .Z(n12626) );
  OR U12931 ( .A(n12624), .B(n12623), .Z(n12625) );
  NAND U12932 ( .A(n12626), .B(n12625), .Z(n12793) );
  OR U12933 ( .A(n12628), .B(n12627), .Z(n12632) );
  OR U12934 ( .A(n12630), .B(n12629), .Z(n12631) );
  AND U12935 ( .A(n12632), .B(n12631), .Z(n12790) );
  OR U12936 ( .A(n12634), .B(n12633), .Z(n12638) );
  NANDN U12937 ( .A(n12636), .B(n12635), .Z(n12637) );
  AND U12938 ( .A(n12638), .B(n12637), .Z(n12791) );
  XOR U12939 ( .A(n12790), .B(n12791), .Z(n12792) );
  XNOR U12940 ( .A(n12793), .B(n12792), .Z(n12712) );
  OR U12941 ( .A(n12639), .B(n12774), .Z(n12643) );
  OR U12942 ( .A(n12641), .B(n12640), .Z(n12642) );
  AND U12943 ( .A(n12643), .B(n12642), .Z(n12749) );
  NAND U12944 ( .A(x[128]), .B(y[784]), .Z(n12784) );
  NAND U12945 ( .A(x[144]), .B(y[768]), .Z(n12783) );
  XOR U12946 ( .A(n12784), .B(n12783), .Z(n12786) );
  AND U12947 ( .A(y[769]), .B(x[143]), .Z(n12771) );
  XOR U12948 ( .A(o[144]), .B(n12771), .Z(n12785) );
  NAND U12949 ( .A(x[135]), .B(y[777]), .Z(n12644) );
  XOR U12950 ( .A(n12645), .B(n12644), .Z(n12776) );
  NAND U12951 ( .A(x[138]), .B(y[774]), .Z(n12775) );
  XNOR U12952 ( .A(n12776), .B(n12775), .Z(n12762) );
  XOR U12953 ( .A(n12761), .B(n12762), .Z(n12764) );
  ANDN U12954 ( .B(y[779]), .A(n161), .Z(n13347) );
  NANDN U12955 ( .A(n12646), .B(n13347), .Z(n12649) );
  NANDN U12956 ( .A(n12647), .B(n13048), .Z(n12648) );
  AND U12957 ( .A(n12649), .B(n12648), .Z(n12763) );
  XNOR U12958 ( .A(n12764), .B(n12763), .Z(n12740) );
  NAND U12959 ( .A(x[136]), .B(y[782]), .Z(n13588) );
  NANDN U12960 ( .A(n13588), .B(n12650), .Z(n12654) );
  NANDN U12961 ( .A(n12652), .B(n12651), .Z(n12653) );
  AND U12962 ( .A(n12654), .B(n12653), .Z(n12737) );
  AND U12963 ( .A(y[783]), .B(x[143]), .Z(n14788) );
  NAND U12964 ( .A(n12655), .B(n14788), .Z(n12659) );
  OR U12965 ( .A(n12657), .B(n12656), .Z(n12658) );
  AND U12966 ( .A(n12659), .B(n12658), .Z(n12738) );
  XOR U12967 ( .A(n12737), .B(n12738), .Z(n12739) );
  XNOR U12968 ( .A(n12740), .B(n12739), .Z(n12750) );
  XOR U12969 ( .A(n12749), .B(n12750), .Z(n12751) );
  NANDN U12970 ( .A(n12660), .B(o[143]), .Z(n12780) );
  NAND U12971 ( .A(x[129]), .B(y[783]), .Z(n12661) );
  XOR U12972 ( .A(n12662), .B(n12661), .Z(n12779) );
  XNOR U12973 ( .A(n12780), .B(n12779), .Z(n12757) );
  AND U12974 ( .A(y[773]), .B(x[139]), .Z(n12664) );
  NAND U12975 ( .A(x[142]), .B(y[770]), .Z(n12663) );
  XOR U12976 ( .A(n12664), .B(n12663), .Z(n12728) );
  NAND U12977 ( .A(x[132]), .B(y[780]), .Z(n12727) );
  XOR U12978 ( .A(n12728), .B(n12727), .Z(n12756) );
  ANDN U12979 ( .B(y[781]), .A(n160), .Z(n13417) );
  NAND U12980 ( .A(n12665), .B(n13417), .Z(n12669) );
  OR U12981 ( .A(n12667), .B(n12666), .Z(n12668) );
  NAND U12982 ( .A(n12669), .B(n12668), .Z(n12755) );
  XNOR U12983 ( .A(n12756), .B(n12755), .Z(n12758) );
  XOR U12984 ( .A(n12757), .B(n12758), .Z(n12752) );
  XOR U12985 ( .A(n12751), .B(n12752), .Z(n12744) );
  NANDN U12986 ( .A(n12671), .B(n12670), .Z(n12675) );
  NANDN U12987 ( .A(n12673), .B(n12672), .Z(n12674) );
  AND U12988 ( .A(n12675), .B(n12674), .Z(n12743) );
  XOR U12989 ( .A(n12744), .B(n12743), .Z(n12745) );
  ANDN U12990 ( .B(y[772]), .A(n163), .Z(n13421) );
  AND U12991 ( .A(x[141]), .B(y[771]), .Z(n12677) );
  NAND U12992 ( .A(x[133]), .B(y[779]), .Z(n12676) );
  XNOR U12993 ( .A(n12677), .B(n12676), .Z(n12768) );
  XNOR U12994 ( .A(n13421), .B(n12768), .Z(n12732) );
  NAND U12995 ( .A(x[130]), .B(y[782]), .Z(n12678) );
  XOR U12996 ( .A(n12679), .B(n12678), .Z(n12723) );
  NAND U12997 ( .A(x[131]), .B(y[781]), .Z(n12722) );
  XNOR U12998 ( .A(n12723), .B(n12722), .Z(n12731) );
  XOR U12999 ( .A(n12732), .B(n12731), .Z(n12733) );
  NAND U13000 ( .A(n12680), .B(n13421), .Z(n12684) );
  OR U13001 ( .A(n12682), .B(n12681), .Z(n12683) );
  AND U13002 ( .A(n12684), .B(n12683), .Z(n12734) );
  OR U13003 ( .A(n12686), .B(n12685), .Z(n12690) );
  NANDN U13004 ( .A(n12688), .B(n12687), .Z(n12689) );
  NAND U13005 ( .A(n12690), .B(n12689), .Z(n12715) );
  XNOR U13006 ( .A(n12716), .B(n12715), .Z(n12718) );
  NANDN U13007 ( .A(n12692), .B(n12691), .Z(n12696) );
  NANDN U13008 ( .A(n12694), .B(n12693), .Z(n12695) );
  NAND U13009 ( .A(n12696), .B(n12695), .Z(n12717) );
  XOR U13010 ( .A(n12718), .B(n12717), .Z(n12746) );
  XNOR U13011 ( .A(n12745), .B(n12746), .Z(n12710) );
  NANDN U13012 ( .A(n12698), .B(n12697), .Z(n12702) );
  NANDN U13013 ( .A(n12700), .B(n12699), .Z(n12701) );
  AND U13014 ( .A(n12702), .B(n12701), .Z(n12709) );
  XOR U13015 ( .A(n12710), .B(n12709), .Z(n12711) );
  XNOR U13016 ( .A(n12712), .B(n12711), .Z(n12706) );
  XOR U13017 ( .A(n12705), .B(n12706), .Z(N305) );
  NANDN U13018 ( .A(n12704), .B(n12703), .Z(n12708) );
  NANDN U13019 ( .A(n12706), .B(n12705), .Z(n12707) );
  NAND U13020 ( .A(n12708), .B(n12707), .Z(n12796) );
  OR U13021 ( .A(n12710), .B(n12709), .Z(n12714) );
  NANDN U13022 ( .A(n12712), .B(n12711), .Z(n12713) );
  NAND U13023 ( .A(n12714), .B(n12713), .Z(n12797) );
  XNOR U13024 ( .A(n12796), .B(n12797), .Z(n12798) );
  OR U13025 ( .A(n12716), .B(n12715), .Z(n12720) );
  OR U13026 ( .A(n12718), .B(n12717), .Z(n12719) );
  AND U13027 ( .A(n12720), .B(n12719), .Z(n12894) );
  AND U13028 ( .A(y[778]), .B(x[135]), .Z(n12976) );
  ANDN U13029 ( .B(y[781]), .A(n155), .Z(n12851) );
  ANDN U13030 ( .B(y[774]), .A(n162), .Z(n12849) );
  ANDN U13031 ( .B(y[772]), .A(n164), .Z(n12848) );
  XNOR U13032 ( .A(n12849), .B(n12848), .Z(n12850) );
  XNOR U13033 ( .A(n12851), .B(n12850), .Z(n12871) );
  ANDN U13034 ( .B(y[780]), .A(n156), .Z(n12890) );
  ANDN U13035 ( .B(y[777]), .A(n159), .Z(n12887) );
  XOR U13036 ( .A(n12888), .B(n12887), .Z(n12889) );
  XNOR U13037 ( .A(n12890), .B(n12889), .Z(n12872) );
  XNOR U13038 ( .A(n12871), .B(n12872), .Z(n12873) );
  XOR U13039 ( .A(n12976), .B(n12873), .Z(n12868) );
  AND U13040 ( .A(y[782]), .B(x[137]), .Z(n12721) );
  NAND U13041 ( .A(n12721), .B(n12880), .Z(n12725) );
  OR U13042 ( .A(n12723), .B(n12722), .Z(n12724) );
  NAND U13043 ( .A(n12725), .B(n12724), .Z(n12866) );
  NAND U13044 ( .A(x[139]), .B(y[770]), .Z(n12938) );
  AND U13045 ( .A(y[773]), .B(x[142]), .Z(n12726) );
  NANDN U13046 ( .A(n12938), .B(n12726), .Z(n12730) );
  OR U13047 ( .A(n12728), .B(n12727), .Z(n12729) );
  AND U13048 ( .A(n12730), .B(n12729), .Z(n12865) );
  XNOR U13049 ( .A(n12868), .B(n12867), .Z(n12808) );
  OR U13050 ( .A(n12732), .B(n12731), .Z(n12736) );
  NANDN U13051 ( .A(n12734), .B(n12733), .Z(n12735) );
  AND U13052 ( .A(n12736), .B(n12735), .Z(n12809) );
  XNOR U13053 ( .A(n12808), .B(n12809), .Z(n12811) );
  OR U13054 ( .A(n12738), .B(n12737), .Z(n12742) );
  NANDN U13055 ( .A(n12740), .B(n12739), .Z(n12741) );
  AND U13056 ( .A(n12742), .B(n12741), .Z(n12810) );
  XOR U13057 ( .A(n12811), .B(n12810), .Z(n12893) );
  OR U13058 ( .A(n12744), .B(n12743), .Z(n12748) );
  NANDN U13059 ( .A(n12746), .B(n12745), .Z(n12747) );
  NAND U13060 ( .A(n12748), .B(n12747), .Z(n12895) );
  XOR U13061 ( .A(n12896), .B(n12895), .Z(n12804) );
  OR U13062 ( .A(n12750), .B(n12749), .Z(n12754) );
  NANDN U13063 ( .A(n12752), .B(n12751), .Z(n12753) );
  NAND U13064 ( .A(n12754), .B(n12753), .Z(n12902) );
  OR U13065 ( .A(n12756), .B(n12755), .Z(n12760) );
  NANDN U13066 ( .A(n12758), .B(n12757), .Z(n12759) );
  NAND U13067 ( .A(n12760), .B(n12759), .Z(n12900) );
  NANDN U13068 ( .A(n12762), .B(n12761), .Z(n12766) );
  OR U13069 ( .A(n12764), .B(n12763), .Z(n12765) );
  NAND U13070 ( .A(n12766), .B(n12765), .Z(n12817) );
  ANDN U13071 ( .B(y[779]), .A(n164), .Z(n13689) );
  NAND U13072 ( .A(n13689), .B(n12767), .Z(n12770) );
  NAND U13073 ( .A(n12768), .B(n13421), .Z(n12769) );
  NAND U13074 ( .A(n12770), .B(n12769), .Z(n12834) );
  NAND U13075 ( .A(x[140]), .B(y[773]), .Z(n12861) );
  ANDN U13076 ( .B(y[771]), .A(n165), .Z(n12860) );
  NAND U13077 ( .A(x[143]), .B(y[770]), .Z(n12859) );
  XOR U13078 ( .A(n12860), .B(n12859), .Z(n12862) );
  XNOR U13079 ( .A(n12861), .B(n12862), .Z(n12833) );
  NAND U13080 ( .A(n12771), .B(o[144]), .Z(n12877) );
  AND U13081 ( .A(y[776]), .B(x[137]), .Z(n12773) );
  AND U13082 ( .A(y[784]), .B(x[129]), .Z(n12772) );
  XNOR U13083 ( .A(n12773), .B(n12772), .Z(n12876) );
  XOR U13084 ( .A(n12877), .B(n12876), .Z(n12832) );
  XOR U13085 ( .A(n12833), .B(n12832), .Z(n12835) );
  XNOR U13086 ( .A(n12834), .B(n12835), .Z(n12814) );
  NAND U13087 ( .A(n12976), .B(n12774), .Z(n12778) );
  OR U13088 ( .A(n12776), .B(n12775), .Z(n12777) );
  NAND U13089 ( .A(n12778), .B(n12777), .Z(n12820) );
  NAND U13090 ( .A(x[136]), .B(y[783]), .Z(n13416) );
  ANDN U13091 ( .B(y[776]), .A(n152), .Z(n12963) );
  NANDN U13092 ( .A(n13416), .B(n12963), .Z(n12782) );
  OR U13093 ( .A(n12780), .B(n12779), .Z(n12781) );
  AND U13094 ( .A(n12782), .B(n12781), .Z(n12821) );
  OR U13095 ( .A(n12784), .B(n12783), .Z(n12788) );
  NAND U13096 ( .A(n12786), .B(n12785), .Z(n12787) );
  NAND U13097 ( .A(n12788), .B(n12787), .Z(n12827) );
  AND U13098 ( .A(y[775]), .B(x[138]), .Z(n13445) );
  NAND U13099 ( .A(x[130]), .B(y[783]), .Z(n12789) );
  XOR U13100 ( .A(n13445), .B(n12789), .Z(n12882) );
  AND U13101 ( .A(y[782]), .B(x[131]), .Z(n12881) );
  XNOR U13102 ( .A(n12882), .B(n12881), .Z(n12826) );
  XNOR U13103 ( .A(n12827), .B(n12826), .Z(n12829) );
  AND U13104 ( .A(y[769]), .B(x[144]), .Z(n12854) );
  XNOR U13105 ( .A(o[145]), .B(n12854), .Z(n12839) );
  AND U13106 ( .A(y[768]), .B(x[145]), .Z(n12838) );
  XOR U13107 ( .A(n12839), .B(n12838), .Z(n12841) );
  AND U13108 ( .A(x[128]), .B(y[785]), .Z(n12840) );
  XNOR U13109 ( .A(n12841), .B(n12840), .Z(n12828) );
  XOR U13110 ( .A(n12829), .B(n12828), .Z(n12823) );
  XNOR U13111 ( .A(n12822), .B(n12823), .Z(n12815) );
  XNOR U13112 ( .A(n12814), .B(n12815), .Z(n12816) );
  XOR U13113 ( .A(n12817), .B(n12816), .Z(n12899) );
  XNOR U13114 ( .A(n12900), .B(n12899), .Z(n12901) );
  XNOR U13115 ( .A(n12902), .B(n12901), .Z(n12802) );
  OR U13116 ( .A(n12791), .B(n12790), .Z(n12795) );
  NANDN U13117 ( .A(n12793), .B(n12792), .Z(n12794) );
  AND U13118 ( .A(n12795), .B(n12794), .Z(n12803) );
  XOR U13119 ( .A(n12802), .B(n12803), .Z(n12805) );
  XNOR U13120 ( .A(n12804), .B(n12805), .Z(n12799) );
  XOR U13121 ( .A(n12798), .B(n12799), .Z(N306) );
  NANDN U13122 ( .A(n12797), .B(n12796), .Z(n12801) );
  NANDN U13123 ( .A(n12799), .B(n12798), .Z(n12800) );
  NAND U13124 ( .A(n12801), .B(n12800), .Z(n13009) );
  NANDN U13125 ( .A(n12803), .B(n12802), .Z(n12807) );
  OR U13126 ( .A(n12805), .B(n12804), .Z(n12806) );
  AND U13127 ( .A(n12807), .B(n12806), .Z(n13010) );
  XNOR U13128 ( .A(n13009), .B(n13010), .Z(n13011) );
  OR U13129 ( .A(n12809), .B(n12808), .Z(n12813) );
  OR U13130 ( .A(n12811), .B(n12810), .Z(n12812) );
  NAND U13131 ( .A(n12813), .B(n12812), .Z(n12912) );
  OR U13132 ( .A(n12815), .B(n12814), .Z(n12819) );
  OR U13133 ( .A(n12817), .B(n12816), .Z(n12818) );
  AND U13134 ( .A(n12819), .B(n12818), .Z(n12911) );
  XOR U13135 ( .A(n12912), .B(n12911), .Z(n12914) );
  NANDN U13136 ( .A(n12821), .B(n12820), .Z(n12825) );
  NANDN U13137 ( .A(n12823), .B(n12822), .Z(n12824) );
  NAND U13138 ( .A(n12825), .B(n12824), .Z(n12987) );
  NAND U13139 ( .A(n12827), .B(n12826), .Z(n12831) );
  NANDN U13140 ( .A(n12829), .B(n12828), .Z(n12830) );
  NAND U13141 ( .A(n12831), .B(n12830), .Z(n12985) );
  NANDN U13142 ( .A(n12833), .B(n12832), .Z(n12837) );
  NANDN U13143 ( .A(n12835), .B(n12834), .Z(n12836) );
  AND U13144 ( .A(n12837), .B(n12836), .Z(n12986) );
  XOR U13145 ( .A(n12987), .B(n12988), .Z(n12907) );
  NANDN U13146 ( .A(n12839), .B(n12838), .Z(n12843) );
  NANDN U13147 ( .A(n12841), .B(n12840), .Z(n12842) );
  NAND U13148 ( .A(n12843), .B(n12842), .Z(n12992) );
  NAND U13149 ( .A(x[132]), .B(y[782]), .Z(n12979) );
  AND U13150 ( .A(y[779]), .B(x[135]), .Z(n12844) );
  XNOR U13151 ( .A(n12845), .B(n12844), .Z(n12978) );
  XOR U13152 ( .A(n12979), .B(n12978), .Z(n12924) );
  ANDN U13153 ( .B(y[780]), .A(n157), .Z(n12923) );
  AND U13154 ( .A(x[133]), .B(y[781]), .Z(n13074) );
  XNOR U13155 ( .A(n12923), .B(n13074), .Z(n12925) );
  XNOR U13156 ( .A(n12924), .B(n12925), .Z(n12991) );
  XOR U13157 ( .A(n12992), .B(n12991), .Z(n12993) );
  NAND U13158 ( .A(x[130]), .B(y[784]), .Z(n12940) );
  AND U13159 ( .A(y[775]), .B(x[139]), .Z(n12847) );
  NAND U13160 ( .A(x[144]), .B(y[770]), .Z(n12846) );
  XOR U13161 ( .A(n12847), .B(n12846), .Z(n12939) );
  XOR U13162 ( .A(n12940), .B(n12939), .Z(n12994) );
  XOR U13163 ( .A(n12993), .B(n12994), .Z(n13005) );
  OR U13164 ( .A(n12849), .B(n12848), .Z(n12853) );
  OR U13165 ( .A(n12851), .B(n12850), .Z(n12852) );
  NAND U13166 ( .A(n12853), .B(n12852), .Z(n12946) );
  NAND U13167 ( .A(n12854), .B(o[145]), .Z(n12965) );
  AND U13168 ( .A(y[776]), .B(x[138]), .Z(n12856) );
  AND U13169 ( .A(x[129]), .B(y[785]), .Z(n12855) );
  XNOR U13170 ( .A(n12856), .B(n12855), .Z(n12964) );
  XOR U13171 ( .A(n12965), .B(n12964), .Z(n12943) );
  NAND U13172 ( .A(x[143]), .B(y[771]), .Z(n12930) );
  AND U13173 ( .A(y[772]), .B(x[142]), .Z(n12857) );
  XNOR U13174 ( .A(n12858), .B(n12857), .Z(n12929) );
  XNOR U13175 ( .A(n12930), .B(n12929), .Z(n12944) );
  XOR U13176 ( .A(n12943), .B(n12944), .Z(n12945) );
  XNOR U13177 ( .A(n12946), .B(n12945), .Z(n13004) );
  NANDN U13178 ( .A(n12860), .B(n12859), .Z(n12864) );
  NANDN U13179 ( .A(n12862), .B(n12861), .Z(n12863) );
  AND U13180 ( .A(n12864), .B(n12863), .Z(n13003) );
  XOR U13181 ( .A(n13005), .B(n13006), .Z(n12905) );
  NANDN U13182 ( .A(n12866), .B(n12865), .Z(n12870) );
  NANDN U13183 ( .A(n12868), .B(n12867), .Z(n12869) );
  NAND U13184 ( .A(n12870), .B(n12869), .Z(n12919) );
  NANDN U13185 ( .A(n12872), .B(n12871), .Z(n12875) );
  NAND U13186 ( .A(n12873), .B(n12976), .Z(n12874) );
  NAND U13187 ( .A(n12875), .B(n12874), .Z(n12918) );
  AND U13188 ( .A(y[784]), .B(x[137]), .Z(n13926) );
  NAND U13189 ( .A(n12963), .B(n13926), .Z(n12879) );
  OR U13190 ( .A(n12877), .B(n12876), .Z(n12878) );
  NAND U13191 ( .A(n12879), .B(n12878), .Z(n13000) );
  IV U13192 ( .A(y[783]), .Z(n13574) );
  NOR U13193 ( .A(n161), .B(n13574), .Z(n13925) );
  NAND U13194 ( .A(n13925), .B(n12880), .Z(n12884) );
  NANDN U13195 ( .A(n12882), .B(n12881), .Z(n12883) );
  AND U13196 ( .A(n12884), .B(n12883), .Z(n12952) );
  AND U13197 ( .A(y[769]), .B(x[145]), .Z(n12982) );
  XNOR U13198 ( .A(o[146]), .B(n12982), .Z(n12960) );
  NAND U13199 ( .A(x[128]), .B(y[786]), .Z(n12958) );
  NAND U13200 ( .A(x[146]), .B(y[768]), .Z(n12957) );
  XNOR U13201 ( .A(n12958), .B(n12957), .Z(n12959) );
  XNOR U13202 ( .A(n12960), .B(n12959), .Z(n12950) );
  AND U13203 ( .A(y[774]), .B(x[140]), .Z(n13042) );
  AND U13204 ( .A(x[131]), .B(y[783]), .Z(n12886) );
  AND U13205 ( .A(y[773]), .B(x[141]), .Z(n12885) );
  XNOR U13206 ( .A(n12886), .B(n12885), .Z(n12971) );
  XOR U13207 ( .A(n13042), .B(n12971), .Z(n12949) );
  XOR U13208 ( .A(n12950), .B(n12949), .Z(n12951) );
  XOR U13209 ( .A(n12952), .B(n12951), .Z(n12997) );
  OR U13210 ( .A(n12888), .B(n12887), .Z(n12892) );
  NANDN U13211 ( .A(n12890), .B(n12889), .Z(n12891) );
  AND U13212 ( .A(n12892), .B(n12891), .Z(n12998) );
  XNOR U13213 ( .A(n12997), .B(n12998), .Z(n12999) );
  XNOR U13214 ( .A(n13000), .B(n12999), .Z(n12917) );
  XOR U13215 ( .A(n12918), .B(n12917), .Z(n12920) );
  XOR U13216 ( .A(n12919), .B(n12920), .Z(n12906) );
  XOR U13217 ( .A(n12905), .B(n12906), .Z(n12908) );
  XNOR U13218 ( .A(n12907), .B(n12908), .Z(n12913) );
  XNOR U13219 ( .A(n12914), .B(n12913), .Z(n13018) );
  NANDN U13220 ( .A(n12894), .B(n12893), .Z(n12898) );
  OR U13221 ( .A(n12896), .B(n12895), .Z(n12897) );
  NAND U13222 ( .A(n12898), .B(n12897), .Z(n13016) );
  OR U13223 ( .A(n12900), .B(n12899), .Z(n12904) );
  OR U13224 ( .A(n12902), .B(n12901), .Z(n12903) );
  NAND U13225 ( .A(n12904), .B(n12903), .Z(n13015) );
  XNOR U13226 ( .A(n13016), .B(n13015), .Z(n13017) );
  XNOR U13227 ( .A(n13018), .B(n13017), .Z(n13012) );
  XOR U13228 ( .A(n13011), .B(n13012), .Z(N307) );
  NANDN U13229 ( .A(n12906), .B(n12905), .Z(n12910) );
  NANDN U13230 ( .A(n12908), .B(n12907), .Z(n12909) );
  AND U13231 ( .A(n12910), .B(n12909), .Z(n13027) );
  OR U13232 ( .A(n12912), .B(n12911), .Z(n12916) );
  NAND U13233 ( .A(n12914), .B(n12913), .Z(n12915) );
  AND U13234 ( .A(n12916), .B(n12915), .Z(n13028) );
  XOR U13235 ( .A(n13027), .B(n13028), .Z(n13030) );
  NANDN U13236 ( .A(n12918), .B(n12917), .Z(n12922) );
  NANDN U13237 ( .A(n12920), .B(n12919), .Z(n12921) );
  NAND U13238 ( .A(n12922), .B(n12921), .Z(n13127) );
  OR U13239 ( .A(n12923), .B(n13074), .Z(n12927) );
  OR U13240 ( .A(n12925), .B(n12924), .Z(n12926) );
  AND U13241 ( .A(n12927), .B(n12926), .Z(n13120) );
  AND U13242 ( .A(y[772]), .B(x[137]), .Z(n12928) );
  ANDN U13243 ( .B(y[777]), .A(n165), .Z(n13629) );
  NAND U13244 ( .A(n12928), .B(n13629), .Z(n12932) );
  OR U13245 ( .A(n12930), .B(n12929), .Z(n12931) );
  AND U13246 ( .A(n12932), .B(n12931), .Z(n13063) );
  NAND U13247 ( .A(x[130]), .B(y[785]), .Z(n13045) );
  AND U13248 ( .A(x[141]), .B(y[774]), .Z(n12933) );
  XNOR U13249 ( .A(n12934), .B(n12933), .Z(n13044) );
  XOR U13250 ( .A(n13045), .B(n13044), .Z(n13062) );
  NAND U13251 ( .A(x[129]), .B(y[786]), .Z(n13092) );
  AND U13252 ( .A(y[779]), .B(x[136]), .Z(n12936) );
  NAND U13253 ( .A(x[142]), .B(y[773]), .Z(n12935) );
  XOR U13254 ( .A(n12936), .B(n12935), .Z(n13091) );
  XNOR U13255 ( .A(n13092), .B(n13091), .Z(n13064) );
  XOR U13256 ( .A(n13065), .B(n13064), .Z(n13118) );
  AND U13257 ( .A(y[775]), .B(x[144]), .Z(n12937) );
  NANDN U13258 ( .A(n12938), .B(n12937), .Z(n12942) );
  OR U13259 ( .A(n12940), .B(n12939), .Z(n12941) );
  NAND U13260 ( .A(n12942), .B(n12941), .Z(n13119) );
  XNOR U13261 ( .A(n13118), .B(n13119), .Z(n13121) );
  XOR U13262 ( .A(n13120), .B(n13121), .Z(n13124) );
  NANDN U13263 ( .A(n12944), .B(n12943), .Z(n12948) );
  OR U13264 ( .A(n12946), .B(n12945), .Z(n12947) );
  NAND U13265 ( .A(n12948), .B(n12947), .Z(n13113) );
  OR U13266 ( .A(n12950), .B(n12949), .Z(n12954) );
  NANDN U13267 ( .A(n12952), .B(n12951), .Z(n12953) );
  NAND U13268 ( .A(n12954), .B(n12953), .Z(n13112) );
  XOR U13269 ( .A(n13113), .B(n13112), .Z(n13114) );
  AND U13270 ( .A(y[778]), .B(x[137]), .Z(n12956) );
  NAND U13271 ( .A(x[144]), .B(y[771]), .Z(n12955) );
  XOR U13272 ( .A(n12956), .B(n12955), .Z(n13035) );
  AND U13273 ( .A(y[772]), .B(x[143]), .Z(n13034) );
  XNOR U13274 ( .A(n13035), .B(n13034), .Z(n13068) );
  OR U13275 ( .A(n12958), .B(n12957), .Z(n12962) );
  OR U13276 ( .A(n12960), .B(n12959), .Z(n12961) );
  AND U13277 ( .A(n12962), .B(n12961), .Z(n13069) );
  IV U13278 ( .A(y[785]), .Z(n14329) );
  NOR U13279 ( .A(n161), .B(n14329), .Z(n14231) );
  NAND U13280 ( .A(n14231), .B(n12963), .Z(n12967) );
  OR U13281 ( .A(n12965), .B(n12964), .Z(n12966) );
  AND U13282 ( .A(n12967), .B(n12966), .Z(n13070) );
  XOR U13283 ( .A(n13071), .B(n13070), .Z(n13108) );
  AND U13284 ( .A(y[769]), .B(x[146]), .Z(n13055) );
  XNOR U13285 ( .A(o[147]), .B(n13055), .Z(n13097) );
  AND U13286 ( .A(x[138]), .B(y[777]), .Z(n12969) );
  AND U13287 ( .A(y[770]), .B(x[145]), .Z(n12968) );
  XNOR U13288 ( .A(n12969), .B(n12968), .Z(n13096) );
  XNOR U13289 ( .A(n13097), .B(n13096), .Z(n13103) );
  AND U13290 ( .A(x[141]), .B(y[783]), .Z(n14382) );
  NAND U13291 ( .A(n12970), .B(n14382), .Z(n12973) );
  NANDN U13292 ( .A(n12971), .B(n13042), .Z(n12972) );
  AND U13293 ( .A(n12973), .B(n12972), .Z(n13100) );
  NAND U13294 ( .A(x[131]), .B(y[784]), .Z(n13050) );
  AND U13295 ( .A(y[776]), .B(x[139]), .Z(n12975) );
  NAND U13296 ( .A(x[135]), .B(y[780]), .Z(n12974) );
  XOR U13297 ( .A(n12975), .B(n12974), .Z(n13049) );
  XNOR U13298 ( .A(n13050), .B(n13049), .Z(n13101) );
  XNOR U13299 ( .A(n13100), .B(n13101), .Z(n13102) );
  XOR U13300 ( .A(n13103), .B(n13102), .Z(n13107) );
  NANDN U13301 ( .A(n12977), .B(n12976), .Z(n12981) );
  OR U13302 ( .A(n12979), .B(n12978), .Z(n12980) );
  AND U13303 ( .A(n12981), .B(n12980), .Z(n13059) );
  NAND U13304 ( .A(n12982), .B(o[146]), .Z(n13083) );
  NAND U13305 ( .A(x[147]), .B(y[768]), .Z(n13081) );
  NAND U13306 ( .A(x[128]), .B(y[787]), .Z(n13080) );
  XNOR U13307 ( .A(n13081), .B(n13080), .Z(n13082) );
  XNOR U13308 ( .A(n13083), .B(n13082), .Z(n13057) );
  AND U13309 ( .A(y[783]), .B(x[132]), .Z(n13148) );
  AND U13310 ( .A(y[781]), .B(x[134]), .Z(n12984) );
  AND U13311 ( .A(y[782]), .B(x[133]), .Z(n12983) );
  XNOR U13312 ( .A(n12984), .B(n12983), .Z(n13075) );
  XOR U13313 ( .A(n13148), .B(n13075), .Z(n13056) );
  XOR U13314 ( .A(n13057), .B(n13056), .Z(n13058) );
  XOR U13315 ( .A(n13059), .B(n13058), .Z(n13106) );
  XOR U13316 ( .A(n13107), .B(n13106), .Z(n13109) );
  XNOR U13317 ( .A(n13108), .B(n13109), .Z(n13115) );
  XNOR U13318 ( .A(n13114), .B(n13115), .Z(n13125) );
  XNOR U13319 ( .A(n13124), .B(n13125), .Z(n13126) );
  XNOR U13320 ( .A(n13127), .B(n13126), .Z(n13132) );
  NANDN U13321 ( .A(n12986), .B(n12985), .Z(n12990) );
  NANDN U13322 ( .A(n12988), .B(n12987), .Z(n12989) );
  NAND U13323 ( .A(n12990), .B(n12989), .Z(n13131) );
  OR U13324 ( .A(n12992), .B(n12991), .Z(n12996) );
  NANDN U13325 ( .A(n12994), .B(n12993), .Z(n12995) );
  AND U13326 ( .A(n12996), .B(n12995), .Z(n13139) );
  NANDN U13327 ( .A(n12998), .B(n12997), .Z(n13002) );
  NANDN U13328 ( .A(n13000), .B(n12999), .Z(n13001) );
  AND U13329 ( .A(n13002), .B(n13001), .Z(n13136) );
  NANDN U13330 ( .A(n13004), .B(n13003), .Z(n13008) );
  NANDN U13331 ( .A(n13006), .B(n13005), .Z(n13007) );
  NAND U13332 ( .A(n13008), .B(n13007), .Z(n13137) );
  XNOR U13333 ( .A(n13136), .B(n13137), .Z(n13138) );
  XOR U13334 ( .A(n13139), .B(n13138), .Z(n13130) );
  XOR U13335 ( .A(n13131), .B(n13130), .Z(n13133) );
  XNOR U13336 ( .A(n13132), .B(n13133), .Z(n13029) );
  XNOR U13337 ( .A(n13030), .B(n13029), .Z(n13024) );
  NANDN U13338 ( .A(n13010), .B(n13009), .Z(n13014) );
  NANDN U13339 ( .A(n13012), .B(n13011), .Z(n13013) );
  NAND U13340 ( .A(n13014), .B(n13013), .Z(n13021) );
  OR U13341 ( .A(n13016), .B(n13015), .Z(n13020) );
  OR U13342 ( .A(n13018), .B(n13017), .Z(n13019) );
  AND U13343 ( .A(n13020), .B(n13019), .Z(n13022) );
  XNOR U13344 ( .A(n13021), .B(n13022), .Z(n13023) );
  XOR U13345 ( .A(n13024), .B(n13023), .Z(N308) );
  NANDN U13346 ( .A(n13022), .B(n13021), .Z(n13026) );
  NANDN U13347 ( .A(n13024), .B(n13023), .Z(n13025) );
  NAND U13348 ( .A(n13026), .B(n13025), .Z(n13247) );
  OR U13349 ( .A(n13028), .B(n13027), .Z(n13032) );
  NAND U13350 ( .A(n13030), .B(n13029), .Z(n13031) );
  AND U13351 ( .A(n13032), .B(n13031), .Z(n13248) );
  XNOR U13352 ( .A(n13247), .B(n13248), .Z(n13249) );
  AND U13353 ( .A(y[778]), .B(x[144]), .Z(n13983) );
  NANDN U13354 ( .A(n13033), .B(n13983), .Z(n13037) );
  NANDN U13355 ( .A(n13035), .B(n13034), .Z(n13036) );
  AND U13356 ( .A(n13037), .B(n13036), .Z(n13184) );
  AND U13357 ( .A(y[773]), .B(x[143]), .Z(n13039) );
  NAND U13358 ( .A(x[137]), .B(y[779]), .Z(n13038) );
  XOR U13359 ( .A(n13039), .B(n13038), .Z(n13203) );
  AND U13360 ( .A(x[142]), .B(y[774]), .Z(n13202) );
  XNOR U13361 ( .A(n13203), .B(n13202), .Z(n13171) );
  NAND U13362 ( .A(x[130]), .B(y[786]), .Z(n13162) );
  AND U13363 ( .A(y[778]), .B(x[138]), .Z(n13041) );
  NAND U13364 ( .A(x[144]), .B(y[772]), .Z(n13040) );
  XOR U13365 ( .A(n13041), .B(n13040), .Z(n13161) );
  XNOR U13366 ( .A(n13162), .B(n13161), .Z(n13172) );
  XOR U13367 ( .A(n13171), .B(n13172), .Z(n13174) );
  AND U13368 ( .A(y[775]), .B(x[141]), .Z(n13043) );
  NAND U13369 ( .A(n13043), .B(n13042), .Z(n13047) );
  OR U13370 ( .A(n13045), .B(n13044), .Z(n13046) );
  AND U13371 ( .A(n13047), .B(n13046), .Z(n13173) );
  XOR U13372 ( .A(n13174), .B(n13173), .Z(n13183) );
  ANDN U13373 ( .B(y[780]), .A(n162), .Z(n13595) );
  NAND U13374 ( .A(n13595), .B(n13048), .Z(n13052) );
  OR U13375 ( .A(n13050), .B(n13049), .Z(n13051) );
  AND U13376 ( .A(n13052), .B(n13051), .Z(n13180) );
  AND U13377 ( .A(y[769]), .B(x[147]), .Z(n13206) );
  XNOR U13378 ( .A(o[148]), .B(n13206), .Z(n13214) );
  AND U13379 ( .A(x[139]), .B(y[777]), .Z(n13054) );
  AND U13380 ( .A(y[787]), .B(x[129]), .Z(n13053) );
  XNOR U13381 ( .A(n13054), .B(n13053), .Z(n13213) );
  XNOR U13382 ( .A(n13214), .B(n13213), .Z(n13178) );
  NAND U13383 ( .A(o[147]), .B(n13055), .Z(n13145) );
  NAND U13384 ( .A(x[148]), .B(y[768]), .Z(n13143) );
  NAND U13385 ( .A(x[128]), .B(y[788]), .Z(n13142) );
  XNOR U13386 ( .A(n13143), .B(n13142), .Z(n13144) );
  XNOR U13387 ( .A(n13145), .B(n13144), .Z(n13177) );
  XOR U13388 ( .A(n13178), .B(n13177), .Z(n13179) );
  XOR U13389 ( .A(n13180), .B(n13179), .Z(n13185) );
  XOR U13390 ( .A(n13186), .B(n13185), .Z(n13232) );
  OR U13391 ( .A(n13057), .B(n13056), .Z(n13061) );
  NANDN U13392 ( .A(n13059), .B(n13058), .Z(n13060) );
  NAND U13393 ( .A(n13061), .B(n13060), .Z(n13230) );
  NANDN U13394 ( .A(n13063), .B(n13062), .Z(n13067) );
  OR U13395 ( .A(n13065), .B(n13064), .Z(n13066) );
  NAND U13396 ( .A(n13067), .B(n13066), .Z(n13229) );
  XOR U13397 ( .A(n13230), .B(n13229), .Z(n13231) );
  XOR U13398 ( .A(n13232), .B(n13231), .Z(n13192) );
  NANDN U13399 ( .A(n13069), .B(n13068), .Z(n13073) );
  OR U13400 ( .A(n13071), .B(n13070), .Z(n13072) );
  NAND U13401 ( .A(n13073), .B(n13072), .Z(n13198) );
  ANDN U13402 ( .B(y[782]), .A(n157), .Z(n13217) );
  NAND U13403 ( .A(n13217), .B(n13074), .Z(n13077) );
  NANDN U13404 ( .A(n13075), .B(n13148), .Z(n13076) );
  AND U13405 ( .A(n13077), .B(n13076), .Z(n13224) );
  NAND U13406 ( .A(x[145]), .B(y[771]), .Z(n13209) );
  AND U13407 ( .A(y[776]), .B(x[140]), .Z(n13079) );
  AND U13408 ( .A(y[770]), .B(x[146]), .Z(n13078) );
  XNOR U13409 ( .A(n13079), .B(n13078), .Z(n13208) );
  XOR U13410 ( .A(n13209), .B(n13208), .Z(n13223) );
  OR U13411 ( .A(n13081), .B(n13080), .Z(n13085) );
  OR U13412 ( .A(n13083), .B(n13082), .Z(n13084) );
  AND U13413 ( .A(n13085), .B(n13084), .Z(n13225) );
  XNOR U13414 ( .A(n13226), .B(n13225), .Z(n13195) );
  NAND U13415 ( .A(x[135]), .B(y[781]), .Z(n13150) );
  AND U13416 ( .A(x[133]), .B(y[783]), .Z(n13087) );
  NAND U13417 ( .A(x[132]), .B(y[784]), .Z(n13086) );
  XOR U13418 ( .A(n13087), .B(n13086), .Z(n13149) );
  XNOR U13419 ( .A(n13150), .B(n13149), .Z(n13218) );
  NAND U13420 ( .A(x[136]), .B(y[780]), .Z(n13157) );
  AND U13421 ( .A(x[131]), .B(y[785]), .Z(n13089) );
  NAND U13422 ( .A(x[141]), .B(y[775]), .Z(n13088) );
  XOR U13423 ( .A(n13089), .B(n13088), .Z(n13156) );
  XNOR U13424 ( .A(n13157), .B(n13156), .Z(n13219) );
  XNOR U13425 ( .A(n13220), .B(n13219), .Z(n13167) );
  AND U13426 ( .A(y[779]), .B(x[142]), .Z(n13853) );
  NAND U13427 ( .A(n13853), .B(n13090), .Z(n13094) );
  OR U13428 ( .A(n13092), .B(n13091), .Z(n13093) );
  NAND U13429 ( .A(n13094), .B(n13093), .Z(n13166) );
  AND U13430 ( .A(x[145]), .B(y[777]), .Z(n13998) );
  NANDN U13431 ( .A(n13095), .B(n13998), .Z(n13099) );
  OR U13432 ( .A(n13097), .B(n13096), .Z(n13098) );
  NAND U13433 ( .A(n13099), .B(n13098), .Z(n13165) );
  XNOR U13434 ( .A(n13166), .B(n13165), .Z(n13168) );
  XNOR U13435 ( .A(n13167), .B(n13168), .Z(n13196) );
  XOR U13436 ( .A(n13198), .B(n13197), .Z(n13190) );
  OR U13437 ( .A(n13101), .B(n13100), .Z(n13105) );
  OR U13438 ( .A(n13103), .B(n13102), .Z(n13104) );
  NAND U13439 ( .A(n13105), .B(n13104), .Z(n13189) );
  XNOR U13440 ( .A(n13190), .B(n13189), .Z(n13191) );
  XNOR U13441 ( .A(n13192), .B(n13191), .Z(n13236) );
  NANDN U13442 ( .A(n13107), .B(n13106), .Z(n13111) );
  OR U13443 ( .A(n13109), .B(n13108), .Z(n13110) );
  NAND U13444 ( .A(n13111), .B(n13110), .Z(n13242) );
  OR U13445 ( .A(n13113), .B(n13112), .Z(n13117) );
  NANDN U13446 ( .A(n13115), .B(n13114), .Z(n13116) );
  NAND U13447 ( .A(n13117), .B(n13116), .Z(n13241) );
  XOR U13448 ( .A(n13242), .B(n13241), .Z(n13243) );
  OR U13449 ( .A(n13119), .B(n13118), .Z(n13123) );
  OR U13450 ( .A(n13121), .B(n13120), .Z(n13122) );
  NAND U13451 ( .A(n13123), .B(n13122), .Z(n13244) );
  XNOR U13452 ( .A(n13243), .B(n13244), .Z(n13235) );
  XNOR U13453 ( .A(n13236), .B(n13235), .Z(n13238) );
  OR U13454 ( .A(n13125), .B(n13124), .Z(n13129) );
  OR U13455 ( .A(n13127), .B(n13126), .Z(n13128) );
  NAND U13456 ( .A(n13129), .B(n13128), .Z(n13237) );
  XNOR U13457 ( .A(n13238), .B(n13237), .Z(n13253) );
  NANDN U13458 ( .A(n13131), .B(n13130), .Z(n13135) );
  NANDN U13459 ( .A(n13133), .B(n13132), .Z(n13134) );
  NAND U13460 ( .A(n13135), .B(n13134), .Z(n13254) );
  XOR U13461 ( .A(n13253), .B(n13254), .Z(n13256) );
  OR U13462 ( .A(n13137), .B(n13136), .Z(n13141) );
  OR U13463 ( .A(n13139), .B(n13138), .Z(n13140) );
  NAND U13464 ( .A(n13141), .B(n13140), .Z(n13255) );
  XOR U13465 ( .A(n13256), .B(n13255), .Z(n13250) );
  XOR U13466 ( .A(n13249), .B(n13250), .Z(N309) );
  OR U13467 ( .A(n13143), .B(n13142), .Z(n13147) );
  OR U13468 ( .A(n13145), .B(n13144), .Z(n13146) );
  AND U13469 ( .A(n13147), .B(n13146), .Z(n13295) );
  ANDN U13470 ( .B(y[784]), .A(n156), .Z(n13353) );
  NAND U13471 ( .A(n13148), .B(n13353), .Z(n13152) );
  OR U13472 ( .A(n13150), .B(n13149), .Z(n13151) );
  AND U13473 ( .A(n13152), .B(n13151), .Z(n13296) );
  XOR U13474 ( .A(n13295), .B(n13296), .Z(n13297) );
  ANDN U13475 ( .B(y[783]), .A(n157), .Z(n13333) );
  ANDN U13476 ( .B(y[782]), .A(n158), .Z(n13415) );
  ANDN U13477 ( .B(y[775]), .A(n165), .Z(n13332) );
  XNOR U13478 ( .A(n13415), .B(n13332), .Z(n13334) );
  XNOR U13479 ( .A(n13333), .B(n13334), .Z(n13316) );
  NAND U13480 ( .A(y[781]), .B(x[136]), .Z(n13313) );
  XOR U13481 ( .A(n13314), .B(n13313), .Z(n13315) );
  XNOR U13482 ( .A(n13316), .B(n13315), .Z(n13374) );
  NAND U13483 ( .A(x[132]), .B(y[785]), .Z(n13362) );
  AND U13484 ( .A(y[786]), .B(x[131]), .Z(n13154) );
  AND U13485 ( .A(y[776]), .B(x[141]), .Z(n13153) );
  XNOR U13486 ( .A(n13154), .B(n13153), .Z(n13361) );
  XOR U13487 ( .A(n13362), .B(n13361), .Z(n13371) );
  NAND U13488 ( .A(y[777]), .B(x[140]), .Z(n13321) );
  ANDN U13489 ( .B(y[787]), .A(n153), .Z(n13320) );
  NAND U13490 ( .A(x[145]), .B(y[772]), .Z(n13319) );
  XOR U13491 ( .A(n13320), .B(n13319), .Z(n13322) );
  XNOR U13492 ( .A(n13321), .B(n13322), .Z(n13372) );
  XNOR U13493 ( .A(n13374), .B(n13373), .Z(n13298) );
  AND U13494 ( .A(y[778]), .B(x[139]), .Z(n13715) );
  NAND U13495 ( .A(x[148]), .B(y[769]), .Z(n13359) );
  XOR U13496 ( .A(o[149]), .B(n13359), .Z(n13328) );
  NAND U13497 ( .A(x[147]), .B(y[770]), .Z(n13327) );
  XNOR U13498 ( .A(n13328), .B(n13327), .Z(n13329) );
  ANDN U13499 ( .B(y[788]), .A(n152), .Z(n13345) );
  ANDN U13500 ( .B(y[771]), .A(n169), .Z(n13346) );
  XNOR U13501 ( .A(n13345), .B(n13346), .Z(n13348) );
  XOR U13502 ( .A(n13347), .B(n13348), .Z(n13301) );
  XNOR U13503 ( .A(n13302), .B(n13301), .Z(n13304) );
  AND U13504 ( .A(x[141]), .B(y[785]), .Z(n14489) );
  NAND U13505 ( .A(n14489), .B(n13155), .Z(n13159) );
  OR U13506 ( .A(n13157), .B(n13156), .Z(n13158) );
  AND U13507 ( .A(n13159), .B(n13158), .Z(n13303) );
  XOR U13508 ( .A(n13304), .B(n13303), .Z(n13307) );
  NAND U13509 ( .A(n13983), .B(n13160), .Z(n13164) );
  OR U13510 ( .A(n13162), .B(n13161), .Z(n13163) );
  NAND U13511 ( .A(n13164), .B(n13163), .Z(n13308) );
  XNOR U13512 ( .A(n13307), .B(n13308), .Z(n13310) );
  XNOR U13513 ( .A(n13309), .B(n13310), .Z(n13272) );
  OR U13514 ( .A(n13166), .B(n13165), .Z(n13170) );
  NANDN U13515 ( .A(n13168), .B(n13167), .Z(n13169) );
  AND U13516 ( .A(n13170), .B(n13169), .Z(n13277) );
  NANDN U13517 ( .A(n13172), .B(n13171), .Z(n13176) );
  OR U13518 ( .A(n13174), .B(n13173), .Z(n13175) );
  NAND U13519 ( .A(n13176), .B(n13175), .Z(n13278) );
  XOR U13520 ( .A(n13277), .B(n13278), .Z(n13279) );
  OR U13521 ( .A(n13178), .B(n13177), .Z(n13182) );
  NANDN U13522 ( .A(n13180), .B(n13179), .Z(n13181) );
  NAND U13523 ( .A(n13182), .B(n13181), .Z(n13280) );
  XOR U13524 ( .A(n13272), .B(n13271), .Z(n13274) );
  NANDN U13525 ( .A(n13184), .B(n13183), .Z(n13188) );
  OR U13526 ( .A(n13186), .B(n13185), .Z(n13187) );
  NAND U13527 ( .A(n13188), .B(n13187), .Z(n13273) );
  XOR U13528 ( .A(n13274), .B(n13273), .Z(n13383) );
  OR U13529 ( .A(n13190), .B(n13189), .Z(n13194) );
  OR U13530 ( .A(n13192), .B(n13191), .Z(n13193) );
  NAND U13531 ( .A(n13194), .B(n13193), .Z(n13384) );
  XNOR U13532 ( .A(n13383), .B(n13384), .Z(n13386) );
  NAND U13533 ( .A(n13196), .B(n13195), .Z(n13200) );
  NANDN U13534 ( .A(n13198), .B(n13197), .Z(n13199) );
  NAND U13535 ( .A(n13200), .B(n13199), .Z(n13378) );
  NAND U13536 ( .A(x[144]), .B(y[773]), .Z(n13354) );
  XOR U13537 ( .A(n13353), .B(n13354), .Z(n13356) );
  NAND U13538 ( .A(y[774]), .B(x[143]), .Z(n13355) );
  XOR U13539 ( .A(n13356), .B(n13355), .Z(n13365) );
  AND U13540 ( .A(y[779]), .B(x[143]), .Z(n13989) );
  NAND U13541 ( .A(n13201), .B(n13989), .Z(n13205) );
  NANDN U13542 ( .A(n13203), .B(n13202), .Z(n13204) );
  NAND U13543 ( .A(n13205), .B(n13204), .Z(n13366) );
  XNOR U13544 ( .A(n13365), .B(n13366), .Z(n13368) );
  NAND U13545 ( .A(x[128]), .B(y[789]), .Z(n13342) );
  AND U13546 ( .A(n13206), .B(o[148]), .Z(n13340) );
  NAND U13547 ( .A(x[149]), .B(y[768]), .Z(n13339) );
  XNOR U13548 ( .A(n13340), .B(n13339), .Z(n13341) );
  XNOR U13549 ( .A(n13342), .B(n13341), .Z(n13367) );
  XNOR U13550 ( .A(n13368), .B(n13367), .Z(n13289) );
  AND U13551 ( .A(y[776]), .B(x[146]), .Z(n13995) );
  NAND U13552 ( .A(n13207), .B(n13995), .Z(n13211) );
  OR U13553 ( .A(n13209), .B(n13208), .Z(n13210) );
  AND U13554 ( .A(n13211), .B(n13210), .Z(n13290) );
  XOR U13555 ( .A(n13289), .B(n13290), .Z(n13292) );
  ANDN U13556 ( .B(y[787]), .A(n162), .Z(n14701) );
  NAND U13557 ( .A(n13212), .B(n14701), .Z(n13216) );
  OR U13558 ( .A(n13214), .B(n13213), .Z(n13215) );
  AND U13559 ( .A(n13216), .B(n13215), .Z(n13291) );
  XOR U13560 ( .A(n13292), .B(n13291), .Z(n13283) );
  NANDN U13561 ( .A(n13218), .B(n13217), .Z(n13222) );
  OR U13562 ( .A(n13220), .B(n13219), .Z(n13221) );
  AND U13563 ( .A(n13222), .B(n13221), .Z(n13284) );
  NANDN U13564 ( .A(n13224), .B(n13223), .Z(n13228) );
  OR U13565 ( .A(n13226), .B(n13225), .Z(n13227) );
  AND U13566 ( .A(n13228), .B(n13227), .Z(n13285) );
  XOR U13567 ( .A(n13286), .B(n13285), .Z(n13377) );
  XOR U13568 ( .A(n13378), .B(n13377), .Z(n13380) );
  OR U13569 ( .A(n13230), .B(n13229), .Z(n13234) );
  NANDN U13570 ( .A(n13232), .B(n13231), .Z(n13233) );
  NAND U13571 ( .A(n13234), .B(n13233), .Z(n13379) );
  XNOR U13572 ( .A(n13380), .B(n13379), .Z(n13385) );
  XNOR U13573 ( .A(n13386), .B(n13385), .Z(n13267) );
  OR U13574 ( .A(n13236), .B(n13235), .Z(n13240) );
  OR U13575 ( .A(n13238), .B(n13237), .Z(n13239) );
  AND U13576 ( .A(n13240), .B(n13239), .Z(n13265) );
  OR U13577 ( .A(n13242), .B(n13241), .Z(n13246) );
  NANDN U13578 ( .A(n13244), .B(n13243), .Z(n13245) );
  NAND U13579 ( .A(n13246), .B(n13245), .Z(n13266) );
  XOR U13580 ( .A(n13265), .B(n13266), .Z(n13268) );
  XNOR U13581 ( .A(n13267), .B(n13268), .Z(n13262) );
  NANDN U13582 ( .A(n13248), .B(n13247), .Z(n13252) );
  NANDN U13583 ( .A(n13250), .B(n13249), .Z(n13251) );
  NAND U13584 ( .A(n13252), .B(n13251), .Z(n13259) );
  NANDN U13585 ( .A(n13254), .B(n13253), .Z(n13258) );
  OR U13586 ( .A(n13256), .B(n13255), .Z(n13257) );
  NAND U13587 ( .A(n13258), .B(n13257), .Z(n13260) );
  XNOR U13588 ( .A(n13259), .B(n13260), .Z(n13261) );
  XOR U13589 ( .A(n13262), .B(n13261), .Z(N310) );
  NANDN U13590 ( .A(n13260), .B(n13259), .Z(n13264) );
  NANDN U13591 ( .A(n13262), .B(n13261), .Z(n13263) );
  NAND U13592 ( .A(n13264), .B(n13263), .Z(n13389) );
  OR U13593 ( .A(n13266), .B(n13265), .Z(n13270) );
  NAND U13594 ( .A(n13268), .B(n13267), .Z(n13269) );
  AND U13595 ( .A(n13270), .B(n13269), .Z(n13390) );
  XNOR U13596 ( .A(n13389), .B(n13390), .Z(n13391) );
  NANDN U13597 ( .A(n13272), .B(n13271), .Z(n13276) );
  OR U13598 ( .A(n13274), .B(n13273), .Z(n13275) );
  AND U13599 ( .A(n13276), .B(n13275), .Z(n13518) );
  OR U13600 ( .A(n13278), .B(n13277), .Z(n13282) );
  NANDN U13601 ( .A(n13280), .B(n13279), .Z(n13281) );
  AND U13602 ( .A(n13282), .B(n13281), .Z(n13519) );
  XOR U13603 ( .A(n13518), .B(n13519), .Z(n13520) );
  NANDN U13604 ( .A(n13284), .B(n13283), .Z(n13288) );
  OR U13605 ( .A(n13286), .B(n13285), .Z(n13287) );
  NAND U13606 ( .A(n13288), .B(n13287), .Z(n13402) );
  NANDN U13607 ( .A(n13290), .B(n13289), .Z(n13294) );
  OR U13608 ( .A(n13292), .B(n13291), .Z(n13293) );
  NAND U13609 ( .A(n13294), .B(n13293), .Z(n13491) );
  OR U13610 ( .A(n13296), .B(n13295), .Z(n13300) );
  NANDN U13611 ( .A(n13298), .B(n13297), .Z(n13299) );
  NAND U13612 ( .A(n13300), .B(n13299), .Z(n13489) );
  OR U13613 ( .A(n13302), .B(n13301), .Z(n13306) );
  OR U13614 ( .A(n13304), .B(n13303), .Z(n13305) );
  NAND U13615 ( .A(n13306), .B(n13305), .Z(n13488) );
  XOR U13616 ( .A(n13489), .B(n13488), .Z(n13490) );
  XOR U13617 ( .A(n13402), .B(n13401), .Z(n13404) );
  OR U13618 ( .A(n13308), .B(n13307), .Z(n13312) );
  OR U13619 ( .A(n13310), .B(n13309), .Z(n13311) );
  NAND U13620 ( .A(n13312), .B(n13311), .Z(n13497) );
  NANDN U13621 ( .A(n13314), .B(n13313), .Z(n13318) );
  OR U13622 ( .A(n13316), .B(n13315), .Z(n13317) );
  AND U13623 ( .A(n13318), .B(n13317), .Z(n13514) );
  NANDN U13624 ( .A(n13320), .B(n13319), .Z(n13324) );
  NANDN U13625 ( .A(n13322), .B(n13321), .Z(n13323) );
  NAND U13626 ( .A(n13324), .B(n13323), .Z(n13471) );
  AND U13627 ( .A(y[778]), .B(x[140]), .Z(n13326) );
  NAND U13628 ( .A(x[146]), .B(y[772]), .Z(n13325) );
  XOR U13629 ( .A(n13326), .B(n13325), .Z(n13423) );
  NAND U13630 ( .A(x[132]), .B(y[786]), .Z(n13422) );
  XOR U13631 ( .A(n13423), .B(n13422), .Z(n13468) );
  NAND U13632 ( .A(x[133]), .B(y[785]), .Z(n13439) );
  NAND U13633 ( .A(x[145]), .B(y[773]), .Z(n13438) );
  XOR U13634 ( .A(n13439), .B(n13438), .Z(n13440) );
  NAND U13635 ( .A(y[774]), .B(x[144]), .Z(n13441) );
  XOR U13636 ( .A(n13440), .B(n13441), .Z(n13469) );
  XOR U13637 ( .A(n13471), .B(n13470), .Z(n13512) );
  OR U13638 ( .A(n13328), .B(n13327), .Z(n13331) );
  NANDN U13639 ( .A(n13329), .B(n13715), .Z(n13330) );
  NAND U13640 ( .A(n13331), .B(n13330), .Z(n13513) );
  XNOR U13641 ( .A(n13512), .B(n13513), .Z(n13515) );
  XOR U13642 ( .A(n13514), .B(n13515), .Z(n13494) );
  OR U13643 ( .A(n13332), .B(n13415), .Z(n13336) );
  OR U13644 ( .A(n13334), .B(n13333), .Z(n13335) );
  NAND U13645 ( .A(n13336), .B(n13335), .Z(n13453) );
  AND U13646 ( .A(y[782]), .B(x[136]), .Z(n13338) );
  NAND U13647 ( .A(x[135]), .B(y[783]), .Z(n13337) );
  XNOR U13648 ( .A(n13338), .B(n13337), .Z(n13418) );
  NAND U13649 ( .A(x[128]), .B(y[790]), .Z(n13427) );
  NAND U13650 ( .A(x[150]), .B(y[768]), .Z(n13426) );
  XOR U13651 ( .A(n13427), .B(n13426), .Z(n13428) );
  NAND U13652 ( .A(x[149]), .B(y[769]), .Z(n13444) );
  XOR U13653 ( .A(o[150]), .B(n13444), .Z(n13429) );
  XOR U13654 ( .A(n13428), .B(n13429), .Z(n13451) );
  XOR U13655 ( .A(n13450), .B(n13451), .Z(n13452) );
  XOR U13656 ( .A(n13453), .B(n13452), .Z(n13465) );
  NANDN U13657 ( .A(n13340), .B(n13339), .Z(n13344) );
  NAND U13658 ( .A(n13342), .B(n13341), .Z(n13343) );
  AND U13659 ( .A(n13344), .B(n13343), .Z(n13462) );
  OR U13660 ( .A(n13346), .B(n13345), .Z(n13350) );
  OR U13661 ( .A(n13348), .B(n13347), .Z(n13349) );
  AND U13662 ( .A(n13350), .B(n13349), .Z(n13463) );
  XOR U13663 ( .A(n13462), .B(n13463), .Z(n13464) );
  NAND U13664 ( .A(x[130]), .B(y[788]), .Z(n13433) );
  NAND U13665 ( .A(x[148]), .B(y[770]), .Z(n13432) );
  XOR U13666 ( .A(n13433), .B(n13432), .Z(n13434) );
  NAND U13667 ( .A(x[141]), .B(y[777]), .Z(n13435) );
  XOR U13668 ( .A(n13434), .B(n13435), .Z(n13410) );
  AND U13669 ( .A(y[775]), .B(x[143]), .Z(n13352) );
  NAND U13670 ( .A(x[138]), .B(y[780]), .Z(n13351) );
  XOR U13671 ( .A(n13352), .B(n13351), .Z(n13447) );
  NAND U13672 ( .A(x[134]), .B(y[784]), .Z(n13446) );
  XNOR U13673 ( .A(n13447), .B(n13446), .Z(n13407) );
  NANDN U13674 ( .A(n13354), .B(n13353), .Z(n13358) );
  OR U13675 ( .A(n13356), .B(n13355), .Z(n13357) );
  NAND U13676 ( .A(n13358), .B(n13357), .Z(n13408) );
  XOR U13677 ( .A(n13410), .B(n13409), .Z(n13506) );
  NAND U13678 ( .A(x[142]), .B(y[776]), .Z(n13483) );
  NAND U13679 ( .A(x[131]), .B(y[787]), .Z(n13482) );
  XOR U13680 ( .A(n13483), .B(n13482), .Z(n13484) );
  NAND U13681 ( .A(y[771]), .B(x[147]), .Z(n13485) );
  XOR U13682 ( .A(n13484), .B(n13485), .Z(n13457) );
  NANDN U13683 ( .A(n13359), .B(o[149]), .Z(n13479) );
  NAND U13684 ( .A(x[129]), .B(y[789]), .Z(n13477) );
  XOR U13685 ( .A(n13476), .B(n13477), .Z(n13478) );
  XNOR U13686 ( .A(n13479), .B(n13478), .Z(n13456) );
  XNOR U13687 ( .A(n13457), .B(n13456), .Z(n13459) );
  ANDN U13688 ( .B(y[786]), .A(n164), .Z(n14746) );
  NAND U13689 ( .A(n13360), .B(n14746), .Z(n13364) );
  OR U13690 ( .A(n13362), .B(n13361), .Z(n13363) );
  AND U13691 ( .A(n13364), .B(n13363), .Z(n13458) );
  XNOR U13692 ( .A(n13459), .B(n13458), .Z(n13507) );
  XNOR U13693 ( .A(n13506), .B(n13507), .Z(n13509) );
  XNOR U13694 ( .A(n13508), .B(n13509), .Z(n13502) );
  OR U13695 ( .A(n13366), .B(n13365), .Z(n13370) );
  OR U13696 ( .A(n13368), .B(n13367), .Z(n13369) );
  AND U13697 ( .A(n13370), .B(n13369), .Z(n13500) );
  NANDN U13698 ( .A(n13372), .B(n13371), .Z(n13376) );
  NAND U13699 ( .A(n13374), .B(n13373), .Z(n13375) );
  NAND U13700 ( .A(n13376), .B(n13375), .Z(n13501) );
  XNOR U13701 ( .A(n13500), .B(n13501), .Z(n13503) );
  XNOR U13702 ( .A(n13502), .B(n13503), .Z(n13495) );
  XNOR U13703 ( .A(n13494), .B(n13495), .Z(n13496) );
  XOR U13704 ( .A(n13497), .B(n13496), .Z(n13403) );
  XNOR U13705 ( .A(n13404), .B(n13403), .Z(n13521) );
  XOR U13706 ( .A(n13520), .B(n13521), .Z(n13398) );
  NANDN U13707 ( .A(n13378), .B(n13377), .Z(n13382) );
  OR U13708 ( .A(n13380), .B(n13379), .Z(n13381) );
  NAND U13709 ( .A(n13382), .B(n13381), .Z(n13396) );
  OR U13710 ( .A(n13384), .B(n13383), .Z(n13388) );
  OR U13711 ( .A(n13386), .B(n13385), .Z(n13387) );
  NAND U13712 ( .A(n13388), .B(n13387), .Z(n13395) );
  XNOR U13713 ( .A(n13396), .B(n13395), .Z(n13397) );
  XNOR U13714 ( .A(n13398), .B(n13397), .Z(n13392) );
  XOR U13715 ( .A(n13391), .B(n13392), .Z(N311) );
  NANDN U13716 ( .A(n13390), .B(n13389), .Z(n13394) );
  NANDN U13717 ( .A(n13392), .B(n13391), .Z(n13393) );
  NAND U13718 ( .A(n13394), .B(n13393), .Z(n13524) );
  OR U13719 ( .A(n13396), .B(n13395), .Z(n13400) );
  OR U13720 ( .A(n13398), .B(n13397), .Z(n13399) );
  AND U13721 ( .A(n13400), .B(n13399), .Z(n13525) );
  XNOR U13722 ( .A(n13524), .B(n13525), .Z(n13526) );
  NANDN U13723 ( .A(n13402), .B(n13401), .Z(n13406) );
  OR U13724 ( .A(n13404), .B(n13403), .Z(n13405) );
  AND U13725 ( .A(n13406), .B(n13405), .Z(n13530) );
  NANDN U13726 ( .A(n13408), .B(n13407), .Z(n13412) );
  NAND U13727 ( .A(n13410), .B(n13409), .Z(n13411) );
  NAND U13728 ( .A(n13412), .B(n13411), .Z(n13561) );
  NAND U13729 ( .A(x[128]), .B(y[791]), .Z(n13576) );
  NAND U13730 ( .A(x[151]), .B(y[768]), .Z(n13575) );
  XOR U13731 ( .A(n13576), .B(n13575), .Z(n13578) );
  ANDN U13732 ( .B(y[769]), .A(n173), .Z(n13604) );
  XOR U13733 ( .A(o[151]), .B(n13604), .Z(n13577) );
  AND U13734 ( .A(x[148]), .B(y[771]), .Z(n13414) );
  NAND U13735 ( .A(x[144]), .B(y[775]), .Z(n13413) );
  XOR U13736 ( .A(n13414), .B(n13413), .Z(n13601) );
  NAND U13737 ( .A(x[147]), .B(y[772]), .Z(n13600) );
  XNOR U13738 ( .A(n13601), .B(n13600), .Z(n13659) );
  NANDN U13739 ( .A(n13416), .B(n13415), .Z(n13420) );
  NAND U13740 ( .A(n13418), .B(n13417), .Z(n13419) );
  NAND U13741 ( .A(n13420), .B(n13419), .Z(n13660) );
  AND U13742 ( .A(y[778]), .B(x[146]), .Z(n14368) );
  NAND U13743 ( .A(n14368), .B(n13421), .Z(n13425) );
  OR U13744 ( .A(n13423), .B(n13422), .Z(n13424) );
  NAND U13745 ( .A(n13425), .B(n13424), .Z(n13653) );
  OR U13746 ( .A(n13427), .B(n13426), .Z(n13431) );
  NANDN U13747 ( .A(n13429), .B(n13428), .Z(n13430) );
  AND U13748 ( .A(n13431), .B(n13430), .Z(n13654) );
  XOR U13749 ( .A(n13561), .B(n13560), .Z(n13563) );
  OR U13750 ( .A(n13433), .B(n13432), .Z(n13437) );
  NANDN U13751 ( .A(n13435), .B(n13434), .Z(n13436) );
  NAND U13752 ( .A(n13437), .B(n13436), .Z(n13567) );
  NAND U13753 ( .A(x[141]), .B(y[778]), .Z(n13624) );
  NAND U13754 ( .A(x[130]), .B(y[789]), .Z(n13623) );
  XOR U13755 ( .A(n13624), .B(n13623), .Z(n13625) );
  NAND U13756 ( .A(x[149]), .B(y[770]), .Z(n13626) );
  XOR U13757 ( .A(n13625), .B(n13626), .Z(n13644) );
  OR U13758 ( .A(n13439), .B(n13438), .Z(n13443) );
  NANDN U13759 ( .A(n13441), .B(n13440), .Z(n13442) );
  AND U13760 ( .A(n13443), .B(n13442), .Z(n13641) );
  NANDN U13761 ( .A(n13444), .B(o[150]), .Z(n13584) );
  NAND U13762 ( .A(x[140]), .B(y[779]), .Z(n13582) );
  NAND U13763 ( .A(x[129]), .B(y[790]), .Z(n13581) );
  XOR U13764 ( .A(n13582), .B(n13581), .Z(n13583) );
  XOR U13765 ( .A(n13584), .B(n13583), .Z(n13642) );
  XOR U13766 ( .A(n13641), .B(n13642), .Z(n13643) );
  XNOR U13767 ( .A(n13644), .B(n13643), .Z(n13566) );
  XNOR U13768 ( .A(n13567), .B(n13566), .Z(n13569) );
  AND U13769 ( .A(y[780]), .B(x[143]), .Z(n14225) );
  NAND U13770 ( .A(n13445), .B(n14225), .Z(n13449) );
  OR U13771 ( .A(n13447), .B(n13446), .Z(n13448) );
  AND U13772 ( .A(n13449), .B(n13448), .Z(n13650) );
  NAND U13773 ( .A(y[788]), .B(x[131]), .Z(n13630) );
  XOR U13774 ( .A(n13629), .B(n13630), .Z(n13632) );
  NAND U13775 ( .A(x[132]), .B(y[787]), .Z(n13631) );
  XOR U13776 ( .A(n13632), .B(n13631), .Z(n13648) );
  NAND U13777 ( .A(x[133]), .B(y[786]), .Z(n13618) );
  NAND U13778 ( .A(x[146]), .B(y[773]), .Z(n13617) );
  XOR U13779 ( .A(n13618), .B(n13617), .Z(n13619) );
  NAND U13780 ( .A(y[774]), .B(x[145]), .Z(n13620) );
  XNOR U13781 ( .A(n13619), .B(n13620), .Z(n13647) );
  XNOR U13782 ( .A(n13650), .B(n13649), .Z(n13568) );
  XNOR U13783 ( .A(n13569), .B(n13568), .Z(n13562) );
  XNOR U13784 ( .A(n13563), .B(n13562), .Z(n13548) );
  NANDN U13785 ( .A(n13451), .B(n13450), .Z(n13455) );
  OR U13786 ( .A(n13453), .B(n13452), .Z(n13454) );
  AND U13787 ( .A(n13455), .B(n13454), .Z(n13605) );
  OR U13788 ( .A(n13457), .B(n13456), .Z(n13461) );
  OR U13789 ( .A(n13459), .B(n13458), .Z(n13460) );
  AND U13790 ( .A(n13461), .B(n13460), .Z(n13606) );
  XOR U13791 ( .A(n13605), .B(n13606), .Z(n13607) );
  OR U13792 ( .A(n13463), .B(n13462), .Z(n13467) );
  NANDN U13793 ( .A(n13465), .B(n13464), .Z(n13466) );
  NAND U13794 ( .A(n13467), .B(n13466), .Z(n13608) );
  NANDN U13795 ( .A(n13469), .B(n13468), .Z(n13473) );
  OR U13796 ( .A(n13471), .B(n13470), .Z(n13472) );
  AND U13797 ( .A(n13473), .B(n13472), .Z(n13536) );
  AND U13798 ( .A(x[136]), .B(y[783]), .Z(n13475) );
  NAND U13799 ( .A(x[137]), .B(y[782]), .Z(n13474) );
  XOR U13800 ( .A(n13475), .B(n13474), .Z(n13590) );
  NAND U13801 ( .A(x[135]), .B(y[784]), .Z(n13589) );
  XOR U13802 ( .A(n13590), .B(n13589), .Z(n13635) );
  NAND U13803 ( .A(y[781]), .B(x[138]), .Z(n13636) );
  XNOR U13804 ( .A(n13635), .B(n13636), .Z(n13637) );
  NAND U13805 ( .A(x[134]), .B(y[785]), .Z(n13594) );
  NAND U13806 ( .A(x[143]), .B(y[776]), .Z(n13593) );
  XOR U13807 ( .A(n13594), .B(n13593), .Z(n13596) );
  XNOR U13808 ( .A(n13595), .B(n13596), .Z(n13638) );
  XOR U13809 ( .A(n13637), .B(n13638), .Z(n13614) );
  NANDN U13810 ( .A(n13477), .B(n13476), .Z(n13481) );
  OR U13811 ( .A(n13479), .B(n13478), .Z(n13480) );
  NAND U13812 ( .A(n13481), .B(n13480), .Z(n13612) );
  OR U13813 ( .A(n13483), .B(n13482), .Z(n13487) );
  NANDN U13814 ( .A(n13485), .B(n13484), .Z(n13486) );
  AND U13815 ( .A(n13487), .B(n13486), .Z(n13611) );
  XOR U13816 ( .A(n13614), .B(n13613), .Z(n13537) );
  XOR U13817 ( .A(n13536), .B(n13537), .Z(n13538) );
  XOR U13818 ( .A(n13548), .B(n13549), .Z(n13551) );
  OR U13819 ( .A(n13489), .B(n13488), .Z(n13493) );
  NANDN U13820 ( .A(n13491), .B(n13490), .Z(n13492) );
  NAND U13821 ( .A(n13493), .B(n13492), .Z(n13550) );
  XOR U13822 ( .A(n13551), .B(n13550), .Z(n13556) );
  OR U13823 ( .A(n13495), .B(n13494), .Z(n13499) );
  OR U13824 ( .A(n13497), .B(n13496), .Z(n13498) );
  NAND U13825 ( .A(n13499), .B(n13498), .Z(n13555) );
  OR U13826 ( .A(n13501), .B(n13500), .Z(n13505) );
  NANDN U13827 ( .A(n13503), .B(n13502), .Z(n13504) );
  AND U13828 ( .A(n13505), .B(n13504), .Z(n13544) );
  OR U13829 ( .A(n13507), .B(n13506), .Z(n13511) );
  OR U13830 ( .A(n13509), .B(n13508), .Z(n13510) );
  NAND U13831 ( .A(n13511), .B(n13510), .Z(n13543) );
  OR U13832 ( .A(n13513), .B(n13512), .Z(n13517) );
  OR U13833 ( .A(n13515), .B(n13514), .Z(n13516) );
  AND U13834 ( .A(n13517), .B(n13516), .Z(n13542) );
  XNOR U13835 ( .A(n13543), .B(n13542), .Z(n13545) );
  XNOR U13836 ( .A(n13544), .B(n13545), .Z(n13554) );
  XNOR U13837 ( .A(n13555), .B(n13554), .Z(n13557) );
  XNOR U13838 ( .A(n13556), .B(n13557), .Z(n13531) );
  XOR U13839 ( .A(n13530), .B(n13531), .Z(n13532) );
  OR U13840 ( .A(n13519), .B(n13518), .Z(n13523) );
  NANDN U13841 ( .A(n13521), .B(n13520), .Z(n13522) );
  AND U13842 ( .A(n13523), .B(n13522), .Z(n13533) );
  XOR U13843 ( .A(n13526), .B(n13527), .Z(N312) );
  NANDN U13844 ( .A(n13525), .B(n13524), .Z(n13529) );
  NANDN U13845 ( .A(n13527), .B(n13526), .Z(n13528) );
  NAND U13846 ( .A(n13529), .B(n13528), .Z(n13665) );
  OR U13847 ( .A(n13531), .B(n13530), .Z(n13535) );
  NANDN U13848 ( .A(n13533), .B(n13532), .Z(n13534) );
  AND U13849 ( .A(n13535), .B(n13534), .Z(n13666) );
  XNOR U13850 ( .A(n13665), .B(n13666), .Z(n13667) );
  OR U13851 ( .A(n13537), .B(n13536), .Z(n13541) );
  NANDN U13852 ( .A(n13539), .B(n13538), .Z(n13540) );
  NAND U13853 ( .A(n13541), .B(n13540), .Z(n13800) );
  OR U13854 ( .A(n13543), .B(n13542), .Z(n13547) );
  OR U13855 ( .A(n13545), .B(n13544), .Z(n13546) );
  AND U13856 ( .A(n13547), .B(n13546), .Z(n13799) );
  XOR U13857 ( .A(n13800), .B(n13799), .Z(n13801) );
  NANDN U13858 ( .A(n13549), .B(n13548), .Z(n13553) );
  OR U13859 ( .A(n13551), .B(n13550), .Z(n13552) );
  NAND U13860 ( .A(n13553), .B(n13552), .Z(n13802) );
  OR U13861 ( .A(n13555), .B(n13554), .Z(n13559) );
  OR U13862 ( .A(n13557), .B(n13556), .Z(n13558) );
  AND U13863 ( .A(n13559), .B(n13558), .Z(n13672) );
  NANDN U13864 ( .A(n13561), .B(n13560), .Z(n13565) );
  NANDN U13865 ( .A(n13563), .B(n13562), .Z(n13564) );
  NAND U13866 ( .A(n13565), .B(n13564), .Z(n13680) );
  NAND U13867 ( .A(n13567), .B(n13566), .Z(n13571) );
  NANDN U13868 ( .A(n13569), .B(n13568), .Z(n13570) );
  NAND U13869 ( .A(n13571), .B(n13570), .Z(n13677) );
  AND U13870 ( .A(x[139]), .B(y[781]), .Z(n13573) );
  NAND U13871 ( .A(x[142]), .B(y[778]), .Z(n13572) );
  XOR U13872 ( .A(n13573), .B(n13572), .Z(n13717) );
  ANDN U13873 ( .B(y[784]), .A(n159), .Z(n13716) );
  XNOR U13874 ( .A(n13717), .B(n13716), .Z(n13711) );
  NOR U13875 ( .A(n160), .B(n13574), .Z(n13587) );
  IV U13876 ( .A(n13587), .Z(n13709) );
  NAND U13877 ( .A(x[138]), .B(y[782]), .Z(n13708) );
  XOR U13878 ( .A(n13709), .B(n13708), .Z(n13710) );
  XNOR U13879 ( .A(n13711), .B(n13710), .Z(n13722) );
  OR U13880 ( .A(n13576), .B(n13575), .Z(n13580) );
  NAND U13881 ( .A(n13578), .B(n13577), .Z(n13579) );
  NAND U13882 ( .A(n13580), .B(n13579), .Z(n13720) );
  NAND U13883 ( .A(x[143]), .B(y[777]), .Z(n13727) );
  NAND U13884 ( .A(x[131]), .B(y[789]), .Z(n13726) );
  XOR U13885 ( .A(n13727), .B(n13726), .Z(n13728) );
  NAND U13886 ( .A(y[788]), .B(x[132]), .Z(n13729) );
  XOR U13887 ( .A(n13728), .B(n13729), .Z(n13721) );
  XOR U13888 ( .A(n13722), .B(n13723), .Z(n13740) );
  OR U13889 ( .A(n13582), .B(n13581), .Z(n13586) );
  NANDN U13890 ( .A(n13584), .B(n13583), .Z(n13585) );
  AND U13891 ( .A(n13586), .B(n13585), .Z(n13784) );
  NANDN U13892 ( .A(n13588), .B(n13587), .Z(n13592) );
  OR U13893 ( .A(n13590), .B(n13589), .Z(n13591) );
  AND U13894 ( .A(n13592), .B(n13591), .Z(n13782) );
  NAND U13895 ( .A(x[144]), .B(y[776]), .Z(n13753) );
  NAND U13896 ( .A(x[133]), .B(y[787]), .Z(n13751) );
  NAND U13897 ( .A(x[149]), .B(y[771]), .Z(n13750) );
  XNOR U13898 ( .A(n13751), .B(n13750), .Z(n13752) );
  XNOR U13899 ( .A(n13753), .B(n13752), .Z(n13772) );
  OR U13900 ( .A(n13594), .B(n13593), .Z(n13598) );
  NAND U13901 ( .A(n13596), .B(n13595), .Z(n13597) );
  AND U13902 ( .A(n13598), .B(n13597), .Z(n13769) );
  ANDN U13903 ( .B(y[772]), .A(n171), .Z(n13896) );
  NAND U13904 ( .A(x[147]), .B(y[773]), .Z(n13759) );
  NAND U13905 ( .A(x[134]), .B(y[786]), .Z(n13758) );
  XNOR U13906 ( .A(n13759), .B(n13758), .Z(n13760) );
  XOR U13907 ( .A(n13896), .B(n13760), .Z(n13770) );
  XOR U13908 ( .A(n13769), .B(n13770), .Z(n13771) );
  XNOR U13909 ( .A(n13772), .B(n13771), .Z(n13781) );
  XNOR U13910 ( .A(n13782), .B(n13781), .Z(n13783) );
  XOR U13911 ( .A(n13784), .B(n13783), .Z(n13738) );
  NAND U13912 ( .A(x[130]), .B(y[790]), .Z(n13696) );
  NAND U13913 ( .A(x[150]), .B(y[770]), .Z(n13695) );
  XOR U13914 ( .A(n13696), .B(n13695), .Z(n13698) );
  XNOR U13915 ( .A(n13697), .B(n13698), .Z(n13778) );
  AND U13916 ( .A(y[771]), .B(x[144]), .Z(n13599) );
  ANDN U13917 ( .B(y[775]), .A(n171), .Z(n14159) );
  NAND U13918 ( .A(n13599), .B(n14159), .Z(n13603) );
  OR U13919 ( .A(n13601), .B(n13600), .Z(n13602) );
  AND U13920 ( .A(n13603), .B(n13602), .Z(n13776) );
  NAND U13921 ( .A(n13604), .B(o[151]), .Z(n13692) );
  NAND U13922 ( .A(x[129]), .B(y[791]), .Z(n13690) );
  XOR U13923 ( .A(n13692), .B(n13691), .Z(n13775) );
  XOR U13924 ( .A(n13778), .B(n13777), .Z(n13739) );
  XOR U13925 ( .A(n13738), .B(n13739), .Z(n13741) );
  XOR U13926 ( .A(n13740), .B(n13741), .Z(n13678) );
  XNOR U13927 ( .A(n13680), .B(n13679), .Z(n13808) );
  OR U13928 ( .A(n13606), .B(n13605), .Z(n13610) );
  NANDN U13929 ( .A(n13608), .B(n13607), .Z(n13609) );
  AND U13930 ( .A(n13610), .B(n13609), .Z(n13806) );
  NANDN U13931 ( .A(n13612), .B(n13611), .Z(n13616) );
  NAND U13932 ( .A(n13614), .B(n13613), .Z(n13615) );
  NAND U13933 ( .A(n13616), .B(n13615), .Z(n13685) );
  NAND U13934 ( .A(x[146]), .B(y[774]), .Z(n13705) );
  NAND U13935 ( .A(x[145]), .B(y[775]), .Z(n13703) );
  NAND U13936 ( .A(y[785]), .B(x[135]), .Z(n13702) );
  XOR U13937 ( .A(n13703), .B(n13702), .Z(n13704) );
  XOR U13938 ( .A(n13705), .B(n13704), .Z(n13764) );
  ANDN U13939 ( .B(y[769]), .A(n174), .Z(n13701) );
  XOR U13940 ( .A(o[152]), .B(n13701), .Z(n13734) );
  NAND U13941 ( .A(x[128]), .B(y[792]), .Z(n13733) );
  NAND U13942 ( .A(x[152]), .B(y[768]), .Z(n13732) );
  XOR U13943 ( .A(n13733), .B(n13732), .Z(n13735) );
  XOR U13944 ( .A(n13734), .B(n13735), .Z(n13763) );
  OR U13945 ( .A(n13618), .B(n13617), .Z(n13622) );
  NANDN U13946 ( .A(n13620), .B(n13619), .Z(n13621) );
  AND U13947 ( .A(n13622), .B(n13621), .Z(n13765) );
  XNOR U13948 ( .A(n13766), .B(n13765), .Z(n13790) );
  OR U13949 ( .A(n13624), .B(n13623), .Z(n13628) );
  NANDN U13950 ( .A(n13626), .B(n13625), .Z(n13627) );
  AND U13951 ( .A(n13628), .B(n13627), .Z(n13787) );
  NANDN U13952 ( .A(n13630), .B(n13629), .Z(n13634) );
  OR U13953 ( .A(n13632), .B(n13631), .Z(n13633) );
  AND U13954 ( .A(n13634), .B(n13633), .Z(n13788) );
  XOR U13955 ( .A(n13787), .B(n13788), .Z(n13789) );
  XNOR U13956 ( .A(n13790), .B(n13789), .Z(n13683) );
  NANDN U13957 ( .A(n13636), .B(n13635), .Z(n13640) );
  NANDN U13958 ( .A(n13638), .B(n13637), .Z(n13639) );
  NAND U13959 ( .A(n13640), .B(n13639), .Z(n13684) );
  XNOR U13960 ( .A(n13683), .B(n13684), .Z(n13686) );
  XOR U13961 ( .A(n13685), .B(n13686), .Z(n13796) );
  OR U13962 ( .A(n13642), .B(n13641), .Z(n13646) );
  NANDN U13963 ( .A(n13644), .B(n13643), .Z(n13645) );
  NAND U13964 ( .A(n13646), .B(n13645), .Z(n13793) );
  NAND U13965 ( .A(n13648), .B(n13647), .Z(n13652) );
  NANDN U13966 ( .A(n13650), .B(n13649), .Z(n13651) );
  NAND U13967 ( .A(n13652), .B(n13651), .Z(n13747) );
  NANDN U13968 ( .A(n13654), .B(n13653), .Z(n13658) );
  NAND U13969 ( .A(n13656), .B(n13655), .Z(n13657) );
  NAND U13970 ( .A(n13658), .B(n13657), .Z(n13744) );
  NANDN U13971 ( .A(n13660), .B(n13659), .Z(n13664) );
  NANDN U13972 ( .A(n13662), .B(n13661), .Z(n13663) );
  NAND U13973 ( .A(n13664), .B(n13663), .Z(n13745) );
  XNOR U13974 ( .A(n13747), .B(n13746), .Z(n13794) );
  XOR U13975 ( .A(n13796), .B(n13795), .Z(n13805) );
  XOR U13976 ( .A(n13806), .B(n13805), .Z(n13807) );
  XNOR U13977 ( .A(n13808), .B(n13807), .Z(n13671) );
  XOR U13978 ( .A(n13672), .B(n13671), .Z(n13673) );
  XNOR U13979 ( .A(n13674), .B(n13673), .Z(n13668) );
  XOR U13980 ( .A(n13667), .B(n13668), .Z(N313) );
  NANDN U13981 ( .A(n13666), .B(n13665), .Z(n13670) );
  NANDN U13982 ( .A(n13668), .B(n13667), .Z(n13669) );
  NAND U13983 ( .A(n13670), .B(n13669), .Z(n13811) );
  NANDN U13984 ( .A(n13672), .B(n13671), .Z(n13676) );
  OR U13985 ( .A(n13674), .B(n13673), .Z(n13675) );
  AND U13986 ( .A(n13676), .B(n13675), .Z(n13812) );
  XNOR U13987 ( .A(n13811), .B(n13812), .Z(n13813) );
  NANDN U13988 ( .A(n13678), .B(n13677), .Z(n13682) );
  NAND U13989 ( .A(n13680), .B(n13679), .Z(n13681) );
  NAND U13990 ( .A(n13682), .B(n13681), .Z(n13951) );
  OR U13991 ( .A(n13684), .B(n13683), .Z(n13688) );
  NANDN U13992 ( .A(n13686), .B(n13685), .Z(n13687) );
  NAND U13993 ( .A(n13688), .B(n13687), .Z(n13831) );
  NANDN U13994 ( .A(n13690), .B(n13689), .Z(n13694) );
  OR U13995 ( .A(n13692), .B(n13691), .Z(n13693) );
  NAND U13996 ( .A(n13694), .B(n13693), .Z(n13933) );
  OR U13997 ( .A(n13696), .B(n13695), .Z(n13700) );
  NAND U13998 ( .A(n13698), .B(n13697), .Z(n13699) );
  NAND U13999 ( .A(n13700), .B(n13699), .Z(n13932) );
  NANDN U14000 ( .A(n14329), .B(x[136]), .Z(n13927) );
  XNOR U14001 ( .A(n13927), .B(n13928), .Z(n13916) );
  AND U14002 ( .A(n13701), .B(o[152]), .Z(n13922) );
  AND U14003 ( .A(y[768]), .B(x[153]), .Z(n13919) );
  AND U14004 ( .A(y[793]), .B(x[128]), .Z(n13920) );
  XNOR U14005 ( .A(n13919), .B(n13920), .Z(n13921) );
  XNOR U14006 ( .A(n13922), .B(n13921), .Z(n13915) );
  XOR U14007 ( .A(n13916), .B(n13915), .Z(n13918) );
  OR U14008 ( .A(n13703), .B(n13702), .Z(n13707) );
  NANDN U14009 ( .A(n13705), .B(n13704), .Z(n13706) );
  AND U14010 ( .A(n13707), .B(n13706), .Z(n13917) );
  XOR U14011 ( .A(n13918), .B(n13917), .Z(n13931) );
  XNOR U14012 ( .A(n13932), .B(n13931), .Z(n13934) );
  XOR U14013 ( .A(n13933), .B(n13934), .Z(n13939) );
  NAND U14014 ( .A(n13709), .B(n13708), .Z(n13713) );
  NANDN U14015 ( .A(n13711), .B(n13710), .Z(n13712) );
  AND U14016 ( .A(n13713), .B(n13712), .Z(n13937) );
  NANDN U14017 ( .A(n162), .B(y[782]), .Z(n13874) );
  NANDN U14018 ( .A(n13714), .B(x[140]), .Z(n13872) );
  NANDN U14019 ( .A(n158), .B(y[786]), .Z(n13873) );
  XNOR U14020 ( .A(n13872), .B(n13873), .Z(n13875) );
  XNOR U14021 ( .A(n13874), .B(n13875), .Z(n13865) );
  AND U14022 ( .A(x[142]), .B(y[781]), .Z(n14216) );
  NAND U14023 ( .A(n13715), .B(n14216), .Z(n13719) );
  NANDN U14024 ( .A(n13717), .B(n13716), .Z(n13718) );
  AND U14025 ( .A(n13719), .B(n13718), .Z(n13866) );
  XNOR U14026 ( .A(n13865), .B(n13866), .Z(n13868) );
  NAND U14027 ( .A(x[141]), .B(y[780]), .Z(n13860) );
  AND U14028 ( .A(y[792]), .B(x[129]), .Z(n13859) );
  XNOR U14029 ( .A(n13860), .B(n13859), .Z(n13862) );
  ANDN U14030 ( .B(y[769]), .A(n175), .Z(n13871) );
  XOR U14031 ( .A(o[153]), .B(n13871), .Z(n13861) );
  XOR U14032 ( .A(n13868), .B(n13867), .Z(n13938) );
  XNOR U14033 ( .A(n13937), .B(n13938), .Z(n13940) );
  XNOR U14034 ( .A(n13939), .B(n13940), .Z(n13837) );
  NANDN U14035 ( .A(n13721), .B(n13720), .Z(n13725) );
  OR U14036 ( .A(n13723), .B(n13722), .Z(n13724) );
  NAND U14037 ( .A(n13725), .B(n13724), .Z(n13835) );
  OR U14038 ( .A(n13727), .B(n13726), .Z(n13731) );
  NANDN U14039 ( .A(n13729), .B(n13728), .Z(n13730) );
  AND U14040 ( .A(n13731), .B(n13730), .Z(n13913) );
  OR U14041 ( .A(n13733), .B(n13732), .Z(n13737) );
  NAND U14042 ( .A(n13735), .B(n13734), .Z(n13736) );
  AND U14043 ( .A(n13737), .B(n13736), .Z(n13911) );
  NAND U14044 ( .A(x[130]), .B(y[791]), .Z(n13856) );
  NAND U14045 ( .A(x[131]), .B(y[790]), .Z(n13854) );
  XNOR U14046 ( .A(n13853), .B(n13854), .Z(n13855) );
  XOR U14047 ( .A(n13856), .B(n13855), .Z(n13912) );
  XOR U14048 ( .A(n13911), .B(n13912), .Z(n13914) );
  XOR U14049 ( .A(n13913), .B(n13914), .Z(n13836) );
  XOR U14050 ( .A(n13837), .B(n13838), .Z(n13830) );
  NANDN U14051 ( .A(n13739), .B(n13738), .Z(n13743) );
  OR U14052 ( .A(n13741), .B(n13740), .Z(n13742) );
  AND U14053 ( .A(n13743), .B(n13742), .Z(n13829) );
  XNOR U14054 ( .A(n13830), .B(n13829), .Z(n13832) );
  XOR U14055 ( .A(n13831), .B(n13832), .Z(n13949) );
  NANDN U14056 ( .A(n13745), .B(n13744), .Z(n13749) );
  NAND U14057 ( .A(n13747), .B(n13746), .Z(n13748) );
  NAND U14058 ( .A(n13749), .B(n13748), .Z(n13824) );
  OR U14059 ( .A(n13751), .B(n13750), .Z(n13755) );
  OR U14060 ( .A(n13753), .B(n13752), .Z(n13754) );
  AND U14061 ( .A(n13755), .B(n13754), .Z(n13909) );
  ANDN U14062 ( .B(y[771]), .A(n173), .Z(n13880) );
  ANDN U14063 ( .B(y[788]), .A(n156), .Z(n13878) );
  ANDN U14064 ( .B(y[776]), .A(n168), .Z(n13879) );
  XNOR U14065 ( .A(n13878), .B(n13879), .Z(n13881) );
  XOR U14066 ( .A(n13880), .B(n13881), .Z(n13908) );
  NAND U14067 ( .A(x[147]), .B(y[774]), .Z(n13898) );
  AND U14068 ( .A(y[772]), .B(x[149]), .Z(n13757) );
  AND U14069 ( .A(y[773]), .B(x[148]), .Z(n13756) );
  XNOR U14070 ( .A(n13757), .B(n13756), .Z(n13897) );
  XOR U14071 ( .A(n13898), .B(n13897), .Z(n13907) );
  XOR U14072 ( .A(n13908), .B(n13907), .Z(n13910) );
  XOR U14073 ( .A(n13909), .B(n13910), .Z(n13944) );
  ANDN U14074 ( .B(y[770]), .A(n174), .Z(n13886) );
  ANDN U14075 ( .B(y[789]), .A(n155), .Z(n13884) );
  ANDN U14076 ( .B(y[777]), .A(n167), .Z(n13885) );
  XNOR U14077 ( .A(n13884), .B(n13885), .Z(n13887) );
  XOR U14078 ( .A(n13886), .B(n13887), .Z(n13904) );
  ANDN U14079 ( .B(y[778]), .A(n166), .Z(n13892) );
  ANDN U14080 ( .B(y[775]), .A(n169), .Z(n13890) );
  ANDN U14081 ( .B(y[787]), .A(n157), .Z(n13891) );
  XNOR U14082 ( .A(n13890), .B(n13891), .Z(n13893) );
  XOR U14083 ( .A(n13892), .B(n13893), .Z(n13902) );
  OR U14084 ( .A(n13759), .B(n13758), .Z(n13762) );
  NANDN U14085 ( .A(n13760), .B(n13896), .Z(n13761) );
  NAND U14086 ( .A(n13762), .B(n13761), .Z(n13901) );
  XOR U14087 ( .A(n13902), .B(n13901), .Z(n13903) );
  XOR U14088 ( .A(n13904), .B(n13903), .Z(n13943) );
  XNOR U14089 ( .A(n13944), .B(n13943), .Z(n13946) );
  NANDN U14090 ( .A(n13764), .B(n13763), .Z(n13768) );
  OR U14091 ( .A(n13766), .B(n13765), .Z(n13767) );
  AND U14092 ( .A(n13768), .B(n13767), .Z(n13945) );
  XOR U14093 ( .A(n13946), .B(n13945), .Z(n13847) );
  OR U14094 ( .A(n13770), .B(n13769), .Z(n13774) );
  NANDN U14095 ( .A(n13772), .B(n13771), .Z(n13773) );
  AND U14096 ( .A(n13774), .B(n13773), .Z(n13848) );
  NANDN U14097 ( .A(n13776), .B(n13775), .Z(n13780) );
  OR U14098 ( .A(n13778), .B(n13777), .Z(n13779) );
  AND U14099 ( .A(n13780), .B(n13779), .Z(n13849) );
  XOR U14100 ( .A(n13850), .B(n13849), .Z(n13844) );
  NANDN U14101 ( .A(n13782), .B(n13781), .Z(n13786) );
  NANDN U14102 ( .A(n13784), .B(n13783), .Z(n13785) );
  NAND U14103 ( .A(n13786), .B(n13785), .Z(n13842) );
  OR U14104 ( .A(n13788), .B(n13787), .Z(n13792) );
  NANDN U14105 ( .A(n13790), .B(n13789), .Z(n13791) );
  AND U14106 ( .A(n13792), .B(n13791), .Z(n13841) );
  XOR U14107 ( .A(n13844), .B(n13843), .Z(n13823) );
  XNOR U14108 ( .A(n13824), .B(n13823), .Z(n13826) );
  NANDN U14109 ( .A(n13794), .B(n13793), .Z(n13798) );
  NAND U14110 ( .A(n13796), .B(n13795), .Z(n13797) );
  NAND U14111 ( .A(n13798), .B(n13797), .Z(n13825) );
  XOR U14112 ( .A(n13826), .B(n13825), .Z(n13950) );
  XOR U14113 ( .A(n13949), .B(n13950), .Z(n13952) );
  XNOR U14114 ( .A(n13951), .B(n13952), .Z(n13820) );
  OR U14115 ( .A(n13800), .B(n13799), .Z(n13804) );
  NANDN U14116 ( .A(n13802), .B(n13801), .Z(n13803) );
  AND U14117 ( .A(n13804), .B(n13803), .Z(n13817) );
  NANDN U14118 ( .A(n13806), .B(n13805), .Z(n13810) );
  OR U14119 ( .A(n13808), .B(n13807), .Z(n13809) );
  NAND U14120 ( .A(n13810), .B(n13809), .Z(n13818) );
  XOR U14121 ( .A(n13817), .B(n13818), .Z(n13819) );
  XOR U14122 ( .A(n13820), .B(n13819), .Z(n13814) );
  XOR U14123 ( .A(n13813), .B(n13814), .Z(N314) );
  NANDN U14124 ( .A(n13812), .B(n13811), .Z(n13816) );
  NANDN U14125 ( .A(n13814), .B(n13813), .Z(n13815) );
  NAND U14126 ( .A(n13816), .B(n13815), .Z(n13955) );
  OR U14127 ( .A(n13818), .B(n13817), .Z(n13822) );
  NANDN U14128 ( .A(n13820), .B(n13819), .Z(n13821) );
  AND U14129 ( .A(n13822), .B(n13821), .Z(n13956) );
  XNOR U14130 ( .A(n13955), .B(n13956), .Z(n13957) );
  OR U14131 ( .A(n13824), .B(n13823), .Z(n13828) );
  OR U14132 ( .A(n13826), .B(n13825), .Z(n13827) );
  NAND U14133 ( .A(n13828), .B(n13827), .Z(n13964) );
  OR U14134 ( .A(n13830), .B(n13829), .Z(n13834) );
  NANDN U14135 ( .A(n13832), .B(n13831), .Z(n13833) );
  NAND U14136 ( .A(n13834), .B(n13833), .Z(n14090) );
  NANDN U14137 ( .A(n13836), .B(n13835), .Z(n13840) );
  OR U14138 ( .A(n13838), .B(n13837), .Z(n13839) );
  NAND U14139 ( .A(n13840), .B(n13839), .Z(n14091) );
  NANDN U14140 ( .A(n13842), .B(n13841), .Z(n13846) );
  NANDN U14141 ( .A(n13844), .B(n13843), .Z(n13845) );
  AND U14142 ( .A(n13846), .B(n13845), .Z(n14096) );
  NANDN U14143 ( .A(n13848), .B(n13847), .Z(n13852) );
  OR U14144 ( .A(n13850), .B(n13849), .Z(n13851) );
  AND U14145 ( .A(n13852), .B(n13851), .Z(n14010) );
  NANDN U14146 ( .A(n13854), .B(n13853), .Z(n13858) );
  NANDN U14147 ( .A(n13856), .B(n13855), .Z(n13857) );
  NAND U14148 ( .A(n13858), .B(n13857), .Z(n14002) );
  NANDN U14149 ( .A(n13860), .B(n13859), .Z(n13864) );
  NAND U14150 ( .A(n13862), .B(n13861), .Z(n13863) );
  NAND U14151 ( .A(n13864), .B(n13863), .Z(n14001) );
  XNOR U14152 ( .A(n14002), .B(n14001), .Z(n14003) );
  ANDN U14153 ( .B(y[785]), .A(n160), .Z(n14078) );
  ANDN U14154 ( .B(y[788]), .A(n157), .Z(n14076) );
  ANDN U14155 ( .B(y[786]), .A(n159), .Z(n14077) );
  XNOR U14156 ( .A(n14076), .B(n14077), .Z(n14079) );
  XNOR U14157 ( .A(n14078), .B(n14079), .Z(n14056) );
  NANDN U14158 ( .A(n158), .B(y[787]), .Z(n14053) );
  ANDN U14159 ( .B(y[784]), .A(n161), .Z(n14031) );
  ANDN U14160 ( .B(y[782]), .A(n163), .Z(n14029) );
  ANDN U14161 ( .B(y[789]), .A(n156), .Z(n14030) );
  XNOR U14162 ( .A(n14029), .B(n14030), .Z(n14032) );
  XNOR U14163 ( .A(n14031), .B(n14032), .Z(n14054) );
  XOR U14164 ( .A(n14053), .B(n14054), .Z(n14055) );
  XNOR U14165 ( .A(n14056), .B(n14055), .Z(n14004) );
  XNOR U14166 ( .A(n14003), .B(n14004), .Z(n14041) );
  OR U14167 ( .A(n13866), .B(n13865), .Z(n13870) );
  OR U14168 ( .A(n13868), .B(n13867), .Z(n13869) );
  AND U14169 ( .A(n13870), .B(n13869), .Z(n14042) );
  XOR U14170 ( .A(n14041), .B(n14042), .Z(n14044) );
  NAND U14171 ( .A(x[128]), .B(y[794]), .Z(n14036) );
  AND U14172 ( .A(y[768]), .B(x[154]), .Z(n14035) );
  XNOR U14173 ( .A(n14036), .B(n14035), .Z(n14037) );
  ANDN U14174 ( .B(y[769]), .A(n14372), .Z(n14075) );
  XNOR U14175 ( .A(o[154]), .B(n14075), .Z(n14038) );
  AND U14176 ( .A(n13871), .B(o[153]), .Z(n14068) );
  AND U14177 ( .A(y[780]), .B(x[142]), .Z(n14065) );
  AND U14178 ( .A(y[793]), .B(x[129]), .Z(n14066) );
  XNOR U14179 ( .A(n14065), .B(n14066), .Z(n14067) );
  XOR U14180 ( .A(n14068), .B(n14067), .Z(n14023) );
  NAND U14181 ( .A(n13873), .B(n13872), .Z(n13877) );
  NANDN U14182 ( .A(n13875), .B(n13874), .Z(n13876) );
  NAND U14183 ( .A(n13877), .B(n13876), .Z(n14024) );
  XOR U14184 ( .A(n14023), .B(n14024), .Z(n14025) );
  OR U14185 ( .A(n13879), .B(n13878), .Z(n13883) );
  OR U14186 ( .A(n13881), .B(n13880), .Z(n13882) );
  AND U14187 ( .A(n13883), .B(n13882), .Z(n13973) );
  OR U14188 ( .A(n13885), .B(n13884), .Z(n13889) );
  OR U14189 ( .A(n13887), .B(n13886), .Z(n13888) );
  AND U14190 ( .A(n13889), .B(n13888), .Z(n13974) );
  XNOR U14191 ( .A(n13973), .B(n13974), .Z(n13976) );
  XNOR U14192 ( .A(n13975), .B(n13976), .Z(n14016) );
  ANDN U14193 ( .B(y[790]), .A(n155), .Z(n13996) );
  XOR U14194 ( .A(n13995), .B(n13996), .Z(n13997) );
  XNOR U14195 ( .A(n13998), .B(n13997), .Z(n13979) );
  OR U14196 ( .A(n13891), .B(n13890), .Z(n13895) );
  OR U14197 ( .A(n13893), .B(n13892), .Z(n13894) );
  NAND U14198 ( .A(n13895), .B(n13894), .Z(n13980) );
  XOR U14199 ( .A(n13979), .B(n13980), .Z(n13982) );
  NAND U14200 ( .A(x[147]), .B(y[775]), .Z(n14060) );
  ANDN U14201 ( .B(y[783]), .A(n162), .Z(n14059) );
  XNOR U14202 ( .A(n14060), .B(n14059), .Z(n14062) );
  ANDN U14203 ( .B(y[791]), .A(n154), .Z(n14061) );
  XNOR U14204 ( .A(n14062), .B(n14061), .Z(n13981) );
  XOR U14205 ( .A(n13982), .B(n13981), .Z(n14013) );
  AND U14206 ( .A(y[773]), .B(x[149]), .Z(n14070) );
  NAND U14207 ( .A(n13896), .B(n14070), .Z(n13900) );
  OR U14208 ( .A(n13898), .B(n13897), .Z(n13899) );
  NAND U14209 ( .A(n13900), .B(n13899), .Z(n13968) );
  NAND U14210 ( .A(x[150]), .B(y[772]), .Z(n13986) );
  AND U14211 ( .A(x[151]), .B(y[771]), .Z(n13984) );
  XNOR U14212 ( .A(n13986), .B(n13985), .Z(n13967) );
  XNOR U14213 ( .A(n13968), .B(n13967), .Z(n13970) );
  NANDN U14214 ( .A(n150), .B(x[148]), .Z(n14071) );
  XNOR U14215 ( .A(n14070), .B(n14069), .Z(n14072) );
  XOR U14216 ( .A(n14071), .B(n14072), .Z(n13969) );
  XOR U14217 ( .A(n13970), .B(n13969), .Z(n14014) );
  XOR U14218 ( .A(n14013), .B(n14014), .Z(n14015) );
  XNOR U14219 ( .A(n14016), .B(n14015), .Z(n14043) );
  XOR U14220 ( .A(n14044), .B(n14043), .Z(n14008) );
  NANDN U14221 ( .A(n13902), .B(n13901), .Z(n13906) );
  OR U14222 ( .A(n13904), .B(n13903), .Z(n13905) );
  NAND U14223 ( .A(n13906), .B(n13905), .Z(n14087) );
  XOR U14224 ( .A(n14087), .B(n14086), .Z(n14088) );
  XNOR U14225 ( .A(n14088), .B(n14089), .Z(n14007) );
  XOR U14226 ( .A(n14008), .B(n14007), .Z(n14009) );
  XNOR U14227 ( .A(n14010), .B(n14009), .Z(n14097) );
  XNOR U14228 ( .A(n14096), .B(n14097), .Z(n14099) );
  NAND U14229 ( .A(x[130]), .B(y[792]), .Z(n13990) );
  XOR U14230 ( .A(n13990), .B(n13989), .Z(n13992) );
  AND U14231 ( .A(y[770]), .B(x[152]), .Z(n13991) );
  XOR U14232 ( .A(n13992), .B(n13991), .Z(n14018) );
  OR U14233 ( .A(n13920), .B(n13919), .Z(n13924) );
  OR U14234 ( .A(n13922), .B(n13921), .Z(n13923) );
  NAND U14235 ( .A(n13924), .B(n13923), .Z(n14017) );
  XNOR U14236 ( .A(n14018), .B(n14017), .Z(n14020) );
  OR U14237 ( .A(n13926), .B(n13925), .Z(n13930) );
  NANDN U14238 ( .A(n13928), .B(n13927), .Z(n13929) );
  NAND U14239 ( .A(n13930), .B(n13929), .Z(n14019) );
  XNOR U14240 ( .A(n14020), .B(n14019), .Z(n14083) );
  XOR U14241 ( .A(n14082), .B(n14083), .Z(n14085) );
  NAND U14242 ( .A(n13932), .B(n13931), .Z(n13936) );
  NANDN U14243 ( .A(n13934), .B(n13933), .Z(n13935) );
  AND U14244 ( .A(n13936), .B(n13935), .Z(n14084) );
  XOR U14245 ( .A(n14085), .B(n14084), .Z(n14049) );
  OR U14246 ( .A(n13938), .B(n13937), .Z(n13942) );
  NANDN U14247 ( .A(n13940), .B(n13939), .Z(n13941) );
  AND U14248 ( .A(n13942), .B(n13941), .Z(n14047) );
  NAND U14249 ( .A(n13944), .B(n13943), .Z(n13948) );
  OR U14250 ( .A(n13946), .B(n13945), .Z(n13947) );
  NAND U14251 ( .A(n13948), .B(n13947), .Z(n14048) );
  XNOR U14252 ( .A(n14047), .B(n14048), .Z(n14050) );
  XOR U14253 ( .A(n14049), .B(n14050), .Z(n14098) );
  XNOR U14254 ( .A(n14099), .B(n14098), .Z(n14093) );
  XOR U14255 ( .A(n14092), .B(n14093), .Z(n13961) );
  NANDN U14256 ( .A(n13950), .B(n13949), .Z(n13954) );
  NANDN U14257 ( .A(n13952), .B(n13951), .Z(n13953) );
  AND U14258 ( .A(n13954), .B(n13953), .Z(n13962) );
  XNOR U14259 ( .A(n13964), .B(n13963), .Z(n13958) );
  XOR U14260 ( .A(n13957), .B(n13958), .Z(N315) );
  NANDN U14261 ( .A(n13956), .B(n13955), .Z(n13960) );
  NANDN U14262 ( .A(n13958), .B(n13957), .Z(n13959) );
  NAND U14263 ( .A(n13960), .B(n13959), .Z(n14102) );
  NANDN U14264 ( .A(n13962), .B(n13961), .Z(n13966) );
  NANDN U14265 ( .A(n13964), .B(n13963), .Z(n13965) );
  NAND U14266 ( .A(n13966), .B(n13965), .Z(n14103) );
  XNOR U14267 ( .A(n14102), .B(n14103), .Z(n14104) );
  OR U14268 ( .A(n13968), .B(n13967), .Z(n13972) );
  OR U14269 ( .A(n13970), .B(n13969), .Z(n13971) );
  NAND U14270 ( .A(n13972), .B(n13971), .Z(n14125) );
  OR U14271 ( .A(n13974), .B(n13973), .Z(n13978) );
  NANDN U14272 ( .A(n13976), .B(n13975), .Z(n13977) );
  AND U14273 ( .A(n13978), .B(n13977), .Z(n14131) );
  OR U14274 ( .A(n13984), .B(n13983), .Z(n13988) );
  NAND U14275 ( .A(n13986), .B(n13985), .Z(n13987) );
  AND U14276 ( .A(n13988), .B(n13987), .Z(n14201) );
  NANDN U14277 ( .A(n13990), .B(n13989), .Z(n13994) );
  NANDN U14278 ( .A(n13992), .B(n13991), .Z(n13993) );
  NAND U14279 ( .A(n13994), .B(n13993), .Z(n14202) );
  XNOR U14280 ( .A(n14201), .B(n14202), .Z(n14204) );
  OR U14281 ( .A(n13996), .B(n13995), .Z(n14000) );
  NANDN U14282 ( .A(n13998), .B(n13997), .Z(n13999) );
  AND U14283 ( .A(n14000), .B(n13999), .Z(n14195) );
  ANDN U14284 ( .B(y[786]), .A(n160), .Z(n14154) );
  ANDN U14285 ( .B(y[777]), .A(n169), .Z(n14152) );
  ANDN U14286 ( .B(y[774]), .A(n172), .Z(n14153) );
  XNOR U14287 ( .A(n14152), .B(n14153), .Z(n14155) );
  XNOR U14288 ( .A(n14154), .B(n14155), .Z(n14196) );
  XNOR U14289 ( .A(n14195), .B(n14196), .Z(n14198) );
  ANDN U14290 ( .B(y[795]), .A(n151), .Z(n14142) );
  NAND U14291 ( .A(x[154]), .B(y[769]), .Z(n14158) );
  XNOR U14292 ( .A(n14158), .B(o[155]), .Z(n14140) );
  ANDN U14293 ( .B(y[768]), .A(n177), .Z(n14141) );
  XNOR U14294 ( .A(n14140), .B(n14141), .Z(n14143) );
  XNOR U14295 ( .A(n14142), .B(n14143), .Z(n14197) );
  XOR U14296 ( .A(n14198), .B(n14197), .Z(n14203) );
  XNOR U14297 ( .A(n14129), .B(n14128), .Z(n14130) );
  XOR U14298 ( .A(n14131), .B(n14130), .Z(n14124) );
  XOR U14299 ( .A(n14125), .B(n14124), .Z(n14127) );
  OR U14300 ( .A(n14002), .B(n14001), .Z(n14006) );
  OR U14301 ( .A(n14004), .B(n14003), .Z(n14005) );
  NAND U14302 ( .A(n14006), .B(n14005), .Z(n14126) );
  XOR U14303 ( .A(n14127), .B(n14126), .Z(n14251) );
  OR U14304 ( .A(n14008), .B(n14007), .Z(n14012) );
  NANDN U14305 ( .A(n14010), .B(n14009), .Z(n14011) );
  AND U14306 ( .A(n14012), .B(n14011), .Z(n14252) );
  OR U14307 ( .A(n14018), .B(n14017), .Z(n14022) );
  OR U14308 ( .A(n14020), .B(n14019), .Z(n14021) );
  AND U14309 ( .A(n14022), .B(n14021), .Z(n14136) );
  OR U14310 ( .A(n14024), .B(n14023), .Z(n14028) );
  NANDN U14311 ( .A(n14026), .B(n14025), .Z(n14027) );
  AND U14312 ( .A(n14028), .B(n14027), .Z(n14135) );
  ANDN U14313 ( .B(y[783]), .A(n163), .Z(n14219) );
  ANDN U14314 ( .B(y[782]), .A(n164), .Z(n14220) );
  XNOR U14315 ( .A(n14219), .B(n14220), .Z(n14222) );
  ANDN U14316 ( .B(y[784]), .A(n162), .Z(n14233) );
  ANDN U14317 ( .B(y[779]), .A(n167), .Z(n14232) );
  XNOR U14318 ( .A(n14231), .B(n14232), .Z(n14234) );
  XNOR U14319 ( .A(n14233), .B(n14234), .Z(n14221) );
  XOR U14320 ( .A(n14222), .B(n14221), .Z(n14179) );
  NAND U14321 ( .A(x[131]), .B(y[792]), .Z(n14228) );
  ANDN U14322 ( .B(y[793]), .A(n153), .Z(n14226) );
  XOR U14323 ( .A(n14225), .B(n14226), .Z(n14227) );
  XNOR U14324 ( .A(n14228), .B(n14227), .Z(n14177) );
  NAND U14325 ( .A(x[134]), .B(y[789]), .Z(n14167) );
  ANDN U14326 ( .B(y[770]), .A(n14372), .Z(n14165) );
  ANDN U14327 ( .B(y[776]), .A(n170), .Z(n14166) );
  XNOR U14328 ( .A(n14165), .B(n14166), .Z(n14168) );
  XNOR U14329 ( .A(n14167), .B(n14168), .Z(n14178) );
  XOR U14330 ( .A(n14177), .B(n14178), .Z(n14180) );
  XNOR U14331 ( .A(n14179), .B(n14180), .Z(n14209) );
  OR U14332 ( .A(n14030), .B(n14029), .Z(n14034) );
  OR U14333 ( .A(n14032), .B(n14031), .Z(n14033) );
  AND U14334 ( .A(n14034), .B(n14033), .Z(n14207) );
  NANDN U14335 ( .A(n14036), .B(n14035), .Z(n14040) );
  NANDN U14336 ( .A(n14038), .B(n14037), .Z(n14039) );
  NAND U14337 ( .A(n14040), .B(n14039), .Z(n14208) );
  XNOR U14338 ( .A(n14207), .B(n14208), .Z(n14210) );
  XOR U14339 ( .A(n14209), .B(n14210), .Z(n14134) );
  XOR U14340 ( .A(n14135), .B(n14134), .Z(n14137) );
  XNOR U14341 ( .A(n14136), .B(n14137), .Z(n14121) );
  XOR U14342 ( .A(n14120), .B(n14121), .Z(n14122) );
  NANDN U14343 ( .A(n14042), .B(n14041), .Z(n14046) );
  NANDN U14344 ( .A(n14044), .B(n14043), .Z(n14045) );
  AND U14345 ( .A(n14046), .B(n14045), .Z(n14123) );
  XNOR U14346 ( .A(n14122), .B(n14123), .Z(n14253) );
  XOR U14347 ( .A(n14254), .B(n14253), .Z(n14247) );
  OR U14348 ( .A(n14048), .B(n14047), .Z(n14052) );
  NANDN U14349 ( .A(n14050), .B(n14049), .Z(n14051) );
  AND U14350 ( .A(n14052), .B(n14051), .Z(n14245) );
  NANDN U14351 ( .A(n14054), .B(n14053), .Z(n14058) );
  OR U14352 ( .A(n14056), .B(n14055), .Z(n14057) );
  AND U14353 ( .A(n14058), .B(n14057), .Z(n14116) );
  NANDN U14354 ( .A(n14060), .B(n14059), .Z(n14064) );
  NAND U14355 ( .A(n14062), .B(n14061), .Z(n14063) );
  AND U14356 ( .A(n14064), .B(n14063), .Z(n14185) );
  NAND U14357 ( .A(x[150]), .B(y[773]), .Z(n14237) );
  ANDN U14358 ( .B(y[772]), .A(n174), .Z(n14235) );
  ANDN U14359 ( .B(y[787]), .A(n159), .Z(n14236) );
  XNOR U14360 ( .A(n14235), .B(n14236), .Z(n14238) );
  XOR U14361 ( .A(n14237), .B(n14238), .Z(n14183) );
  NAND U14362 ( .A(y[788]), .B(x[135]), .Z(n14161) );
  ANDN U14363 ( .B(y[771]), .A(n175), .Z(n14160) );
  XNOR U14364 ( .A(n14159), .B(n14160), .Z(n14162) );
  XNOR U14365 ( .A(n14161), .B(n14162), .Z(n14184) );
  XOR U14366 ( .A(n14183), .B(n14184), .Z(n14186) );
  XOR U14367 ( .A(n14185), .B(n14186), .Z(n14114) );
  OR U14368 ( .A(n14070), .B(n14069), .Z(n14074) );
  NANDN U14369 ( .A(n14072), .B(n14071), .Z(n14073) );
  NAND U14370 ( .A(n14074), .B(n14073), .Z(n14171) );
  XNOR U14371 ( .A(n14172), .B(n14171), .Z(n14174) );
  AND U14372 ( .A(n14075), .B(o[154]), .Z(n14213) );
  ANDN U14373 ( .B(y[794]), .A(n152), .Z(n14214) );
  XNOR U14374 ( .A(n14213), .B(n14214), .Z(n14215) );
  XOR U14375 ( .A(n14216), .B(n14215), .Z(n14189) );
  NAND U14376 ( .A(x[145]), .B(y[778]), .Z(n14147) );
  AND U14377 ( .A(y[791]), .B(x[132]), .Z(n14146) );
  XOR U14378 ( .A(n14147), .B(n14146), .Z(n14149) );
  AND U14379 ( .A(y[790]), .B(x[133]), .Z(n14148) );
  XOR U14380 ( .A(n14149), .B(n14148), .Z(n14190) );
  XNOR U14381 ( .A(n14189), .B(n14190), .Z(n14192) );
  OR U14382 ( .A(n14077), .B(n14076), .Z(n14081) );
  OR U14383 ( .A(n14079), .B(n14078), .Z(n14080) );
  NAND U14384 ( .A(n14081), .B(n14080), .Z(n14191) );
  XNOR U14385 ( .A(n14192), .B(n14191), .Z(n14173) );
  XOR U14386 ( .A(n14174), .B(n14173), .Z(n14115) );
  XNOR U14387 ( .A(n14114), .B(n14115), .Z(n14117) );
  XOR U14388 ( .A(n14116), .B(n14117), .Z(n14241) );
  XNOR U14389 ( .A(n14241), .B(n14242), .Z(n14244) );
  XOR U14390 ( .A(n14244), .B(n14243), .Z(n14246) );
  XNOR U14391 ( .A(n14245), .B(n14246), .Z(n14248) );
  XNOR U14392 ( .A(n14247), .B(n14248), .Z(n14111) );
  NANDN U14393 ( .A(n14091), .B(n14090), .Z(n14095) );
  NANDN U14394 ( .A(n14093), .B(n14092), .Z(n14094) );
  NAND U14395 ( .A(n14095), .B(n14094), .Z(n14109) );
  OR U14396 ( .A(n14097), .B(n14096), .Z(n14101) );
  OR U14397 ( .A(n14099), .B(n14098), .Z(n14100) );
  AND U14398 ( .A(n14101), .B(n14100), .Z(n14108) );
  XNOR U14399 ( .A(n14111), .B(n14110), .Z(n14105) );
  XOR U14400 ( .A(n14104), .B(n14105), .Z(N316) );
  NANDN U14401 ( .A(n14103), .B(n14102), .Z(n14107) );
  NANDN U14402 ( .A(n14105), .B(n14104), .Z(n14106) );
  NAND U14403 ( .A(n14107), .B(n14106), .Z(n14257) );
  NANDN U14404 ( .A(n14109), .B(n14108), .Z(n14113) );
  NANDN U14405 ( .A(n14111), .B(n14110), .Z(n14112) );
  NAND U14406 ( .A(n14113), .B(n14112), .Z(n14258) );
  XNOR U14407 ( .A(n14257), .B(n14258), .Z(n14259) );
  OR U14408 ( .A(n14115), .B(n14114), .Z(n14119) );
  OR U14409 ( .A(n14117), .B(n14116), .Z(n14118) );
  AND U14410 ( .A(n14119), .B(n14118), .Z(n14419) );
  XOR U14411 ( .A(n14417), .B(n14416), .Z(n14418) );
  XNOR U14412 ( .A(n14419), .B(n14418), .Z(n14424) );
  NANDN U14413 ( .A(n14129), .B(n14128), .Z(n14133) );
  NANDN U14414 ( .A(n14131), .B(n14130), .Z(n14132) );
  AND U14415 ( .A(n14133), .B(n14132), .Z(n14404) );
  NANDN U14416 ( .A(n14135), .B(n14134), .Z(n14139) );
  OR U14417 ( .A(n14137), .B(n14136), .Z(n14138) );
  NAND U14418 ( .A(n14139), .B(n14138), .Z(n14405) );
  XNOR U14419 ( .A(n14404), .B(n14405), .Z(n14407) );
  OR U14420 ( .A(n14141), .B(n14140), .Z(n14145) );
  OR U14421 ( .A(n14143), .B(n14142), .Z(n14144) );
  AND U14422 ( .A(n14145), .B(n14144), .Z(n14287) );
  NANDN U14423 ( .A(n14147), .B(n14146), .Z(n14151) );
  NANDN U14424 ( .A(n14149), .B(n14148), .Z(n14150) );
  NAND U14425 ( .A(n14151), .B(n14150), .Z(n14288) );
  XNOR U14426 ( .A(n14287), .B(n14288), .Z(n14290) );
  OR U14427 ( .A(n14153), .B(n14152), .Z(n14157) );
  OR U14428 ( .A(n14155), .B(n14154), .Z(n14156) );
  AND U14429 ( .A(n14157), .B(n14156), .Z(n14317) );
  ANDN U14430 ( .B(y[787]), .A(n160), .Z(n14330) );
  ANDN U14431 ( .B(y[788]), .A(n159), .Z(n14331) );
  XNOR U14432 ( .A(n14330), .B(n14331), .Z(n14333) );
  ANDN U14433 ( .B(y[786]), .A(n161), .Z(n14332) );
  XNOR U14434 ( .A(n14333), .B(n14332), .Z(n14318) );
  XOR U14435 ( .A(n14317), .B(n14318), .Z(n14319) );
  ANDN U14436 ( .B(o[155]), .A(n14158), .Z(n14336) );
  ANDN U14437 ( .B(y[768]), .A(n14373), .Z(n14337) );
  XNOR U14438 ( .A(n14336), .B(n14337), .Z(n14339) );
  ANDN U14439 ( .B(y[796]), .A(n151), .Z(n14338) );
  XNOR U14440 ( .A(n14339), .B(n14338), .Z(n14320) );
  XOR U14441 ( .A(n14319), .B(n14320), .Z(n14289) );
  XOR U14442 ( .A(n14290), .B(n14289), .Z(n14271) );
  ANDN U14443 ( .B(y[795]), .A(n152), .Z(n14355) );
  NAND U14444 ( .A(y[771]), .B(x[153]), .Z(n14354) );
  XOR U14445 ( .A(n14355), .B(n14354), .Z(n14357) );
  XNOR U14446 ( .A(n14356), .B(n14357), .Z(n14283) );
  NAND U14447 ( .A(x[144]), .B(y[780]), .Z(n14344) );
  ANDN U14448 ( .B(y[794]), .A(n153), .Z(n14343) );
  NAND U14449 ( .A(x[152]), .B(y[772]), .Z(n14342) );
  XOR U14450 ( .A(n14343), .B(n14342), .Z(n14345) );
  XNOR U14451 ( .A(n14344), .B(n14345), .Z(n14281) );
  OR U14452 ( .A(n14160), .B(n14159), .Z(n14164) );
  NANDN U14453 ( .A(n14162), .B(n14161), .Z(n14163) );
  NAND U14454 ( .A(n14164), .B(n14163), .Z(n14282) );
  XOR U14455 ( .A(n14281), .B(n14282), .Z(n14284) );
  XOR U14456 ( .A(n14283), .B(n14284), .Z(n14269) );
  ANDN U14457 ( .B(y[773]), .A(n174), .Z(n14381) );
  NAND U14458 ( .A(x[131]), .B(y[793]), .Z(n14380) );
  XOR U14459 ( .A(n14381), .B(n14380), .Z(n14383) );
  XNOR U14460 ( .A(n14382), .B(n14383), .Z(n14295) );
  NAND U14461 ( .A(x[133]), .B(y[791]), .Z(n14362) );
  ANDN U14462 ( .B(y[776]), .A(n171), .Z(n14361) );
  NAND U14463 ( .A(x[149]), .B(y[775]), .Z(n14360) );
  XOR U14464 ( .A(n14361), .B(n14360), .Z(n14363) );
  XNOR U14465 ( .A(n14362), .B(n14363), .Z(n14293) );
  OR U14466 ( .A(n14166), .B(n14165), .Z(n14170) );
  NANDN U14467 ( .A(n14168), .B(n14167), .Z(n14169) );
  NAND U14468 ( .A(n14170), .B(n14169), .Z(n14294) );
  XOR U14469 ( .A(n14293), .B(n14294), .Z(n14296) );
  XOR U14470 ( .A(n14295), .B(n14296), .Z(n14270) );
  XNOR U14471 ( .A(n14269), .B(n14270), .Z(n14272) );
  OR U14472 ( .A(n14172), .B(n14171), .Z(n14176) );
  OR U14473 ( .A(n14174), .B(n14173), .Z(n14175) );
  NAND U14474 ( .A(n14176), .B(n14175), .Z(n14308) );
  NANDN U14475 ( .A(n14178), .B(n14177), .Z(n14182) );
  OR U14476 ( .A(n14180), .B(n14179), .Z(n14181) );
  NAND U14477 ( .A(n14182), .B(n14181), .Z(n14306) );
  NANDN U14478 ( .A(n14184), .B(n14183), .Z(n14188) );
  OR U14479 ( .A(n14186), .B(n14185), .Z(n14187) );
  NAND U14480 ( .A(n14188), .B(n14187), .Z(n14305) );
  XNOR U14481 ( .A(n14306), .B(n14305), .Z(n14307) );
  XNOR U14482 ( .A(n14308), .B(n14307), .Z(n14410) );
  XNOR U14483 ( .A(n14411), .B(n14410), .Z(n14413) );
  OR U14484 ( .A(n14190), .B(n14189), .Z(n14194) );
  OR U14485 ( .A(n14192), .B(n14191), .Z(n14193) );
  AND U14486 ( .A(n14194), .B(n14193), .Z(n14299) );
  OR U14487 ( .A(n14196), .B(n14195), .Z(n14200) );
  OR U14488 ( .A(n14198), .B(n14197), .Z(n14199) );
  NAND U14489 ( .A(n14200), .B(n14199), .Z(n14300) );
  XNOR U14490 ( .A(n14299), .B(n14300), .Z(n14302) );
  OR U14491 ( .A(n14202), .B(n14201), .Z(n14206) );
  NANDN U14492 ( .A(n14204), .B(n14203), .Z(n14205) );
  NAND U14493 ( .A(n14206), .B(n14205), .Z(n14301) );
  XOR U14494 ( .A(n14302), .B(n14301), .Z(n14401) );
  OR U14495 ( .A(n14208), .B(n14207), .Z(n14212) );
  NANDN U14496 ( .A(n14210), .B(n14209), .Z(n14211) );
  AND U14497 ( .A(n14212), .B(n14211), .Z(n14398) );
  OR U14498 ( .A(n14214), .B(n14213), .Z(n14218) );
  OR U14499 ( .A(n14216), .B(n14215), .Z(n14217) );
  AND U14500 ( .A(n14218), .B(n14217), .Z(n14314) );
  OR U14501 ( .A(n14220), .B(n14219), .Z(n14224) );
  OR U14502 ( .A(n14222), .B(n14221), .Z(n14223) );
  AND U14503 ( .A(n14224), .B(n14223), .Z(n14311) );
  OR U14504 ( .A(n14226), .B(n14225), .Z(n14230) );
  NAND U14505 ( .A(n14228), .B(n14227), .Z(n14229) );
  AND U14506 ( .A(n14230), .B(n14229), .Z(n14312) );
  XOR U14507 ( .A(n14311), .B(n14312), .Z(n14313) );
  NAND U14508 ( .A(x[154]), .B(y[770]), .Z(n14387) );
  AND U14509 ( .A(x[143]), .B(y[781]), .Z(n14386) );
  XNOR U14510 ( .A(n14387), .B(n14386), .Z(n14389) );
  NAND U14511 ( .A(x[155]), .B(y[769]), .Z(n14543) );
  XNOR U14512 ( .A(n14543), .B(o[156]), .Z(n14388) );
  XNOR U14513 ( .A(n14389), .B(n14388), .Z(n14377) );
  ANDN U14514 ( .B(y[789]), .A(n158), .Z(n14350) );
  ANDN U14515 ( .B(y[785]), .A(n162), .Z(n14348) );
  ANDN U14516 ( .B(y[784]), .A(n163), .Z(n14349) );
  XNOR U14517 ( .A(n14348), .B(n14349), .Z(n14351) );
  XOR U14518 ( .A(n14350), .B(n14351), .Z(n14374) );
  XNOR U14519 ( .A(n14375), .B(n14374), .Z(n14376) );
  XOR U14520 ( .A(n14377), .B(n14376), .Z(n14275) );
  OR U14521 ( .A(n14236), .B(n14235), .Z(n14240) );
  NANDN U14522 ( .A(n14238), .B(n14237), .Z(n14239) );
  AND U14523 ( .A(n14240), .B(n14239), .Z(n14392) );
  ANDN U14524 ( .B(y[790]), .A(n157), .Z(n14370) );
  ANDN U14525 ( .B(y[777]), .A(n170), .Z(n14369) );
  XNOR U14526 ( .A(n14368), .B(n14369), .Z(n14371) );
  XNOR U14527 ( .A(n14370), .B(n14371), .Z(n14393) );
  XOR U14528 ( .A(n14392), .B(n14393), .Z(n14395) );
  NAND U14529 ( .A(x[145]), .B(y[779]), .Z(n14325) );
  ANDN U14530 ( .B(y[792]), .A(n155), .Z(n14324) );
  NAND U14531 ( .A(y[774]), .B(x[150]), .Z(n14323) );
  XOR U14532 ( .A(n14324), .B(n14323), .Z(n14326) );
  XNOR U14533 ( .A(n14325), .B(n14326), .Z(n14394) );
  XNOR U14534 ( .A(n14395), .B(n14394), .Z(n14276) );
  XOR U14535 ( .A(n14275), .B(n14276), .Z(n14277) );
  XOR U14536 ( .A(n14398), .B(n14399), .Z(n14400) );
  XOR U14537 ( .A(n14413), .B(n14412), .Z(n14406) );
  XNOR U14538 ( .A(n14407), .B(n14406), .Z(n14422) );
  XNOR U14539 ( .A(n14422), .B(n14423), .Z(n14425) );
  XNOR U14540 ( .A(n14424), .B(n14425), .Z(n14263) );
  OR U14541 ( .A(n14246), .B(n14245), .Z(n14250) );
  NANDN U14542 ( .A(n14248), .B(n14247), .Z(n14249) );
  AND U14543 ( .A(n14250), .B(n14249), .Z(n14264) );
  XOR U14544 ( .A(n14263), .B(n14264), .Z(n14266) );
  NANDN U14545 ( .A(n14252), .B(n14251), .Z(n14256) );
  NANDN U14546 ( .A(n14254), .B(n14253), .Z(n14255) );
  NAND U14547 ( .A(n14256), .B(n14255), .Z(n14265) );
  XOR U14548 ( .A(n14266), .B(n14265), .Z(n14260) );
  XNOR U14549 ( .A(n14259), .B(n14260), .Z(N317) );
  NANDN U14550 ( .A(n14258), .B(n14257), .Z(n14262) );
  NAND U14551 ( .A(n14260), .B(n14259), .Z(n14261) );
  NAND U14552 ( .A(n14262), .B(n14261), .Z(n14428) );
  NANDN U14553 ( .A(n14264), .B(n14263), .Z(n14268) );
  OR U14554 ( .A(n14266), .B(n14265), .Z(n14267) );
  AND U14555 ( .A(n14268), .B(n14267), .Z(n14429) );
  XNOR U14556 ( .A(n14428), .B(n14429), .Z(n14430) );
  OR U14557 ( .A(n14270), .B(n14269), .Z(n14274) );
  NANDN U14558 ( .A(n14272), .B(n14271), .Z(n14273) );
  NAND U14559 ( .A(n14274), .B(n14273), .Z(n14446) );
  OR U14560 ( .A(n14276), .B(n14275), .Z(n14280) );
  NANDN U14561 ( .A(n14278), .B(n14277), .Z(n14279) );
  NAND U14562 ( .A(n14280), .B(n14279), .Z(n14451) );
  OR U14563 ( .A(n14282), .B(n14281), .Z(n14286) );
  NAND U14564 ( .A(n14284), .B(n14283), .Z(n14285) );
  NAND U14565 ( .A(n14286), .B(n14285), .Z(n14514) );
  OR U14566 ( .A(n14288), .B(n14287), .Z(n14292) );
  OR U14567 ( .A(n14290), .B(n14289), .Z(n14291) );
  AND U14568 ( .A(n14292), .B(n14291), .Z(n14511) );
  OR U14569 ( .A(n14294), .B(n14293), .Z(n14298) );
  NAND U14570 ( .A(n14296), .B(n14295), .Z(n14297) );
  NAND U14571 ( .A(n14298), .B(n14297), .Z(n14512) );
  XNOR U14572 ( .A(n14511), .B(n14512), .Z(n14513) );
  XOR U14573 ( .A(n14514), .B(n14513), .Z(n14450) );
  XNOR U14574 ( .A(n14451), .B(n14450), .Z(n14453) );
  OR U14575 ( .A(n14300), .B(n14299), .Z(n14304) );
  OR U14576 ( .A(n14302), .B(n14301), .Z(n14303) );
  AND U14577 ( .A(n14304), .B(n14303), .Z(n14452) );
  XOR U14578 ( .A(n14453), .B(n14452), .Z(n14444) );
  OR U14579 ( .A(n14306), .B(n14305), .Z(n14310) );
  OR U14580 ( .A(n14308), .B(n14307), .Z(n14309) );
  AND U14581 ( .A(n14310), .B(n14309), .Z(n14445) );
  XOR U14582 ( .A(n14444), .B(n14445), .Z(n14447) );
  OR U14583 ( .A(n14312), .B(n14311), .Z(n14316) );
  NANDN U14584 ( .A(n14314), .B(n14313), .Z(n14315) );
  AND U14585 ( .A(n14316), .B(n14315), .Z(n14507) );
  OR U14586 ( .A(n14318), .B(n14317), .Z(n14322) );
  NANDN U14587 ( .A(n14320), .B(n14319), .Z(n14321) );
  AND U14588 ( .A(n14322), .B(n14321), .Z(n14505) );
  NANDN U14589 ( .A(n14324), .B(n14323), .Z(n14328) );
  NANDN U14590 ( .A(n14326), .B(n14325), .Z(n14327) );
  AND U14591 ( .A(n14328), .B(n14327), .Z(n14499) );
  ANDN U14592 ( .B(y[775]), .A(n173), .Z(n14573) );
  ANDN U14593 ( .B(y[796]), .A(n152), .Z(n14574) );
  XNOR U14594 ( .A(n14573), .B(n14574), .Z(n14575) );
  NOR U14595 ( .A(n163), .B(n14329), .Z(n14703) );
  XNOR U14596 ( .A(n14575), .B(n14703), .Z(n14471) );
  OR U14597 ( .A(n14331), .B(n14330), .Z(n14335) );
  OR U14598 ( .A(n14333), .B(n14332), .Z(n14334) );
  AND U14599 ( .A(n14335), .B(n14334), .Z(n14469) );
  ANDN U14600 ( .B(y[777]), .A(n171), .Z(n14576) );
  ANDN U14601 ( .B(y[776]), .A(n172), .Z(n14708) );
  XNOR U14602 ( .A(n14576), .B(n14708), .Z(n14578) );
  ANDN U14603 ( .B(y[782]), .A(n166), .Z(n14577) );
  XOR U14604 ( .A(n14578), .B(n14577), .Z(n14468) );
  XOR U14605 ( .A(n14469), .B(n14468), .Z(n14470) );
  XNOR U14606 ( .A(n14471), .B(n14470), .Z(n14500) );
  XOR U14607 ( .A(n14499), .B(n14500), .Z(n14501) );
  OR U14608 ( .A(n14337), .B(n14336), .Z(n14341) );
  OR U14609 ( .A(n14339), .B(n14338), .Z(n14340) );
  AND U14610 ( .A(n14341), .B(n14340), .Z(n14502) );
  XNOR U14611 ( .A(n14505), .B(n14506), .Z(n14508) );
  XOR U14612 ( .A(n14507), .B(n14508), .Z(n14465) );
  NANDN U14613 ( .A(n14343), .B(n14342), .Z(n14347) );
  NANDN U14614 ( .A(n14345), .B(n14344), .Z(n14346) );
  AND U14615 ( .A(n14347), .B(n14346), .Z(n14474) );
  ANDN U14616 ( .B(y[774]), .A(n174), .Z(n14554) );
  ANDN U14617 ( .B(y[773]), .A(n175), .Z(n14785) );
  XNOR U14618 ( .A(n14554), .B(n14785), .Z(n14556) );
  ANDN U14619 ( .B(y[784]), .A(n164), .Z(n14555) );
  XNOR U14620 ( .A(n14556), .B(n14555), .Z(n14526) );
  OR U14621 ( .A(n14349), .B(n14348), .Z(n14353) );
  OR U14622 ( .A(n14351), .B(n14350), .Z(n14352) );
  AND U14623 ( .A(n14353), .B(n14352), .Z(n14524) );
  ANDN U14624 ( .B(y[786]), .A(n162), .Z(n14548) );
  ANDN U14625 ( .B(y[780]), .A(n168), .Z(n14549) );
  XNOR U14626 ( .A(n14548), .B(n14549), .Z(n14551) );
  ANDN U14627 ( .B(y[794]), .A(n154), .Z(n14550) );
  XOR U14628 ( .A(n14551), .B(n14550), .Z(n14523) );
  XOR U14629 ( .A(n14524), .B(n14523), .Z(n14525) );
  XNOR U14630 ( .A(n14526), .B(n14525), .Z(n14475) );
  XOR U14631 ( .A(n14474), .B(n14475), .Z(n14476) );
  NANDN U14632 ( .A(n14355), .B(n14354), .Z(n14359) );
  OR U14633 ( .A(n14357), .B(n14356), .Z(n14358) );
  AND U14634 ( .A(n14359), .B(n14358), .Z(n14477) );
  ANDN U14635 ( .B(y[779]), .A(n169), .Z(n14535) );
  ANDN U14636 ( .B(y[778]), .A(n170), .Z(n14536) );
  XNOR U14637 ( .A(n14535), .B(n14536), .Z(n14538) );
  ANDN U14638 ( .B(y[795]), .A(n153), .Z(n14537) );
  XNOR U14639 ( .A(n14538), .B(n14537), .Z(n14570) );
  NANDN U14640 ( .A(n14361), .B(n14360), .Z(n14365) );
  NANDN U14641 ( .A(n14363), .B(n14362), .Z(n14364) );
  AND U14642 ( .A(n14365), .B(n14364), .Z(n14568) );
  NAND U14643 ( .A(y[769]), .B(o[156]), .Z(n14366) );
  XNOR U14644 ( .A(y[770]), .B(n14366), .Z(n14367) );
  NAND U14645 ( .A(x[155]), .B(n14367), .Z(n14542) );
  ANDN U14646 ( .B(y[781]), .A(n167), .Z(n14541) );
  XOR U14647 ( .A(n14542), .B(n14541), .Z(n14567) );
  XOR U14648 ( .A(n14568), .B(n14567), .Z(n14569) );
  XNOR U14649 ( .A(n14570), .B(n14569), .Z(n14597) );
  ANDN U14650 ( .B(y[772]), .A(n14372), .Z(n14584) );
  ANDN U14651 ( .B(y[771]), .A(n176), .Z(n14585) );
  XNOR U14652 ( .A(n14584), .B(n14585), .Z(n14587) );
  ANDN U14653 ( .B(y[783]), .A(n165), .Z(n14586) );
  XOR U14654 ( .A(n14587), .B(n14586), .Z(n14480) );
  NAND U14655 ( .A(x[128]), .B(y[797]), .Z(n14496) );
  ANDN U14656 ( .B(y[769]), .A(n14373), .Z(n14583) );
  XOR U14657 ( .A(o[157]), .B(n14583), .Z(n14494) );
  NAND U14658 ( .A(x[157]), .B(y[768]), .Z(n14493) );
  XNOR U14659 ( .A(n14494), .B(n14493), .Z(n14495) );
  XOR U14660 ( .A(n14496), .B(n14495), .Z(n14481) );
  XNOR U14661 ( .A(n14480), .B(n14481), .Z(n14482) );
  XOR U14662 ( .A(n14483), .B(n14482), .Z(n14596) );
  XNOR U14663 ( .A(n14597), .B(n14596), .Z(n14598) );
  XOR U14664 ( .A(n14599), .B(n14598), .Z(n14593) );
  OR U14665 ( .A(n14375), .B(n14374), .Z(n14379) );
  OR U14666 ( .A(n14377), .B(n14376), .Z(n14378) );
  AND U14667 ( .A(n14379), .B(n14378), .Z(n14590) );
  NANDN U14668 ( .A(n14381), .B(n14380), .Z(n14385) );
  OR U14669 ( .A(n14383), .B(n14382), .Z(n14384) );
  AND U14670 ( .A(n14385), .B(n14384), .Z(n14517) );
  NANDN U14671 ( .A(n14387), .B(n14386), .Z(n14391) );
  NAND U14672 ( .A(n14389), .B(n14388), .Z(n14390) );
  NAND U14673 ( .A(n14391), .B(n14390), .Z(n14518) );
  XOR U14674 ( .A(n14517), .B(n14518), .Z(n14519) );
  ANDN U14675 ( .B(y[792]), .A(n156), .Z(n14529) );
  ANDN U14676 ( .B(y[787]), .A(n161), .Z(n14530) );
  XNOR U14677 ( .A(n14529), .B(n14530), .Z(n14532) );
  ANDN U14678 ( .B(y[793]), .A(n155), .Z(n14531) );
  XNOR U14679 ( .A(n14532), .B(n14531), .Z(n14486) );
  XNOR U14680 ( .A(n14696), .B(n14486), .Z(n14488) );
  ANDN U14681 ( .B(y[789]), .A(n159), .Z(n14559) );
  ANDN U14682 ( .B(y[790]), .A(n158), .Z(n14560) );
  XNOR U14683 ( .A(n14559), .B(n14560), .Z(n14562) );
  ANDN U14684 ( .B(y[791]), .A(n157), .Z(n14561) );
  XOR U14685 ( .A(n14562), .B(n14561), .Z(n14487) );
  XOR U14686 ( .A(n14488), .B(n14487), .Z(n14520) );
  XNOR U14687 ( .A(n14519), .B(n14520), .Z(n14591) );
  XOR U14688 ( .A(n14590), .B(n14591), .Z(n14592) );
  XOR U14689 ( .A(n14593), .B(n14592), .Z(n14463) );
  OR U14690 ( .A(n14393), .B(n14392), .Z(n14397) );
  NAND U14691 ( .A(n14395), .B(n14394), .Z(n14396) );
  NAND U14692 ( .A(n14397), .B(n14396), .Z(n14462) );
  XOR U14693 ( .A(n14463), .B(n14462), .Z(n14464) );
  XOR U14694 ( .A(n14465), .B(n14464), .Z(n14457) );
  OR U14695 ( .A(n14399), .B(n14398), .Z(n14403) );
  NANDN U14696 ( .A(n14401), .B(n14400), .Z(n14402) );
  NAND U14697 ( .A(n14403), .B(n14402), .Z(n14456) );
  XNOR U14698 ( .A(n14457), .B(n14456), .Z(n14459) );
  XOR U14699 ( .A(n14458), .B(n14459), .Z(n14440) );
  OR U14700 ( .A(n14405), .B(n14404), .Z(n14409) );
  NANDN U14701 ( .A(n14407), .B(n14406), .Z(n14408) );
  AND U14702 ( .A(n14409), .B(n14408), .Z(n14438) );
  OR U14703 ( .A(n14411), .B(n14410), .Z(n14415) );
  OR U14704 ( .A(n14413), .B(n14412), .Z(n14414) );
  AND U14705 ( .A(n14415), .B(n14414), .Z(n14439) );
  XNOR U14706 ( .A(n14438), .B(n14439), .Z(n14441) );
  XNOR U14707 ( .A(n14440), .B(n14441), .Z(n14437) );
  OR U14708 ( .A(n14417), .B(n14416), .Z(n14421) );
  NANDN U14709 ( .A(n14419), .B(n14418), .Z(n14420) );
  NAND U14710 ( .A(n14421), .B(n14420), .Z(n14435) );
  OR U14711 ( .A(n14423), .B(n14422), .Z(n14427) );
  OR U14712 ( .A(n14425), .B(n14424), .Z(n14426) );
  NAND U14713 ( .A(n14427), .B(n14426), .Z(n14434) );
  XOR U14714 ( .A(n14435), .B(n14434), .Z(n14436) );
  XOR U14715 ( .A(n14437), .B(n14436), .Z(n14431) );
  XNOR U14716 ( .A(n14430), .B(n14431), .Z(N318) );
  NANDN U14717 ( .A(n14429), .B(n14428), .Z(n14433) );
  NAND U14718 ( .A(n14431), .B(n14430), .Z(n14432) );
  NAND U14719 ( .A(n14433), .B(n14432), .Z(n14603) );
  XNOR U14720 ( .A(n14603), .B(n14602), .Z(n14605) );
  OR U14721 ( .A(n14439), .B(n14438), .Z(n14443) );
  OR U14722 ( .A(n14441), .B(n14440), .Z(n14442) );
  AND U14723 ( .A(n14443), .B(n14442), .Z(n14897) );
  OR U14724 ( .A(n14445), .B(n14444), .Z(n14449) );
  NAND U14725 ( .A(n14447), .B(n14446), .Z(n14448) );
  NAND U14726 ( .A(n14449), .B(n14448), .Z(n14609) );
  OR U14727 ( .A(n14451), .B(n14450), .Z(n14455) );
  OR U14728 ( .A(n14453), .B(n14452), .Z(n14454) );
  AND U14729 ( .A(n14455), .B(n14454), .Z(n14608) );
  XOR U14730 ( .A(n14609), .B(n14608), .Z(n14610) );
  OR U14731 ( .A(n14457), .B(n14456), .Z(n14461) );
  OR U14732 ( .A(n14459), .B(n14458), .Z(n14460) );
  AND U14733 ( .A(n14461), .B(n14460), .Z(n14611) );
  OR U14734 ( .A(n14463), .B(n14462), .Z(n14467) );
  NANDN U14735 ( .A(n14465), .B(n14464), .Z(n14466) );
  AND U14736 ( .A(n14467), .B(n14466), .Z(n14881) );
  NANDN U14737 ( .A(n14469), .B(n14468), .Z(n14473) );
  OR U14738 ( .A(n14471), .B(n14470), .Z(n14472) );
  AND U14739 ( .A(n14473), .B(n14472), .Z(n14630) );
  OR U14740 ( .A(n14475), .B(n14474), .Z(n14479) );
  NANDN U14741 ( .A(n14477), .B(n14476), .Z(n14478) );
  AND U14742 ( .A(n14479), .B(n14478), .Z(n14631) );
  XOR U14743 ( .A(n14630), .B(n14631), .Z(n14628) );
  OR U14744 ( .A(n14481), .B(n14480), .Z(n14485) );
  OR U14745 ( .A(n14483), .B(n14482), .Z(n14484) );
  NAND U14746 ( .A(n14485), .B(n14484), .Z(n14629) );
  XNOR U14747 ( .A(n14628), .B(n14629), .Z(n14862) );
  NAND U14748 ( .A(x[155]), .B(y[771]), .Z(n14791) );
  NAND U14749 ( .A(x[129]), .B(y[797]), .Z(n14790) );
  XNOR U14750 ( .A(n14791), .B(n14790), .Z(n14789) );
  XNOR U14751 ( .A(n14788), .B(n14789), .Z(n14662) );
  AND U14752 ( .A(y[786]), .B(x[140]), .Z(n14490) );
  XNOR U14753 ( .A(n14490), .B(n14489), .Z(n14702) );
  XNOR U14754 ( .A(n14701), .B(n14702), .Z(n14694) );
  AND U14755 ( .A(x[138]), .B(y[788]), .Z(n14492) );
  AND U14756 ( .A(y[789]), .B(x[137]), .Z(n14491) );
  XNOR U14757 ( .A(n14492), .B(n14491), .Z(n14695) );
  XNOR U14758 ( .A(n14694), .B(n14695), .Z(n14664) );
  NANDN U14759 ( .A(n14494), .B(n14493), .Z(n14498) );
  NAND U14760 ( .A(n14496), .B(n14495), .Z(n14497) );
  AND U14761 ( .A(n14498), .B(n14497), .Z(n14665) );
  XNOR U14762 ( .A(n14664), .B(n14665), .Z(n14663) );
  XOR U14763 ( .A(n14662), .B(n14663), .Z(n14638) );
  XNOR U14764 ( .A(n14639), .B(n14638), .Z(n14637) );
  OR U14765 ( .A(n14500), .B(n14499), .Z(n14504) );
  NANDN U14766 ( .A(n14502), .B(n14501), .Z(n14503) );
  NAND U14767 ( .A(n14504), .B(n14503), .Z(n14636) );
  XOR U14768 ( .A(n14637), .B(n14636), .Z(n14863) );
  XOR U14769 ( .A(n14862), .B(n14863), .Z(n14864) );
  OR U14770 ( .A(n14506), .B(n14505), .Z(n14510) );
  OR U14771 ( .A(n14508), .B(n14507), .Z(n14509) );
  NAND U14772 ( .A(n14510), .B(n14509), .Z(n14865) );
  XOR U14773 ( .A(n14864), .B(n14865), .Z(n14880) );
  OR U14774 ( .A(n14512), .B(n14511), .Z(n14516) );
  OR U14775 ( .A(n14514), .B(n14513), .Z(n14515) );
  NAND U14776 ( .A(n14516), .B(n14515), .Z(n14885) );
  OR U14777 ( .A(n14518), .B(n14517), .Z(n14522) );
  NANDN U14778 ( .A(n14520), .B(n14519), .Z(n14521) );
  AND U14779 ( .A(n14522), .B(n14521), .Z(n14856) );
  NANDN U14780 ( .A(n14524), .B(n14523), .Z(n14528) );
  OR U14781 ( .A(n14526), .B(n14525), .Z(n14527) );
  AND U14782 ( .A(n14528), .B(n14527), .Z(n14859) );
  OR U14783 ( .A(n14530), .B(n14529), .Z(n14534) );
  OR U14784 ( .A(n14532), .B(n14531), .Z(n14533) );
  AND U14785 ( .A(n14534), .B(n14533), .Z(n14655) );
  NAND U14786 ( .A(x[134]), .B(y[792]), .Z(n14833) );
  NAND U14787 ( .A(x[133]), .B(y[793]), .Z(n14835) );
  NAND U14788 ( .A(x[147]), .B(y[779]), .Z(n14834) );
  XNOR U14789 ( .A(n14835), .B(n14834), .Z(n14832) );
  XNOR U14790 ( .A(n14833), .B(n14832), .Z(n14674) );
  OR U14791 ( .A(n14536), .B(n14535), .Z(n14540) );
  OR U14792 ( .A(n14538), .B(n14537), .Z(n14539) );
  AND U14793 ( .A(n14540), .B(n14539), .Z(n14676) );
  NAND U14794 ( .A(x[132]), .B(y[794]), .Z(n14827) );
  NAND U14795 ( .A(x[131]), .B(y[795]), .Z(n14829) );
  AND U14796 ( .A(y[780]), .B(x[146]), .Z(n14828) );
  XNOR U14797 ( .A(n14829), .B(n14828), .Z(n14826) );
  XNOR U14798 ( .A(n14827), .B(n14826), .Z(n14677) );
  XOR U14799 ( .A(n14676), .B(n14677), .Z(n14675) );
  XNOR U14800 ( .A(n14674), .B(n14675), .Z(n14654) );
  XOR U14801 ( .A(n14655), .B(n14654), .Z(n14657) );
  OR U14802 ( .A(n14542), .B(n14541), .Z(n14547) );
  NANDN U14803 ( .A(n14543), .B(o[156]), .Z(n14545) );
  NAND U14804 ( .A(x[155]), .B(y[770]), .Z(n14544) );
  AND U14805 ( .A(n14545), .B(n14544), .Z(n14546) );
  ANDN U14806 ( .B(n14547), .A(n14546), .Z(n14656) );
  XNOR U14807 ( .A(n14859), .B(n14858), .Z(n14857) );
  XNOR U14808 ( .A(n14856), .B(n14857), .Z(n14617) );
  OR U14809 ( .A(n14549), .B(n14548), .Z(n14553) );
  OR U14810 ( .A(n14551), .B(n14550), .Z(n14552) );
  NAND U14811 ( .A(n14553), .B(n14552), .Z(n14683) );
  NAND U14812 ( .A(x[148]), .B(y[778]), .Z(n14714) );
  AND U14813 ( .A(y[784]), .B(x[142]), .Z(n14713) );
  XOR U14814 ( .A(n14714), .B(n14713), .Z(n14712) );
  AND U14815 ( .A(y[790]), .B(x[136]), .Z(n14711) );
  XOR U14816 ( .A(n14712), .B(n14711), .Z(n14685) );
  NAND U14817 ( .A(y[768]), .B(x[158]), .Z(n14691) );
  NAND U14818 ( .A(x[157]), .B(y[769]), .Z(n14743) );
  XNOR U14819 ( .A(o[158]), .B(n14743), .Z(n14690) );
  XOR U14820 ( .A(n14691), .B(n14690), .Z(n14689) );
  AND U14821 ( .A(y[798]), .B(x[128]), .Z(n14688) );
  XNOR U14822 ( .A(n14689), .B(n14688), .Z(n14684) );
  XOR U14823 ( .A(n14683), .B(n14682), .Z(n14644) );
  OR U14824 ( .A(n14785), .B(n14554), .Z(n14558) );
  OR U14825 ( .A(n14556), .B(n14555), .Z(n14557) );
  AND U14826 ( .A(n14558), .B(n14557), .Z(n14645) );
  XNOR U14827 ( .A(n14644), .B(n14645), .Z(n14643) );
  OR U14828 ( .A(n14560), .B(n14559), .Z(n14564) );
  OR U14829 ( .A(n14562), .B(n14561), .Z(n14563) );
  AND U14830 ( .A(n14564), .B(n14563), .Z(n14738) );
  NAND U14831 ( .A(x[145]), .B(y[781]), .Z(n14819) );
  NAND U14832 ( .A(x[130]), .B(y[796]), .Z(n14821) );
  NAND U14833 ( .A(x[154]), .B(y[772]), .Z(n14820) );
  XNOR U14834 ( .A(n14821), .B(n14820), .Z(n14818) );
  XNOR U14835 ( .A(n14819), .B(n14818), .Z(n14739) );
  NAND U14836 ( .A(x[135]), .B(y[791]), .Z(n14707) );
  AND U14837 ( .A(y[776]), .B(x[150]), .Z(n14566) );
  AND U14838 ( .A(x[149]), .B(y[777]), .Z(n14565) );
  XNOR U14839 ( .A(n14566), .B(n14565), .Z(n14706) );
  XOR U14840 ( .A(n14707), .B(n14706), .Z(n14740) );
  XNOR U14841 ( .A(n14739), .B(n14740), .Z(n14737) );
  XOR U14842 ( .A(n14738), .B(n14737), .Z(n14642) );
  XNOR U14843 ( .A(n14643), .B(n14642), .Z(n14622) );
  NANDN U14844 ( .A(n14568), .B(n14567), .Z(n14572) );
  OR U14845 ( .A(n14570), .B(n14569), .Z(n14571) );
  NAND U14846 ( .A(n14572), .B(n14571), .Z(n14625) );
  OR U14847 ( .A(n14708), .B(n14576), .Z(n14580) );
  OR U14848 ( .A(n14578), .B(n14577), .Z(n14579) );
  AND U14849 ( .A(n14580), .B(n14579), .Z(n14668) );
  NAND U14850 ( .A(x[151]), .B(y[775]), .Z(n14784) );
  AND U14851 ( .A(y[773]), .B(x[153]), .Z(n14582) );
  AND U14852 ( .A(x[152]), .B(y[774]), .Z(n14581) );
  XNOR U14853 ( .A(n14582), .B(n14581), .Z(n14783) );
  XOR U14854 ( .A(n14784), .B(n14783), .Z(n14670) );
  NAND U14855 ( .A(n14583), .B(o[157]), .Z(n14813) );
  NAND U14856 ( .A(x[156]), .B(y[770]), .Z(n14815) );
  AND U14857 ( .A(y[782]), .B(x[144]), .Z(n14814) );
  XNOR U14858 ( .A(n14815), .B(n14814), .Z(n14812) );
  XNOR U14859 ( .A(n14813), .B(n14812), .Z(n14671) );
  XNOR U14860 ( .A(n14670), .B(n14671), .Z(n14669) );
  XOR U14861 ( .A(n14668), .B(n14669), .Z(n14650) );
  OR U14862 ( .A(n14585), .B(n14584), .Z(n14589) );
  OR U14863 ( .A(n14587), .B(n14586), .Z(n14588) );
  AND U14864 ( .A(n14589), .B(n14588), .Z(n14648) );
  XOR U14865 ( .A(n14649), .B(n14648), .Z(n14624) );
  XNOR U14866 ( .A(n14625), .B(n14624), .Z(n14623) );
  OR U14867 ( .A(n14591), .B(n14590), .Z(n14595) );
  NANDN U14868 ( .A(n14593), .B(n14592), .Z(n14594) );
  NAND U14869 ( .A(n14595), .B(n14594), .Z(n14618) );
  XNOR U14870 ( .A(n14619), .B(n14618), .Z(n14616) );
  XOR U14871 ( .A(n14617), .B(n14616), .Z(n14884) );
  XNOR U14872 ( .A(n14885), .B(n14884), .Z(n14887) );
  OR U14873 ( .A(n14597), .B(n14596), .Z(n14601) );
  OR U14874 ( .A(n14599), .B(n14598), .Z(n14600) );
  NAND U14875 ( .A(n14601), .B(n14600), .Z(n14886) );
  XOR U14876 ( .A(n14887), .B(n14886), .Z(n14878) );
  XNOR U14877 ( .A(n14879), .B(n14878), .Z(n14899) );
  XOR U14878 ( .A(n14898), .B(n14899), .Z(n14896) );
  XOR U14879 ( .A(n14897), .B(n14896), .Z(n14604) );
  XOR U14880 ( .A(n14605), .B(n14604), .Z(N319) );
  ANDN U14881 ( .B(n14603), .A(n14602), .Z(n14607) );
  ANDN U14882 ( .B(n14605), .A(n14604), .Z(n14606) );
  NOR U14883 ( .A(n14607), .B(n14606), .Z(n14615) );
  OR U14884 ( .A(n14609), .B(n14608), .Z(n14613) );
  NANDN U14885 ( .A(n14611), .B(n14610), .Z(n14612) );
  AND U14886 ( .A(n14613), .B(n14612), .Z(n14614) );
  XNOR U14887 ( .A(n14615), .B(n14614), .Z(n14895) );
  OR U14888 ( .A(n14617), .B(n14616), .Z(n14621) );
  OR U14889 ( .A(n14619), .B(n14618), .Z(n14620) );
  AND U14890 ( .A(n14621), .B(n14620), .Z(n14877) );
  NANDN U14891 ( .A(n14623), .B(n14622), .Z(n14627) );
  OR U14892 ( .A(n14625), .B(n14624), .Z(n14626) );
  AND U14893 ( .A(n14627), .B(n14626), .Z(n14635) );
  NANDN U14894 ( .A(n14629), .B(n14628), .Z(n14633) );
  OR U14895 ( .A(n14631), .B(n14630), .Z(n14632) );
  NAND U14896 ( .A(n14633), .B(n14632), .Z(n14634) );
  XNOR U14897 ( .A(n14635), .B(n14634), .Z(n14875) );
  OR U14898 ( .A(n14637), .B(n14636), .Z(n14641) );
  OR U14899 ( .A(n14639), .B(n14638), .Z(n14640) );
  AND U14900 ( .A(n14641), .B(n14640), .Z(n14873) );
  OR U14901 ( .A(n14643), .B(n14642), .Z(n14647) );
  OR U14902 ( .A(n14645), .B(n14644), .Z(n14646) );
  AND U14903 ( .A(n14647), .B(n14646), .Z(n14855) );
  OR U14904 ( .A(n14649), .B(n14648), .Z(n14653) );
  NANDN U14905 ( .A(n14651), .B(n14650), .Z(n14652) );
  AND U14906 ( .A(n14653), .B(n14652), .Z(n14661) );
  NOR U14907 ( .A(n14655), .B(n14654), .Z(n14659) );
  ANDN U14908 ( .B(n14657), .A(n14656), .Z(n14658) );
  OR U14909 ( .A(n14659), .B(n14658), .Z(n14660) );
  XNOR U14910 ( .A(n14661), .B(n14660), .Z(n14853) );
  OR U14911 ( .A(n14663), .B(n14662), .Z(n14667) );
  OR U14912 ( .A(n14665), .B(n14664), .Z(n14666) );
  AND U14913 ( .A(n14667), .B(n14666), .Z(n14851) );
  OR U14914 ( .A(n14669), .B(n14668), .Z(n14673) );
  OR U14915 ( .A(n14671), .B(n14670), .Z(n14672) );
  AND U14916 ( .A(n14673), .B(n14672), .Z(n14681) );
  NAND U14917 ( .A(n14675), .B(n14674), .Z(n14679) );
  OR U14918 ( .A(n14677), .B(n14676), .Z(n14678) );
  NAND U14919 ( .A(n14679), .B(n14678), .Z(n14680) );
  XNOR U14920 ( .A(n14681), .B(n14680), .Z(n14849) );
  OR U14921 ( .A(n14683), .B(n14682), .Z(n14687) );
  NANDN U14922 ( .A(n14685), .B(n14684), .Z(n14686) );
  AND U14923 ( .A(n14687), .B(n14686), .Z(n14847) );
  NANDN U14924 ( .A(n14689), .B(n14688), .Z(n14693) );
  NANDN U14925 ( .A(n14691), .B(n14690), .Z(n14692) );
  AND U14926 ( .A(n14693), .B(n14692), .Z(n14700) );
  NANDN U14927 ( .A(n14695), .B(n14694), .Z(n14698) );
  NAND U14928 ( .A(x[138]), .B(y[789]), .Z(n14745) );
  NANDN U14929 ( .A(n14745), .B(n14696), .Z(n14697) );
  NAND U14930 ( .A(n14698), .B(n14697), .Z(n14699) );
  XNOR U14931 ( .A(n14700), .B(n14699), .Z(n14845) );
  NANDN U14932 ( .A(n14702), .B(n14701), .Z(n14705) );
  NAND U14933 ( .A(n14703), .B(n14746), .Z(n14704) );
  AND U14934 ( .A(n14705), .B(n14704), .Z(n14736) );
  OR U14935 ( .A(n14707), .B(n14706), .Z(n14710) );
  NAND U14936 ( .A(x[150]), .B(y[777]), .Z(n14744) );
  NANDN U14937 ( .A(n14744), .B(n14708), .Z(n14709) );
  AND U14938 ( .A(n14710), .B(n14709), .Z(n14718) );
  NANDN U14939 ( .A(n14712), .B(n14711), .Z(n14716) );
  NANDN U14940 ( .A(n14714), .B(n14713), .Z(n14715) );
  NAND U14941 ( .A(n14716), .B(n14715), .Z(n14717) );
  XNOR U14942 ( .A(n14718), .B(n14717), .Z(n14734) );
  AND U14943 ( .A(y[782]), .B(x[145]), .Z(n14720) );
  NAND U14944 ( .A(x[130]), .B(y[797]), .Z(n14719) );
  XNOR U14945 ( .A(n14720), .B(n14719), .Z(n14724) );
  AND U14946 ( .A(x[146]), .B(y[781]), .Z(n14722) );
  NAND U14947 ( .A(x[133]), .B(y[794]), .Z(n14721) );
  XNOR U14948 ( .A(n14722), .B(n14721), .Z(n14723) );
  XOR U14949 ( .A(n14724), .B(n14723), .Z(n14732) );
  AND U14950 ( .A(x[159]), .B(y[768]), .Z(n14726) );
  NAND U14951 ( .A(x[132]), .B(y[795]), .Z(n14725) );
  XNOR U14952 ( .A(n14726), .B(n14725), .Z(n14730) );
  AND U14953 ( .A(y[793]), .B(x[134]), .Z(n14728) );
  NAND U14954 ( .A(x[152]), .B(y[775]), .Z(n14727) );
  XNOR U14955 ( .A(n14728), .B(n14727), .Z(n14729) );
  XNOR U14956 ( .A(n14730), .B(n14729), .Z(n14731) );
  XNOR U14957 ( .A(n14732), .B(n14731), .Z(n14733) );
  XNOR U14958 ( .A(n14734), .B(n14733), .Z(n14735) );
  XNOR U14959 ( .A(n14736), .B(n14735), .Z(n14811) );
  NANDN U14960 ( .A(n14738), .B(n14737), .Z(n14742) );
  NANDN U14961 ( .A(n14740), .B(n14739), .Z(n14741) );
  AND U14962 ( .A(n14742), .B(n14741), .Z(n14809) );
  AND U14963 ( .A(y[778]), .B(x[149]), .Z(n14752) );
  ANDN U14964 ( .B(o[158]), .A(n14743), .Z(n14750) );
  XNOR U14965 ( .A(n14744), .B(o[159]), .Z(n14748) );
  XOR U14966 ( .A(n14746), .B(n14745), .Z(n14747) );
  XNOR U14967 ( .A(n14748), .B(n14747), .Z(n14749) );
  XNOR U14968 ( .A(n14750), .B(n14749), .Z(n14751) );
  XNOR U14969 ( .A(n14752), .B(n14751), .Z(n14760) );
  AND U14970 ( .A(y[776]), .B(x[151]), .Z(n14754) );
  NAND U14971 ( .A(x[155]), .B(y[772]), .Z(n14753) );
  XNOR U14972 ( .A(n14754), .B(n14753), .Z(n14758) );
  AND U14973 ( .A(y[780]), .B(x[147]), .Z(n14756) );
  NAND U14974 ( .A(x[136]), .B(y[791]), .Z(n14755) );
  XNOR U14975 ( .A(n14756), .B(n14755), .Z(n14757) );
  XNOR U14976 ( .A(n14758), .B(n14757), .Z(n14759) );
  XNOR U14977 ( .A(n14760), .B(n14759), .Z(n14807) );
  AND U14978 ( .A(y[796]), .B(x[131]), .Z(n14762) );
  NAND U14979 ( .A(x[135]), .B(y[792]), .Z(n14761) );
  XNOR U14980 ( .A(n14762), .B(n14761), .Z(n14766) );
  AND U14981 ( .A(y[787]), .B(x[140]), .Z(n14764) );
  NAND U14982 ( .A(x[154]), .B(y[773]), .Z(n14763) );
  XNOR U14983 ( .A(n14764), .B(n14763), .Z(n14765) );
  XOR U14984 ( .A(n14766), .B(n14765), .Z(n14774) );
  AND U14985 ( .A(x[158]), .B(y[769]), .Z(n14768) );
  NAND U14986 ( .A(x[139]), .B(y[788]), .Z(n14767) );
  XNOR U14987 ( .A(n14768), .B(n14767), .Z(n14772) );
  AND U14988 ( .A(y[770]), .B(x[157]), .Z(n14770) );
  NAND U14989 ( .A(x[148]), .B(y[779]), .Z(n14769) );
  XNOR U14990 ( .A(n14770), .B(n14769), .Z(n14771) );
  XNOR U14991 ( .A(n14772), .B(n14771), .Z(n14773) );
  XNOR U14992 ( .A(n14774), .B(n14773), .Z(n14782) );
  AND U14993 ( .A(y[790]), .B(x[137]), .Z(n14776) );
  NAND U14994 ( .A(x[144]), .B(y[783]), .Z(n14775) );
  XNOR U14995 ( .A(n14776), .B(n14775), .Z(n14780) );
  AND U14996 ( .A(y[798]), .B(x[129]), .Z(n14778) );
  NAND U14997 ( .A(x[142]), .B(y[785]), .Z(n14777) );
  XNOR U14998 ( .A(n14778), .B(n14777), .Z(n14779) );
  XNOR U14999 ( .A(n14780), .B(n14779), .Z(n14781) );
  XNOR U15000 ( .A(n14782), .B(n14781), .Z(n14797) );
  OR U15001 ( .A(n14784), .B(n14783), .Z(n14787) );
  NAND U15002 ( .A(x[153]), .B(y[774]), .Z(n14803) );
  NANDN U15003 ( .A(n14803), .B(n14785), .Z(n14786) );
  AND U15004 ( .A(n14787), .B(n14786), .Z(n14795) );
  NANDN U15005 ( .A(n14789), .B(n14788), .Z(n14793) );
  OR U15006 ( .A(n14791), .B(n14790), .Z(n14792) );
  NAND U15007 ( .A(n14793), .B(n14792), .Z(n14794) );
  XNOR U15008 ( .A(n14795), .B(n14794), .Z(n14796) );
  XOR U15009 ( .A(n14797), .B(n14796), .Z(n14805) );
  AND U15010 ( .A(x[156]), .B(y[771]), .Z(n14799) );
  NAND U15011 ( .A(x[128]), .B(y[799]), .Z(n14798) );
  XNOR U15012 ( .A(n14799), .B(n14798), .Z(n14801) );
  NAND U15013 ( .A(x[143]), .B(y[784]), .Z(n14800) );
  XNOR U15014 ( .A(n14801), .B(n14800), .Z(n14802) );
  XOR U15015 ( .A(n14803), .B(n14802), .Z(n14804) );
  XNOR U15016 ( .A(n14805), .B(n14804), .Z(n14806) );
  XNOR U15017 ( .A(n14807), .B(n14806), .Z(n14808) );
  XNOR U15018 ( .A(n14809), .B(n14808), .Z(n14810) );
  XOR U15019 ( .A(n14811), .B(n14810), .Z(n14843) );
  NANDN U15020 ( .A(n14813), .B(n14812), .Z(n14817) );
  NANDN U15021 ( .A(n14815), .B(n14814), .Z(n14816) );
  AND U15022 ( .A(n14817), .B(n14816), .Z(n14825) );
  OR U15023 ( .A(n14819), .B(n14818), .Z(n14823) );
  OR U15024 ( .A(n14821), .B(n14820), .Z(n14822) );
  NAND U15025 ( .A(n14823), .B(n14822), .Z(n14824) );
  XNOR U15026 ( .A(n14825), .B(n14824), .Z(n14841) );
  NANDN U15027 ( .A(n14827), .B(n14826), .Z(n14831) );
  NANDN U15028 ( .A(n14829), .B(n14828), .Z(n14830) );
  AND U15029 ( .A(n14831), .B(n14830), .Z(n14839) );
  OR U15030 ( .A(n14833), .B(n14832), .Z(n14837) );
  OR U15031 ( .A(n14835), .B(n14834), .Z(n14836) );
  NAND U15032 ( .A(n14837), .B(n14836), .Z(n14838) );
  XNOR U15033 ( .A(n14839), .B(n14838), .Z(n14840) );
  XNOR U15034 ( .A(n14841), .B(n14840), .Z(n14842) );
  XNOR U15035 ( .A(n14843), .B(n14842), .Z(n14844) );
  XNOR U15036 ( .A(n14845), .B(n14844), .Z(n14846) );
  XNOR U15037 ( .A(n14847), .B(n14846), .Z(n14848) );
  XNOR U15038 ( .A(n14849), .B(n14848), .Z(n14850) );
  XNOR U15039 ( .A(n14851), .B(n14850), .Z(n14852) );
  XNOR U15040 ( .A(n14853), .B(n14852), .Z(n14854) );
  XNOR U15041 ( .A(n14855), .B(n14854), .Z(n14871) );
  OR U15042 ( .A(n14857), .B(n14856), .Z(n14861) );
  NOR U15043 ( .A(n14859), .B(n14858), .Z(n14860) );
  ANDN U15044 ( .B(n14861), .A(n14860), .Z(n14869) );
  ANDN U15045 ( .B(n14863), .A(n14862), .Z(n14867) );
  NOR U15046 ( .A(n14865), .B(n14864), .Z(n14866) );
  OR U15047 ( .A(n14867), .B(n14866), .Z(n14868) );
  XNOR U15048 ( .A(n14869), .B(n14868), .Z(n14870) );
  XNOR U15049 ( .A(n14871), .B(n14870), .Z(n14872) );
  XNOR U15050 ( .A(n14873), .B(n14872), .Z(n14874) );
  XNOR U15051 ( .A(n14875), .B(n14874), .Z(n14876) );
  XNOR U15052 ( .A(n14877), .B(n14876), .Z(n14893) );
  NANDN U15053 ( .A(n14879), .B(n14878), .Z(n14883) );
  NANDN U15054 ( .A(n14881), .B(n14880), .Z(n14882) );
  AND U15055 ( .A(n14883), .B(n14882), .Z(n14891) );
  OR U15056 ( .A(n14885), .B(n14884), .Z(n14889) );
  OR U15057 ( .A(n14887), .B(n14886), .Z(n14888) );
  AND U15058 ( .A(n14889), .B(n14888), .Z(n14890) );
  XNOR U15059 ( .A(n14891), .B(n14890), .Z(n14892) );
  XNOR U15060 ( .A(n14893), .B(n14892), .Z(n14894) );
  XNOR U15061 ( .A(n14895), .B(n14894), .Z(n14903) );
  NANDN U15062 ( .A(n14897), .B(n14896), .Z(n14901) );
  OR U15063 ( .A(n14899), .B(n14898), .Z(n14900) );
  NAND U15064 ( .A(n14901), .B(n14900), .Z(n14902) );
  XNOR U15065 ( .A(n14903), .B(n14902), .Z(N320) );
endmodule

