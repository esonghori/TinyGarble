
module matrixMult_N_M_3_N16_M32 ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;
  wire   N33, N34, N35, N40, N41, N42, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N57, N58, N59, N61, N62, N63, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470;

  DFF \o_reg[31]  ( .D(n12494), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \o_reg[30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \o_reg[29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \o_reg[28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \o_reg[27]  ( .D(n6253), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \o_reg[26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \o_reg[25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \o_reg[24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \o_reg[23]  ( .D(n6254), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \o_reg[22]  ( .D(n12495), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \o_reg[21]  ( .D(n6255), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \o_reg[20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \o_reg[19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \o_reg[18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \o_reg[17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \o_reg[16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \o_reg[15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \o_reg[14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \o_reg[13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \o_reg[12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \o_reg[11]  ( .D(n12496), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \o_reg[10]  ( .D(n6256), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \o_reg[9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \o_reg[8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \o_reg[7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \o_reg[6]  ( .D(n6257), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \o_reg[5]  ( .D(n12497), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \o_reg[4]  ( .D(n6258), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \o_reg[3]  ( .D(n6259), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \o_reg[2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \o_reg[1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \o_reg[0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  XNOR U6573 ( .A(n15135), .B(n15134), .Z(n15123) );
  XNOR U6574 ( .A(n13035), .B(n13034), .Z(n13036) );
  XNOR U6575 ( .A(n15121), .B(n15120), .Z(n15122) );
  XNOR U6576 ( .A(n15014), .B(n15013), .Z(n15135) );
  XNOR U6577 ( .A(n15187), .B(n15186), .Z(n15446) );
  XNOR U6578 ( .A(n13072), .B(n13071), .Z(n13074) );
  NAND U6579 ( .A(n14284), .B(n14285), .Z(n12498) );
  NANDN U6580 ( .A(n14283), .B(n14282), .Z(n12499) );
  AND U6581 ( .A(n12498), .B(n12499), .Z(n14423) );
  NAND U6582 ( .A(n13767), .B(n13036), .Z(n12500) );
  NANDN U6583 ( .A(n13035), .B(n13034), .Z(n12501) );
  AND U6584 ( .A(n12500), .B(n12501), .Z(n13139) );
  XNOR U6585 ( .A(n13282), .B(n13281), .Z(n13283) );
  XNOR U6586 ( .A(n14863), .B(n14862), .Z(n14865) );
  XNOR U6587 ( .A(n15133), .B(n15132), .Z(n15134) );
  XNOR U6588 ( .A(n15039), .B(n15038), .Z(n15043) );
  XNOR U6589 ( .A(n14948), .B(n14947), .Z(n14941) );
  XNOR U6590 ( .A(n13567), .B(n13566), .Z(n13569) );
  NAND U6591 ( .A(n14205), .B(n14204), .Z(n12502) );
  NAND U6592 ( .A(n14202), .B(n14203), .Z(n12503) );
  AND U6593 ( .A(n12502), .B(n12503), .Z(n14481) );
  XNOR U6594 ( .A(n15444), .B(n15443), .Z(n15440) );
  XNOR U6595 ( .A(n15278), .B(n15277), .Z(n15410) );
  NAND U6596 ( .A(n13463), .B(n13462), .Z(n12504) );
  NAND U6597 ( .A(n13460), .B(n13461), .Z(n12505) );
  NAND U6598 ( .A(n12504), .B(n12505), .Z(n13572) );
  XNOR U6599 ( .A(n13605), .B(n13604), .Z(n13610) );
  XNOR U6600 ( .A(n14307), .B(n14306), .Z(n14308) );
  NAND U6601 ( .A(n14281), .B(n14280), .Z(n12506) );
  NAND U6602 ( .A(n14278), .B(n14279), .Z(n12507) );
  AND U6603 ( .A(n12506), .B(n12507), .Z(n14424) );
  NAND U6604 ( .A(n13074), .B(n13073), .Z(n12508) );
  NANDN U6605 ( .A(n13072), .B(n13071), .Z(n12509) );
  AND U6606 ( .A(n12508), .B(n12509), .Z(n13130) );
  NAND U6607 ( .A(n13194), .B(n13193), .Z(n12510) );
  NANDN U6608 ( .A(n13192), .B(n13191), .Z(n12511) );
  AND U6609 ( .A(n12510), .B(n12511), .Z(n13324) );
  XNOR U6610 ( .A(n13220), .B(n13219), .Z(n13221) );
  NAND U6611 ( .A(n13384), .B(n13385), .Z(n12512) );
  NAND U6612 ( .A(n14438), .B(n13524), .Z(n12513) );
  NAND U6613 ( .A(n12512), .B(n12513), .Z(n13551) );
  NAND U6614 ( .A(n14436), .B(n14435), .Z(n12514) );
  NANDN U6615 ( .A(n14434), .B(n14433), .Z(n12515) );
  AND U6616 ( .A(n12514), .B(n12515), .Z(n14509) );
  NAND U6617 ( .A(n12818), .B(n12817), .Z(n12516) );
  NANDN U6618 ( .A(n12816), .B(n12815), .Z(n12517) );
  NAND U6619 ( .A(n12516), .B(n12517), .Z(n12865) );
  NAND U6620 ( .A(n13136), .B(n13137), .Z(n12518) );
  NANDN U6621 ( .A(n13139), .B(n13138), .Z(n12519) );
  AND U6622 ( .A(n12518), .B(n12519), .Z(n13246) );
  XOR U6623 ( .A(n13284), .B(n13283), .Z(n13275) );
  XNOR U6624 ( .A(n13349), .B(n13348), .Z(n13350) );
  XOR U6625 ( .A(n14928), .B(n14927), .Z(n14930) );
  XNOR U6626 ( .A(n15057), .B(n15056), .Z(n15059) );
  XOR U6627 ( .A(n14804), .B(n14803), .Z(n14806) );
  NAND U6628 ( .A(n12716), .B(n12655), .Z(n12520) );
  NANDN U6629 ( .A(n12657), .B(n12656), .Z(n12521) );
  AND U6630 ( .A(n12520), .B(n12521), .Z(n12691) );
  XNOR U6631 ( .A(n13449), .B(n13448), .Z(n13450) );
  XNOR U6632 ( .A(n15223), .B(n15222), .Z(n15221) );
  XOR U6633 ( .A(n15215), .B(n15214), .Z(n15213) );
  XNOR U6634 ( .A(n15141), .B(n15140), .Z(n15000) );
  XNOR U6635 ( .A(n14936), .B(n14935), .Z(n14948) );
  NAND U6636 ( .A(n13565), .B(n13564), .Z(n12522) );
  NANDN U6637 ( .A(n13563), .B(n13562), .Z(n12523) );
  NAND U6638 ( .A(n12522), .B(n12523), .Z(n13582) );
  NAND U6639 ( .A(n13983), .B(n13984), .Z(n12524) );
  NANDN U6640 ( .A(n14116), .B(n14117), .Z(n12525) );
  AND U6641 ( .A(n12524), .B(n12525), .Z(n14203) );
  XNOR U6642 ( .A(n14331), .B(n14330), .Z(n14333) );
  NAND U6643 ( .A(n14768), .B(n14769), .Z(n12526) );
  XOR U6644 ( .A(n14768), .B(n14769), .Z(n12527) );
  NANDN U6645 ( .A(n14767), .B(n12527), .Z(n12528) );
  NAND U6646 ( .A(n12526), .B(n12528), .Z(n14782) );
  XNOR U6647 ( .A(n15446), .B(n15445), .Z(n15443) );
  XNOR U6648 ( .A(n15425), .B(n15426), .Z(n15428) );
  XNOR U6649 ( .A(n15410), .B(n15409), .Z(n15408) );
  NAND U6650 ( .A(n13573), .B(n13572), .Z(n12529) );
  XOR U6651 ( .A(n13573), .B(n13572), .Z(n12530) );
  NANDN U6652 ( .A(n13574), .B(n12530), .Z(n12531) );
  NAND U6653 ( .A(n12529), .B(n12531), .Z(n13577) );
  XOR U6654 ( .A(n15462), .B(n15461), .Z(n15464) );
  XNOR U6655 ( .A(n13798), .B(n13745), .Z(n13836) );
  NAND U6656 ( .A(n13639), .B(n13638), .Z(n12532) );
  NANDN U6657 ( .A(n13637), .B(n13636), .Z(n12533) );
  AND U6658 ( .A(n12532), .B(n12533), .Z(n13928) );
  NAND U6659 ( .A(n12895), .B(n12894), .Z(n12534) );
  NANDN U6660 ( .A(n12893), .B(n12892), .Z(n12535) );
  AND U6661 ( .A(n12534), .B(n12535), .Z(n12964) );
  NAND U6662 ( .A(n13062), .B(n13063), .Z(n12536) );
  NANDN U6663 ( .A(n13065), .B(n13064), .Z(n12537) );
  AND U6664 ( .A(n12536), .B(n12537), .Z(n13106) );
  NAND U6665 ( .A(n13873), .B(n13068), .Z(n12538) );
  NANDN U6666 ( .A(n13070), .B(n13069), .Z(n12539) );
  AND U6667 ( .A(n12538), .B(n12539), .Z(n13131) );
  NAND U6668 ( .A(n13525), .B(n13526), .Z(n12540) );
  NAND U6669 ( .A(n14549), .B(n13524), .Z(n12541) );
  AND U6670 ( .A(n12540), .B(n12541), .Z(n13628) );
  NAND U6671 ( .A(n13610), .B(n13611), .Z(n12542) );
  NANDN U6672 ( .A(n13613), .B(n13612), .Z(n12543) );
  AND U6673 ( .A(n12542), .B(n12543), .Z(n14127) );
  NAND U6674 ( .A(n13711), .B(n13828), .Z(n12544) );
  NANDN U6675 ( .A(n13784), .B(n13785), .Z(n12545) );
  NAND U6676 ( .A(n12544), .B(n12545), .Z(n13713) );
  XOR U6677 ( .A(n14297), .B(n14296), .Z(n14264) );
  NAND U6678 ( .A(n14234), .B(n14235), .Z(n12546) );
  NANDN U6679 ( .A(n14237), .B(n14236), .Z(n12547) );
  AND U6680 ( .A(n12546), .B(n12547), .Z(n14349) );
  XOR U6681 ( .A(n14529), .B(n14528), .Z(n14507) );
  NAND U6682 ( .A(n14429), .B(n14430), .Z(n12548) );
  NANDN U6683 ( .A(n14432), .B(n14431), .Z(n12549) );
  AND U6684 ( .A(n12548), .B(n12549), .Z(n14688) );
  NAND U6685 ( .A(n12756), .B(n12755), .Z(n12550) );
  NAND U6686 ( .A(n13508), .B(n12754), .Z(n12551) );
  AND U6687 ( .A(n12550), .B(n12551), .Z(n12918) );
  XOR U6688 ( .A(n12871), .B(n12870), .Z(n12883) );
  NAND U6689 ( .A(n13161), .B(n13160), .Z(n12552) );
  NAND U6690 ( .A(n13159), .B(n13158), .Z(n12553) );
  AND U6691 ( .A(n12552), .B(n12553), .Z(n13253) );
  XNOR U6692 ( .A(n13351), .B(n13350), .Z(n13319) );
  NAND U6693 ( .A(n13534), .B(n13535), .Z(n12554) );
  NANDN U6694 ( .A(n13537), .B(n13536), .Z(n12555) );
  AND U6695 ( .A(n12554), .B(n12555), .Z(n13677) );
  XNOR U6696 ( .A(n15390), .B(n15389), .Z(n15388) );
  XNOR U6697 ( .A(n15285), .B(n15286), .Z(n15284) );
  XNOR U6698 ( .A(n14592), .B(n14591), .Z(n14538) );
  XNOR U6699 ( .A(n14598), .B(n14597), .Z(n14504) );
  NAND U6700 ( .A(n13165), .B(n13164), .Z(n12556) );
  NAND U6701 ( .A(n13162), .B(n13163), .Z(n12557) );
  AND U6702 ( .A(n12556), .B(n12557), .Z(n13178) );
  XNOR U6703 ( .A(n13455), .B(n13454), .Z(n13456) );
  NAND U6704 ( .A(n14607), .B(n14608), .Z(n12558) );
  NAND U6705 ( .A(n14548), .B(n14857), .Z(n12559) );
  AND U6706 ( .A(n12558), .B(n12559), .Z(n14876) );
  XOR U6707 ( .A(n14871), .B(n14870), .Z(n14818) );
  XNOR U6708 ( .A(n15043), .B(n15042), .Z(n15045) );
  XNOR U6709 ( .A(n15280), .B(n15279), .Z(n15277) );
  XNOR U6710 ( .A(n14946), .B(n14945), .Z(n14947) );
  XNOR U6711 ( .A(n13025), .B(n13024), .Z(n12956) );
  XOR U6712 ( .A(n13451), .B(n13450), .Z(n13465) );
  XOR U6713 ( .A(n14778), .B(n14777), .Z(n12560) );
  NANDN U6714 ( .A(n14776), .B(n12560), .Z(n12561) );
  NAND U6715 ( .A(n14778), .B(n14777), .Z(n12562) );
  AND U6716 ( .A(n12561), .B(n12562), .Z(n14791) );
  XNOR U6717 ( .A(n15123), .B(n15122), .Z(n15139) );
  XNOR U6718 ( .A(n15440), .B(n15439), .Z(n15438) );
  XNOR U6719 ( .A(n15422), .B(n15421), .Z(n15420) );
  XNOR U6720 ( .A(n15183), .B(n15182), .Z(n15181) );
  XNOR U6721 ( .A(n14982), .B(n14981), .Z(n14984) );
  XOR U6722 ( .A(n12605), .B(n12606), .Z(n12563) );
  NANDN U6723 ( .A(n12607), .B(n12563), .Z(n12564) );
  NAND U6724 ( .A(n12605), .B(n12606), .Z(n12565) );
  AND U6725 ( .A(n12564), .B(n12565), .Z(n15159) );
  NAND U6726 ( .A(n15155), .B(n15152), .Z(n12566) );
  NANDN U6727 ( .A(n15155), .B(n12658), .Z(n12567) );
  NANDN U6728 ( .A(n15153), .B(n12567), .Z(n12568) );
  NAND U6729 ( .A(n12566), .B(n12568), .Z(n12734) );
  XOR U6730 ( .A(n13577), .B(n13576), .Z(n12569) );
  NANDN U6731 ( .A(n13578), .B(n12569), .Z(n12570) );
  NAND U6732 ( .A(n13577), .B(n13576), .Z(n12571) );
  AND U6733 ( .A(n12570), .B(n12571), .Z(n14185) );
  NAND U6734 ( .A(n14483), .B(n14482), .Z(n12572) );
  NAND U6735 ( .A(n14480), .B(n14481), .Z(n12573) );
  AND U6736 ( .A(n12572), .B(n12573), .Z(n14767) );
  XNOR U6737 ( .A(n15171), .B(n15170), .Z(n15169) );
  AND U6738 ( .A(y[0]), .B(x[0]), .Z(n13115) );
  XOR U6739 ( .A(n13115), .B(o[0]), .Z(N33) );
  NAND U6740 ( .A(o[0]), .B(x[0]), .Z(n12574) );
  XNOR U6741 ( .A(x[1]), .B(n12574), .Z(n12575) );
  AND U6742 ( .A(y[0]), .B(n12575), .Z(n12579) );
  AND U6743 ( .A(y[1]), .B(x[0]), .Z(n12582) );
  XNOR U6744 ( .A(n12582), .B(o[1]), .Z(n12578) );
  XNOR U6745 ( .A(n12579), .B(n12578), .Z(N34) );
  NAND U6746 ( .A(n13115), .B(o[0]), .Z(n12577) );
  NAND U6747 ( .A(x[1]), .B(y[0]), .Z(n12576) );
  AND U6748 ( .A(n12577), .B(n12576), .Z(n12581) );
  NAND U6749 ( .A(n12579), .B(n12578), .Z(n12580) );
  NANDN U6750 ( .A(n12581), .B(n12580), .Z(n12607) );
  AND U6751 ( .A(x[2]), .B(y[0]), .Z(n12599) );
  AND U6752 ( .A(y[1]), .B(x[1]), .Z(n12600) );
  XOR U6753 ( .A(n12599), .B(n12600), .Z(n12602) );
  AND U6754 ( .A(n12582), .B(o[1]), .Z(n12601) );
  XOR U6755 ( .A(n12602), .B(n12601), .Z(n12605) );
  AND U6756 ( .A(y[2]), .B(x[0]), .Z(n12589) );
  XOR U6757 ( .A(n12589), .B(o[2]), .Z(n12606) );
  XOR U6758 ( .A(n12605), .B(n12606), .Z(n12583) );
  XNOR U6759 ( .A(n12607), .B(n12583), .Z(N35) );
  AND U6760 ( .A(x[0]), .B(y[4]), .Z(n12585) );
  NAND U6761 ( .A(y[0]), .B(x[4]), .Z(n12584) );
  XNOR U6762 ( .A(n12585), .B(n12584), .Z(n12629) );
  NAND U6763 ( .A(y[1]), .B(x[2]), .Z(n12594) );
  ANDN U6764 ( .B(o[3]), .A(n12594), .Z(n12628) );
  XOR U6765 ( .A(n12629), .B(n12628), .Z(n12618) );
  NAND U6766 ( .A(y[1]), .B(x[3]), .Z(n12623) );
  XNOR U6767 ( .A(o[4]), .B(n12623), .Z(n12625) );
  AND U6768 ( .A(y[3]), .B(x[1]), .Z(n12781) );
  NAND U6769 ( .A(x[2]), .B(y[2]), .Z(n12586) );
  XNOR U6770 ( .A(n12781), .B(n12586), .Z(n12624) );
  XNOR U6771 ( .A(n12625), .B(n12624), .Z(n12617) );
  XNOR U6772 ( .A(n12618), .B(n12617), .Z(n12619) );
  AND U6773 ( .A(x[3]), .B(y[3]), .Z(n12639) );
  NAND U6774 ( .A(n13115), .B(n12639), .Z(n12591) );
  AND U6775 ( .A(y[3]), .B(x[0]), .Z(n12588) );
  NAND U6776 ( .A(y[0]), .B(x[3]), .Z(n12587) );
  XOR U6777 ( .A(n12588), .B(n12587), .Z(n12592) );
  AND U6778 ( .A(n12589), .B(o[2]), .Z(n12593) );
  NANDN U6779 ( .A(n12592), .B(n12593), .Z(n12590) );
  NAND U6780 ( .A(n12591), .B(n12590), .Z(n12620) );
  XOR U6781 ( .A(n12619), .B(n12620), .Z(n12613) );
  XOR U6782 ( .A(n12593), .B(n12592), .Z(n12595) );
  XNOR U6783 ( .A(o[3]), .B(n12594), .Z(n12596) );
  NANDN U6784 ( .A(n12595), .B(n12596), .Z(n12598) );
  XOR U6785 ( .A(n12596), .B(n12595), .Z(n12609) );
  AND U6786 ( .A(y[2]), .B(x[1]), .Z(n12703) );
  NANDN U6787 ( .A(n12609), .B(n12703), .Z(n12597) );
  AND U6788 ( .A(n12598), .B(n12597), .Z(n12614) );
  NANDN U6789 ( .A(n12613), .B(n12614), .Z(n12616) );
  NAND U6790 ( .A(n12600), .B(n12599), .Z(n12604) );
  NAND U6791 ( .A(n12602), .B(n12601), .Z(n12603) );
  AND U6792 ( .A(n12604), .B(n12603), .Z(n12608) );
  IV U6793 ( .A(n12608), .Z(n15158) );
  NANDN U6794 ( .A(n15158), .B(n15159), .Z(n12612) );
  NOR U6795 ( .A(n12608), .B(n15159), .Z(n12610) );
  XNOR U6796 ( .A(n12703), .B(n12609), .Z(n15161) );
  OR U6797 ( .A(n12610), .B(n15161), .Z(n12611) );
  AND U6798 ( .A(n12612), .B(n12611), .Z(n15157) );
  XNOR U6799 ( .A(n12614), .B(n12613), .Z(n15156) );
  NANDN U6800 ( .A(n15157), .B(n15156), .Z(n12615) );
  NAND U6801 ( .A(n12616), .B(n12615), .Z(n12632) );
  NANDN U6802 ( .A(n12618), .B(n12617), .Z(n12622) );
  NANDN U6803 ( .A(n12620), .B(n12619), .Z(n12621) );
  AND U6804 ( .A(n12622), .B(n12621), .Z(n12633) );
  NANDN U6805 ( .A(n12632), .B(n12633), .Z(n12635) );
  AND U6806 ( .A(y[5]), .B(x[0]), .Z(n12643) );
  NAND U6807 ( .A(y[0]), .B(x[5]), .Z(n12644) );
  XNOR U6808 ( .A(n12643), .B(n12644), .Z(n12646) );
  ANDN U6809 ( .B(o[4]), .A(n12623), .Z(n12645) );
  XOR U6810 ( .A(n12646), .B(n12645), .Z(n12657) );
  NAND U6811 ( .A(x[2]), .B(y[3]), .Z(n12716) );
  AND U6812 ( .A(y[2]), .B(x[3]), .Z(n12650) );
  AND U6813 ( .A(y[4]), .B(x[1]), .Z(n12649) );
  XOR U6814 ( .A(n12650), .B(n12649), .Z(n12652) );
  NAND U6815 ( .A(x[4]), .B(y[1]), .Z(n12642) );
  XNOR U6816 ( .A(o[5]), .B(n12642), .Z(n12651) );
  XNOR U6817 ( .A(n12652), .B(n12651), .Z(n12655) );
  XOR U6818 ( .A(n12716), .B(n12655), .Z(n12656) );
  XOR U6819 ( .A(n12657), .B(n12656), .Z(n12661) );
  NANDN U6820 ( .A(n12716), .B(n12703), .Z(n12627) );
  NAND U6821 ( .A(n12625), .B(n12624), .Z(n12626) );
  NAND U6822 ( .A(n12627), .B(n12626), .Z(n12660) );
  AND U6823 ( .A(x[4]), .B(y[4]), .Z(n13425) );
  NAND U6824 ( .A(n13425), .B(n13115), .Z(n12631) );
  NAND U6825 ( .A(n12629), .B(n12628), .Z(n12630) );
  NAND U6826 ( .A(n12631), .B(n12630), .Z(n12659) );
  XOR U6827 ( .A(n12660), .B(n12659), .Z(n12662) );
  XOR U6828 ( .A(n12661), .B(n12662), .Z(n15163) );
  XNOR U6829 ( .A(n12633), .B(n12632), .Z(n15162) );
  NAND U6830 ( .A(n15163), .B(n15162), .Z(n12634) );
  AND U6831 ( .A(n12635), .B(n12634), .Z(n12658) );
  IV U6832 ( .A(n12658), .Z(n15152) );
  AND U6833 ( .A(x[1]), .B(y[5]), .Z(n12637) );
  NAND U6834 ( .A(y[2]), .B(x[4]), .Z(n12636) );
  XNOR U6835 ( .A(n12637), .B(n12636), .Z(n12670) );
  NAND U6836 ( .A(y[1]), .B(x[5]), .Z(n12667) );
  XOR U6837 ( .A(o[6]), .B(n12667), .Z(n12671) );
  XNOR U6838 ( .A(n12670), .B(n12671), .Z(n12677) );
  NAND U6839 ( .A(x[2]), .B(y[4]), .Z(n12638) );
  XNOR U6840 ( .A(n12639), .B(n12638), .Z(n12676) );
  XOR U6841 ( .A(n12677), .B(n12676), .Z(n12687) );
  AND U6842 ( .A(y[0]), .B(x[6]), .Z(n12641) );
  NAND U6843 ( .A(x[0]), .B(y[6]), .Z(n12640) );
  XNOR U6844 ( .A(n12641), .B(n12640), .Z(n12682) );
  ANDN U6845 ( .B(o[5]), .A(n12642), .Z(n12681) );
  XOR U6846 ( .A(n12682), .B(n12681), .Z(n12686) );
  NANDN U6847 ( .A(n12644), .B(n12643), .Z(n12648) );
  NAND U6848 ( .A(n12646), .B(n12645), .Z(n12647) );
  AND U6849 ( .A(n12648), .B(n12647), .Z(n12685) );
  XOR U6850 ( .A(n12686), .B(n12685), .Z(n12688) );
  XOR U6851 ( .A(n12687), .B(n12688), .Z(n12694) );
  NAND U6852 ( .A(n12650), .B(n12649), .Z(n12654) );
  NAND U6853 ( .A(n12652), .B(n12651), .Z(n12653) );
  AND U6854 ( .A(n12654), .B(n12653), .Z(n12692) );
  XNOR U6855 ( .A(n12692), .B(n12691), .Z(n12693) );
  XOR U6856 ( .A(n12694), .B(n12693), .Z(n15153) );
  NAND U6857 ( .A(n12660), .B(n12659), .Z(n12664) );
  NAND U6858 ( .A(n12662), .B(n12661), .Z(n12663) );
  NAND U6859 ( .A(n12664), .B(n12663), .Z(n15155) );
  AND U6860 ( .A(y[7]), .B(x[0]), .Z(n12666) );
  NAND U6861 ( .A(y[0]), .B(x[7]), .Z(n12665) );
  XNOR U6862 ( .A(n12666), .B(n12665), .Z(n12722) );
  ANDN U6863 ( .B(o[6]), .A(n12667), .Z(n12721) );
  XOR U6864 ( .A(n12722), .B(n12721), .Z(n12711) );
  AND U6865 ( .A(x[2]), .B(y[5]), .Z(n12669) );
  NAND U6866 ( .A(y[3]), .B(x[4]), .Z(n12668) );
  XNOR U6867 ( .A(n12669), .B(n12668), .Z(n12718) );
  AND U6868 ( .A(y[4]), .B(x[3]), .Z(n12717) );
  XNOR U6869 ( .A(n12718), .B(n12717), .Z(n12710) );
  XNOR U6870 ( .A(n12711), .B(n12710), .Z(n12713) );
  AND U6871 ( .A(x[4]), .B(y[5]), .Z(n13186) );
  NAND U6872 ( .A(n13186), .B(n12703), .Z(n12673) );
  NANDN U6873 ( .A(n12671), .B(n12670), .Z(n12672) );
  AND U6874 ( .A(n12673), .B(n12672), .Z(n12712) );
  XOR U6875 ( .A(n12713), .B(n12712), .Z(n12698) );
  AND U6876 ( .A(x[5]), .B(y[2]), .Z(n12675) );
  NAND U6877 ( .A(x[1]), .B(y[6]), .Z(n12674) );
  XNOR U6878 ( .A(n12675), .B(n12674), .Z(n12706) );
  NAND U6879 ( .A(x[6]), .B(y[1]), .Z(n12709) );
  XNOR U6880 ( .A(o[7]), .B(n12709), .Z(n12705) );
  XOR U6881 ( .A(n12706), .B(n12705), .Z(n12726) );
  NANDN U6882 ( .A(n12716), .B(n12717), .Z(n12679) );
  NAND U6883 ( .A(n12677), .B(n12676), .Z(n12678) );
  AND U6884 ( .A(n12679), .B(n12678), .Z(n12725) );
  XNOR U6885 ( .A(n12726), .B(n12725), .Z(n12728) );
  AND U6886 ( .A(y[6]), .B(x[6]), .Z(n12680) );
  NAND U6887 ( .A(n13115), .B(n12680), .Z(n12684) );
  NAND U6888 ( .A(n12682), .B(n12681), .Z(n12683) );
  AND U6889 ( .A(n12684), .B(n12683), .Z(n12727) );
  XNOR U6890 ( .A(n12728), .B(n12727), .Z(n12697) );
  XNOR U6891 ( .A(n12698), .B(n12697), .Z(n12700) );
  NANDN U6892 ( .A(n12686), .B(n12685), .Z(n12690) );
  OR U6893 ( .A(n12688), .B(n12687), .Z(n12689) );
  AND U6894 ( .A(n12690), .B(n12689), .Z(n12699) );
  XOR U6895 ( .A(n12700), .B(n12699), .Z(n12732) );
  NANDN U6896 ( .A(n12692), .B(n12691), .Z(n12696) );
  NANDN U6897 ( .A(n12694), .B(n12693), .Z(n12695) );
  AND U6898 ( .A(n12696), .B(n12695), .Z(n12731) );
  XNOR U6899 ( .A(n12732), .B(n12731), .Z(n12733) );
  XOR U6900 ( .A(n12734), .B(n12733), .Z(N40) );
  NANDN U6901 ( .A(n12698), .B(n12697), .Z(n12702) );
  NAND U6902 ( .A(n12700), .B(n12699), .Z(n12701) );
  AND U6903 ( .A(n12702), .B(n12701), .Z(n12776) );
  AND U6904 ( .A(y[6]), .B(x[5]), .Z(n12704) );
  NAND U6905 ( .A(n12704), .B(n12703), .Z(n12708) );
  NAND U6906 ( .A(n12706), .B(n12705), .Z(n12707) );
  AND U6907 ( .A(n12708), .B(n12707), .Z(n12764) );
  ANDN U6908 ( .B(o[7]), .A(n12709), .Z(n12738) );
  NAND U6909 ( .A(x[5]), .B(y[3]), .Z(n13310) );
  NAND U6910 ( .A(x[1]), .B(y[7]), .Z(n12737) );
  XOR U6911 ( .A(n13310), .B(n12737), .Z(n12739) );
  XNOR U6912 ( .A(n12738), .B(n12739), .Z(n12756) );
  NAND U6913 ( .A(y[5]), .B(x[3]), .Z(n13508) );
  AND U6914 ( .A(y[6]), .B(x[2]), .Z(n13603) );
  AND U6915 ( .A(x[6]), .B(y[2]), .Z(n12750) );
  XOR U6916 ( .A(n13603), .B(n12750), .Z(n12751) );
  XNOR U6917 ( .A(n13425), .B(n12751), .Z(n12754) );
  XOR U6918 ( .A(n13508), .B(n12754), .Z(n12755) );
  XNOR U6919 ( .A(n12756), .B(n12755), .Z(n12763) );
  XNOR U6920 ( .A(n12764), .B(n12763), .Z(n12766) );
  NANDN U6921 ( .A(n12711), .B(n12710), .Z(n12715) );
  NAND U6922 ( .A(n12713), .B(n12712), .Z(n12714) );
  AND U6923 ( .A(n12715), .B(n12714), .Z(n12765) );
  XOR U6924 ( .A(n12766), .B(n12765), .Z(n12771) );
  NANDN U6925 ( .A(n12716), .B(n13186), .Z(n12720) );
  NAND U6926 ( .A(n12718), .B(n12717), .Z(n12719) );
  AND U6927 ( .A(n12720), .B(n12719), .Z(n12759) );
  AND U6928 ( .A(x[7]), .B(y[7]), .Z(n13041) );
  NAND U6929 ( .A(n13041), .B(n13115), .Z(n12724) );
  NAND U6930 ( .A(n12722), .B(n12721), .Z(n12723) );
  AND U6931 ( .A(n12724), .B(n12723), .Z(n12758) );
  NAND U6932 ( .A(x[7]), .B(y[1]), .Z(n12743) );
  XNOR U6933 ( .A(o[8]), .B(n12743), .Z(n12746) );
  AND U6934 ( .A(x[0]), .B(y[8]), .Z(n12744) );
  NAND U6935 ( .A(x[8]), .B(y[0]), .Z(n12745) );
  XOR U6936 ( .A(n12744), .B(n12745), .Z(n12747) );
  XNOR U6937 ( .A(n12746), .B(n12747), .Z(n12757) );
  XOR U6938 ( .A(n12758), .B(n12757), .Z(n12760) );
  XOR U6939 ( .A(n12759), .B(n12760), .Z(n12770) );
  NANDN U6940 ( .A(n12726), .B(n12725), .Z(n12730) );
  NAND U6941 ( .A(n12728), .B(n12727), .Z(n12729) );
  NAND U6942 ( .A(n12730), .B(n12729), .Z(n12769) );
  XOR U6943 ( .A(n12770), .B(n12769), .Z(n12772) );
  XNOR U6944 ( .A(n12771), .B(n12772), .Z(n12775) );
  XNOR U6945 ( .A(n12776), .B(n12775), .Z(n12778) );
  NANDN U6946 ( .A(n12732), .B(n12731), .Z(n12736) );
  NANDN U6947 ( .A(n12734), .B(n12733), .Z(n12735) );
  AND U6948 ( .A(n12736), .B(n12735), .Z(n12777) );
  XOR U6949 ( .A(n12778), .B(n12777), .Z(N41) );
  NAND U6950 ( .A(n13310), .B(n12737), .Z(n12741) );
  ANDN U6951 ( .B(n12739), .A(n12738), .Z(n12740) );
  ANDN U6952 ( .B(n12741), .A(n12740), .Z(n12852) );
  AND U6953 ( .A(y[8]), .B(x[1]), .Z(n13524) );
  NAND U6954 ( .A(y[3]), .B(x[6]), .Z(n12742) );
  XNOR U6955 ( .A(n13524), .B(n12742), .Z(n12782) );
  XOR U6956 ( .A(n13186), .B(n12782), .Z(n12839) );
  AND U6957 ( .A(x[2]), .B(y[7]), .Z(n13372) );
  NAND U6958 ( .A(y[6]), .B(x[3]), .Z(n13121) );
  XNOR U6959 ( .A(n13372), .B(n13121), .Z(n12840) );
  XNOR U6960 ( .A(n12839), .B(n12840), .Z(n12851) );
  XNOR U6961 ( .A(n12852), .B(n12851), .Z(n12854) );
  AND U6962 ( .A(x[7]), .B(y[2]), .Z(n13151) );
  NAND U6963 ( .A(y[4]), .B(x[5]), .Z(n12794) );
  XNOR U6964 ( .A(n13151), .B(n12794), .Z(n12796) );
  ANDN U6965 ( .B(o[8]), .A(n12743), .Z(n12795) );
  XOR U6966 ( .A(n12796), .B(n12795), .Z(n12844) );
  AND U6967 ( .A(y[9]), .B(x[0]), .Z(n12786) );
  NAND U6968 ( .A(y[0]), .B(x[9]), .Z(n12787) );
  XNOR U6969 ( .A(n12786), .B(n12787), .Z(n12789) );
  NAND U6970 ( .A(x[8]), .B(y[1]), .Z(n12785) );
  XNOR U6971 ( .A(o[9]), .B(n12785), .Z(n12788) );
  XNOR U6972 ( .A(n12789), .B(n12788), .Z(n12843) );
  XNOR U6973 ( .A(n12844), .B(n12843), .Z(n12845) );
  NANDN U6974 ( .A(n12745), .B(n12744), .Z(n12749) );
  NANDN U6975 ( .A(n12747), .B(n12746), .Z(n12748) );
  NAND U6976 ( .A(n12749), .B(n12748), .Z(n12846) );
  XNOR U6977 ( .A(n12845), .B(n12846), .Z(n12853) );
  XOR U6978 ( .A(n12854), .B(n12853), .Z(n12920) );
  NAND U6979 ( .A(n13603), .B(n12750), .Z(n12753) );
  NAND U6980 ( .A(n13425), .B(n12751), .Z(n12752) );
  AND U6981 ( .A(n12753), .B(n12752), .Z(n12919) );
  XOR U6982 ( .A(n12919), .B(n12918), .Z(n12921) );
  XOR U6983 ( .A(n12920), .B(n12921), .Z(n12930) );
  NANDN U6984 ( .A(n12758), .B(n12757), .Z(n12762) );
  OR U6985 ( .A(n12760), .B(n12759), .Z(n12761) );
  AND U6986 ( .A(n12762), .B(n12761), .Z(n12928) );
  NANDN U6987 ( .A(n12764), .B(n12763), .Z(n12768) );
  NAND U6988 ( .A(n12766), .B(n12765), .Z(n12767) );
  NAND U6989 ( .A(n12768), .B(n12767), .Z(n12929) );
  XOR U6990 ( .A(n12928), .B(n12929), .Z(n12931) );
  XOR U6991 ( .A(n12930), .B(n12931), .Z(n12937) );
  NANDN U6992 ( .A(n12770), .B(n12769), .Z(n12774) );
  OR U6993 ( .A(n12772), .B(n12771), .Z(n12773) );
  AND U6994 ( .A(n12774), .B(n12773), .Z(n12936) );
  XNOR U6995 ( .A(n12937), .B(n12936), .Z(n12939) );
  NANDN U6996 ( .A(n12776), .B(n12775), .Z(n12780) );
  NAND U6997 ( .A(n12778), .B(n12777), .Z(n12779) );
  NAND U6998 ( .A(n12780), .B(n12779), .Z(n12938) );
  XOR U6999 ( .A(n12939), .B(n12938), .Z(N42) );
  NAND U7000 ( .A(x[6]), .B(y[8]), .Z(n13158) );
  NANDN U7001 ( .A(n13158), .B(n12781), .Z(n12784) );
  NAND U7002 ( .A(n13186), .B(n12782), .Z(n12783) );
  AND U7003 ( .A(n12784), .B(n12783), .Z(n12804) );
  AND U7004 ( .A(x[3]), .B(y[7]), .Z(n13789) );
  AND U7005 ( .A(y[9]), .B(x[1]), .Z(n13822) );
  XOR U7006 ( .A(n13789), .B(n13822), .Z(n12829) );
  NAND U7007 ( .A(x[2]), .B(y[8]), .Z(n12830) );
  XNOR U7008 ( .A(n12829), .B(n12830), .Z(n12803) );
  XNOR U7009 ( .A(n12804), .B(n12803), .Z(n12806) );
  AND U7010 ( .A(y[10]), .B(x[0]), .Z(n12815) );
  NAND U7011 ( .A(x[10]), .B(y[0]), .Z(n12816) );
  XNOR U7012 ( .A(n12815), .B(n12816), .Z(n12818) );
  ANDN U7013 ( .B(o[9]), .A(n12785), .Z(n12817) );
  XOR U7014 ( .A(n12818), .B(n12817), .Z(n12805) );
  XOR U7015 ( .A(n12806), .B(n12805), .Z(n12800) );
  NANDN U7016 ( .A(n12787), .B(n12786), .Z(n12791) );
  NAND U7017 ( .A(n12789), .B(n12788), .Z(n12790) );
  AND U7018 ( .A(n12791), .B(n12790), .Z(n12799) );
  NANDN U7019 ( .A(n12800), .B(n12799), .Z(n12802) );
  AND U7020 ( .A(y[3]), .B(x[7]), .Z(n12793) );
  NAND U7021 ( .A(y[6]), .B(x[4]), .Z(n12792) );
  XNOR U7022 ( .A(n12793), .B(n12792), .Z(n12811) );
  AND U7023 ( .A(x[6]), .B(y[4]), .Z(n12810) );
  XOR U7024 ( .A(n12811), .B(n12810), .Z(n12820) );
  NAND U7025 ( .A(y[1]), .B(x[9]), .Z(n12814) );
  XNOR U7026 ( .A(o[10]), .B(n12814), .Z(n12833) );
  NAND U7027 ( .A(x[8]), .B(y[2]), .Z(n12834) );
  XNOR U7028 ( .A(n12833), .B(n12834), .Z(n12836) );
  AND U7029 ( .A(y[5]), .B(x[5]), .Z(n12835) );
  XNOR U7030 ( .A(n12836), .B(n12835), .Z(n12819) );
  XNOR U7031 ( .A(n12820), .B(n12819), .Z(n12821) );
  NANDN U7032 ( .A(n12794), .B(n13151), .Z(n12798) );
  NAND U7033 ( .A(n12796), .B(n12795), .Z(n12797) );
  NAND U7034 ( .A(n12798), .B(n12797), .Z(n12822) );
  XNOR U7035 ( .A(n12821), .B(n12822), .Z(n12927) );
  XNOR U7036 ( .A(n12800), .B(n12799), .Z(n12926) );
  NAND U7037 ( .A(n12927), .B(n12926), .Z(n12801) );
  AND U7038 ( .A(n12802), .B(n12801), .Z(n12860) );
  NANDN U7039 ( .A(n12804), .B(n12803), .Z(n12808) );
  NAND U7040 ( .A(n12806), .B(n12805), .Z(n12807) );
  AND U7041 ( .A(n12808), .B(n12807), .Z(n12877) );
  NAND U7042 ( .A(y[6]), .B(x[7]), .Z(n13072) );
  AND U7043 ( .A(x[4]), .B(y[3]), .Z(n12809) );
  NANDN U7044 ( .A(n13072), .B(n12809), .Z(n12813) );
  NAND U7045 ( .A(n12811), .B(n12810), .Z(n12812) );
  AND U7046 ( .A(n12813), .B(n12812), .Z(n12875) );
  AND U7047 ( .A(x[10]), .B(y[1]), .Z(n12887) );
  XOR U7048 ( .A(n12887), .B(o[11]), .Z(n12909) );
  AND U7049 ( .A(y[10]), .B(x[1]), .Z(n12907) );
  NAND U7050 ( .A(x[6]), .B(y[5]), .Z(n12906) );
  XNOR U7051 ( .A(n12907), .B(n12906), .Z(n12908) );
  XOR U7052 ( .A(n12909), .B(n12908), .Z(n12863) );
  AND U7053 ( .A(y[11]), .B(x[0]), .Z(n12892) );
  NAND U7054 ( .A(x[11]), .B(y[0]), .Z(n12893) );
  XNOR U7055 ( .A(n12892), .B(n12893), .Z(n12895) );
  ANDN U7056 ( .B(o[10]), .A(n12814), .Z(n12894) );
  XOR U7057 ( .A(n12895), .B(n12894), .Z(n12864) );
  XOR U7058 ( .A(n12863), .B(n12864), .Z(n12866) );
  XOR U7059 ( .A(n12866), .B(n12865), .Z(n12874) );
  XNOR U7060 ( .A(n12875), .B(n12874), .Z(n12876) );
  XNOR U7061 ( .A(n12877), .B(n12876), .Z(n12915) );
  NANDN U7062 ( .A(n12820), .B(n12819), .Z(n12824) );
  NANDN U7063 ( .A(n12822), .B(n12821), .Z(n12823) );
  AND U7064 ( .A(n12824), .B(n12823), .Z(n12912) );
  AND U7065 ( .A(x[9]), .B(y[2]), .Z(n12826) );
  NAND U7066 ( .A(x[7]), .B(y[4]), .Z(n12825) );
  XNOR U7067 ( .A(n12826), .B(n12825), .Z(n12888) );
  NAND U7068 ( .A(x[8]), .B(y[3]), .Z(n12889) );
  XOR U7069 ( .A(n12888), .B(n12889), .Z(n12870) );
  NAND U7070 ( .A(x[3]), .B(y[8]), .Z(n13689) );
  AND U7071 ( .A(x[2]), .B(y[9]), .Z(n12828) );
  NAND U7072 ( .A(x[5]), .B(y[6]), .Z(n12827) );
  XNOR U7073 ( .A(n12828), .B(n12827), .Z(n12902) );
  NAND U7074 ( .A(x[4]), .B(y[7]), .Z(n12903) );
  XOR U7075 ( .A(n12902), .B(n12903), .Z(n12869) );
  XNOR U7076 ( .A(n13689), .B(n12869), .Z(n12871) );
  NAND U7077 ( .A(n13822), .B(n13789), .Z(n12832) );
  NANDN U7078 ( .A(n12830), .B(n12829), .Z(n12831) );
  AND U7079 ( .A(n12832), .B(n12831), .Z(n12881) );
  NANDN U7080 ( .A(n12834), .B(n12833), .Z(n12838) );
  NAND U7081 ( .A(n12836), .B(n12835), .Z(n12837) );
  NAND U7082 ( .A(n12838), .B(n12837), .Z(n12880) );
  XNOR U7083 ( .A(n12881), .B(n12880), .Z(n12882) );
  XNOR U7084 ( .A(n12883), .B(n12882), .Z(n12913) );
  XNOR U7085 ( .A(n12912), .B(n12913), .Z(n12914) );
  XNOR U7086 ( .A(n12915), .B(n12914), .Z(n12859) );
  NANDN U7087 ( .A(n12860), .B(n12859), .Z(n12862) );
  NANDN U7088 ( .A(n13372), .B(n13121), .Z(n12842) );
  ANDN U7089 ( .B(n12840), .A(n12839), .Z(n12841) );
  ANDN U7090 ( .B(n12842), .A(n12841), .Z(n12850) );
  NANDN U7091 ( .A(n12844), .B(n12843), .Z(n12848) );
  NANDN U7092 ( .A(n12846), .B(n12845), .Z(n12847) );
  NAND U7093 ( .A(n12848), .B(n12847), .Z(n12849) );
  NANDN U7094 ( .A(n12850), .B(n12849), .Z(n12858) );
  XOR U7095 ( .A(n12850), .B(n12849), .Z(n12924) );
  NANDN U7096 ( .A(n12852), .B(n12851), .Z(n12856) );
  NAND U7097 ( .A(n12854), .B(n12853), .Z(n12855) );
  AND U7098 ( .A(n12856), .B(n12855), .Z(n12925) );
  OR U7099 ( .A(n12924), .B(n12925), .Z(n12857) );
  AND U7100 ( .A(n12858), .B(n12857), .Z(n12953) );
  XNOR U7101 ( .A(n12860), .B(n12859), .Z(n12952) );
  NANDN U7102 ( .A(n12953), .B(n12952), .Z(n12861) );
  AND U7103 ( .A(n12862), .B(n12861), .Z(n12957) );
  NAND U7104 ( .A(n12864), .B(n12863), .Z(n12868) );
  NAND U7105 ( .A(n12866), .B(n12865), .Z(n12867) );
  AND U7106 ( .A(n12868), .B(n12867), .Z(n13018) );
  NAND U7107 ( .A(n13689), .B(n12869), .Z(n12873) );
  NANDN U7108 ( .A(n12871), .B(n12870), .Z(n12872) );
  AND U7109 ( .A(n12873), .B(n12872), .Z(n13017) );
  NANDN U7110 ( .A(n12875), .B(n12874), .Z(n12879) );
  NANDN U7111 ( .A(n12877), .B(n12876), .Z(n12878) );
  AND U7112 ( .A(n12879), .B(n12878), .Z(n13016) );
  XOR U7113 ( .A(n13017), .B(n13016), .Z(n13019) );
  XNOR U7114 ( .A(n13018), .B(n13019), .Z(n13024) );
  NANDN U7115 ( .A(n12881), .B(n12880), .Z(n12885) );
  NAND U7116 ( .A(n12883), .B(n12882), .Z(n12884) );
  AND U7117 ( .A(n12885), .B(n12884), .Z(n13013) );
  AND U7118 ( .A(x[1]), .B(y[11]), .Z(n13646) );
  NAND U7119 ( .A(x[6]), .B(y[6]), .Z(n12886) );
  XNOR U7120 ( .A(n13646), .B(n12886), .Z(n12979) );
  AND U7121 ( .A(n12887), .B(o[11]), .Z(n12978) );
  XOR U7122 ( .A(n12979), .B(n12978), .Z(n12963) );
  NAND U7123 ( .A(y[4]), .B(x[9]), .Z(n13035) );
  NANDN U7124 ( .A(n13035), .B(n13151), .Z(n12891) );
  NANDN U7125 ( .A(n12889), .B(n12888), .Z(n12890) );
  AND U7126 ( .A(n12891), .B(n12890), .Z(n12962) );
  XNOR U7127 ( .A(n12963), .B(n12962), .Z(n12965) );
  XOR U7128 ( .A(n12965), .B(n12964), .Z(n13011) );
  AND U7129 ( .A(y[4]), .B(x[8]), .Z(n12897) );
  NAND U7130 ( .A(x[2]), .B(y[10]), .Z(n12896) );
  XNOR U7131 ( .A(n12897), .B(n12896), .Z(n13006) );
  AND U7132 ( .A(y[9]), .B(x[3]), .Z(n13005) );
  XOR U7133 ( .A(n13006), .B(n13005), .Z(n12999) );
  AND U7134 ( .A(x[0]), .B(y[12]), .Z(n12899) );
  NAND U7135 ( .A(y[0]), .B(x[12]), .Z(n12898) );
  XNOR U7136 ( .A(n12899), .B(n12898), .Z(n12983) );
  NAND U7137 ( .A(x[11]), .B(y[1]), .Z(n13009) );
  XNOR U7138 ( .A(o[12]), .B(n13009), .Z(n12982) );
  XNOR U7139 ( .A(n12983), .B(n12982), .Z(n12998) );
  XNOR U7140 ( .A(n12999), .B(n12998), .Z(n13001) );
  AND U7141 ( .A(x[9]), .B(y[3]), .Z(n13598) );
  AND U7142 ( .A(y[2]), .B(x[10]), .Z(n12901) );
  NAND U7143 ( .A(y[8]), .B(x[4]), .Z(n12900) );
  XOR U7144 ( .A(n12901), .B(n12900), .Z(n12970) );
  XOR U7145 ( .A(n13598), .B(n12970), .Z(n12994) );
  NAND U7146 ( .A(x[5]), .B(y[7]), .Z(n12993) );
  NAND U7147 ( .A(y[5]), .B(x[7]), .Z(n12992) );
  XOR U7148 ( .A(n12993), .B(n12992), .Z(n12995) );
  XOR U7149 ( .A(n12994), .B(n12995), .Z(n13000) );
  XOR U7150 ( .A(n13001), .B(n13000), .Z(n12989) );
  AND U7151 ( .A(y[9]), .B(x[5]), .Z(n13379) );
  NAND U7152 ( .A(n13603), .B(n13379), .Z(n12905) );
  NANDN U7153 ( .A(n12903), .B(n12902), .Z(n12904) );
  AND U7154 ( .A(n12905), .B(n12904), .Z(n12987) );
  NANDN U7155 ( .A(n12907), .B(n12906), .Z(n12911) );
  NANDN U7156 ( .A(n12909), .B(n12908), .Z(n12910) );
  AND U7157 ( .A(n12911), .B(n12910), .Z(n12986) );
  XNOR U7158 ( .A(n12987), .B(n12986), .Z(n12988) );
  XNOR U7159 ( .A(n12989), .B(n12988), .Z(n13010) );
  XNOR U7160 ( .A(n13011), .B(n13010), .Z(n13012) );
  XOR U7161 ( .A(n13013), .B(n13012), .Z(n13022) );
  NANDN U7162 ( .A(n12913), .B(n12912), .Z(n12917) );
  NAND U7163 ( .A(n12915), .B(n12914), .Z(n12916) );
  AND U7164 ( .A(n12917), .B(n12916), .Z(n13023) );
  XNOR U7165 ( .A(n13022), .B(n13023), .Z(n13025) );
  XNOR U7166 ( .A(n12957), .B(n12956), .Z(n12959) );
  NANDN U7167 ( .A(n12919), .B(n12918), .Z(n12923) );
  OR U7168 ( .A(n12921), .B(n12920), .Z(n12922) );
  AND U7169 ( .A(n12923), .B(n12922), .Z(n12946) );
  XOR U7170 ( .A(n12925), .B(n12924), .Z(n12945) );
  XNOR U7171 ( .A(n12927), .B(n12926), .Z(n12944) );
  XOR U7172 ( .A(n12945), .B(n12944), .Z(n12947) );
  XOR U7173 ( .A(n12946), .B(n12947), .Z(n12935) );
  NANDN U7174 ( .A(n12929), .B(n12928), .Z(n12933) );
  OR U7175 ( .A(n12931), .B(n12930), .Z(n12932) );
  NAND U7176 ( .A(n12933), .B(n12932), .Z(n12934) );
  NANDN U7177 ( .A(n12935), .B(n12934), .Z(n12943) );
  XNOR U7178 ( .A(n12935), .B(n12934), .Z(n15151) );
  NANDN U7179 ( .A(n12937), .B(n12936), .Z(n12941) );
  NAND U7180 ( .A(n12939), .B(n12938), .Z(n12940) );
  AND U7181 ( .A(n12941), .B(n12940), .Z(n15150) );
  NAND U7182 ( .A(n15151), .B(n15150), .Z(n12942) );
  AND U7183 ( .A(n12943), .B(n12942), .Z(n12951) );
  NANDN U7184 ( .A(n12945), .B(n12944), .Z(n12949) );
  OR U7185 ( .A(n12947), .B(n12946), .Z(n12948) );
  AND U7186 ( .A(n12949), .B(n12948), .Z(n12950) );
  NANDN U7187 ( .A(n12951), .B(n12950), .Z(n12955) );
  XNOR U7188 ( .A(n12951), .B(n12950), .Z(n15165) );
  XNOR U7189 ( .A(n12953), .B(n12952), .Z(n15164) );
  NAND U7190 ( .A(n15165), .B(n15164), .Z(n12954) );
  NAND U7191 ( .A(n12955), .B(n12954), .Z(n12958) );
  XNOR U7192 ( .A(n12959), .B(n12958), .Z(N45) );
  NANDN U7193 ( .A(n12957), .B(n12956), .Z(n12961) );
  NAND U7194 ( .A(n12959), .B(n12958), .Z(n12960) );
  AND U7195 ( .A(n12961), .B(n12960), .Z(n13093) );
  NANDN U7196 ( .A(n12963), .B(n12962), .Z(n12967) );
  NAND U7197 ( .A(n12965), .B(n12964), .Z(n12966) );
  AND U7198 ( .A(n12967), .B(n12966), .Z(n13031) );
  AND U7199 ( .A(x[10]), .B(y[8]), .Z(n12969) );
  AND U7200 ( .A(x[4]), .B(y[2]), .Z(n12968) );
  NAND U7201 ( .A(n12969), .B(n12968), .Z(n12972) );
  NANDN U7202 ( .A(n12970), .B(n13598), .Z(n12971) );
  AND U7203 ( .A(n12972), .B(n12971), .Z(n13052) );
  AND U7204 ( .A(y[8]), .B(x[5]), .Z(n12974) );
  NAND U7205 ( .A(x[3]), .B(y[10]), .Z(n12973) );
  XNOR U7206 ( .A(n12974), .B(n12973), .Z(n13042) );
  NAND U7207 ( .A(x[4]), .B(y[9]), .Z(n13043) );
  XNOR U7208 ( .A(n13042), .B(n13043), .Z(n13050) );
  AND U7209 ( .A(x[12]), .B(y[1]), .Z(n13039) );
  XOR U7210 ( .A(o[13]), .B(n13039), .Z(n13046) );
  AND U7211 ( .A(y[0]), .B(x[13]), .Z(n12976) );
  NAND U7212 ( .A(x[0]), .B(y[13]), .Z(n12975) );
  XOR U7213 ( .A(n12976), .B(n12975), .Z(n13047) );
  XOR U7214 ( .A(n13046), .B(n13047), .Z(n13051) );
  XOR U7215 ( .A(n13050), .B(n13051), .Z(n13053) );
  XOR U7216 ( .A(n13052), .B(n13053), .Z(n13029) );
  AND U7217 ( .A(y[11]), .B(x[6]), .Z(n13380) );
  AND U7218 ( .A(y[6]), .B(x[1]), .Z(n12977) );
  NAND U7219 ( .A(n13380), .B(n12977), .Z(n12981) );
  NAND U7220 ( .A(n12979), .B(n12978), .Z(n12980) );
  AND U7221 ( .A(n12981), .B(n12980), .Z(n13058) );
  NAND U7222 ( .A(x[12]), .B(y[12]), .Z(n14284) );
  NANDN U7223 ( .A(n14284), .B(n13115), .Z(n12985) );
  NAND U7224 ( .A(n12983), .B(n12982), .Z(n12984) );
  AND U7225 ( .A(n12985), .B(n12984), .Z(n13057) );
  AND U7226 ( .A(x[10]), .B(y[3]), .Z(n13070) );
  NAND U7227 ( .A(x[11]), .B(y[2]), .Z(n13873) );
  NAND U7228 ( .A(x[8]), .B(y[5]), .Z(n13068) );
  XOR U7229 ( .A(n13873), .B(n13068), .Z(n13069) );
  XOR U7230 ( .A(n13070), .B(n13069), .Z(n13056) );
  XOR U7231 ( .A(n13057), .B(n13056), .Z(n13059) );
  XNOR U7232 ( .A(n13058), .B(n13059), .Z(n13028) );
  XNOR U7233 ( .A(n13029), .B(n13028), .Z(n13030) );
  XNOR U7234 ( .A(n13031), .B(n13030), .Z(n13084) );
  NANDN U7235 ( .A(n12987), .B(n12986), .Z(n12991) );
  NANDN U7236 ( .A(n12989), .B(n12988), .Z(n12990) );
  AND U7237 ( .A(n12991), .B(n12990), .Z(n13081) );
  NAND U7238 ( .A(n12993), .B(n12992), .Z(n12997) );
  NAND U7239 ( .A(n12995), .B(n12994), .Z(n12996) );
  AND U7240 ( .A(n12997), .B(n12996), .Z(n13078) );
  NANDN U7241 ( .A(n12999), .B(n12998), .Z(n13003) );
  NAND U7242 ( .A(n13001), .B(n13000), .Z(n13002) );
  AND U7243 ( .A(n13003), .B(n13002), .Z(n13076) );
  AND U7244 ( .A(x[8]), .B(y[10]), .Z(n14273) );
  AND U7245 ( .A(y[4]), .B(x[2]), .Z(n13004) );
  NAND U7246 ( .A(n14273), .B(n13004), .Z(n13008) );
  NAND U7247 ( .A(n13006), .B(n13005), .Z(n13007) );
  AND U7248 ( .A(n13008), .B(n13007), .Z(n13065) );
  AND U7249 ( .A(x[6]), .B(y[7]), .Z(n13767) );
  AND U7250 ( .A(y[11]), .B(x[2]), .Z(n13034) );
  XOR U7251 ( .A(n13767), .B(n13036), .Z(n13063) );
  AND U7252 ( .A(y[12]), .B(x[1]), .Z(n13071) );
  ANDN U7253 ( .B(o[12]), .A(n13009), .Z(n13073) );
  XOR U7254 ( .A(n13074), .B(n13073), .Z(n13062) );
  XOR U7255 ( .A(n13063), .B(n13062), .Z(n13064) );
  XOR U7256 ( .A(n13065), .B(n13064), .Z(n13075) );
  XNOR U7257 ( .A(n13076), .B(n13075), .Z(n13077) );
  XOR U7258 ( .A(n13078), .B(n13077), .Z(n13082) );
  XNOR U7259 ( .A(n13081), .B(n13082), .Z(n13083) );
  XOR U7260 ( .A(n13084), .B(n13083), .Z(n13088) );
  NANDN U7261 ( .A(n13011), .B(n13010), .Z(n13015) );
  NANDN U7262 ( .A(n13013), .B(n13012), .Z(n13014) );
  NAND U7263 ( .A(n13015), .B(n13014), .Z(n13087) );
  XNOR U7264 ( .A(n13088), .B(n13087), .Z(n13089) );
  NANDN U7265 ( .A(n13017), .B(n13016), .Z(n13021) );
  NANDN U7266 ( .A(n13019), .B(n13018), .Z(n13020) );
  NAND U7267 ( .A(n13021), .B(n13020), .Z(n13090) );
  XOR U7268 ( .A(n13089), .B(n13090), .Z(n13094) );
  XNOR U7269 ( .A(n13093), .B(n13094), .Z(n13096) );
  NAND U7270 ( .A(n13023), .B(n13022), .Z(n13027) );
  NANDN U7271 ( .A(n13025), .B(n13024), .Z(n13026) );
  AND U7272 ( .A(n13027), .B(n13026), .Z(n13095) );
  XOR U7273 ( .A(n13096), .B(n13095), .Z(N46) );
  NANDN U7274 ( .A(n13029), .B(n13028), .Z(n13033) );
  NANDN U7275 ( .A(n13031), .B(n13030), .Z(n13032) );
  AND U7276 ( .A(n13033), .B(n13032), .Z(n13101) );
  AND U7277 ( .A(y[0]), .B(x[14]), .Z(n13038) );
  NAND U7278 ( .A(x[0]), .B(y[14]), .Z(n13037) );
  XNOR U7279 ( .A(n13038), .B(n13037), .Z(n13117) );
  AND U7280 ( .A(o[13]), .B(n13039), .Z(n13116) );
  XOR U7281 ( .A(n13117), .B(n13116), .Z(n13137) );
  NAND U7282 ( .A(y[1]), .B(x[13]), .Z(n13157) );
  XNOR U7283 ( .A(o[14]), .B(n13157), .Z(n13152) );
  NAND U7284 ( .A(y[2]), .B(x[12]), .Z(n13040) );
  XNOR U7285 ( .A(n13041), .B(n13040), .Z(n13153) );
  XOR U7286 ( .A(n13152), .B(n13153), .Z(n13136) );
  XOR U7287 ( .A(n13137), .B(n13136), .Z(n13138) );
  XOR U7288 ( .A(n13139), .B(n13138), .Z(n13162) );
  AND U7289 ( .A(y[10]), .B(x[5]), .Z(n13210) );
  NANDN U7290 ( .A(n13689), .B(n13210), .Z(n13045) );
  NANDN U7291 ( .A(n13043), .B(n13042), .Z(n13044) );
  AND U7292 ( .A(n13045), .B(n13044), .Z(n13142) );
  NAND U7293 ( .A(y[13]), .B(x[1]), .Z(n13160) );
  NAND U7294 ( .A(x[11]), .B(y[3]), .Z(n13159) );
  XOR U7295 ( .A(n13158), .B(n13159), .Z(n13161) );
  XOR U7296 ( .A(n13160), .B(n13161), .Z(n13140) );
  NAND U7297 ( .A(y[13]), .B(x[13]), .Z(n14622) );
  NANDN U7298 ( .A(n14622), .B(n13115), .Z(n13049) );
  NANDN U7299 ( .A(n13047), .B(n13046), .Z(n13048) );
  NAND U7300 ( .A(n13049), .B(n13048), .Z(n13141) );
  XOR U7301 ( .A(n13140), .B(n13141), .Z(n13143) );
  XNOR U7302 ( .A(n13142), .B(n13143), .Z(n13163) );
  XOR U7303 ( .A(n13162), .B(n13163), .Z(n13165) );
  NANDN U7304 ( .A(n13051), .B(n13050), .Z(n13055) );
  OR U7305 ( .A(n13053), .B(n13052), .Z(n13054) );
  AND U7306 ( .A(n13055), .B(n13054), .Z(n13164) );
  XOR U7307 ( .A(n13165), .B(n13164), .Z(n13100) );
  NANDN U7308 ( .A(n13057), .B(n13056), .Z(n13061) );
  OR U7309 ( .A(n13059), .B(n13058), .Z(n13060) );
  AND U7310 ( .A(n13061), .B(n13060), .Z(n13108) );
  AND U7311 ( .A(x[4]), .B(y[10]), .Z(n13515) );
  AND U7312 ( .A(x[3]), .B(y[11]), .Z(n13067) );
  NAND U7313 ( .A(x[8]), .B(y[6]), .Z(n13066) );
  XOR U7314 ( .A(n13067), .B(n13066), .Z(n13122) );
  XOR U7315 ( .A(n13379), .B(n13122), .Z(n13125) );
  XNOR U7316 ( .A(n13515), .B(n13125), .Z(n13126) );
  AND U7317 ( .A(y[4]), .B(x[10]), .Z(n13882) );
  AND U7318 ( .A(y[12]), .B(x[2]), .Z(n13146) );
  XOR U7319 ( .A(n13882), .B(n13146), .Z(n13148) );
  AND U7320 ( .A(y[5]), .B(x[9]), .Z(n13147) );
  XOR U7321 ( .A(n13148), .B(n13147), .Z(n13127) );
  XOR U7322 ( .A(n13126), .B(n13127), .Z(n13132) );
  XOR U7323 ( .A(n13131), .B(n13130), .Z(n13133) );
  XNOR U7324 ( .A(n13132), .B(n13133), .Z(n13105) );
  XNOR U7325 ( .A(n13106), .B(n13105), .Z(n13107) );
  XNOR U7326 ( .A(n13108), .B(n13107), .Z(n13099) );
  XOR U7327 ( .A(n13100), .B(n13099), .Z(n13102) );
  XOR U7328 ( .A(n13101), .B(n13102), .Z(n13174) );
  NANDN U7329 ( .A(n13076), .B(n13075), .Z(n13080) );
  NANDN U7330 ( .A(n13078), .B(n13077), .Z(n13079) );
  NAND U7331 ( .A(n13080), .B(n13079), .Z(n13173) );
  NANDN U7332 ( .A(n13082), .B(n13081), .Z(n13086) );
  NAND U7333 ( .A(n13084), .B(n13083), .Z(n13085) );
  NAND U7334 ( .A(n13086), .B(n13085), .Z(n13172) );
  XOR U7335 ( .A(n13173), .B(n13172), .Z(n13175) );
  XOR U7336 ( .A(n13174), .B(n13175), .Z(n13166) );
  NANDN U7337 ( .A(n13088), .B(n13087), .Z(n13092) );
  NANDN U7338 ( .A(n13090), .B(n13089), .Z(n13091) );
  NAND U7339 ( .A(n13092), .B(n13091), .Z(n13167) );
  XNOR U7340 ( .A(n13166), .B(n13167), .Z(n13169) );
  NANDN U7341 ( .A(n13094), .B(n13093), .Z(n13098) );
  NAND U7342 ( .A(n13096), .B(n13095), .Z(n13097) );
  AND U7343 ( .A(n13098), .B(n13097), .Z(n13168) );
  XNOR U7344 ( .A(n13169), .B(n13168), .Z(N47) );
  NANDN U7345 ( .A(n13100), .B(n13099), .Z(n13104) );
  NANDN U7346 ( .A(n13102), .B(n13101), .Z(n13103) );
  AND U7347 ( .A(n13104), .B(n13103), .Z(n13181) );
  NANDN U7348 ( .A(n13106), .B(n13105), .Z(n13110) );
  NANDN U7349 ( .A(n13108), .B(n13107), .Z(n13109) );
  AND U7350 ( .A(n13110), .B(n13109), .Z(n13242) );
  AND U7351 ( .A(x[6]), .B(y[9]), .Z(n13301) );
  AND U7352 ( .A(x[10]), .B(y[5]), .Z(n13112) );
  NAND U7353 ( .A(y[11]), .B(x[4]), .Z(n13111) );
  XNOR U7354 ( .A(n13112), .B(n13111), .Z(n13187) );
  NAND U7355 ( .A(x[7]), .B(y[8]), .Z(n13188) );
  XNOR U7356 ( .A(n13187), .B(n13188), .Z(n13208) );
  XOR U7357 ( .A(n13301), .B(n13208), .Z(n13209) );
  XOR U7358 ( .A(n13209), .B(n13210), .Z(n13222) );
  AND U7359 ( .A(y[1]), .B(x[14]), .Z(n13207) );
  XOR U7360 ( .A(n13207), .B(o[15]), .Z(n13197) );
  AND U7361 ( .A(y[14]), .B(x[1]), .Z(n13196) );
  NAND U7362 ( .A(x[8]), .B(y[7]), .Z(n13195) );
  XOR U7363 ( .A(n13196), .B(n13195), .Z(n13198) );
  XOR U7364 ( .A(n13197), .B(n13198), .Z(n13220) );
  AND U7365 ( .A(x[2]), .B(y[13]), .Z(n13114) );
  NAND U7366 ( .A(x[9]), .B(y[6]), .Z(n13113) );
  XNOR U7367 ( .A(n13114), .B(n13113), .Z(n13201) );
  AND U7368 ( .A(y[12]), .B(x[3]), .Z(n13202) );
  XOR U7369 ( .A(n13201), .B(n13202), .Z(n13219) );
  XNOR U7370 ( .A(n13222), .B(n13221), .Z(n13216) );
  AND U7371 ( .A(y[14]), .B(x[14]), .Z(n14892) );
  NAND U7372 ( .A(n14892), .B(n13115), .Z(n13119) );
  NAND U7373 ( .A(n13117), .B(n13116), .Z(n13118) );
  AND U7374 ( .A(n13119), .B(n13118), .Z(n13213) );
  AND U7375 ( .A(y[11]), .B(x[8]), .Z(n13120) );
  NANDN U7376 ( .A(n13121), .B(n13120), .Z(n13124) );
  NANDN U7377 ( .A(n13122), .B(n13379), .Z(n13123) );
  AND U7378 ( .A(n13124), .B(n13123), .Z(n13214) );
  XOR U7379 ( .A(n13213), .B(n13214), .Z(n13215) );
  XNOR U7380 ( .A(n13216), .B(n13215), .Z(n13258) );
  NANDN U7381 ( .A(n13125), .B(n13515), .Z(n13129) );
  NAND U7382 ( .A(n13127), .B(n13126), .Z(n13128) );
  NAND U7383 ( .A(n13129), .B(n13128), .Z(n13257) );
  XOR U7384 ( .A(n13258), .B(n13257), .Z(n13260) );
  NANDN U7385 ( .A(n13131), .B(n13130), .Z(n13135) );
  OR U7386 ( .A(n13133), .B(n13132), .Z(n13134) );
  AND U7387 ( .A(n13135), .B(n13134), .Z(n13259) );
  XOR U7388 ( .A(n13260), .B(n13259), .Z(n13240) );
  NANDN U7389 ( .A(n13141), .B(n13140), .Z(n13145) );
  NANDN U7390 ( .A(n13143), .B(n13142), .Z(n13144) );
  AND U7391 ( .A(n13145), .B(n13144), .Z(n13245) );
  XNOR U7392 ( .A(n13246), .B(n13245), .Z(n13248) );
  AND U7393 ( .A(n13882), .B(n13146), .Z(n13150) );
  NAND U7394 ( .A(n13148), .B(n13147), .Z(n13149) );
  NANDN U7395 ( .A(n13150), .B(n13149), .Z(n13251) );
  NAND U7396 ( .A(x[12]), .B(y[7]), .Z(n13605) );
  NANDN U7397 ( .A(n13605), .B(n13151), .Z(n13155) );
  NAND U7398 ( .A(n13153), .B(n13152), .Z(n13154) );
  NAND U7399 ( .A(n13155), .B(n13154), .Z(n13228) );
  AND U7400 ( .A(x[13]), .B(y[2]), .Z(n13772) );
  NAND U7401 ( .A(x[11]), .B(y[4]), .Z(n13156) );
  XNOR U7402 ( .A(n13772), .B(n13156), .Z(n13231) );
  NAND U7403 ( .A(x[12]), .B(y[3]), .Z(n13232) );
  XNOR U7404 ( .A(n13231), .B(n13232), .Z(n13226) );
  AND U7405 ( .A(x[15]), .B(y[0]), .Z(n13191) );
  NAND U7406 ( .A(y[15]), .B(x[0]), .Z(n13192) );
  XNOR U7407 ( .A(n13191), .B(n13192), .Z(n13194) );
  ANDN U7408 ( .B(o[14]), .A(n13157), .Z(n13193) );
  XOR U7409 ( .A(n13194), .B(n13193), .Z(n13225) );
  XOR U7410 ( .A(n13226), .B(n13225), .Z(n13227) );
  XOR U7411 ( .A(n13228), .B(n13227), .Z(n13252) );
  XOR U7412 ( .A(n13251), .B(n13252), .Z(n13254) );
  XOR U7413 ( .A(n13254), .B(n13253), .Z(n13247) );
  XNOR U7414 ( .A(n13248), .B(n13247), .Z(n13239) );
  XNOR U7415 ( .A(n13240), .B(n13239), .Z(n13241) );
  XOR U7416 ( .A(n13242), .B(n13241), .Z(n13179) );
  XNOR U7417 ( .A(n13179), .B(n13178), .Z(n13180) );
  XNOR U7418 ( .A(n13181), .B(n13180), .Z(n13263) );
  NANDN U7419 ( .A(n13167), .B(n13166), .Z(n13171) );
  NAND U7420 ( .A(n13169), .B(n13168), .Z(n13170) );
  NAND U7421 ( .A(n13171), .B(n13170), .Z(n13264) );
  XNOR U7422 ( .A(n13263), .B(n13264), .Z(n13266) );
  NAND U7423 ( .A(n13173), .B(n13172), .Z(n13177) );
  NAND U7424 ( .A(n13175), .B(n13174), .Z(n13176) );
  AND U7425 ( .A(n13177), .B(n13176), .Z(n13265) );
  XOR U7426 ( .A(n13266), .B(n13265), .Z(N48) );
  NANDN U7427 ( .A(n13179), .B(n13178), .Z(n13183) );
  NANDN U7428 ( .A(n13181), .B(n13180), .Z(n13182) );
  AND U7429 ( .A(n13183), .B(n13182), .Z(n13361) );
  AND U7430 ( .A(x[7]), .B(y[9]), .Z(n13185) );
  NAND U7431 ( .A(x[6]), .B(y[10]), .Z(n13184) );
  XNOR U7432 ( .A(n13185), .B(n13184), .Z(n13303) );
  AND U7433 ( .A(y[6]), .B(x[10]), .Z(n13302) );
  XOR U7434 ( .A(n13303), .B(n13302), .Z(n13288) );
  NAND U7435 ( .A(y[1]), .B(x[15]), .Z(n13316) );
  XNOR U7436 ( .A(o[16]), .B(n13316), .Z(n13298) );
  AND U7437 ( .A(x[16]), .B(y[0]), .Z(n13295) );
  NAND U7438 ( .A(y[16]), .B(x[0]), .Z(n13296) );
  XNOR U7439 ( .A(n13295), .B(n13296), .Z(n13297) );
  XNOR U7440 ( .A(n13298), .B(n13297), .Z(n13287) );
  XNOR U7441 ( .A(n13288), .B(n13287), .Z(n13290) );
  NAND U7442 ( .A(y[11]), .B(x[10]), .Z(n13711) );
  NANDN U7443 ( .A(n13711), .B(n13186), .Z(n13190) );
  NANDN U7444 ( .A(n13188), .B(n13187), .Z(n13189) );
  AND U7445 ( .A(n13190), .B(n13189), .Z(n13289) );
  XOR U7446 ( .A(n13290), .B(n13289), .Z(n13325) );
  NANDN U7447 ( .A(n13196), .B(n13195), .Z(n13200) );
  OR U7448 ( .A(n13198), .B(n13197), .Z(n13199) );
  AND U7449 ( .A(n13200), .B(n13199), .Z(n13323) );
  XOR U7450 ( .A(n13324), .B(n13323), .Z(n13326) );
  XNOR U7451 ( .A(n13325), .B(n13326), .Z(n13278) );
  AND U7452 ( .A(y[13]), .B(x[9]), .Z(n13868) );
  NAND U7453 ( .A(n13868), .B(n13603), .Z(n13204) );
  NAND U7454 ( .A(n13202), .B(n13201), .Z(n13203) );
  AND U7455 ( .A(n13204), .B(n13203), .Z(n13284) );
  AND U7456 ( .A(x[4]), .B(y[12]), .Z(n13340) );
  AND U7457 ( .A(y[2]), .B(x[14]), .Z(n13339) );
  NAND U7458 ( .A(y[5]), .B(x[11]), .Z(n13338) );
  XOR U7459 ( .A(n13339), .B(n13338), .Z(n13341) );
  XOR U7460 ( .A(n13340), .B(n13341), .Z(n13282) );
  AND U7461 ( .A(x[1]), .B(y[15]), .Z(n13206) );
  NAND U7462 ( .A(y[8]), .B(x[8]), .Z(n13205) );
  XNOR U7463 ( .A(n13206), .B(n13205), .Z(n13306) );
  NAND U7464 ( .A(n13207), .B(o[15]), .Z(n13307) );
  XNOR U7465 ( .A(n13306), .B(n13307), .Z(n13281) );
  NAND U7466 ( .A(n13208), .B(n13301), .Z(n13212) );
  NAND U7467 ( .A(n13210), .B(n13209), .Z(n13211) );
  AND U7468 ( .A(n13212), .B(n13211), .Z(n13276) );
  XOR U7469 ( .A(n13275), .B(n13276), .Z(n13277) );
  XNOR U7470 ( .A(n13278), .B(n13277), .Z(n13317) );
  NAND U7471 ( .A(n13214), .B(n13213), .Z(n13218) );
  NAND U7472 ( .A(n13216), .B(n13215), .Z(n13217) );
  AND U7473 ( .A(n13218), .B(n13217), .Z(n13318) );
  XOR U7474 ( .A(n13317), .B(n13318), .Z(n13320) );
  NANDN U7475 ( .A(n13220), .B(n13219), .Z(n13224) );
  NAND U7476 ( .A(n13222), .B(n13221), .Z(n13223) );
  AND U7477 ( .A(n13224), .B(n13223), .Z(n13351) );
  NAND U7478 ( .A(n13226), .B(n13225), .Z(n13230) );
  NAND U7479 ( .A(n13228), .B(n13227), .Z(n13229) );
  AND U7480 ( .A(n13230), .B(n13229), .Z(n13349) );
  AND U7481 ( .A(y[4]), .B(x[13]), .Z(n13337) );
  NANDN U7482 ( .A(n13873), .B(n13337), .Z(n13234) );
  NANDN U7483 ( .A(n13232), .B(n13231), .Z(n13233) );
  AND U7484 ( .A(n13234), .B(n13233), .Z(n13332) );
  AND U7485 ( .A(y[7]), .B(x[9]), .Z(n13236) );
  NAND U7486 ( .A(x[2]), .B(y[14]), .Z(n13235) );
  XNOR U7487 ( .A(n13236), .B(n13235), .Z(n13344) );
  NAND U7488 ( .A(y[13]), .B(x[3]), .Z(n13345) );
  XNOR U7489 ( .A(n13344), .B(n13345), .Z(n13329) );
  AND U7490 ( .A(y[4]), .B(x[12]), .Z(n13752) );
  AND U7491 ( .A(y[3]), .B(x[13]), .Z(n13238) );
  NAND U7492 ( .A(x[5]), .B(y[11]), .Z(n13237) );
  XOR U7493 ( .A(n13238), .B(n13237), .Z(n13311) );
  XOR U7494 ( .A(n13752), .B(n13311), .Z(n13330) );
  XNOR U7495 ( .A(n13329), .B(n13330), .Z(n13331) );
  XNOR U7496 ( .A(n13332), .B(n13331), .Z(n13348) );
  XOR U7497 ( .A(n13320), .B(n13319), .Z(n13271) );
  NANDN U7498 ( .A(n13240), .B(n13239), .Z(n13244) );
  NAND U7499 ( .A(n13242), .B(n13241), .Z(n13243) );
  AND U7500 ( .A(n13244), .B(n13243), .Z(n13270) );
  NANDN U7501 ( .A(n13246), .B(n13245), .Z(n13250) );
  NAND U7502 ( .A(n13248), .B(n13247), .Z(n13249) );
  AND U7503 ( .A(n13250), .B(n13249), .Z(n13357) );
  NAND U7504 ( .A(n13252), .B(n13251), .Z(n13256) );
  NAND U7505 ( .A(n13254), .B(n13253), .Z(n13255) );
  AND U7506 ( .A(n13256), .B(n13255), .Z(n13355) );
  NAND U7507 ( .A(n13258), .B(n13257), .Z(n13262) );
  NAND U7508 ( .A(n13260), .B(n13259), .Z(n13261) );
  AND U7509 ( .A(n13262), .B(n13261), .Z(n13354) );
  XOR U7510 ( .A(n13355), .B(n13354), .Z(n13356) );
  XOR U7511 ( .A(n13357), .B(n13356), .Z(n13269) );
  XOR U7512 ( .A(n13270), .B(n13269), .Z(n13272) );
  XNOR U7513 ( .A(n13271), .B(n13272), .Z(n13360) );
  XNOR U7514 ( .A(n13361), .B(n13360), .Z(n13363) );
  NANDN U7515 ( .A(n13264), .B(n13263), .Z(n13268) );
  NAND U7516 ( .A(n13266), .B(n13265), .Z(n13267) );
  NAND U7517 ( .A(n13268), .B(n13267), .Z(n13362) );
  XOR U7518 ( .A(n13363), .B(n13362), .Z(N49) );
  NANDN U7519 ( .A(n13270), .B(n13269), .Z(n13274) );
  OR U7520 ( .A(n13272), .B(n13271), .Z(n13273) );
  AND U7521 ( .A(n13274), .B(n13273), .Z(n13461) );
  NAND U7522 ( .A(n13276), .B(n13275), .Z(n13280) );
  NAND U7523 ( .A(n13278), .B(n13277), .Z(n13279) );
  AND U7524 ( .A(n13280), .B(n13279), .Z(n13451) );
  NANDN U7525 ( .A(n13282), .B(n13281), .Z(n13286) );
  NANDN U7526 ( .A(n13284), .B(n13283), .Z(n13285) );
  AND U7527 ( .A(n13286), .B(n13285), .Z(n13448) );
  NANDN U7528 ( .A(n13288), .B(n13287), .Z(n13292) );
  NAND U7529 ( .A(n13290), .B(n13289), .Z(n13291) );
  AND U7530 ( .A(n13292), .B(n13291), .Z(n13445) );
  AND U7531 ( .A(x[2]), .B(y[15]), .Z(n13294) );
  NAND U7532 ( .A(y[7]), .B(x[10]), .Z(n13293) );
  XNOR U7533 ( .A(n13294), .B(n13293), .Z(n13374) );
  AND U7534 ( .A(y[14]), .B(x[3]), .Z(n13373) );
  XOR U7535 ( .A(n13374), .B(n13373), .Z(n13406) );
  NAND U7536 ( .A(x[16]), .B(y[1]), .Z(n13422) );
  XNOR U7537 ( .A(o[17]), .B(n13422), .Z(n13415) );
  AND U7538 ( .A(y[17]), .B(x[0]), .Z(n13412) );
  NAND U7539 ( .A(x[17]), .B(y[0]), .Z(n13413) );
  XNOR U7540 ( .A(n13412), .B(n13413), .Z(n13414) );
  XOR U7541 ( .A(n13415), .B(n13414), .Z(n13405) );
  NANDN U7542 ( .A(n13296), .B(n13295), .Z(n13300) );
  NAND U7543 ( .A(n13298), .B(n13297), .Z(n13299) );
  AND U7544 ( .A(n13300), .B(n13299), .Z(n13404) );
  XOR U7545 ( .A(n13405), .B(n13404), .Z(n13407) );
  XOR U7546 ( .A(n13406), .B(n13407), .Z(n13394) );
  AND U7547 ( .A(y[10]), .B(x[7]), .Z(n13367) );
  NAND U7548 ( .A(n13367), .B(n13301), .Z(n13305) );
  NAND U7549 ( .A(n13303), .B(n13302), .Z(n13304) );
  AND U7550 ( .A(n13305), .B(n13304), .Z(n13393) );
  AND U7551 ( .A(x[8]), .B(y[15]), .Z(n14071) );
  NAND U7552 ( .A(n14071), .B(n13524), .Z(n13309) );
  NANDN U7553 ( .A(n13307), .B(n13306), .Z(n13308) );
  NAND U7554 ( .A(n13309), .B(n13308), .Z(n13392) );
  XOR U7555 ( .A(n13393), .B(n13392), .Z(n13395) );
  XOR U7556 ( .A(n13394), .B(n13395), .Z(n13443) );
  AND U7557 ( .A(y[11]), .B(x[13]), .Z(n14279) );
  NANDN U7558 ( .A(n13310), .B(n14279), .Z(n13313) );
  NANDN U7559 ( .A(n13311), .B(n13752), .Z(n13312) );
  AND U7560 ( .A(n13313), .B(n13312), .Z(n13399) );
  AND U7561 ( .A(y[2]), .B(x[15]), .Z(n13430) );
  NAND U7562 ( .A(y[5]), .B(x[12]), .Z(n13431) );
  XNOR U7563 ( .A(n13430), .B(n13431), .Z(n13432) );
  NAND U7564 ( .A(x[14]), .B(y[3]), .Z(n13433) );
  XNOR U7565 ( .A(n13432), .B(n13433), .Z(n13398) );
  XNOR U7566 ( .A(n13399), .B(n13398), .Z(n13401) );
  AND U7567 ( .A(y[8]), .B(x[9]), .Z(n13315) );
  NAND U7568 ( .A(x[1]), .B(y[16]), .Z(n13314) );
  XNOR U7569 ( .A(n13315), .B(n13314), .Z(n13385) );
  ANDN U7570 ( .B(o[16]), .A(n13316), .Z(n13384) );
  XOR U7571 ( .A(n13385), .B(n13384), .Z(n13400) );
  XNOR U7572 ( .A(n13401), .B(n13400), .Z(n13442) );
  XNOR U7573 ( .A(n13443), .B(n13442), .Z(n13444) );
  XOR U7574 ( .A(n13445), .B(n13444), .Z(n13449) );
  NAND U7575 ( .A(n13318), .B(n13317), .Z(n13322) );
  NAND U7576 ( .A(n13320), .B(n13319), .Z(n13321) );
  AND U7577 ( .A(n13322), .B(n13321), .Z(n13457) );
  NANDN U7578 ( .A(n13324), .B(n13323), .Z(n13328) );
  OR U7579 ( .A(n13326), .B(n13325), .Z(n13327) );
  AND U7580 ( .A(n13328), .B(n13327), .Z(n13438) );
  NANDN U7581 ( .A(n13330), .B(n13329), .Z(n13334) );
  NANDN U7582 ( .A(n13332), .B(n13331), .Z(n13333) );
  AND U7583 ( .A(n13334), .B(n13333), .Z(n13437) );
  AND U7584 ( .A(x[5]), .B(y[12]), .Z(n13477) );
  NAND U7585 ( .A(x[8]), .B(y[9]), .Z(n13335) );
  XNOR U7586 ( .A(n13477), .B(n13335), .Z(n13381) );
  XOR U7587 ( .A(n13381), .B(n13380), .Z(n13366) );
  XOR U7588 ( .A(n13367), .B(n13366), .Z(n13369) );
  NAND U7589 ( .A(y[13]), .B(x[4]), .Z(n13336) );
  XNOR U7590 ( .A(n13337), .B(n13336), .Z(n13426) );
  NAND U7591 ( .A(y[6]), .B(x[11]), .Z(n13427) );
  XNOR U7592 ( .A(n13426), .B(n13427), .Z(n13368) );
  XOR U7593 ( .A(n13369), .B(n13368), .Z(n13388) );
  NANDN U7594 ( .A(n13339), .B(n13338), .Z(n13343) );
  OR U7595 ( .A(n13341), .B(n13340), .Z(n13342) );
  AND U7596 ( .A(n13343), .B(n13342), .Z(n13387) );
  AND U7597 ( .A(x[9]), .B(y[14]), .Z(n14268) );
  NAND U7598 ( .A(n13372), .B(n14268), .Z(n13347) );
  NANDN U7599 ( .A(n13345), .B(n13344), .Z(n13346) );
  AND U7600 ( .A(n13347), .B(n13346), .Z(n13386) );
  XOR U7601 ( .A(n13387), .B(n13386), .Z(n13389) );
  XNOR U7602 ( .A(n13388), .B(n13389), .Z(n13436) );
  XOR U7603 ( .A(n13437), .B(n13436), .Z(n13439) );
  XOR U7604 ( .A(n13438), .B(n13439), .Z(n13455) );
  NANDN U7605 ( .A(n13349), .B(n13348), .Z(n13353) );
  NANDN U7606 ( .A(n13351), .B(n13350), .Z(n13352) );
  AND U7607 ( .A(n13353), .B(n13352), .Z(n13454) );
  XNOR U7608 ( .A(n13457), .B(n13456), .Z(n13464) );
  XOR U7609 ( .A(n13465), .B(n13464), .Z(n13467) );
  NAND U7610 ( .A(n13355), .B(n13354), .Z(n13359) );
  NAND U7611 ( .A(n13357), .B(n13356), .Z(n13358) );
  AND U7612 ( .A(n13359), .B(n13358), .Z(n13466) );
  XOR U7613 ( .A(n13467), .B(n13466), .Z(n13460) );
  XOR U7614 ( .A(n13461), .B(n13460), .Z(n13463) );
  NANDN U7615 ( .A(n13361), .B(n13360), .Z(n13365) );
  NAND U7616 ( .A(n13363), .B(n13362), .Z(n13364) );
  NAND U7617 ( .A(n13365), .B(n13364), .Z(n13462) );
  XOR U7618 ( .A(n13463), .B(n13462), .Z(N50) );
  NAND U7619 ( .A(n13367), .B(n13366), .Z(n13371) );
  NAND U7620 ( .A(n13369), .B(n13368), .Z(n13370) );
  AND U7621 ( .A(n13371), .B(n13370), .Z(n13537) );
  AND U7622 ( .A(x[10]), .B(y[15]), .Z(n14292) );
  IV U7623 ( .A(n14292), .Z(n14437) );
  NANDN U7624 ( .A(n14437), .B(n13372), .Z(n13376) );
  NAND U7625 ( .A(n13374), .B(n13373), .Z(n13375) );
  NAND U7626 ( .A(n13376), .B(n13375), .Z(n13498) );
  AND U7627 ( .A(x[3]), .B(y[15]), .Z(n13378) );
  NAND U7628 ( .A(x[13]), .B(y[5]), .Z(n13377) );
  XNOR U7629 ( .A(n13378), .B(n13377), .Z(n13509) );
  NAND U7630 ( .A(y[6]), .B(x[12]), .Z(n13510) );
  XNOR U7631 ( .A(n13509), .B(n13510), .Z(n13497) );
  NAND U7632 ( .A(x[17]), .B(y[1]), .Z(n13521) );
  XNOR U7633 ( .A(o[18]), .B(n13521), .Z(n13529) );
  AND U7634 ( .A(x[0]), .B(y[18]), .Z(n13527) );
  NAND U7635 ( .A(x[18]), .B(y[0]), .Z(n13528) );
  XOR U7636 ( .A(n13527), .B(n13528), .Z(n13530) );
  XNOR U7637 ( .A(n13529), .B(n13530), .Z(n13496) );
  XOR U7638 ( .A(n13497), .B(n13496), .Z(n13499) );
  XNOR U7639 ( .A(n13498), .B(n13499), .Z(n13552) );
  AND U7640 ( .A(x[8]), .B(y[12]), .Z(n13867) );
  NAND U7641 ( .A(n13867), .B(n13379), .Z(n13383) );
  NAND U7642 ( .A(n13381), .B(n13380), .Z(n13382) );
  AND U7643 ( .A(n13383), .B(n13382), .Z(n13550) );
  AND U7644 ( .A(y[16]), .B(x[9]), .Z(n14438) );
  XOR U7645 ( .A(n13550), .B(n13551), .Z(n13553) );
  XOR U7646 ( .A(n13552), .B(n13553), .Z(n13534) );
  NANDN U7647 ( .A(n13387), .B(n13386), .Z(n13391) );
  OR U7648 ( .A(n13389), .B(n13388), .Z(n13390) );
  AND U7649 ( .A(n13391), .B(n13390), .Z(n13535) );
  XOR U7650 ( .A(n13534), .B(n13535), .Z(n13536) );
  XOR U7651 ( .A(n13537), .B(n13536), .Z(n13473) );
  NANDN U7652 ( .A(n13393), .B(n13392), .Z(n13397) );
  OR U7653 ( .A(n13395), .B(n13394), .Z(n13396) );
  AND U7654 ( .A(n13397), .B(n13396), .Z(n13558) );
  NANDN U7655 ( .A(n13399), .B(n13398), .Z(n13403) );
  NAND U7656 ( .A(n13401), .B(n13400), .Z(n13402) );
  AND U7657 ( .A(n13403), .B(n13402), .Z(n13557) );
  NANDN U7658 ( .A(n13405), .B(n13404), .Z(n13409) );
  OR U7659 ( .A(n13407), .B(n13406), .Z(n13408) );
  AND U7660 ( .A(n13409), .B(n13408), .Z(n13556) );
  XOR U7661 ( .A(n13557), .B(n13556), .Z(n13559) );
  XOR U7662 ( .A(n13558), .B(n13559), .Z(n13472) );
  AND U7663 ( .A(x[5]), .B(y[13]), .Z(n13632) );
  NAND U7664 ( .A(y[12]), .B(x[6]), .Z(n13410) );
  XNOR U7665 ( .A(n13632), .B(n13410), .Z(n13480) );
  NAND U7666 ( .A(y[14]), .B(x[4]), .Z(n13411) );
  XNOR U7667 ( .A(n14273), .B(n13411), .Z(n13518) );
  AND U7668 ( .A(y[11]), .B(x[7]), .Z(n13517) );
  XOR U7669 ( .A(n13518), .B(n13517), .Z(n13479) );
  XOR U7670 ( .A(n13480), .B(n13479), .Z(n13541) );
  NANDN U7671 ( .A(n13413), .B(n13412), .Z(n13417) );
  NAND U7672 ( .A(n13415), .B(n13414), .Z(n13416) );
  AND U7673 ( .A(n13417), .B(n13416), .Z(n13539) );
  AND U7674 ( .A(y[7]), .B(x[11]), .Z(n13419) );
  NAND U7675 ( .A(y[2]), .B(x[16]), .Z(n13418) );
  XNOR U7676 ( .A(n13419), .B(n13418), .Z(n13485) );
  AND U7677 ( .A(y[16]), .B(x[2]), .Z(n13484) );
  XOR U7678 ( .A(n13485), .B(n13484), .Z(n13538) );
  XNOR U7679 ( .A(n13539), .B(n13538), .Z(n13540) );
  XOR U7680 ( .A(n13541), .B(n13540), .Z(n13547) );
  AND U7681 ( .A(x[1]), .B(y[17]), .Z(n13421) );
  NAND U7682 ( .A(y[8]), .B(x[10]), .Z(n13420) );
  XNOR U7683 ( .A(n13421), .B(n13420), .Z(n13526) );
  ANDN U7684 ( .B(o[17]), .A(n13422), .Z(n13525) );
  XNOR U7685 ( .A(n13526), .B(n13525), .Z(n13503) );
  AND U7686 ( .A(y[3]), .B(x[15]), .Z(n13424) );
  NAND U7687 ( .A(x[9]), .B(y[9]), .Z(n13423) );
  XNOR U7688 ( .A(n13424), .B(n13423), .Z(n13489) );
  AND U7689 ( .A(y[4]), .B(x[14]), .Z(n13488) );
  XNOR U7690 ( .A(n13489), .B(n13488), .Z(n13502) );
  XOR U7691 ( .A(n13503), .B(n13502), .Z(n13505) );
  NANDN U7692 ( .A(n14622), .B(n13425), .Z(n13429) );
  NANDN U7693 ( .A(n13427), .B(n13426), .Z(n13428) );
  AND U7694 ( .A(n13429), .B(n13428), .Z(n13504) );
  XOR U7695 ( .A(n13505), .B(n13504), .Z(n13544) );
  NANDN U7696 ( .A(n13431), .B(n13430), .Z(n13435) );
  NANDN U7697 ( .A(n13433), .B(n13432), .Z(n13434) );
  NAND U7698 ( .A(n13435), .B(n13434), .Z(n13545) );
  XNOR U7699 ( .A(n13544), .B(n13545), .Z(n13546) );
  XNOR U7700 ( .A(n13547), .B(n13546), .Z(n13471) );
  XOR U7701 ( .A(n13472), .B(n13471), .Z(n13474) );
  XOR U7702 ( .A(n13473), .B(n13474), .Z(n13564) );
  NANDN U7703 ( .A(n13437), .B(n13436), .Z(n13441) );
  OR U7704 ( .A(n13439), .B(n13438), .Z(n13440) );
  AND U7705 ( .A(n13441), .B(n13440), .Z(n13563) );
  NANDN U7706 ( .A(n13443), .B(n13442), .Z(n13447) );
  NANDN U7707 ( .A(n13445), .B(n13444), .Z(n13446) );
  AND U7708 ( .A(n13447), .B(n13446), .Z(n13562) );
  XNOR U7709 ( .A(n13563), .B(n13562), .Z(n13565) );
  XOR U7710 ( .A(n13564), .B(n13565), .Z(n13566) );
  NANDN U7711 ( .A(n13449), .B(n13448), .Z(n13453) );
  NANDN U7712 ( .A(n13451), .B(n13450), .Z(n13452) );
  NAND U7713 ( .A(n13453), .B(n13452), .Z(n13567) );
  NANDN U7714 ( .A(n13455), .B(n13454), .Z(n13459) );
  NAND U7715 ( .A(n13457), .B(n13456), .Z(n13458) );
  AND U7716 ( .A(n13459), .B(n13458), .Z(n13568) );
  XNOR U7717 ( .A(n13569), .B(n13568), .Z(n13574) );
  NAND U7718 ( .A(n13465), .B(n13464), .Z(n13469) );
  NAND U7719 ( .A(n13467), .B(n13466), .Z(n13468) );
  NAND U7720 ( .A(n13469), .B(n13468), .Z(n13573) );
  XOR U7721 ( .A(n13572), .B(n13573), .Z(n13470) );
  XNOR U7722 ( .A(n13574), .B(n13470), .Z(N51) );
  NANDN U7723 ( .A(n13472), .B(n13471), .Z(n13476) );
  NANDN U7724 ( .A(n13474), .B(n13473), .Z(n13475) );
  AND U7725 ( .A(n13476), .B(n13475), .Z(n13580) );
  AND U7726 ( .A(x[6]), .B(y[13]), .Z(n13478) );
  NAND U7727 ( .A(n13478), .B(n13477), .Z(n13482) );
  NAND U7728 ( .A(n13480), .B(n13479), .Z(n13481) );
  NAND U7729 ( .A(n13482), .B(n13481), .Z(n13671) );
  AND U7730 ( .A(x[16]), .B(y[7]), .Z(n13483) );
  NANDN U7731 ( .A(n13873), .B(n13483), .Z(n13487) );
  NAND U7732 ( .A(n13485), .B(n13484), .Z(n13486) );
  NAND U7733 ( .A(n13487), .B(n13486), .Z(n13669) );
  NAND U7734 ( .A(y[9]), .B(x[15]), .Z(n14307) );
  NANDN U7735 ( .A(n14307), .B(n13598), .Z(n13491) );
  NAND U7736 ( .A(n13489), .B(n13488), .Z(n13490) );
  AND U7737 ( .A(n13491), .B(n13490), .Z(n13613) );
  AND U7738 ( .A(y[18]), .B(x[1]), .Z(n13493) );
  NAND U7739 ( .A(x[8]), .B(y[11]), .Z(n13492) );
  XNOR U7740 ( .A(n13493), .B(n13492), .Z(n13647) );
  NAND U7741 ( .A(y[5]), .B(x[14]), .Z(n13648) );
  XNOR U7742 ( .A(n13647), .B(n13648), .Z(n13611) );
  AND U7743 ( .A(x[2]), .B(y[17]), .Z(n13495) );
  NAND U7744 ( .A(x[13]), .B(y[6]), .Z(n13494) );
  XNOR U7745 ( .A(n13495), .B(n13494), .Z(n13604) );
  XOR U7746 ( .A(n13611), .B(n13610), .Z(n13612) );
  XNOR U7747 ( .A(n13613), .B(n13612), .Z(n13670) );
  XOR U7748 ( .A(n13669), .B(n13670), .Z(n13672) );
  XNOR U7749 ( .A(n13671), .B(n13672), .Z(n13676) );
  NAND U7750 ( .A(n13497), .B(n13496), .Z(n13501) );
  NAND U7751 ( .A(n13499), .B(n13498), .Z(n13500) );
  NAND U7752 ( .A(n13501), .B(n13500), .Z(n13663) );
  NAND U7753 ( .A(n13503), .B(n13502), .Z(n13507) );
  NAND U7754 ( .A(n13505), .B(n13504), .Z(n13506) );
  AND U7755 ( .A(n13507), .B(n13506), .Z(n13664) );
  XOR U7756 ( .A(n13663), .B(n13664), .Z(n13666) );
  AND U7757 ( .A(x[13]), .B(y[15]), .Z(n14923) );
  NANDN U7758 ( .A(n13508), .B(n14923), .Z(n13512) );
  NANDN U7759 ( .A(n13510), .B(n13509), .Z(n13511) );
  AND U7760 ( .A(n13512), .B(n13511), .Z(n13622) );
  AND U7761 ( .A(y[8]), .B(x[11]), .Z(n13514) );
  NAND U7762 ( .A(x[3]), .B(y[16]), .Z(n13513) );
  XNOR U7763 ( .A(n13514), .B(n13513), .Z(n13592) );
  AND U7764 ( .A(x[7]), .B(y[12]), .Z(n13591) );
  XOR U7765 ( .A(n13592), .B(n13591), .Z(n13621) );
  AND U7766 ( .A(x[18]), .B(y[1]), .Z(n13595) );
  XOR U7767 ( .A(n13595), .B(o[19]), .Z(n13652) );
  NAND U7768 ( .A(x[17]), .B(y[2]), .Z(n13653) );
  NAND U7769 ( .A(y[9]), .B(x[10]), .Z(n13654) );
  XOR U7770 ( .A(n13653), .B(n13654), .Z(n13651) );
  XNOR U7771 ( .A(n13652), .B(n13651), .Z(n13620) );
  XOR U7772 ( .A(n13621), .B(n13620), .Z(n13623) );
  XOR U7773 ( .A(n13622), .B(n13623), .Z(n13657) );
  AND U7774 ( .A(x[8]), .B(y[14]), .Z(n13516) );
  NAND U7775 ( .A(n13516), .B(n13515), .Z(n13520) );
  NAND U7776 ( .A(n13518), .B(n13517), .Z(n13519) );
  AND U7777 ( .A(n13520), .B(n13519), .Z(n13617) );
  AND U7778 ( .A(y[19]), .B(x[0]), .Z(n13636) );
  NAND U7779 ( .A(x[19]), .B(y[0]), .Z(n13637) );
  XNOR U7780 ( .A(n13636), .B(n13637), .Z(n13639) );
  ANDN U7781 ( .B(o[18]), .A(n13521), .Z(n13638) );
  XOR U7782 ( .A(n13639), .B(n13638), .Z(n13614) );
  AND U7783 ( .A(x[4]), .B(y[15]), .Z(n13797) );
  AND U7784 ( .A(x[5]), .B(y[14]), .Z(n13523) );
  NAND U7785 ( .A(y[13]), .B(x[6]), .Z(n13522) );
  XOR U7786 ( .A(n13523), .B(n13522), .Z(n13633) );
  XOR U7787 ( .A(n13797), .B(n13633), .Z(n13615) );
  XNOR U7788 ( .A(n13614), .B(n13615), .Z(n13616) );
  XNOR U7789 ( .A(n13617), .B(n13616), .Z(n13658) );
  XOR U7790 ( .A(n13657), .B(n13658), .Z(n13660) );
  AND U7791 ( .A(x[10]), .B(y[17]), .Z(n14549) );
  NANDN U7792 ( .A(n13528), .B(n13527), .Z(n13532) );
  NANDN U7793 ( .A(n13530), .B(n13529), .Z(n13531) );
  AND U7794 ( .A(n13532), .B(n13531), .Z(n13627) );
  AND U7795 ( .A(y[3]), .B(x[16]), .Z(n14224) );
  NAND U7796 ( .A(x[9]), .B(y[10]), .Z(n13533) );
  XNOR U7797 ( .A(n14224), .B(n13533), .Z(n13599) );
  NAND U7798 ( .A(y[4]), .B(x[15]), .Z(n13600) );
  XNOR U7799 ( .A(n13599), .B(n13600), .Z(n13626) );
  XOR U7800 ( .A(n13627), .B(n13626), .Z(n13629) );
  XOR U7801 ( .A(n13628), .B(n13629), .Z(n13659) );
  XOR U7802 ( .A(n13660), .B(n13659), .Z(n13665) );
  XNOR U7803 ( .A(n13666), .B(n13665), .Z(n13675) );
  XOR U7804 ( .A(n13676), .B(n13675), .Z(n13678) );
  XOR U7805 ( .A(n13678), .B(n13677), .Z(n13683) );
  NANDN U7806 ( .A(n13539), .B(n13538), .Z(n13543) );
  NAND U7807 ( .A(n13541), .B(n13540), .Z(n13542) );
  AND U7808 ( .A(n13543), .B(n13542), .Z(n13586) );
  NANDN U7809 ( .A(n13545), .B(n13544), .Z(n13549) );
  NANDN U7810 ( .A(n13547), .B(n13546), .Z(n13548) );
  NAND U7811 ( .A(n13549), .B(n13548), .Z(n13585) );
  XOR U7812 ( .A(n13586), .B(n13585), .Z(n13588) );
  NANDN U7813 ( .A(n13551), .B(n13550), .Z(n13555) );
  NANDN U7814 ( .A(n13553), .B(n13552), .Z(n13554) );
  NAND U7815 ( .A(n13555), .B(n13554), .Z(n13587) );
  XOR U7816 ( .A(n13588), .B(n13587), .Z(n13682) );
  NANDN U7817 ( .A(n13557), .B(n13556), .Z(n13561) );
  OR U7818 ( .A(n13559), .B(n13558), .Z(n13560) );
  NAND U7819 ( .A(n13561), .B(n13560), .Z(n13681) );
  XOR U7820 ( .A(n13682), .B(n13681), .Z(n13684) );
  XNOR U7821 ( .A(n13683), .B(n13684), .Z(n13579) );
  XNOR U7822 ( .A(n13580), .B(n13579), .Z(n13581) );
  XNOR U7823 ( .A(n13581), .B(n13582), .Z(n13578) );
  NANDN U7824 ( .A(n13567), .B(n13566), .Z(n13571) );
  NAND U7825 ( .A(n13569), .B(n13568), .Z(n13570) );
  NAND U7826 ( .A(n13571), .B(n13570), .Z(n13576) );
  XOR U7827 ( .A(n13576), .B(n13577), .Z(n13575) );
  XNOR U7828 ( .A(n13578), .B(n13575), .Z(N52) );
  NANDN U7829 ( .A(n13580), .B(n13579), .Z(n13584) );
  NANDN U7830 ( .A(n13582), .B(n13581), .Z(n13583) );
  AND U7831 ( .A(n13584), .B(n13583), .Z(n14183) );
  NAND U7832 ( .A(n13586), .B(n13585), .Z(n13590) );
  NAND U7833 ( .A(n13588), .B(n13587), .Z(n13589) );
  AND U7834 ( .A(n13590), .B(n13589), .Z(n14163) );
  AND U7835 ( .A(y[16]), .B(x[11]), .Z(n14551) );
  NANDN U7836 ( .A(n13689), .B(n14551), .Z(n13594) );
  NAND U7837 ( .A(n13592), .B(n13591), .Z(n13593) );
  AND U7838 ( .A(n13594), .B(n13593), .Z(n13958) );
  AND U7839 ( .A(n13595), .B(o[19]), .Z(n13805) );
  AND U7840 ( .A(x[0]), .B(y[20]), .Z(n13804) );
  NAND U7841 ( .A(y[0]), .B(x[20]), .Z(n13803) );
  XOR U7842 ( .A(n13804), .B(n13803), .Z(n13806) );
  XOR U7843 ( .A(n13805), .B(n13806), .Z(n13956) );
  NAND U7844 ( .A(x[19]), .B(y[1]), .Z(n13706) );
  XNOR U7845 ( .A(o[20]), .B(n13706), .Z(n13823) );
  AND U7846 ( .A(x[1]), .B(y[19]), .Z(n13597) );
  NAND U7847 ( .A(x[11]), .B(y[9]), .Z(n13596) );
  XOR U7848 ( .A(n13597), .B(n13596), .Z(n13824) );
  XNOR U7849 ( .A(n13823), .B(n13824), .Z(n13955) );
  XNOR U7850 ( .A(n13956), .B(n13955), .Z(n13957) );
  XNOR U7851 ( .A(n13958), .B(n13957), .Z(n13965) );
  AND U7852 ( .A(y[10]), .B(x[16]), .Z(n14520) );
  NAND U7853 ( .A(n14520), .B(n13598), .Z(n13602) );
  NANDN U7854 ( .A(n13600), .B(n13599), .Z(n13601) );
  AND U7855 ( .A(n13602), .B(n13601), .Z(n13964) );
  AND U7856 ( .A(y[17]), .B(x[13]), .Z(n15286) );
  NAND U7857 ( .A(n15286), .B(n13603), .Z(n13607) );
  NANDN U7858 ( .A(n13605), .B(n13604), .Z(n13606) );
  AND U7859 ( .A(n13607), .B(n13606), .Z(n13952) );
  AND U7860 ( .A(y[6]), .B(x[14]), .Z(n13839) );
  AND U7861 ( .A(y[11]), .B(x[9]), .Z(n13838) );
  NAND U7862 ( .A(y[5]), .B(x[15]), .Z(n13837) );
  XOR U7863 ( .A(n13838), .B(n13837), .Z(n13840) );
  XOR U7864 ( .A(n13839), .B(n13840), .Z(n13950) );
  AND U7865 ( .A(x[16]), .B(y[4]), .Z(n13609) );
  NAND U7866 ( .A(x[10]), .B(y[10]), .Z(n13608) );
  XNOR U7867 ( .A(n13609), .B(n13608), .Z(n13883) );
  NAND U7868 ( .A(x[2]), .B(y[18]), .Z(n13884) );
  XNOR U7869 ( .A(n13883), .B(n13884), .Z(n13949) );
  XNOR U7870 ( .A(n13950), .B(n13949), .Z(n13951) );
  XNOR U7871 ( .A(n13952), .B(n13951), .Z(n13963) );
  XOR U7872 ( .A(n13964), .B(n13963), .Z(n13966) );
  XNOR U7873 ( .A(n13965), .B(n13966), .Z(n14129) );
  NANDN U7874 ( .A(n13615), .B(n13614), .Z(n13619) );
  NANDN U7875 ( .A(n13617), .B(n13616), .Z(n13618) );
  NAND U7876 ( .A(n13619), .B(n13618), .Z(n14126) );
  XNOR U7877 ( .A(n14127), .B(n14126), .Z(n14128) );
  XOR U7878 ( .A(n14129), .B(n14128), .Z(n14143) );
  NANDN U7879 ( .A(n13621), .B(n13620), .Z(n13625) );
  NANDN U7880 ( .A(n13623), .B(n13622), .Z(n13624) );
  AND U7881 ( .A(n13625), .B(n13624), .Z(n14141) );
  NANDN U7882 ( .A(n13627), .B(n13626), .Z(n13631) );
  OR U7883 ( .A(n13629), .B(n13628), .Z(n13630) );
  AND U7884 ( .A(n13631), .B(n13630), .Z(n14122) );
  AND U7885 ( .A(x[6]), .B(y[14]), .Z(n13920) );
  NAND U7886 ( .A(n13920), .B(n13632), .Z(n13635) );
  NANDN U7887 ( .A(n13633), .B(n13797), .Z(n13634) );
  AND U7888 ( .A(n13635), .B(n13634), .Z(n13929) );
  AND U7889 ( .A(y[2]), .B(x[18]), .Z(n13641) );
  NAND U7890 ( .A(y[3]), .B(x[17]), .Z(n13640) );
  XNOR U7891 ( .A(n13641), .B(n13640), .Z(n13829) );
  NAND U7892 ( .A(x[12]), .B(y[8]), .Z(n13830) );
  XNOR U7893 ( .A(n13829), .B(n13830), .Z(n13927) );
  XOR U7894 ( .A(n13928), .B(n13927), .Z(n13930) );
  XOR U7895 ( .A(n13929), .B(n13930), .Z(n14121) );
  AND U7896 ( .A(y[7]), .B(x[13]), .Z(n13643) );
  NAND U7897 ( .A(x[3]), .B(y[17]), .Z(n13642) );
  XNOR U7898 ( .A(n13643), .B(n13642), .Z(n13790) );
  XOR U7899 ( .A(n13867), .B(n13790), .Z(n13921) );
  AND U7900 ( .A(x[5]), .B(y[15]), .Z(n13645) );
  NAND U7901 ( .A(y[16]), .B(x[4]), .Z(n13644) );
  XNOR U7902 ( .A(n13645), .B(n13644), .Z(n13800) );
  AND U7903 ( .A(x[7]), .B(y[13]), .Z(n13799) );
  XNOR U7904 ( .A(n13800), .B(n13799), .Z(n13919) );
  XOR U7905 ( .A(n13920), .B(n13919), .Z(n13922) );
  XOR U7906 ( .A(n13921), .B(n13922), .Z(n13945) );
  AND U7907 ( .A(x[8]), .B(y[18]), .Z(n14355) );
  NAND U7908 ( .A(n14355), .B(n13646), .Z(n13650) );
  NANDN U7909 ( .A(n13648), .B(n13647), .Z(n13649) );
  AND U7910 ( .A(n13650), .B(n13649), .Z(n13944) );
  NANDN U7911 ( .A(n13652), .B(n13651), .Z(n13656) );
  IV U7912 ( .A(n13653), .Z(n13827) );
  ANDN U7913 ( .B(n13654), .A(n13827), .Z(n13655) );
  ANDN U7914 ( .B(n13656), .A(n13655), .Z(n13943) );
  XOR U7915 ( .A(n13944), .B(n13943), .Z(n13946) );
  XNOR U7916 ( .A(n13945), .B(n13946), .Z(n14120) );
  XOR U7917 ( .A(n14121), .B(n14120), .Z(n14123) );
  XNOR U7918 ( .A(n14122), .B(n14123), .Z(n14140) );
  XNOR U7919 ( .A(n14141), .B(n14140), .Z(n14142) );
  XOR U7920 ( .A(n14143), .B(n14142), .Z(n14172) );
  NAND U7921 ( .A(n13658), .B(n13657), .Z(n13662) );
  NAND U7922 ( .A(n13660), .B(n13659), .Z(n13661) );
  NAND U7923 ( .A(n13662), .B(n13661), .Z(n14167) );
  NAND U7924 ( .A(n13664), .B(n13663), .Z(n13668) );
  NAND U7925 ( .A(n13666), .B(n13665), .Z(n13667) );
  NAND U7926 ( .A(n13668), .B(n13667), .Z(n14166) );
  XOR U7927 ( .A(n14167), .B(n14166), .Z(n14169) );
  NAND U7928 ( .A(n13670), .B(n13669), .Z(n13674) );
  NAND U7929 ( .A(n13672), .B(n13671), .Z(n13673) );
  NAND U7930 ( .A(n13674), .B(n13673), .Z(n14168) );
  XOR U7931 ( .A(n14169), .B(n14168), .Z(n14173) );
  XOR U7932 ( .A(n14172), .B(n14173), .Z(n14175) );
  NAND U7933 ( .A(n13676), .B(n13675), .Z(n13680) );
  NAND U7934 ( .A(n13678), .B(n13677), .Z(n13679) );
  AND U7935 ( .A(n13680), .B(n13679), .Z(n14174) );
  XOR U7936 ( .A(n14175), .B(n14174), .Z(n14161) );
  NANDN U7937 ( .A(n13682), .B(n13681), .Z(n13686) );
  OR U7938 ( .A(n13684), .B(n13683), .Z(n13685) );
  AND U7939 ( .A(n13686), .B(n13685), .Z(n14160) );
  XNOR U7940 ( .A(n14161), .B(n14160), .Z(n14162) );
  XNOR U7941 ( .A(n14163), .B(n14162), .Z(n14182) );
  XNOR U7942 ( .A(n14183), .B(n14182), .Z(n14184) );
  XNOR U7943 ( .A(n14185), .B(n14184), .Z(N53) );
  AND U7944 ( .A(y[1]), .B(x[20]), .Z(n13786) );
  AND U7945 ( .A(o[21]), .B(n13786), .Z(n13725) );
  AND U7946 ( .A(y[21]), .B(x[1]), .Z(n13726) );
  XOR U7947 ( .A(n13725), .B(n13726), .Z(n13727) );
  AND U7948 ( .A(y[11]), .B(x[11]), .Z(n13728) );
  XOR U7949 ( .A(n13727), .B(n13728), .Z(n13688) );
  AND U7950 ( .A(y[19]), .B(x[3]), .Z(n13719) );
  AND U7951 ( .A(x[14]), .B(y[8]), .Z(n13720) );
  XOR U7952 ( .A(n13719), .B(n13720), .Z(n13722) );
  AND U7953 ( .A(x[19]), .B(y[3]), .Z(n13721) );
  XOR U7954 ( .A(n13722), .B(n13721), .Z(n13687) );
  NAND U7955 ( .A(n13688), .B(n13687), .Z(n13695) );
  XOR U7956 ( .A(n13688), .B(n13687), .Z(n13861) );
  AND U7957 ( .A(x[13]), .B(y[18]), .Z(n15349) );
  NANDN U7958 ( .A(n13689), .B(n15349), .Z(n13693) );
  AND U7959 ( .A(y[18]), .B(x[3]), .Z(n13691) );
  NAND U7960 ( .A(y[8]), .B(x[13]), .Z(n13690) );
  XNOR U7961 ( .A(n13691), .B(n13690), .Z(n13812) );
  AND U7962 ( .A(x[4]), .B(y[17]), .Z(n13811) );
  NAND U7963 ( .A(n13812), .B(n13811), .Z(n13692) );
  NAND U7964 ( .A(n13693), .B(n13692), .Z(n13862) );
  NAND U7965 ( .A(n13861), .B(n13862), .Z(n13694) );
  NAND U7966 ( .A(n13695), .B(n13694), .Z(n14040) );
  AND U7967 ( .A(y[1]), .B(x[21]), .Z(n13783) );
  XNOR U7968 ( .A(n13783), .B(o[22]), .Z(n13760) );
  NAND U7969 ( .A(x[22]), .B(y[0]), .Z(n13758) );
  NAND U7970 ( .A(y[22]), .B(x[0]), .Z(n13757) );
  XOR U7971 ( .A(n13758), .B(n13757), .Z(n13759) );
  XNOR U7972 ( .A(n13760), .B(n13759), .Z(n13698) );
  AND U7973 ( .A(y[15]), .B(x[7]), .Z(n13697) );
  NAND U7974 ( .A(y[14]), .B(x[8]), .Z(n13696) );
  XNOR U7975 ( .A(n13697), .B(n13696), .Z(n13763) );
  XOR U7976 ( .A(n13868), .B(n13763), .Z(n13699) );
  NAND U7977 ( .A(n13698), .B(n13699), .Z(n13705) );
  XOR U7978 ( .A(n13699), .B(n13698), .Z(n13714) );
  AND U7979 ( .A(y[15]), .B(x[14]), .Z(n15070) );
  NAND U7980 ( .A(n15070), .B(n13767), .Z(n13703) );
  AND U7981 ( .A(x[7]), .B(y[14]), .Z(n14069) );
  AND U7982 ( .A(y[7]), .B(x[14]), .Z(n13701) );
  AND U7983 ( .A(y[15]), .B(x[6]), .Z(n13700) );
  XOR U7984 ( .A(n13701), .B(n13700), .Z(n13817) );
  NAND U7985 ( .A(n14069), .B(n13817), .Z(n13702) );
  NAND U7986 ( .A(n13703), .B(n13702), .Z(n13715) );
  NAND U7987 ( .A(n13714), .B(n13715), .Z(n13704) );
  NAND U7988 ( .A(n13705), .B(n13704), .Z(n14039) );
  XOR U7989 ( .A(n14040), .B(n14039), .Z(n14042) );
  AND U7990 ( .A(y[21]), .B(x[0]), .Z(n13708) );
  AND U7991 ( .A(y[0]), .B(x[21]), .Z(n13707) );
  NAND U7992 ( .A(n13708), .B(n13707), .Z(n13710) );
  ANDN U7993 ( .B(o[20]), .A(n13706), .Z(n13834) );
  XOR U7994 ( .A(n13708), .B(n13707), .Z(n13833) );
  NAND U7995 ( .A(n13834), .B(n13833), .Z(n13709) );
  AND U7996 ( .A(n13710), .B(n13709), .Z(n13712) );
  NAND U7997 ( .A(x[18]), .B(y[3]), .Z(n13828) );
  XNOR U7998 ( .A(n13711), .B(n13828), .Z(n13784) );
  NAND U7999 ( .A(x[1]), .B(y[20]), .Z(n13785) );
  NAND U8000 ( .A(n13712), .B(n13713), .Z(n13717) );
  XOR U8001 ( .A(n13713), .B(n13712), .Z(n13865) );
  XNOR U8002 ( .A(n13715), .B(n13714), .Z(n13866) );
  NAND U8003 ( .A(n13865), .B(n13866), .Z(n13716) );
  AND U8004 ( .A(n13717), .B(n13716), .Z(n14041) );
  XNOR U8005 ( .A(n14042), .B(n14041), .Z(n14101) );
  AND U8006 ( .A(x[15]), .B(y[8]), .Z(n14063) );
  NAND U8007 ( .A(x[6]), .B(y[17]), .Z(n14064) );
  XNOR U8008 ( .A(n14063), .B(n14064), .Z(n14066) );
  AND U8009 ( .A(x[11]), .B(y[12]), .Z(n14065) );
  XNOR U8010 ( .A(n14066), .B(n14065), .Z(n14012) );
  NAND U8011 ( .A(x[10]), .B(y[13]), .Z(n14010) );
  NAND U8012 ( .A(x[7]), .B(y[16]), .Z(n13718) );
  XNOR U8013 ( .A(n14268), .B(n13718), .Z(n14070) );
  XNOR U8014 ( .A(n14071), .B(n14070), .Z(n14009) );
  XOR U8015 ( .A(n14010), .B(n14009), .Z(n14011) );
  XNOR U8016 ( .A(n14012), .B(n14011), .Z(n13987) );
  NAND U8017 ( .A(n13720), .B(n13719), .Z(n13724) );
  NAND U8018 ( .A(n13722), .B(n13721), .Z(n13723) );
  NAND U8019 ( .A(n13724), .B(n13723), .Z(n13986) );
  NAND U8020 ( .A(n13726), .B(n13725), .Z(n13730) );
  NAND U8021 ( .A(n13728), .B(n13727), .Z(n13729) );
  NAND U8022 ( .A(n13730), .B(n13729), .Z(n13985) );
  XOR U8023 ( .A(n13986), .B(n13985), .Z(n13988) );
  XNOR U8024 ( .A(n13987), .B(n13988), .Z(n14099) );
  AND U8025 ( .A(x[17]), .B(y[5]), .Z(n13777) );
  AND U8026 ( .A(y[17]), .B(x[5]), .Z(n13778) );
  XOR U8027 ( .A(n13777), .B(n13778), .Z(n13779) );
  AND U8028 ( .A(y[6]), .B(x[16]), .Z(n13780) );
  XOR U8029 ( .A(n13779), .B(n13780), .Z(n13734) );
  AND U8030 ( .A(y[4]), .B(x[18]), .Z(n13732) );
  NAND U8031 ( .A(x[12]), .B(y[10]), .Z(n13731) );
  XNOR U8032 ( .A(n13732), .B(n13731), .Z(n13754) );
  AND U8033 ( .A(x[4]), .B(y[18]), .Z(n13753) );
  XOR U8034 ( .A(n13754), .B(n13753), .Z(n13733) );
  NAND U8035 ( .A(n13734), .B(n13733), .Z(n13740) );
  XOR U8036 ( .A(n13734), .B(n13733), .Z(n13878) );
  AND U8037 ( .A(x[17]), .B(y[9]), .Z(n14515) );
  NAND U8038 ( .A(n14515), .B(n13752), .Z(n13738) );
  AND U8039 ( .A(x[12]), .B(y[9]), .Z(n13736) );
  NAND U8040 ( .A(y[4]), .B(x[17]), .Z(n13735) );
  XNOR U8041 ( .A(n13736), .B(n13735), .Z(n13814) );
  AND U8042 ( .A(y[19]), .B(x[2]), .Z(n13813) );
  NAND U8043 ( .A(n13814), .B(n13813), .Z(n13737) );
  NAND U8044 ( .A(n13738), .B(n13737), .Z(n13879) );
  NAND U8045 ( .A(n13878), .B(n13879), .Z(n13739) );
  AND U8046 ( .A(n13740), .B(n13739), .Z(n14098) );
  XOR U8047 ( .A(n14099), .B(n14098), .Z(n14100) );
  XNOR U8048 ( .A(n14101), .B(n14100), .Z(n14093) );
  AND U8049 ( .A(y[7]), .B(x[15]), .Z(n13742) );
  NAND U8050 ( .A(y[16]), .B(x[6]), .Z(n13741) );
  XNOR U8051 ( .A(n13742), .B(n13741), .Z(n13768) );
  AND U8052 ( .A(x[10]), .B(y[12]), .Z(n13769) );
  XOR U8053 ( .A(n13768), .B(n13769), .Z(n13749) );
  AND U8054 ( .A(x[20]), .B(y[2]), .Z(n13744) );
  NAND U8055 ( .A(x[13]), .B(y[9]), .Z(n13743) );
  XNOR U8056 ( .A(n13744), .B(n13743), .Z(n13773) );
  AND U8057 ( .A(x[2]), .B(y[20]), .Z(n13774) );
  XOR U8058 ( .A(n13773), .B(n13774), .Z(n13748) );
  NAND U8059 ( .A(n13749), .B(n13748), .Z(n13751) );
  NAND U8060 ( .A(y[16]), .B(x[5]), .Z(n13798) );
  AND U8061 ( .A(y[5]), .B(x[16]), .Z(n13745) );
  NANDN U8062 ( .A(n13798), .B(n13745), .Z(n13747) );
  AND U8063 ( .A(y[6]), .B(x[15]), .Z(n13835) );
  NAND U8064 ( .A(n13836), .B(n13835), .Z(n13746) );
  AND U8065 ( .A(n13747), .B(n13746), .Z(n13864) );
  XOR U8066 ( .A(n13749), .B(n13748), .Z(n13863) );
  NANDN U8067 ( .A(n13864), .B(n13863), .Z(n13750) );
  NAND U8068 ( .A(n13751), .B(n13750), .Z(n14046) );
  AND U8069 ( .A(y[10]), .B(x[18]), .Z(n15101) );
  NAND U8070 ( .A(n15101), .B(n13752), .Z(n13756) );
  NAND U8071 ( .A(n13754), .B(n13753), .Z(n13755) );
  NAND U8072 ( .A(n13756), .B(n13755), .Z(n14022) );
  NAND U8073 ( .A(n13758), .B(n13757), .Z(n13762) );
  NAND U8074 ( .A(n13760), .B(n13759), .Z(n13761) );
  AND U8075 ( .A(n13762), .B(n13761), .Z(n14021) );
  XOR U8076 ( .A(n14022), .B(n14021), .Z(n14024) );
  NAND U8077 ( .A(n14069), .B(n14071), .Z(n13765) );
  NAND U8078 ( .A(n13763), .B(n13868), .Z(n13764) );
  NAND U8079 ( .A(n13765), .B(n13764), .Z(n14028) );
  AND U8080 ( .A(x[23]), .B(y[0]), .Z(n14055) );
  AND U8081 ( .A(x[0]), .B(y[23]), .Z(n14056) );
  XOR U8082 ( .A(n14055), .B(n14056), .Z(n14057) );
  NAND U8083 ( .A(x[22]), .B(y[1]), .Z(n14085) );
  XNOR U8084 ( .A(o[23]), .B(n14085), .Z(n14058) );
  XOR U8085 ( .A(n14057), .B(n14058), .Z(n14027) );
  XOR U8086 ( .A(n14028), .B(n14027), .Z(n14029) );
  AND U8087 ( .A(y[3]), .B(x[20]), .Z(n14639) );
  NAND U8088 ( .A(y[7]), .B(x[16]), .Z(n13766) );
  XNOR U8089 ( .A(n14639), .B(n13766), .Z(n14081) );
  NAND U8090 ( .A(x[19]), .B(y[4]), .Z(n14082) );
  XNOR U8091 ( .A(n14081), .B(n14082), .Z(n14030) );
  XOR U8092 ( .A(n14029), .B(n14030), .Z(n14023) );
  XOR U8093 ( .A(n14024), .B(n14023), .Z(n14045) );
  XOR U8094 ( .A(n14046), .B(n14045), .Z(n14048) );
  AND U8095 ( .A(y[16]), .B(x[15]), .Z(n15350) );
  NAND U8096 ( .A(n15350), .B(n13767), .Z(n13771) );
  NAND U8097 ( .A(n13769), .B(n13768), .Z(n13770) );
  NAND U8098 ( .A(n13771), .B(n13770), .Z(n14036) );
  AND U8099 ( .A(y[9]), .B(x[14]), .Z(n13991) );
  AND U8100 ( .A(x[3]), .B(y[20]), .Z(n13992) );
  XOR U8101 ( .A(n13991), .B(n13992), .Z(n13993) );
  AND U8102 ( .A(x[4]), .B(y[19]), .Z(n13994) );
  XOR U8103 ( .A(n13993), .B(n13994), .Z(n14033) );
  AND U8104 ( .A(x[5]), .B(y[18]), .Z(n14003) );
  NAND U8105 ( .A(x[18]), .B(y[5]), .Z(n14004) );
  XNOR U8106 ( .A(n14003), .B(n14004), .Z(n14005) );
  NAND U8107 ( .A(y[6]), .B(x[17]), .Z(n14006) );
  XNOR U8108 ( .A(n14005), .B(n14006), .Z(n14034) );
  XOR U8109 ( .A(n14033), .B(n14034), .Z(n14035) );
  XOR U8110 ( .A(n14036), .B(n14035), .Z(n14089) );
  AND U8111 ( .A(y[9]), .B(x[20]), .Z(n15058) );
  NAND U8112 ( .A(n15058), .B(n13772), .Z(n13776) );
  NAND U8113 ( .A(n13774), .B(n13773), .Z(n13775) );
  NAND U8114 ( .A(n13776), .B(n13775), .Z(n14087) );
  NAND U8115 ( .A(n13778), .B(n13777), .Z(n13782) );
  NAND U8116 ( .A(n13780), .B(n13779), .Z(n13781) );
  NAND U8117 ( .A(n13782), .B(n13781), .Z(n14018) );
  NAND U8118 ( .A(n13783), .B(o[22]), .Z(n14077) );
  NAND U8119 ( .A(y[22]), .B(x[1]), .Z(n14075) );
  NAND U8120 ( .A(y[11]), .B(x[12]), .Z(n14074) );
  XOR U8121 ( .A(n14075), .B(n14074), .Z(n14076) );
  XNOR U8122 ( .A(n14077), .B(n14076), .Z(n14015) );
  AND U8123 ( .A(y[21]), .B(x[2]), .Z(n13997) );
  AND U8124 ( .A(y[10]), .B(x[13]), .Z(n13998) );
  XOR U8125 ( .A(n13997), .B(n13998), .Z(n13999) );
  AND U8126 ( .A(y[2]), .B(x[21]), .Z(n14000) );
  XOR U8127 ( .A(n13999), .B(n14000), .Z(n14016) );
  XOR U8128 ( .A(n14015), .B(n14016), .Z(n14017) );
  XOR U8129 ( .A(n14018), .B(n14017), .Z(n14086) );
  XOR U8130 ( .A(n14087), .B(n14086), .Z(n14088) );
  XOR U8131 ( .A(n14089), .B(n14088), .Z(n14047) );
  XOR U8132 ( .A(n14048), .B(n14047), .Z(n14092) );
  XOR U8133 ( .A(n14093), .B(n14092), .Z(n14095) );
  XOR U8134 ( .A(n13785), .B(n13784), .Z(n13794) );
  XOR U8135 ( .A(o[21]), .B(n13786), .Z(n13875) );
  AND U8136 ( .A(y[2]), .B(x[19]), .Z(n13788) );
  AND U8137 ( .A(x[11]), .B(y[10]), .Z(n13787) );
  XOR U8138 ( .A(n13788), .B(n13787), .Z(n13874) );
  XOR U8139 ( .A(n13875), .B(n13874), .Z(n13793) );
  NAND U8140 ( .A(n13794), .B(n13793), .Z(n13796) );
  NAND U8141 ( .A(n15286), .B(n13789), .Z(n13792) );
  NAND U8142 ( .A(n13867), .B(n13790), .Z(n13791) );
  AND U8143 ( .A(n13792), .B(n13791), .Z(n13888) );
  XOR U8144 ( .A(n13794), .B(n13793), .Z(n13887) );
  NANDN U8145 ( .A(n13888), .B(n13887), .Z(n13795) );
  AND U8146 ( .A(n13796), .B(n13795), .Z(n13821) );
  NANDN U8147 ( .A(n13798), .B(n13797), .Z(n13802) );
  NAND U8148 ( .A(n13800), .B(n13799), .Z(n13801) );
  AND U8149 ( .A(n13802), .B(n13801), .Z(n13810) );
  NANDN U8150 ( .A(n13804), .B(n13803), .Z(n13808) );
  OR U8151 ( .A(n13806), .B(n13805), .Z(n13807) );
  AND U8152 ( .A(n13808), .B(n13807), .Z(n13809) );
  NANDN U8153 ( .A(n13810), .B(n13809), .Z(n13819) );
  XOR U8154 ( .A(n13810), .B(n13809), .Z(n13891) );
  XOR U8155 ( .A(n13812), .B(n13811), .Z(n13850) );
  XOR U8156 ( .A(n13814), .B(n13813), .Z(n13849) );
  XOR U8157 ( .A(n13850), .B(n13849), .Z(n13852) );
  AND U8158 ( .A(x[9]), .B(y[12]), .Z(n13816) );
  NAND U8159 ( .A(y[13]), .B(x[8]), .Z(n13815) );
  XNOR U8160 ( .A(n13816), .B(n13815), .Z(n13870) );
  XOR U8161 ( .A(n14069), .B(n13817), .Z(n13869) );
  XOR U8162 ( .A(n13870), .B(n13869), .Z(n13851) );
  XOR U8163 ( .A(n13852), .B(n13851), .Z(n13892) );
  NANDN U8164 ( .A(n13891), .B(n13892), .Z(n13818) );
  AND U8165 ( .A(n13819), .B(n13818), .Z(n13820) );
  NAND U8166 ( .A(n13821), .B(n13820), .Z(n13848) );
  XOR U8167 ( .A(n13821), .B(n13820), .Z(n13916) );
  NAND U8168 ( .A(y[19]), .B(x[11]), .Z(n15285) );
  NANDN U8169 ( .A(n15285), .B(n13822), .Z(n13826) );
  NANDN U8170 ( .A(n13824), .B(n13823), .Z(n13825) );
  NAND U8171 ( .A(n13826), .B(n13825), .Z(n13844) );
  NANDN U8172 ( .A(n13828), .B(n13827), .Z(n13832) );
  NANDN U8173 ( .A(n13830), .B(n13829), .Z(n13831) );
  NAND U8174 ( .A(n13832), .B(n13831), .Z(n13843) );
  NAND U8175 ( .A(n13844), .B(n13843), .Z(n13846) );
  XOR U8176 ( .A(n13834), .B(n13833), .Z(n13856) );
  XOR U8177 ( .A(n13836), .B(n13835), .Z(n13855) );
  XOR U8178 ( .A(n13856), .B(n13855), .Z(n13858) );
  NANDN U8179 ( .A(n13838), .B(n13837), .Z(n13842) );
  OR U8180 ( .A(n13840), .B(n13839), .Z(n13841) );
  AND U8181 ( .A(n13842), .B(n13841), .Z(n13857) );
  XOR U8182 ( .A(n13858), .B(n13857), .Z(n13918) );
  XOR U8183 ( .A(n13844), .B(n13843), .Z(n13917) );
  NAND U8184 ( .A(n13918), .B(n13917), .Z(n13845) );
  AND U8185 ( .A(n13846), .B(n13845), .Z(n13915) );
  NAND U8186 ( .A(n13916), .B(n13915), .Z(n13847) );
  AND U8187 ( .A(n13848), .B(n13847), .Z(n14094) );
  XNOR U8188 ( .A(n14095), .B(n14094), .Z(n14113) );
  NAND U8189 ( .A(n13850), .B(n13849), .Z(n13854) );
  NAND U8190 ( .A(n13852), .B(n13851), .Z(n13853) );
  NAND U8191 ( .A(n13854), .B(n13853), .Z(n13911) );
  NAND U8192 ( .A(n13856), .B(n13855), .Z(n13860) );
  NAND U8193 ( .A(n13858), .B(n13857), .Z(n13859) );
  NAND U8194 ( .A(n13860), .B(n13859), .Z(n13909) );
  XNOR U8195 ( .A(n13862), .B(n13861), .Z(n13898) );
  XOR U8196 ( .A(n13864), .B(n13863), .Z(n13897) );
  XOR U8197 ( .A(n13898), .B(n13897), .Z(n13899) );
  XNOR U8198 ( .A(n13866), .B(n13865), .Z(n13900) );
  XOR U8199 ( .A(n13899), .B(n13900), .Z(n13910) );
  XNOR U8200 ( .A(n13909), .B(n13910), .Z(n13912) );
  XOR U8201 ( .A(n13911), .B(n13912), .Z(n13880) );
  NAND U8202 ( .A(n13868), .B(n13867), .Z(n13872) );
  NAND U8203 ( .A(n13870), .B(n13869), .Z(n13871) );
  NAND U8204 ( .A(n13872), .B(n13871), .Z(n13905) );
  AND U8205 ( .A(y[10]), .B(x[19]), .Z(n14905) );
  NANDN U8206 ( .A(n13873), .B(n14905), .Z(n13877) );
  NAND U8207 ( .A(n13875), .B(n13874), .Z(n13876) );
  NAND U8208 ( .A(n13877), .B(n13876), .Z(n13903) );
  XOR U8209 ( .A(n13879), .B(n13878), .Z(n13904) );
  XOR U8210 ( .A(n13903), .B(n13904), .Z(n13906) );
  XOR U8211 ( .A(n13905), .B(n13906), .Z(n13881) );
  NANDN U8212 ( .A(n13880), .B(n13881), .Z(n13896) );
  XNOR U8213 ( .A(n13881), .B(n13880), .Z(n13937) );
  NAND U8214 ( .A(n14520), .B(n13882), .Z(n13886) );
  NANDN U8215 ( .A(n13884), .B(n13883), .Z(n13885) );
  AND U8216 ( .A(n13886), .B(n13885), .Z(n13890) );
  XNOR U8217 ( .A(n13888), .B(n13887), .Z(n13889) );
  NANDN U8218 ( .A(n13890), .B(n13889), .Z(n13894) );
  XNOR U8219 ( .A(n13890), .B(n13889), .Z(n13942) );
  XNOR U8220 ( .A(n13892), .B(n13891), .Z(n13941) );
  NAND U8221 ( .A(n13942), .B(n13941), .Z(n13893) );
  NAND U8222 ( .A(n13894), .B(n13893), .Z(n13938) );
  NAND U8223 ( .A(n13937), .B(n13938), .Z(n13895) );
  AND U8224 ( .A(n13896), .B(n13895), .Z(n14111) );
  NAND U8225 ( .A(n13898), .B(n13897), .Z(n13902) );
  NANDN U8226 ( .A(n13900), .B(n13899), .Z(n13901) );
  NAND U8227 ( .A(n13902), .B(n13901), .Z(n14104) );
  NAND U8228 ( .A(n13904), .B(n13903), .Z(n13908) );
  NAND U8229 ( .A(n13906), .B(n13905), .Z(n13907) );
  AND U8230 ( .A(n13908), .B(n13907), .Z(n14105) );
  XOR U8231 ( .A(n14104), .B(n14105), .Z(n14107) );
  NAND U8232 ( .A(n13910), .B(n13909), .Z(n13914) );
  NANDN U8233 ( .A(n13912), .B(n13911), .Z(n13913) );
  AND U8234 ( .A(n13914), .B(n13913), .Z(n14106) );
  XOR U8235 ( .A(n14107), .B(n14106), .Z(n14110) );
  XOR U8236 ( .A(n14111), .B(n14110), .Z(n14112) );
  XOR U8237 ( .A(n14113), .B(n14112), .Z(n13983) );
  XOR U8238 ( .A(n13916), .B(n13915), .Z(n13936) );
  XOR U8239 ( .A(n13918), .B(n13917), .Z(n13926) );
  NANDN U8240 ( .A(n13920), .B(n13919), .Z(n13924) );
  OR U8241 ( .A(n13922), .B(n13921), .Z(n13923) );
  NAND U8242 ( .A(n13924), .B(n13923), .Z(n13925) );
  NANDN U8243 ( .A(n13926), .B(n13925), .Z(n13934) );
  XOR U8244 ( .A(n13926), .B(n13925), .Z(n14134) );
  NANDN U8245 ( .A(n13928), .B(n13927), .Z(n13932) );
  OR U8246 ( .A(n13930), .B(n13929), .Z(n13931) );
  AND U8247 ( .A(n13932), .B(n13931), .Z(n14135) );
  NANDN U8248 ( .A(n14134), .B(n14135), .Z(n13933) );
  AND U8249 ( .A(n13934), .B(n13933), .Z(n13935) );
  NANDN U8250 ( .A(n13936), .B(n13935), .Z(n13940) );
  XOR U8251 ( .A(n13936), .B(n13935), .Z(n13977) );
  XOR U8252 ( .A(n13938), .B(n13937), .Z(n13978) );
  NANDN U8253 ( .A(n13977), .B(n13978), .Z(n13939) );
  AND U8254 ( .A(n13940), .B(n13939), .Z(n13984) );
  XOR U8255 ( .A(n13942), .B(n13941), .Z(n13962) );
  NANDN U8256 ( .A(n13944), .B(n13943), .Z(n13948) );
  OR U8257 ( .A(n13946), .B(n13945), .Z(n13947) );
  NAND U8258 ( .A(n13948), .B(n13947), .Z(n13973) );
  NANDN U8259 ( .A(n13950), .B(n13949), .Z(n13954) );
  NANDN U8260 ( .A(n13952), .B(n13951), .Z(n13953) );
  NAND U8261 ( .A(n13954), .B(n13953), .Z(n13972) );
  NANDN U8262 ( .A(n13956), .B(n13955), .Z(n13960) );
  NANDN U8263 ( .A(n13958), .B(n13957), .Z(n13959) );
  NAND U8264 ( .A(n13960), .B(n13959), .Z(n13971) );
  XNOR U8265 ( .A(n13972), .B(n13971), .Z(n13974) );
  XOR U8266 ( .A(n13973), .B(n13974), .Z(n13961) );
  NANDN U8267 ( .A(n13962), .B(n13961), .Z(n13970) );
  XNOR U8268 ( .A(n13962), .B(n13961), .Z(n14139) );
  NANDN U8269 ( .A(n13964), .B(n13963), .Z(n13968) );
  NANDN U8270 ( .A(n13966), .B(n13965), .Z(n13967) );
  AND U8271 ( .A(n13968), .B(n13967), .Z(n14138) );
  NAND U8272 ( .A(n14139), .B(n14138), .Z(n13969) );
  AND U8273 ( .A(n13970), .B(n13969), .Z(n13980) );
  NAND U8274 ( .A(n13972), .B(n13971), .Z(n13976) );
  NANDN U8275 ( .A(n13974), .B(n13973), .Z(n13975) );
  NAND U8276 ( .A(n13976), .B(n13975), .Z(n13979) );
  NAND U8277 ( .A(n13980), .B(n13979), .Z(n13982) );
  XOR U8278 ( .A(n13978), .B(n13977), .Z(n14118) );
  XOR U8279 ( .A(n13980), .B(n13979), .Z(n14119) );
  NANDN U8280 ( .A(n14118), .B(n14119), .Z(n13981) );
  NAND U8281 ( .A(n13982), .B(n13981), .Z(n14116) );
  XOR U8282 ( .A(n13984), .B(n13983), .Z(n14117) );
  NAND U8283 ( .A(n13986), .B(n13985), .Z(n13990) );
  NAND U8284 ( .A(n13988), .B(n13987), .Z(n13989) );
  NAND U8285 ( .A(n13990), .B(n13989), .Z(n14315) );
  NAND U8286 ( .A(n13992), .B(n13991), .Z(n13996) );
  NAND U8287 ( .A(n13994), .B(n13993), .Z(n13995) );
  AND U8288 ( .A(n13996), .B(n13995), .Z(n14245) );
  NAND U8289 ( .A(n13998), .B(n13997), .Z(n14002) );
  NAND U8290 ( .A(n14000), .B(n13999), .Z(n14001) );
  AND U8291 ( .A(n14002), .B(n14001), .Z(n14244) );
  XOR U8292 ( .A(n14245), .B(n14244), .Z(n14247) );
  NANDN U8293 ( .A(n14004), .B(n14003), .Z(n14008) );
  NANDN U8294 ( .A(n14006), .B(n14005), .Z(n14007) );
  AND U8295 ( .A(n14008), .B(n14007), .Z(n14220) );
  AND U8296 ( .A(y[17]), .B(x[7]), .Z(n14286) );
  NAND U8297 ( .A(y[6]), .B(x[18]), .Z(n14287) );
  XNOR U8298 ( .A(n14286), .B(n14287), .Z(n14289) );
  AND U8299 ( .A(x[17]), .B(y[7]), .Z(n14288) );
  XOR U8300 ( .A(n14289), .B(n14288), .Z(n14219) );
  NAND U8301 ( .A(x[23]), .B(y[1]), .Z(n14293) );
  XNOR U8302 ( .A(o[24]), .B(n14293), .Z(n14303) );
  AND U8303 ( .A(y[0]), .B(x[24]), .Z(n14300) );
  NAND U8304 ( .A(y[24]), .B(x[0]), .Z(n14301) );
  XNOR U8305 ( .A(n14300), .B(n14301), .Z(n14302) );
  XNOR U8306 ( .A(n14303), .B(n14302), .Z(n14218) );
  XOR U8307 ( .A(n14219), .B(n14218), .Z(n14221) );
  XNOR U8308 ( .A(n14220), .B(n14221), .Z(n14246) );
  XNOR U8309 ( .A(n14247), .B(n14246), .Z(n14313) );
  NAND U8310 ( .A(n14010), .B(n14009), .Z(n14014) );
  NAND U8311 ( .A(n14012), .B(n14011), .Z(n14013) );
  AND U8312 ( .A(n14014), .B(n14013), .Z(n14312) );
  XOR U8313 ( .A(n14313), .B(n14312), .Z(n14314) );
  XOR U8314 ( .A(n14315), .B(n14314), .Z(n14259) );
  NAND U8315 ( .A(n14016), .B(n14015), .Z(n14020) );
  NAND U8316 ( .A(n14018), .B(n14017), .Z(n14019) );
  NAND U8317 ( .A(n14020), .B(n14019), .Z(n14257) );
  NAND U8318 ( .A(n14022), .B(n14021), .Z(n14026) );
  NAND U8319 ( .A(n14024), .B(n14023), .Z(n14025) );
  NAND U8320 ( .A(n14026), .B(n14025), .Z(n14215) );
  NAND U8321 ( .A(n14028), .B(n14027), .Z(n14032) );
  NAND U8322 ( .A(n14030), .B(n14029), .Z(n14031) );
  NAND U8323 ( .A(n14032), .B(n14031), .Z(n14213) );
  NAND U8324 ( .A(n14034), .B(n14033), .Z(n14038) );
  NAND U8325 ( .A(n14036), .B(n14035), .Z(n14037) );
  NAND U8326 ( .A(n14038), .B(n14037), .Z(n14212) );
  XOR U8327 ( .A(n14213), .B(n14212), .Z(n14214) );
  XOR U8328 ( .A(n14215), .B(n14214), .Z(n14256) );
  XOR U8329 ( .A(n14257), .B(n14256), .Z(n14258) );
  XNOR U8330 ( .A(n14259), .B(n14258), .Z(n14207) );
  NAND U8331 ( .A(n14040), .B(n14039), .Z(n14044) );
  NAND U8332 ( .A(n14042), .B(n14041), .Z(n14043) );
  AND U8333 ( .A(n14044), .B(n14043), .Z(n14206) );
  XOR U8334 ( .A(n14207), .B(n14206), .Z(n14209) );
  NAND U8335 ( .A(n14046), .B(n14045), .Z(n14050) );
  NAND U8336 ( .A(n14048), .B(n14047), .Z(n14049) );
  AND U8337 ( .A(n14050), .B(n14049), .Z(n14321) );
  AND U8338 ( .A(y[16]), .B(x[8]), .Z(n14052) );
  NAND U8339 ( .A(x[14]), .B(y[10]), .Z(n14051) );
  XNOR U8340 ( .A(n14052), .B(n14051), .Z(n14274) );
  NAND U8341 ( .A(x[11]), .B(y[13]), .Z(n14275) );
  XNOR U8342 ( .A(n14274), .B(n14275), .Z(n14269) );
  AND U8343 ( .A(x[9]), .B(y[15]), .Z(n14054) );
  NAND U8344 ( .A(y[14]), .B(x[10]), .Z(n14053) );
  XOR U8345 ( .A(n14054), .B(n14053), .Z(n14270) );
  XOR U8346 ( .A(n14269), .B(n14270), .Z(n14296) );
  AND U8347 ( .A(y[21]), .B(x[3]), .Z(n14306) );
  NAND U8348 ( .A(x[4]), .B(y[20]), .Z(n14309) );
  XOR U8349 ( .A(n14308), .B(n14309), .Z(n14294) );
  NAND U8350 ( .A(n14056), .B(n14055), .Z(n14060) );
  NAND U8351 ( .A(n14058), .B(n14057), .Z(n14059) );
  AND U8352 ( .A(n14060), .B(n14059), .Z(n14295) );
  XNOR U8353 ( .A(n14294), .B(n14295), .Z(n14297) );
  AND U8354 ( .A(x[6]), .B(y[18]), .Z(n14582) );
  AND U8355 ( .A(y[4]), .B(x[20]), .Z(n14229) );
  XOR U8356 ( .A(n14582), .B(n14229), .Z(n14231) );
  AND U8357 ( .A(x[19]), .B(y[5]), .Z(n14230) );
  XOR U8358 ( .A(n14231), .B(n14230), .Z(n14239) );
  AND U8359 ( .A(y[3]), .B(x[21]), .Z(n14062) );
  NAND U8360 ( .A(y[8]), .B(x[16]), .Z(n14061) );
  XNOR U8361 ( .A(n14062), .B(n14061), .Z(n14226) );
  AND U8362 ( .A(y[19]), .B(x[5]), .Z(n14225) );
  XNOR U8363 ( .A(n14226), .B(n14225), .Z(n14238) );
  XNOR U8364 ( .A(n14239), .B(n14238), .Z(n14240) );
  NANDN U8365 ( .A(n14064), .B(n14063), .Z(n14068) );
  NAND U8366 ( .A(n14066), .B(n14065), .Z(n14067) );
  NAND U8367 ( .A(n14068), .B(n14067), .Z(n14241) );
  XOR U8368 ( .A(n14240), .B(n14241), .Z(n14252) );
  NAND U8369 ( .A(n14438), .B(n14069), .Z(n14073) );
  NAND U8370 ( .A(n14071), .B(n14070), .Z(n14072) );
  NAND U8371 ( .A(n14073), .B(n14072), .Z(n14250) );
  NAND U8372 ( .A(n14075), .B(n14074), .Z(n14079) );
  NAND U8373 ( .A(n14077), .B(n14076), .Z(n14078) );
  AND U8374 ( .A(n14079), .B(n14078), .Z(n14251) );
  XOR U8375 ( .A(n14250), .B(n14251), .Z(n14253) );
  XOR U8376 ( .A(n14252), .B(n14253), .Z(n14262) );
  AND U8377 ( .A(y[7]), .B(x[20]), .Z(n14080) );
  NAND U8378 ( .A(n14080), .B(n14224), .Z(n14084) );
  NANDN U8379 ( .A(n14082), .B(n14081), .Z(n14083) );
  AND U8380 ( .A(n14084), .B(n14083), .Z(n14237) );
  AND U8381 ( .A(y[22]), .B(x[2]), .Z(n14283) );
  NAND U8382 ( .A(x[22]), .B(y[2]), .Z(n14285) );
  XOR U8383 ( .A(n14284), .B(n14285), .Z(n14282) );
  XOR U8384 ( .A(n14283), .B(n14282), .Z(n14234) );
  AND U8385 ( .A(x[1]), .B(y[23]), .Z(n14278) );
  XOR U8386 ( .A(n14279), .B(n14278), .Z(n14281) );
  ANDN U8387 ( .B(o[23]), .A(n14085), .Z(n14280) );
  XOR U8388 ( .A(n14281), .B(n14280), .Z(n14235) );
  XOR U8389 ( .A(n14234), .B(n14235), .Z(n14236) );
  XNOR U8390 ( .A(n14237), .B(n14236), .Z(n14263) );
  XOR U8391 ( .A(n14262), .B(n14263), .Z(n14265) );
  XNOR U8392 ( .A(n14264), .B(n14265), .Z(n14318) );
  NAND U8393 ( .A(n14087), .B(n14086), .Z(n14091) );
  NAND U8394 ( .A(n14089), .B(n14088), .Z(n14090) );
  AND U8395 ( .A(n14091), .B(n14090), .Z(n14319) );
  XOR U8396 ( .A(n14318), .B(n14319), .Z(n14320) );
  XOR U8397 ( .A(n14321), .B(n14320), .Z(n14208) );
  XOR U8398 ( .A(n14209), .B(n14208), .Z(n14331) );
  NAND U8399 ( .A(n14093), .B(n14092), .Z(n14097) );
  NAND U8400 ( .A(n14095), .B(n14094), .Z(n14096) );
  NAND U8401 ( .A(n14097), .B(n14096), .Z(n14326) );
  NAND U8402 ( .A(n14099), .B(n14098), .Z(n14103) );
  NAND U8403 ( .A(n14101), .B(n14100), .Z(n14102) );
  AND U8404 ( .A(n14103), .B(n14102), .Z(n14325) );
  NAND U8405 ( .A(n14105), .B(n14104), .Z(n14109) );
  NAND U8406 ( .A(n14107), .B(n14106), .Z(n14108) );
  AND U8407 ( .A(n14109), .B(n14108), .Z(n14324) );
  XOR U8408 ( .A(n14325), .B(n14324), .Z(n14327) );
  XOR U8409 ( .A(n14326), .B(n14327), .Z(n14330) );
  NAND U8410 ( .A(n14111), .B(n14110), .Z(n14115) );
  NAND U8411 ( .A(n14113), .B(n14112), .Z(n14114) );
  AND U8412 ( .A(n14115), .B(n14114), .Z(n14332) );
  XOR U8413 ( .A(n14333), .B(n14332), .Z(n14202) );
  XOR U8414 ( .A(n14203), .B(n14202), .Z(n14205) );
  XOR U8415 ( .A(n14117), .B(n14116), .Z(n14156) );
  XOR U8416 ( .A(n14119), .B(n14118), .Z(n14152) );
  NANDN U8417 ( .A(n14121), .B(n14120), .Z(n14125) );
  NANDN U8418 ( .A(n14123), .B(n14122), .Z(n14124) );
  AND U8419 ( .A(n14125), .B(n14124), .Z(n14133) );
  NANDN U8420 ( .A(n14127), .B(n14126), .Z(n14131) );
  NAND U8421 ( .A(n14129), .B(n14128), .Z(n14130) );
  AND U8422 ( .A(n14131), .B(n14130), .Z(n14132) );
  NANDN U8423 ( .A(n14133), .B(n14132), .Z(n14137) );
  XNOR U8424 ( .A(n14133), .B(n14132), .Z(n14149) );
  XNOR U8425 ( .A(n14135), .B(n14134), .Z(n14148) );
  NAND U8426 ( .A(n14149), .B(n14148), .Z(n14136) );
  AND U8427 ( .A(n14137), .B(n14136), .Z(n14153) );
  NANDN U8428 ( .A(n14152), .B(n14153), .Z(n14155) );
  XOR U8429 ( .A(n14139), .B(n14138), .Z(n14147) );
  NANDN U8430 ( .A(n14141), .B(n14140), .Z(n14145) );
  NANDN U8431 ( .A(n14143), .B(n14142), .Z(n14144) );
  AND U8432 ( .A(n14145), .B(n14144), .Z(n14146) );
  NANDN U8433 ( .A(n14147), .B(n14146), .Z(n14151) );
  XOR U8434 ( .A(n14147), .B(n14146), .Z(n14178) );
  XOR U8435 ( .A(n14149), .B(n14148), .Z(n14179) );
  OR U8436 ( .A(n14178), .B(n14179), .Z(n14150) );
  AND U8437 ( .A(n14151), .B(n14150), .Z(n14159) );
  XNOR U8438 ( .A(n14153), .B(n14152), .Z(n14158) );
  NANDN U8439 ( .A(n14159), .B(n14158), .Z(n14154) );
  AND U8440 ( .A(n14155), .B(n14154), .Z(n14157) );
  NANDN U8441 ( .A(n14156), .B(n14157), .Z(n14201) );
  XNOR U8442 ( .A(n14157), .B(n14156), .Z(n15147) );
  XOR U8443 ( .A(n14159), .B(n14158), .Z(n14190) );
  NANDN U8444 ( .A(n14161), .B(n14160), .Z(n14165) );
  NANDN U8445 ( .A(n14163), .B(n14162), .Z(n14164) );
  AND U8446 ( .A(n14165), .B(n14164), .Z(n14181) );
  NAND U8447 ( .A(n14167), .B(n14166), .Z(n14171) );
  NAND U8448 ( .A(n14169), .B(n14168), .Z(n14170) );
  NAND U8449 ( .A(n14171), .B(n14170), .Z(n14194) );
  NAND U8450 ( .A(n14173), .B(n14172), .Z(n14177) );
  NAND U8451 ( .A(n14175), .B(n14174), .Z(n14176) );
  NAND U8452 ( .A(n14177), .B(n14176), .Z(n14192) );
  XOR U8453 ( .A(n14179), .B(n14178), .Z(n14193) );
  XNOR U8454 ( .A(n14192), .B(n14193), .Z(n14195) );
  XOR U8455 ( .A(n14194), .B(n14195), .Z(n14180) );
  NANDN U8456 ( .A(n14181), .B(n14180), .Z(n14189) );
  XNOR U8457 ( .A(n14181), .B(n14180), .Z(n15149) );
  NANDN U8458 ( .A(n14183), .B(n14182), .Z(n14187) );
  NAND U8459 ( .A(n14185), .B(n14184), .Z(n14186) );
  NAND U8460 ( .A(n14187), .B(n14186), .Z(n15148) );
  NAND U8461 ( .A(n15149), .B(n15148), .Z(n14188) );
  AND U8462 ( .A(n14189), .B(n14188), .Z(n14191) );
  NANDN U8463 ( .A(n14190), .B(n14191), .Z(n14199) );
  XNOR U8464 ( .A(n14191), .B(n14190), .Z(n15167) );
  NAND U8465 ( .A(n14193), .B(n14192), .Z(n14197) );
  NANDN U8466 ( .A(n14195), .B(n14194), .Z(n14196) );
  NAND U8467 ( .A(n14197), .B(n14196), .Z(n15166) );
  NAND U8468 ( .A(n15167), .B(n15166), .Z(n14198) );
  AND U8469 ( .A(n14199), .B(n14198), .Z(n15146) );
  NAND U8470 ( .A(n15147), .B(n15146), .Z(n14200) );
  AND U8471 ( .A(n14201), .B(n14200), .Z(n14204) );
  XOR U8472 ( .A(n14205), .B(n14204), .Z(N57) );
  NAND U8473 ( .A(n14207), .B(n14206), .Z(n14211) );
  NAND U8474 ( .A(n14209), .B(n14208), .Z(n14210) );
  NAND U8475 ( .A(n14211), .B(n14210), .Z(n14337) );
  NAND U8476 ( .A(n14213), .B(n14212), .Z(n14217) );
  NAND U8477 ( .A(n14215), .B(n14214), .Z(n14216) );
  AND U8478 ( .A(n14217), .B(n14216), .Z(n14469) );
  NANDN U8479 ( .A(n14219), .B(n14218), .Z(n14223) );
  NANDN U8480 ( .A(n14221), .B(n14220), .Z(n14222) );
  NAND U8481 ( .A(n14223), .B(n14222), .Z(n14450) );
  NAND U8482 ( .A(x[21]), .B(y[8]), .Z(n15057) );
  NANDN U8483 ( .A(n15057), .B(n14224), .Z(n14228) );
  NAND U8484 ( .A(n14226), .B(n14225), .Z(n14227) );
  AND U8485 ( .A(n14228), .B(n14227), .Z(n14419) );
  AND U8486 ( .A(y[6]), .B(x[19]), .Z(n14395) );
  AND U8487 ( .A(y[5]), .B(x[20]), .Z(n14394) );
  NAND U8488 ( .A(y[4]), .B(x[21]), .Z(n14393) );
  XOR U8489 ( .A(n14394), .B(n14393), .Z(n14396) );
  XOR U8490 ( .A(n14395), .B(n14396), .Z(n14418) );
  AND U8491 ( .A(x[22]), .B(y[3]), .Z(n14376) );
  AND U8492 ( .A(x[17]), .B(y[8]), .Z(n14375) );
  NAND U8493 ( .A(x[5]), .B(y[20]), .Z(n14374) );
  XOR U8494 ( .A(n14375), .B(n14374), .Z(n14377) );
  XNOR U8495 ( .A(n14376), .B(n14377), .Z(n14417) );
  XOR U8496 ( .A(n14418), .B(n14417), .Z(n14420) );
  XNOR U8497 ( .A(n14419), .B(n14420), .Z(n14449) );
  XOR U8498 ( .A(n14450), .B(n14449), .Z(n14452) );
  NAND U8499 ( .A(n14582), .B(n14229), .Z(n14233) );
  AND U8500 ( .A(n14231), .B(n14230), .Z(n14232) );
  ANDN U8501 ( .B(n14233), .A(n14232), .Z(n14413) );
  AND U8502 ( .A(x[23]), .B(y[2]), .Z(n14382) );
  AND U8503 ( .A(y[9]), .B(x[16]), .Z(n14381) );
  NAND U8504 ( .A(x[4]), .B(y[21]), .Z(n14380) );
  XOR U8505 ( .A(n14381), .B(n14380), .Z(n14383) );
  XOR U8506 ( .A(n14382), .B(n14383), .Z(n14412) );
  AND U8507 ( .A(y[10]), .B(x[15]), .Z(n14401) );
  AND U8508 ( .A(x[6]), .B(y[19]), .Z(n14400) );
  NAND U8509 ( .A(x[18]), .B(y[7]), .Z(n14399) );
  XOR U8510 ( .A(n14400), .B(n14399), .Z(n14402) );
  XNOR U8511 ( .A(n14401), .B(n14402), .Z(n14411) );
  XOR U8512 ( .A(n14412), .B(n14411), .Z(n14414) );
  XNOR U8513 ( .A(n14413), .B(n14414), .Z(n14451) );
  XOR U8514 ( .A(n14452), .B(n14451), .Z(n14350) );
  NANDN U8515 ( .A(n14239), .B(n14238), .Z(n14243) );
  NANDN U8516 ( .A(n14241), .B(n14240), .Z(n14242) );
  AND U8517 ( .A(n14243), .B(n14242), .Z(n14348) );
  XOR U8518 ( .A(n14349), .B(n14348), .Z(n14351) );
  XNOR U8519 ( .A(n14350), .B(n14351), .Z(n14345) );
  NAND U8520 ( .A(n14245), .B(n14244), .Z(n14249) );
  NAND U8521 ( .A(n14247), .B(n14246), .Z(n14248) );
  NAND U8522 ( .A(n14249), .B(n14248), .Z(n14343) );
  NAND U8523 ( .A(n14251), .B(n14250), .Z(n14255) );
  NAND U8524 ( .A(n14253), .B(n14252), .Z(n14254) );
  AND U8525 ( .A(n14255), .B(n14254), .Z(n14342) );
  XOR U8526 ( .A(n14343), .B(n14342), .Z(n14344) );
  XOR U8527 ( .A(n14345), .B(n14344), .Z(n14468) );
  XOR U8528 ( .A(n14469), .B(n14468), .Z(n14471) );
  NAND U8529 ( .A(n14257), .B(n14256), .Z(n14261) );
  NAND U8530 ( .A(n14259), .B(n14258), .Z(n14260) );
  AND U8531 ( .A(n14261), .B(n14260), .Z(n14470) );
  XOR U8532 ( .A(n14471), .B(n14470), .Z(n14477) );
  NAND U8533 ( .A(n14263), .B(n14262), .Z(n14267) );
  NAND U8534 ( .A(n14265), .B(n14264), .Z(n14266) );
  AND U8535 ( .A(n14267), .B(n14266), .Z(n14456) );
  NANDN U8536 ( .A(n14437), .B(n14268), .Z(n14272) );
  NANDN U8537 ( .A(n14270), .B(n14269), .Z(n14271) );
  AND U8538 ( .A(n14272), .B(n14271), .Z(n14444) );
  NAND U8539 ( .A(y[16]), .B(x[14]), .Z(n15390) );
  NANDN U8540 ( .A(n15390), .B(n14273), .Z(n14277) );
  NANDN U8541 ( .A(n14275), .B(n14274), .Z(n14276) );
  AND U8542 ( .A(n14277), .B(n14276), .Z(n14371) );
  AND U8543 ( .A(x[11]), .B(y[14]), .Z(n14389) );
  AND U8544 ( .A(x[12]), .B(y[13]), .Z(n14388) );
  NAND U8545 ( .A(x[7]), .B(y[18]), .Z(n14387) );
  XOR U8546 ( .A(n14388), .B(n14387), .Z(n14390) );
  XOR U8547 ( .A(n14389), .B(n14390), .Z(n14369) );
  NAND U8548 ( .A(x[13]), .B(y[12]), .Z(n14364) );
  NAND U8549 ( .A(y[24]), .B(x[1]), .Z(n14363) );
  NAND U8550 ( .A(y[1]), .B(x[24]), .Z(n14386) );
  XOR U8551 ( .A(o[25]), .B(n14386), .Z(n14362) );
  XNOR U8552 ( .A(n14363), .B(n14362), .Z(n14365) );
  XOR U8553 ( .A(n14364), .B(n14365), .Z(n14368) );
  XNOR U8554 ( .A(n14369), .B(n14368), .Z(n14370) );
  XNOR U8555 ( .A(n14371), .B(n14370), .Z(n14443) );
  XNOR U8556 ( .A(n14444), .B(n14443), .Z(n14445) );
  XNOR U8557 ( .A(n14424), .B(n14423), .Z(n14425) );
  NANDN U8558 ( .A(n14287), .B(n14286), .Z(n14291) );
  NAND U8559 ( .A(n14289), .B(n14288), .Z(n14290) );
  AND U8560 ( .A(n14291), .B(n14290), .Z(n14432) );
  AND U8561 ( .A(x[8]), .B(y[17]), .Z(n14440) );
  XOR U8562 ( .A(n14438), .B(n14292), .Z(n14439) );
  XOR U8563 ( .A(n14440), .B(n14439), .Z(n14429) );
  AND U8564 ( .A(x[25]), .B(y[0]), .Z(n14433) );
  NAND U8565 ( .A(y[25]), .B(x[0]), .Z(n14434) );
  XNOR U8566 ( .A(n14433), .B(n14434), .Z(n14436) );
  ANDN U8567 ( .B(o[24]), .A(n14293), .Z(n14435) );
  XOR U8568 ( .A(n14436), .B(n14435), .Z(n14430) );
  XOR U8569 ( .A(n14429), .B(n14430), .Z(n14431) );
  XOR U8570 ( .A(n14432), .B(n14431), .Z(n14426) );
  XOR U8571 ( .A(n14425), .B(n14426), .Z(n14446) );
  XOR U8572 ( .A(n14445), .B(n14446), .Z(n14463) );
  NAND U8573 ( .A(n14295), .B(n14294), .Z(n14299) );
  NANDN U8574 ( .A(n14297), .B(n14296), .Z(n14298) );
  NAND U8575 ( .A(n14299), .B(n14298), .Z(n14461) );
  AND U8576 ( .A(y[22]), .B(x[3]), .Z(n14356) );
  NAND U8577 ( .A(y[11]), .B(x[14]), .Z(n14357) );
  XNOR U8578 ( .A(n14356), .B(n14357), .Z(n14359) );
  AND U8579 ( .A(x[2]), .B(y[23]), .Z(n14358) );
  XOR U8580 ( .A(n14359), .B(n14358), .Z(n14406) );
  NANDN U8581 ( .A(n14301), .B(n14300), .Z(n14305) );
  NAND U8582 ( .A(n14303), .B(n14302), .Z(n14304) );
  AND U8583 ( .A(n14305), .B(n14304), .Z(n14405) );
  XNOR U8584 ( .A(n14406), .B(n14405), .Z(n14407) );
  NANDN U8585 ( .A(n14307), .B(n14306), .Z(n14311) );
  NANDN U8586 ( .A(n14309), .B(n14308), .Z(n14310) );
  NAND U8587 ( .A(n14311), .B(n14310), .Z(n14408) );
  XNOR U8588 ( .A(n14407), .B(n14408), .Z(n14462) );
  XOR U8589 ( .A(n14461), .B(n14462), .Z(n14464) );
  XOR U8590 ( .A(n14463), .B(n14464), .Z(n14455) );
  XOR U8591 ( .A(n14456), .B(n14455), .Z(n14458) );
  NAND U8592 ( .A(n14313), .B(n14312), .Z(n14317) );
  NAND U8593 ( .A(n14315), .B(n14314), .Z(n14316) );
  AND U8594 ( .A(n14317), .B(n14316), .Z(n14457) );
  XNOR U8595 ( .A(n14458), .B(n14457), .Z(n14475) );
  NAND U8596 ( .A(n14319), .B(n14318), .Z(n14323) );
  NAND U8597 ( .A(n14321), .B(n14320), .Z(n14322) );
  AND U8598 ( .A(n14323), .B(n14322), .Z(n14474) );
  XOR U8599 ( .A(n14475), .B(n14474), .Z(n14476) );
  XOR U8600 ( .A(n14477), .B(n14476), .Z(n14336) );
  XOR U8601 ( .A(n14337), .B(n14336), .Z(n14339) );
  NAND U8602 ( .A(n14325), .B(n14324), .Z(n14329) );
  NAND U8603 ( .A(n14327), .B(n14326), .Z(n14328) );
  AND U8604 ( .A(n14329), .B(n14328), .Z(n14338) );
  XOR U8605 ( .A(n14339), .B(n14338), .Z(n14480) );
  XOR U8606 ( .A(n14481), .B(n14480), .Z(n14483) );
  NANDN U8607 ( .A(n14331), .B(n14330), .Z(n14335) );
  NAND U8608 ( .A(n14333), .B(n14332), .Z(n14334) );
  AND U8609 ( .A(n14335), .B(n14334), .Z(n14482) );
  XNOR U8610 ( .A(n14483), .B(n14482), .Z(N58) );
  NAND U8611 ( .A(n14337), .B(n14336), .Z(n14341) );
  NAND U8612 ( .A(n14339), .B(n14338), .Z(n14340) );
  NAND U8613 ( .A(n14341), .B(n14340), .Z(n14769) );
  NAND U8614 ( .A(n14343), .B(n14342), .Z(n14347) );
  NAND U8615 ( .A(n14345), .B(n14344), .Z(n14346) );
  AND U8616 ( .A(n14347), .B(n14346), .Z(n14773) );
  NANDN U8617 ( .A(n14349), .B(n14348), .Z(n14353) );
  OR U8618 ( .A(n14351), .B(n14350), .Z(n14352) );
  AND U8619 ( .A(n14353), .B(n14352), .Z(n14746) );
  AND U8620 ( .A(x[12]), .B(y[14]), .Z(n14556) );
  AND U8621 ( .A(y[21]), .B(x[5]), .Z(n14487) );
  XOR U8622 ( .A(n14556), .B(n14487), .Z(n14488) );
  NAND U8623 ( .A(x[10]), .B(y[16]), .Z(n14489) );
  XNOR U8624 ( .A(n14488), .B(n14489), .Z(n14680) );
  NAND U8625 ( .A(y[20]), .B(x[6]), .Z(n14354) );
  XNOR U8626 ( .A(n14355), .B(n14354), .Z(n14584) );
  AND U8627 ( .A(y[17]), .B(x[9]), .Z(n14583) );
  XOR U8628 ( .A(n14584), .B(n14583), .Z(n14678) );
  AND U8629 ( .A(y[19]), .B(x[7]), .Z(n14677) );
  XOR U8630 ( .A(n14678), .B(n14677), .Z(n14679) );
  XOR U8631 ( .A(n14680), .B(n14679), .Z(n14706) );
  NANDN U8632 ( .A(n14357), .B(n14356), .Z(n14361) );
  NAND U8633 ( .A(n14359), .B(n14358), .Z(n14360) );
  NAND U8634 ( .A(n14361), .B(n14360), .Z(n14703) );
  NAND U8635 ( .A(n14363), .B(n14362), .Z(n14367) );
  NANDN U8636 ( .A(n14365), .B(n14364), .Z(n14366) );
  AND U8637 ( .A(n14367), .B(n14366), .Z(n14704) );
  XOR U8638 ( .A(n14703), .B(n14704), .Z(n14705) );
  XOR U8639 ( .A(n14706), .B(n14705), .Z(n14730) );
  NANDN U8640 ( .A(n14369), .B(n14368), .Z(n14373) );
  NANDN U8641 ( .A(n14371), .B(n14370), .Z(n14372) );
  AND U8642 ( .A(n14373), .B(n14372), .Z(n14729) );
  XNOR U8643 ( .A(n14730), .B(n14729), .Z(n14732) );
  NANDN U8644 ( .A(n14375), .B(n14374), .Z(n14379) );
  OR U8645 ( .A(n14377), .B(n14376), .Z(n14378) );
  NAND U8646 ( .A(n14379), .B(n14378), .Z(n14542) );
  NANDN U8647 ( .A(n14381), .B(n14380), .Z(n14385) );
  OR U8648 ( .A(n14383), .B(n14382), .Z(n14384) );
  NAND U8649 ( .A(n14385), .B(n14384), .Z(n14541) );
  NAND U8650 ( .A(y[26]), .B(x[0]), .Z(n14494) );
  NAND U8651 ( .A(x[26]), .B(y[0]), .Z(n14492) );
  AND U8652 ( .A(y[1]), .B(x[25]), .Z(n14569) );
  XNOR U8653 ( .A(o[26]), .B(n14569), .Z(n14493) );
  XNOR U8654 ( .A(n14492), .B(n14493), .Z(n14495) );
  XOR U8655 ( .A(n14494), .B(n14495), .Z(n14499) );
  ANDN U8656 ( .B(o[25]), .A(n14386), .Z(n14628) );
  AND U8657 ( .A(y[12]), .B(x[14]), .Z(n14627) );
  XOR U8658 ( .A(n14628), .B(n14627), .Z(n14630) );
  AND U8659 ( .A(y[25]), .B(x[1]), .Z(n14629) );
  XOR U8660 ( .A(n14630), .B(n14629), .Z(n14498) );
  XOR U8661 ( .A(n14499), .B(n14498), .Z(n14501) );
  NANDN U8662 ( .A(n14388), .B(n14387), .Z(n14392) );
  OR U8663 ( .A(n14390), .B(n14389), .Z(n14391) );
  AND U8664 ( .A(n14392), .B(n14391), .Z(n14500) );
  XNOR U8665 ( .A(n14501), .B(n14500), .Z(n14540) );
  XOR U8666 ( .A(n14541), .B(n14540), .Z(n14543) );
  XOR U8667 ( .A(n14542), .B(n14543), .Z(n14723) );
  NAND U8668 ( .A(y[6]), .B(x[20]), .Z(n14623) );
  NAND U8669 ( .A(y[5]), .B(x[21]), .Z(n14621) );
  XOR U8670 ( .A(n14621), .B(n14622), .Z(n14624) );
  XNOR U8671 ( .A(n14623), .B(n14624), .Z(n14698) );
  AND U8672 ( .A(x[23]), .B(y[3]), .Z(n14521) );
  XOR U8673 ( .A(n14521), .B(n14520), .Z(n14523) );
  AND U8674 ( .A(x[22]), .B(y[4]), .Z(n14522) );
  XOR U8675 ( .A(n14523), .B(n14522), .Z(n14697) );
  XOR U8676 ( .A(n14698), .B(n14697), .Z(n14700) );
  NANDN U8677 ( .A(n14394), .B(n14393), .Z(n14398) );
  OR U8678 ( .A(n14396), .B(n14395), .Z(n14397) );
  AND U8679 ( .A(n14398), .B(n14397), .Z(n14699) );
  XOR U8680 ( .A(n14700), .B(n14699), .Z(n14722) );
  AND U8681 ( .A(x[11]), .B(y[15]), .Z(n14614) );
  AND U8682 ( .A(x[3]), .B(y[23]), .Z(n14613) );
  XOR U8683 ( .A(n14614), .B(n14613), .Z(n14616) );
  AND U8684 ( .A(x[19]), .B(y[7]), .Z(n14615) );
  XOR U8685 ( .A(n14616), .B(n14615), .Z(n14533) );
  AND U8686 ( .A(x[4]), .B(y[22]), .Z(n14514) );
  XOR U8687 ( .A(n14515), .B(n14514), .Z(n14517) );
  AND U8688 ( .A(x[18]), .B(y[8]), .Z(n14516) );
  XOR U8689 ( .A(n14517), .B(n14516), .Z(n14532) );
  XOR U8690 ( .A(n14533), .B(n14532), .Z(n14535) );
  NANDN U8691 ( .A(n14400), .B(n14399), .Z(n14404) );
  OR U8692 ( .A(n14402), .B(n14401), .Z(n14403) );
  AND U8693 ( .A(n14404), .B(n14403), .Z(n14534) );
  XNOR U8694 ( .A(n14535), .B(n14534), .Z(n14721) );
  XOR U8695 ( .A(n14722), .B(n14721), .Z(n14724) );
  XNOR U8696 ( .A(n14723), .B(n14724), .Z(n14731) );
  XOR U8697 ( .A(n14732), .B(n14731), .Z(n14744) );
  NANDN U8698 ( .A(n14406), .B(n14405), .Z(n14410) );
  NANDN U8699 ( .A(n14408), .B(n14407), .Z(n14409) );
  AND U8700 ( .A(n14410), .B(n14409), .Z(n14673) );
  NANDN U8701 ( .A(n14412), .B(n14411), .Z(n14416) );
  OR U8702 ( .A(n14414), .B(n14413), .Z(n14415) );
  AND U8703 ( .A(n14416), .B(n14415), .Z(n14672) );
  NANDN U8704 ( .A(n14418), .B(n14417), .Z(n14422) );
  OR U8705 ( .A(n14420), .B(n14419), .Z(n14421) );
  NAND U8706 ( .A(n14422), .B(n14421), .Z(n14671) );
  XOR U8707 ( .A(n14672), .B(n14671), .Z(n14674) );
  XNOR U8708 ( .A(n14673), .B(n14674), .Z(n14743) );
  XNOR U8709 ( .A(n14744), .B(n14743), .Z(n14745) );
  XNOR U8710 ( .A(n14746), .B(n14745), .Z(n14771) );
  NANDN U8711 ( .A(n14424), .B(n14423), .Z(n14428) );
  NANDN U8712 ( .A(n14426), .B(n14425), .Z(n14427) );
  AND U8713 ( .A(n14428), .B(n14427), .Z(n14690) );
  NAND U8714 ( .A(y[2]), .B(x[24]), .Z(n14528) );
  NAND U8715 ( .A(y[24]), .B(x[2]), .Z(n14527) );
  NAND U8716 ( .A(y[11]), .B(x[15]), .Z(n14526) );
  XNOR U8717 ( .A(n14527), .B(n14526), .Z(n14529) );
  NANDN U8718 ( .A(n14438), .B(n14437), .Z(n14442) );
  NANDN U8719 ( .A(n14440), .B(n14439), .Z(n14441) );
  AND U8720 ( .A(n14442), .B(n14441), .Z(n14506) );
  XOR U8721 ( .A(n14507), .B(n14506), .Z(n14508) );
  XNOR U8722 ( .A(n14509), .B(n14508), .Z(n14687) );
  XNOR U8723 ( .A(n14688), .B(n14687), .Z(n14689) );
  XNOR U8724 ( .A(n14690), .B(n14689), .Z(n14755) );
  NANDN U8725 ( .A(n14444), .B(n14443), .Z(n14448) );
  NANDN U8726 ( .A(n14446), .B(n14445), .Z(n14447) );
  AND U8727 ( .A(n14448), .B(n14447), .Z(n14754) );
  NAND U8728 ( .A(n14450), .B(n14449), .Z(n14454) );
  NAND U8729 ( .A(n14452), .B(n14451), .Z(n14453) );
  AND U8730 ( .A(n14454), .B(n14453), .Z(n14753) );
  XOR U8731 ( .A(n14754), .B(n14753), .Z(n14756) );
  XNOR U8732 ( .A(n14755), .B(n14756), .Z(n14770) );
  XOR U8733 ( .A(n14771), .B(n14770), .Z(n14772) );
  XOR U8734 ( .A(n14773), .B(n14772), .Z(n14778) );
  NAND U8735 ( .A(n14456), .B(n14455), .Z(n14460) );
  NAND U8736 ( .A(n14458), .B(n14457), .Z(n14459) );
  NAND U8737 ( .A(n14460), .B(n14459), .Z(n14776) );
  NAND U8738 ( .A(n14462), .B(n14461), .Z(n14466) );
  NAND U8739 ( .A(n14464), .B(n14463), .Z(n14465) );
  AND U8740 ( .A(n14466), .B(n14465), .Z(n14777) );
  XOR U8741 ( .A(n14776), .B(n14777), .Z(n14467) );
  XOR U8742 ( .A(n14778), .B(n14467), .Z(n14785) );
  NAND U8743 ( .A(n14469), .B(n14468), .Z(n14473) );
  NAND U8744 ( .A(n14471), .B(n14470), .Z(n14472) );
  NAND U8745 ( .A(n14473), .B(n14472), .Z(n14783) );
  NAND U8746 ( .A(n14475), .B(n14474), .Z(n14479) );
  NANDN U8747 ( .A(n14477), .B(n14476), .Z(n14478) );
  AND U8748 ( .A(n14479), .B(n14478), .Z(n14784) );
  XOR U8749 ( .A(n14783), .B(n14784), .Z(n14786) );
  XOR U8750 ( .A(n14785), .B(n14786), .Z(n14768) );
  XNOR U8751 ( .A(n14768), .B(n14767), .Z(n14484) );
  XNOR U8752 ( .A(n14769), .B(n14484), .Z(N59) );
  AND U8753 ( .A(x[15]), .B(y[12]), .Z(n14562) );
  AND U8754 ( .A(y[25]), .B(x[2]), .Z(n14561) );
  XOR U8755 ( .A(n14562), .B(n14561), .Z(n14564) );
  AND U8756 ( .A(y[24]), .B(x[3]), .Z(n14563) );
  XOR U8757 ( .A(n14564), .B(n14563), .Z(n14602) );
  AND U8758 ( .A(x[19]), .B(y[8]), .Z(n14645) );
  AND U8759 ( .A(y[2]), .B(x[25]), .Z(n14644) );
  XOR U8760 ( .A(n14645), .B(n14644), .Z(n14647) );
  AND U8761 ( .A(x[6]), .B(y[21]), .Z(n14646) );
  XOR U8762 ( .A(n14647), .B(n14646), .Z(n14601) );
  XOR U8763 ( .A(n14602), .B(n14601), .Z(n14604) );
  AND U8764 ( .A(y[11]), .B(x[16]), .Z(n14550) );
  XOR U8765 ( .A(n14550), .B(n14549), .Z(n14552) );
  XOR U8766 ( .A(n14552), .B(n14551), .Z(n14558) );
  AND U8767 ( .A(y[14]), .B(x[13]), .Z(n14486) );
  NAND U8768 ( .A(y[15]), .B(x[12]), .Z(n14485) );
  XNOR U8769 ( .A(n14486), .B(n14485), .Z(n14557) );
  XOR U8770 ( .A(n14558), .B(n14557), .Z(n14603) );
  XOR U8771 ( .A(n14604), .B(n14603), .Z(n14597) );
  AND U8772 ( .A(n14556), .B(n14487), .Z(n14491) );
  NANDN U8773 ( .A(n14489), .B(n14488), .Z(n14490) );
  NANDN U8774 ( .A(n14491), .B(n14490), .Z(n14595) );
  NAND U8775 ( .A(n14493), .B(n14492), .Z(n14497) );
  NANDN U8776 ( .A(n14495), .B(n14494), .Z(n14496) );
  AND U8777 ( .A(n14497), .B(n14496), .Z(n14596) );
  XNOR U8778 ( .A(n14595), .B(n14596), .Z(n14598) );
  NAND U8779 ( .A(n14499), .B(n14498), .Z(n14503) );
  NAND U8780 ( .A(n14501), .B(n14500), .Z(n14502) );
  NAND U8781 ( .A(n14503), .B(n14502), .Z(n14505) );
  NAND U8782 ( .A(n14504), .B(n14505), .Z(n14513) );
  XOR U8783 ( .A(n14505), .B(n14504), .Z(n14727) );
  NAND U8784 ( .A(n14507), .B(n14506), .Z(n14511) );
  NANDN U8785 ( .A(n14509), .B(n14508), .Z(n14510) );
  NAND U8786 ( .A(n14511), .B(n14510), .Z(n14728) );
  NAND U8787 ( .A(n14727), .B(n14728), .Z(n14512) );
  NAND U8788 ( .A(n14513), .B(n14512), .Z(n14940) );
  AND U8789 ( .A(n14515), .B(n14514), .Z(n14519) );
  NAND U8790 ( .A(n14517), .B(n14516), .Z(n14518) );
  NANDN U8791 ( .A(n14519), .B(n14518), .Z(n14574) );
  AND U8792 ( .A(x[9]), .B(y[18]), .Z(n14651) );
  AND U8793 ( .A(y[6]), .B(x[21]), .Z(n14650) );
  XOR U8794 ( .A(n14651), .B(n14650), .Z(n14653) );
  AND U8795 ( .A(x[18]), .B(y[9]), .Z(n14652) );
  XOR U8796 ( .A(n14653), .B(n14652), .Z(n14573) );
  AND U8797 ( .A(y[1]), .B(x[26]), .Z(n14656) );
  XOR U8798 ( .A(o[27]), .B(n14656), .Z(n14662) );
  AND U8799 ( .A(x[27]), .B(y[0]), .Z(n14660) );
  AND U8800 ( .A(y[27]), .B(x[0]), .Z(n14659) );
  XOR U8801 ( .A(n14660), .B(n14659), .Z(n14661) );
  XOR U8802 ( .A(n14662), .B(n14661), .Z(n14572) );
  XOR U8803 ( .A(n14573), .B(n14572), .Z(n14575) );
  XOR U8804 ( .A(n14574), .B(n14575), .Z(n14591) );
  NAND U8805 ( .A(n14521), .B(n14520), .Z(n14525) );
  NAND U8806 ( .A(n14523), .B(n14522), .Z(n14524) );
  NAND U8807 ( .A(n14525), .B(n14524), .Z(n14589) );
  NAND U8808 ( .A(n14527), .B(n14526), .Z(n14531) );
  NANDN U8809 ( .A(n14529), .B(n14528), .Z(n14530) );
  AND U8810 ( .A(n14531), .B(n14530), .Z(n14590) );
  XNOR U8811 ( .A(n14589), .B(n14590), .Z(n14592) );
  NAND U8812 ( .A(n14533), .B(n14532), .Z(n14537) );
  NAND U8813 ( .A(n14535), .B(n14534), .Z(n14536) );
  NAND U8814 ( .A(n14537), .B(n14536), .Z(n14539) );
  NAND U8815 ( .A(n14538), .B(n14539), .Z(n14547) );
  XOR U8816 ( .A(n14539), .B(n14538), .Z(n14712) );
  NAND U8817 ( .A(n14541), .B(n14540), .Z(n14545) );
  NAND U8818 ( .A(n14543), .B(n14542), .Z(n14544) );
  AND U8819 ( .A(n14545), .B(n14544), .Z(n14711) );
  NAND U8820 ( .A(n14712), .B(n14711), .Z(n14546) );
  NAND U8821 ( .A(n14547), .B(n14546), .Z(n14939) );
  XOR U8822 ( .A(n14940), .B(n14939), .Z(n14942) );
  AND U8823 ( .A(y[24]), .B(x[4]), .Z(n14848) );
  AND U8824 ( .A(y[6]), .B(x[22]), .Z(n14846) );
  AND U8825 ( .A(y[11]), .B(x[17]), .Z(n14845) );
  XOR U8826 ( .A(n14846), .B(n14845), .Z(n14847) );
  XOR U8827 ( .A(n14848), .B(n14847), .Z(n14875) );
  AND U8828 ( .A(x[6]), .B(y[22]), .Z(n15080) );
  AND U8829 ( .A(x[19]), .B(y[9]), .Z(n14906) );
  XOR U8830 ( .A(n15080), .B(n14906), .Z(n14907) );
  XOR U8831 ( .A(n15101), .B(n14907), .Z(n14874) );
  XOR U8832 ( .A(n14875), .B(n14874), .Z(n14877) );
  NAND U8833 ( .A(y[19]), .B(x[8]), .Z(n14857) );
  NAND U8834 ( .A(x[23]), .B(y[4]), .Z(n14548) );
  XOR U8835 ( .A(n14857), .B(n14548), .Z(n14607) );
  NAND U8836 ( .A(x[22]), .B(y[5]), .Z(n14608) );
  XOR U8837 ( .A(n14877), .B(n14876), .Z(n14815) );
  NAND U8838 ( .A(n14550), .B(n14549), .Z(n14554) );
  NAND U8839 ( .A(n14552), .B(n14551), .Z(n14553) );
  NAND U8840 ( .A(n14554), .B(n14553), .Z(n14929) );
  NAND U8841 ( .A(y[17]), .B(x[11]), .Z(n14882) );
  NAND U8842 ( .A(y[16]), .B(x[12]), .Z(n14881) );
  NAND U8843 ( .A(y[21]), .B(x[7]), .Z(n14880) );
  XOR U8844 ( .A(n14881), .B(n14880), .Z(n14883) );
  XOR U8845 ( .A(n14882), .B(n14883), .Z(n14928) );
  NAND U8846 ( .A(x[27]), .B(y[1]), .Z(n14555) );
  XNOR U8847 ( .A(o[28]), .B(n14555), .Z(n14915) );
  AND U8848 ( .A(y[2]), .B(x[26]), .Z(n14914) );
  XOR U8849 ( .A(n14915), .B(n14914), .Z(n14917) );
  AND U8850 ( .A(y[13]), .B(x[15]), .Z(n14916) );
  XOR U8851 ( .A(n14917), .B(n14916), .Z(n14927) );
  XOR U8852 ( .A(n14929), .B(n14930), .Z(n14816) );
  XNOR U8853 ( .A(n14815), .B(n14816), .Z(n14817) );
  NAND U8854 ( .A(n14923), .B(n14556), .Z(n14560) );
  NAND U8855 ( .A(n14558), .B(n14557), .Z(n14559) );
  NAND U8856 ( .A(n14560), .B(n14559), .Z(n14870) );
  NAND U8857 ( .A(n14562), .B(n14561), .Z(n14566) );
  NAND U8858 ( .A(n14564), .B(n14563), .Z(n14565) );
  NAND U8859 ( .A(n14566), .B(n14565), .Z(n14869) );
  AND U8860 ( .A(y[13]), .B(x[14]), .Z(n14568) );
  AND U8861 ( .A(y[26]), .B(x[1]), .Z(n14567) );
  NAND U8862 ( .A(n14568), .B(n14567), .Z(n14571) );
  XOR U8863 ( .A(n14568), .B(n14567), .Z(n14579) );
  AND U8864 ( .A(n14569), .B(o[26]), .Z(n14578) );
  NAND U8865 ( .A(n14579), .B(n14578), .Z(n14570) );
  NAND U8866 ( .A(n14571), .B(n14570), .Z(n14868) );
  XNOR U8867 ( .A(n14869), .B(n14868), .Z(n14871) );
  XNOR U8868 ( .A(n14817), .B(n14818), .Z(n14936) );
  NAND U8869 ( .A(n14573), .B(n14572), .Z(n14577) );
  NAND U8870 ( .A(n14575), .B(n14574), .Z(n14576) );
  AND U8871 ( .A(n14577), .B(n14576), .Z(n14840) );
  AND U8872 ( .A(x[4]), .B(y[23]), .Z(n14666) );
  AND U8873 ( .A(x[17]), .B(y[10]), .Z(n14665) );
  XOR U8874 ( .A(n14666), .B(n14665), .Z(n14668) );
  AND U8875 ( .A(y[22]), .B(x[5]), .Z(n14667) );
  XOR U8876 ( .A(n14668), .B(n14667), .Z(n14581) );
  XOR U8877 ( .A(n14579), .B(n14578), .Z(n14580) );
  NAND U8878 ( .A(n14581), .B(n14580), .Z(n14588) );
  XOR U8879 ( .A(n14581), .B(n14580), .Z(n14635) );
  AND U8880 ( .A(y[20]), .B(x[8]), .Z(n14658) );
  NAND U8881 ( .A(n14658), .B(n14582), .Z(n14586) );
  NAND U8882 ( .A(n14584), .B(n14583), .Z(n14585) );
  NAND U8883 ( .A(n14586), .B(n14585), .Z(n14636) );
  NAND U8884 ( .A(n14635), .B(n14636), .Z(n14587) );
  AND U8885 ( .A(n14588), .B(n14587), .Z(n14839) );
  XOR U8886 ( .A(n14840), .B(n14839), .Z(n14842) );
  NAND U8887 ( .A(n14590), .B(n14589), .Z(n14594) );
  NANDN U8888 ( .A(n14592), .B(n14591), .Z(n14593) );
  AND U8889 ( .A(n14594), .B(n14593), .Z(n14841) );
  XOR U8890 ( .A(n14842), .B(n14841), .Z(n14934) );
  NAND U8891 ( .A(n14596), .B(n14595), .Z(n14600) );
  NANDN U8892 ( .A(n14598), .B(n14597), .Z(n14599) );
  AND U8893 ( .A(n14600), .B(n14599), .Z(n14933) );
  XOR U8894 ( .A(n14934), .B(n14933), .Z(n14935) );
  NAND U8895 ( .A(n14602), .B(n14601), .Z(n14606) );
  NAND U8896 ( .A(n14604), .B(n14603), .Z(n14605) );
  AND U8897 ( .A(n14606), .B(n14605), .Z(n14810) );
  XNOR U8898 ( .A(n14608), .B(n14607), .Z(n14612) );
  AND U8899 ( .A(x[24]), .B(y[3]), .Z(n14610) );
  NAND U8900 ( .A(x[20]), .B(y[7]), .Z(n14609) );
  XNOR U8901 ( .A(n14610), .B(n14609), .Z(n14641) );
  AND U8902 ( .A(x[7]), .B(y[20]), .Z(n14640) );
  XOR U8903 ( .A(n14641), .B(n14640), .Z(n14611) );
  NAND U8904 ( .A(n14612), .B(n14611), .Z(n14620) );
  XNOR U8905 ( .A(n14612), .B(n14611), .Z(n14683) );
  NAND U8906 ( .A(n14614), .B(n14613), .Z(n14618) );
  NAND U8907 ( .A(n14616), .B(n14615), .Z(n14617) );
  NAND U8908 ( .A(n14618), .B(n14617), .Z(n14684) );
  NANDN U8909 ( .A(n14683), .B(n14684), .Z(n14619) );
  AND U8910 ( .A(n14620), .B(n14619), .Z(n14809) );
  XOR U8911 ( .A(n14810), .B(n14809), .Z(n14812) );
  NAND U8912 ( .A(n14622), .B(n14621), .Z(n14626) );
  NAND U8913 ( .A(n14624), .B(n14623), .Z(n14625) );
  AND U8914 ( .A(n14626), .B(n14625), .Z(n14633) );
  NAND U8915 ( .A(n14628), .B(n14627), .Z(n14632) );
  NAND U8916 ( .A(n14630), .B(n14629), .Z(n14631) );
  NAND U8917 ( .A(n14632), .B(n14631), .Z(n14634) );
  NAND U8918 ( .A(n14633), .B(n14634), .Z(n14638) );
  XOR U8919 ( .A(n14634), .B(n14633), .Z(n14686) );
  XOR U8920 ( .A(n14636), .B(n14635), .Z(n14685) );
  NAND U8921 ( .A(n14686), .B(n14685), .Z(n14637) );
  AND U8922 ( .A(n14638), .B(n14637), .Z(n14811) );
  XOR U8923 ( .A(n14812), .B(n14811), .Z(n14946) );
  AND U8924 ( .A(y[7]), .B(x[24]), .Z(n15370) );
  NAND U8925 ( .A(n15370), .B(n14639), .Z(n14643) );
  NAND U8926 ( .A(n14641), .B(n14640), .Z(n14642) );
  NAND U8927 ( .A(n14643), .B(n14642), .Z(n14835) );
  AND U8928 ( .A(x[25]), .B(y[3]), .Z(n15069) );
  XOR U8929 ( .A(n15069), .B(n14892), .Z(n14894) );
  AND U8930 ( .A(x[1]), .B(y[27]), .Z(n14893) );
  XOR U8931 ( .A(n14894), .B(n14893), .Z(n14834) );
  AND U8932 ( .A(x[16]), .B(y[12]), .Z(n14887) );
  AND U8933 ( .A(y[4]), .B(x[24]), .Z(n14886) );
  XOR U8934 ( .A(n14887), .B(n14886), .Z(n14889) );
  AND U8935 ( .A(x[2]), .B(y[26]), .Z(n14888) );
  XOR U8936 ( .A(n14889), .B(n14888), .Z(n14833) );
  XOR U8937 ( .A(n14834), .B(n14833), .Z(n14836) );
  XNOR U8938 ( .A(n14835), .B(n14836), .Z(n14805) );
  NAND U8939 ( .A(n14645), .B(n14644), .Z(n14649) );
  NAND U8940 ( .A(n14647), .B(n14646), .Z(n14648) );
  NAND U8941 ( .A(n14649), .B(n14648), .Z(n14829) );
  AND U8942 ( .A(y[23]), .B(x[5]), .Z(n14898) );
  AND U8943 ( .A(x[21]), .B(y[7]), .Z(n14897) );
  XOR U8944 ( .A(n14898), .B(n14897), .Z(n14900) );
  AND U8945 ( .A(y[8]), .B(x[20]), .Z(n14899) );
  XOR U8946 ( .A(n14900), .B(n14899), .Z(n14828) );
  AND U8947 ( .A(x[23]), .B(y[5]), .Z(n14921) );
  AND U8948 ( .A(y[25]), .B(x[3]), .Z(n14920) );
  XOR U8949 ( .A(n14921), .B(n14920), .Z(n14922) );
  XOR U8950 ( .A(n14923), .B(n14922), .Z(n14827) );
  XOR U8951 ( .A(n14828), .B(n14827), .Z(n14830) );
  XOR U8952 ( .A(n14829), .B(n14830), .Z(n14804) );
  NAND U8953 ( .A(n14651), .B(n14650), .Z(n14655) );
  NAND U8954 ( .A(n14653), .B(n14652), .Z(n14654) );
  NAND U8955 ( .A(n14655), .B(n14654), .Z(n14864) );
  NAND U8956 ( .A(x[0]), .B(y[28]), .Z(n14853) );
  NAND U8957 ( .A(o[27]), .B(n14656), .Z(n14852) );
  NAND U8958 ( .A(y[0]), .B(x[28]), .Z(n14851) );
  XOR U8959 ( .A(n14852), .B(n14851), .Z(n14854) );
  XOR U8960 ( .A(n14853), .B(n14854), .Z(n14863) );
  AND U8961 ( .A(x[10]), .B(y[18]), .Z(n14859) );
  AND U8962 ( .A(x[9]), .B(y[19]), .Z(n14657) );
  XOR U8963 ( .A(n14658), .B(n14657), .Z(n14858) );
  XOR U8964 ( .A(n14859), .B(n14858), .Z(n14862) );
  XOR U8965 ( .A(n14864), .B(n14865), .Z(n14823) );
  NAND U8966 ( .A(n14660), .B(n14659), .Z(n14664) );
  NAND U8967 ( .A(n14662), .B(n14661), .Z(n14663) );
  NAND U8968 ( .A(n14664), .B(n14663), .Z(n14822) );
  NAND U8969 ( .A(n14666), .B(n14665), .Z(n14670) );
  NAND U8970 ( .A(n14668), .B(n14667), .Z(n14669) );
  NAND U8971 ( .A(n14670), .B(n14669), .Z(n14821) );
  XOR U8972 ( .A(n14822), .B(n14821), .Z(n14824) );
  XNOR U8973 ( .A(n14823), .B(n14824), .Z(n14803) );
  XOR U8974 ( .A(n14805), .B(n14806), .Z(n14945) );
  XOR U8975 ( .A(n14942), .B(n14941), .Z(n14958) );
  NANDN U8976 ( .A(n14672), .B(n14671), .Z(n14676) );
  NANDN U8977 ( .A(n14674), .B(n14673), .Z(n14675) );
  AND U8978 ( .A(n14676), .B(n14675), .Z(n14694) );
  NAND U8979 ( .A(n14678), .B(n14677), .Z(n14682) );
  NAND U8980 ( .A(n14680), .B(n14679), .Z(n14681) );
  AND U8981 ( .A(n14682), .B(n14681), .Z(n14718) );
  XOR U8982 ( .A(n14684), .B(n14683), .Z(n14716) );
  XNOR U8983 ( .A(n14686), .B(n14685), .Z(n14715) );
  XOR U8984 ( .A(n14716), .B(n14715), .Z(n14717) );
  XNOR U8985 ( .A(n14718), .B(n14717), .Z(n14693) );
  NANDN U8986 ( .A(n14694), .B(n14693), .Z(n14696) );
  NANDN U8987 ( .A(n14688), .B(n14687), .Z(n14692) );
  NANDN U8988 ( .A(n14690), .B(n14689), .Z(n14691) );
  AND U8989 ( .A(n14692), .B(n14691), .Z(n14764) );
  XNOR U8990 ( .A(n14694), .B(n14693), .Z(n14763) );
  NANDN U8991 ( .A(n14764), .B(n14763), .Z(n14695) );
  AND U8992 ( .A(n14696), .B(n14695), .Z(n14957) );
  XNOR U8993 ( .A(n14958), .B(n14957), .Z(n14960) );
  NAND U8994 ( .A(n14698), .B(n14697), .Z(n14702) );
  NAND U8995 ( .A(n14700), .B(n14699), .Z(n14701) );
  NAND U8996 ( .A(n14702), .B(n14701), .Z(n14709) );
  NAND U8997 ( .A(n14704), .B(n14703), .Z(n14708) );
  NAND U8998 ( .A(n14706), .B(n14705), .Z(n14707) );
  AND U8999 ( .A(n14708), .B(n14707), .Z(n14710) );
  NANDN U9000 ( .A(n14709), .B(n14710), .Z(n14714) );
  XOR U9001 ( .A(n14710), .B(n14709), .Z(n14739) );
  XOR U9002 ( .A(n14712), .B(n14711), .Z(n14740) );
  OR U9003 ( .A(n14739), .B(n14740), .Z(n14713) );
  AND U9004 ( .A(n14714), .B(n14713), .Z(n14954) );
  NAND U9005 ( .A(n14716), .B(n14715), .Z(n14720) );
  NAND U9006 ( .A(n14718), .B(n14717), .Z(n14719) );
  AND U9007 ( .A(n14720), .B(n14719), .Z(n14952) );
  NANDN U9008 ( .A(n14722), .B(n14721), .Z(n14726) );
  NANDN U9009 ( .A(n14724), .B(n14723), .Z(n14725) );
  NAND U9010 ( .A(n14726), .B(n14725), .Z(n14735) );
  XOR U9011 ( .A(n14728), .B(n14727), .Z(n14736) );
  NANDN U9012 ( .A(n14735), .B(n14736), .Z(n14738) );
  NANDN U9013 ( .A(n14730), .B(n14729), .Z(n14734) );
  NAND U9014 ( .A(n14732), .B(n14731), .Z(n14733) );
  NAND U9015 ( .A(n14734), .B(n14733), .Z(n14741) );
  XNOR U9016 ( .A(n14736), .B(n14735), .Z(n14742) );
  NANDN U9017 ( .A(n14741), .B(n14742), .Z(n14737) );
  AND U9018 ( .A(n14738), .B(n14737), .Z(n14951) );
  XNOR U9019 ( .A(n14952), .B(n14951), .Z(n14953) );
  XNOR U9020 ( .A(n14954), .B(n14953), .Z(n14959) );
  XOR U9021 ( .A(n14960), .B(n14959), .Z(n14799) );
  XOR U9022 ( .A(n14740), .B(n14739), .Z(n14750) );
  XNOR U9023 ( .A(n14742), .B(n14741), .Z(n14749) );
  NANDN U9024 ( .A(n14750), .B(n14749), .Z(n14752) );
  NANDN U9025 ( .A(n14744), .B(n14743), .Z(n14748) );
  NANDN U9026 ( .A(n14746), .B(n14745), .Z(n14747) );
  AND U9027 ( .A(n14748), .B(n14747), .Z(n14760) );
  XNOR U9028 ( .A(n14750), .B(n14749), .Z(n14759) );
  NANDN U9029 ( .A(n14760), .B(n14759), .Z(n14751) );
  AND U9030 ( .A(n14752), .B(n14751), .Z(n14798) );
  NANDN U9031 ( .A(n14754), .B(n14753), .Z(n14758) );
  NANDN U9032 ( .A(n14756), .B(n14755), .Z(n14757) );
  AND U9033 ( .A(n14758), .B(n14757), .Z(n14762) );
  XNOR U9034 ( .A(n14760), .B(n14759), .Z(n14761) );
  NANDN U9035 ( .A(n14762), .B(n14761), .Z(n14766) );
  XNOR U9036 ( .A(n14762), .B(n14761), .Z(n14780) );
  XNOR U9037 ( .A(n14764), .B(n14763), .Z(n14779) );
  NAND U9038 ( .A(n14780), .B(n14779), .Z(n14765) );
  NAND U9039 ( .A(n14766), .B(n14765), .Z(n14797) );
  XOR U9040 ( .A(n14798), .B(n14797), .Z(n14800) );
  XOR U9041 ( .A(n14799), .B(n14800), .Z(n14964) );
  NAND U9042 ( .A(n14771), .B(n14770), .Z(n14775) );
  NAND U9043 ( .A(n14773), .B(n14772), .Z(n14774) );
  AND U9044 ( .A(n14775), .B(n14774), .Z(n14792) );
  XOR U9045 ( .A(n14792), .B(n14791), .Z(n14794) );
  XNOR U9046 ( .A(n14780), .B(n14779), .Z(n14793) );
  XNOR U9047 ( .A(n14794), .B(n14793), .Z(n14781) );
  NANDN U9048 ( .A(n14782), .B(n14781), .Z(n14790) );
  XNOR U9049 ( .A(n14782), .B(n14781), .Z(n15145) );
  NAND U9050 ( .A(n14784), .B(n14783), .Z(n14788) );
  NAND U9051 ( .A(n14786), .B(n14785), .Z(n14787) );
  AND U9052 ( .A(n14788), .B(n14787), .Z(n15144) );
  NAND U9053 ( .A(n15145), .B(n15144), .Z(n14789) );
  AND U9054 ( .A(n14790), .B(n14789), .Z(n14963) );
  XNOR U9055 ( .A(n14964), .B(n14963), .Z(n14966) );
  NAND U9056 ( .A(n14792), .B(n14791), .Z(n14796) );
  NAND U9057 ( .A(n14794), .B(n14793), .Z(n14795) );
  NAND U9058 ( .A(n14796), .B(n14795), .Z(n14965) );
  XNOR U9059 ( .A(n14966), .B(n14965), .Z(N61) );
  NANDN U9060 ( .A(n14798), .B(n14797), .Z(n14802) );
  OR U9061 ( .A(n14800), .B(n14799), .Z(n14801) );
  AND U9062 ( .A(n14802), .B(n14801), .Z(n14976) );
  NANDN U9063 ( .A(n14804), .B(n14803), .Z(n14808) );
  NANDN U9064 ( .A(n14806), .B(n14805), .Z(n14807) );
  AND U9065 ( .A(n14808), .B(n14807), .Z(n14994) );
  NAND U9066 ( .A(n14810), .B(n14809), .Z(n14814) );
  NAND U9067 ( .A(n14812), .B(n14811), .Z(n14813) );
  AND U9068 ( .A(n14814), .B(n14813), .Z(n14993) );
  XOR U9069 ( .A(n14994), .B(n14993), .Z(n14996) );
  NANDN U9070 ( .A(n14816), .B(n14815), .Z(n14820) );
  NANDN U9071 ( .A(n14818), .B(n14817), .Z(n14819) );
  NAND U9072 ( .A(n14820), .B(n14819), .Z(n14988) );
  NAND U9073 ( .A(n14822), .B(n14821), .Z(n14826) );
  NAND U9074 ( .A(n14824), .B(n14823), .Z(n14825) );
  NAND U9075 ( .A(n14826), .B(n14825), .Z(n15128) );
  NAND U9076 ( .A(n14828), .B(n14827), .Z(n14832) );
  NAND U9077 ( .A(n14830), .B(n14829), .Z(n14831) );
  NAND U9078 ( .A(n14832), .B(n14831), .Z(n15127) );
  NAND U9079 ( .A(n14834), .B(n14833), .Z(n14838) );
  NAND U9080 ( .A(n14836), .B(n14835), .Z(n14837) );
  NAND U9081 ( .A(n14838), .B(n14837), .Z(n15126) );
  XOR U9082 ( .A(n15127), .B(n15126), .Z(n15129) );
  XOR U9083 ( .A(n15128), .B(n15129), .Z(n14987) );
  XOR U9084 ( .A(n14988), .B(n14987), .Z(n14990) );
  NAND U9085 ( .A(n14840), .B(n14839), .Z(n14844) );
  NAND U9086 ( .A(n14842), .B(n14841), .Z(n14843) );
  AND U9087 ( .A(n14844), .B(n14843), .Z(n14989) );
  XOR U9088 ( .A(n14990), .B(n14989), .Z(n14995) );
  XOR U9089 ( .A(n14996), .B(n14995), .Z(n15002) );
  NAND U9090 ( .A(n14846), .B(n14845), .Z(n14850) );
  NAND U9091 ( .A(n14848), .B(n14847), .Z(n14849) );
  NAND U9092 ( .A(n14850), .B(n14849), .Z(n15036) );
  NAND U9093 ( .A(n14852), .B(n14851), .Z(n14856) );
  NAND U9094 ( .A(n14854), .B(n14853), .Z(n14855) );
  AND U9095 ( .A(n14856), .B(n14855), .Z(n15037) );
  XOR U9096 ( .A(n15036), .B(n15037), .Z(n15038) );
  AND U9097 ( .A(x[9]), .B(y[20]), .Z(n15300) );
  NANDN U9098 ( .A(n14857), .B(n15300), .Z(n14861) );
  NAND U9099 ( .A(n14859), .B(n14858), .Z(n14860) );
  NAND U9100 ( .A(n14861), .B(n14860), .Z(n15007) );
  AND U9101 ( .A(y[17]), .B(x[12]), .Z(n15064) );
  AND U9102 ( .A(x[1]), .B(y[28]), .Z(n15063) );
  XOR U9103 ( .A(n15064), .B(n15063), .Z(n15066) );
  AND U9104 ( .A(x[22]), .B(y[7]), .Z(n15065) );
  XOR U9105 ( .A(n15066), .B(n15065), .Z(n15006) );
  AND U9106 ( .A(x[15]), .B(y[14]), .Z(n15056) );
  XOR U9107 ( .A(n15059), .B(n15058), .Z(n15005) );
  XOR U9108 ( .A(n15006), .B(n15005), .Z(n15008) );
  XNOR U9109 ( .A(n15007), .B(n15008), .Z(n15039) );
  NANDN U9110 ( .A(n14863), .B(n14862), .Z(n14867) );
  NAND U9111 ( .A(n14865), .B(n14864), .Z(n14866) );
  AND U9112 ( .A(n14867), .B(n14866), .Z(n15042) );
  NAND U9113 ( .A(n14869), .B(n14868), .Z(n14873) );
  NANDN U9114 ( .A(n14871), .B(n14870), .Z(n14872) );
  AND U9115 ( .A(n14873), .B(n14872), .Z(n15044) );
  XOR U9116 ( .A(n15045), .B(n15044), .Z(n15141) );
  NAND U9117 ( .A(n14875), .B(n14874), .Z(n14879) );
  NAND U9118 ( .A(n14877), .B(n14876), .Z(n14878) );
  NAND U9119 ( .A(n14879), .B(n14878), .Z(n15138) );
  AND U9120 ( .A(x[3]), .B(y[26]), .Z(n15075) );
  AND U9121 ( .A(x[17]), .B(y[12]), .Z(n15074) );
  XOR U9122 ( .A(n15075), .B(n15074), .Z(n15077) );
  AND U9123 ( .A(x[11]), .B(y[18]), .Z(n15076) );
  XOR U9124 ( .A(n15077), .B(n15076), .Z(n15109) );
  AND U9125 ( .A(y[16]), .B(x[13]), .Z(n15086) );
  AND U9126 ( .A(y[5]), .B(x[24]), .Z(n15085) );
  XOR U9127 ( .A(n15086), .B(n15085), .Z(n15087) );
  AND U9128 ( .A(y[6]), .B(x[23]), .Z(n15369) );
  XOR U9129 ( .A(n15087), .B(n15369), .Z(n15108) );
  XOR U9130 ( .A(n15109), .B(n15108), .Z(n15111) );
  NAND U9131 ( .A(n14881), .B(n14880), .Z(n14885) );
  NAND U9132 ( .A(n14883), .B(n14882), .Z(n14884) );
  AND U9133 ( .A(n14885), .B(n14884), .Z(n15110) );
  XOR U9134 ( .A(n15111), .B(n15110), .Z(n15013) );
  NAND U9135 ( .A(n14887), .B(n14886), .Z(n14891) );
  NAND U9136 ( .A(n14889), .B(n14888), .Z(n14890) );
  NAND U9137 ( .A(n14891), .B(n14890), .Z(n15012) );
  NAND U9138 ( .A(n15069), .B(n14892), .Z(n14896) );
  NAND U9139 ( .A(n14894), .B(n14893), .Z(n14895) );
  NAND U9140 ( .A(n14896), .B(n14895), .Z(n15011) );
  XNOR U9141 ( .A(n15012), .B(n15011), .Z(n15014) );
  NAND U9142 ( .A(n14898), .B(n14897), .Z(n14902) );
  NAND U9143 ( .A(n14900), .B(n14899), .Z(n14901) );
  NAND U9144 ( .A(n14902), .B(n14901), .Z(n15050) );
  AND U9145 ( .A(y[1]), .B(o[28]), .Z(n15092) );
  XOR U9146 ( .A(n15092), .B(y[2]), .Z(n14903) );
  AND U9147 ( .A(x[27]), .B(n14903), .Z(n15091) );
  AND U9148 ( .A(x[16]), .B(y[13]), .Z(n15090) );
  XOR U9149 ( .A(n15091), .B(n15090), .Z(n15049) );
  NAND U9150 ( .A(x[18]), .B(y[11]), .Z(n14904) );
  XNOR U9151 ( .A(n14905), .B(n14904), .Z(n15103) );
  AND U9152 ( .A(x[2]), .B(y[27]), .Z(n15102) );
  XOR U9153 ( .A(n15103), .B(n15102), .Z(n15048) );
  XOR U9154 ( .A(n15049), .B(n15048), .Z(n15051) );
  XOR U9155 ( .A(n15050), .B(n15051), .Z(n15133) );
  AND U9156 ( .A(n15080), .B(n14906), .Z(n14909) );
  NAND U9157 ( .A(n15101), .B(n14907), .Z(n14908) );
  NANDN U9158 ( .A(n14909), .B(n14908), .Z(n15019) );
  AND U9159 ( .A(y[3]), .B(x[26]), .Z(n14911) );
  NAND U9160 ( .A(x[25]), .B(y[4]), .Z(n14910) );
  XNOR U9161 ( .A(n14911), .B(n14910), .Z(n15071) );
  XOR U9162 ( .A(n15071), .B(n15070), .Z(n15018) );
  AND U9163 ( .A(y[1]), .B(x[28]), .Z(n15062) );
  XOR U9164 ( .A(o[29]), .B(n15062), .Z(n15024) );
  AND U9165 ( .A(x[0]), .B(y[29]), .Z(n15023) );
  XOR U9166 ( .A(n15024), .B(n15023), .Z(n15026) );
  AND U9167 ( .A(y[0]), .B(x[29]), .Z(n15025) );
  XOR U9168 ( .A(n15026), .B(n15025), .Z(n15017) );
  XOR U9169 ( .A(n15018), .B(n15017), .Z(n15020) );
  XNOR U9170 ( .A(n15019), .B(n15020), .Z(n15132) );
  AND U9171 ( .A(y[19]), .B(x[10]), .Z(n15097) );
  AND U9172 ( .A(x[4]), .B(y[25]), .Z(n15096) );
  XOR U9173 ( .A(n15097), .B(n15096), .Z(n15098) );
  AND U9174 ( .A(y[24]), .B(x[5]), .Z(n15248) );
  XOR U9175 ( .A(n15098), .B(n15248), .Z(n15032) );
  AND U9176 ( .A(x[7]), .B(y[22]), .Z(n14913) );
  NAND U9177 ( .A(y[23]), .B(x[6]), .Z(n14912) );
  XNOR U9178 ( .A(n14913), .B(n14912), .Z(n15082) );
  AND U9179 ( .A(x[8]), .B(y[21]), .Z(n15081) );
  XOR U9180 ( .A(n15082), .B(n15081), .Z(n15031) );
  XOR U9181 ( .A(n15032), .B(n15031), .Z(n15033) );
  XOR U9182 ( .A(n15300), .B(n15033), .Z(n15117) );
  IV U9183 ( .A(n15117), .Z(n14926) );
  NAND U9184 ( .A(n14915), .B(n14914), .Z(n14919) );
  NAND U9185 ( .A(n14917), .B(n14916), .Z(n14918) );
  AND U9186 ( .A(n14919), .B(n14918), .Z(n15115) );
  NAND U9187 ( .A(n14921), .B(n14920), .Z(n14925) );
  NAND U9188 ( .A(n14923), .B(n14922), .Z(n14924) );
  AND U9189 ( .A(n14925), .B(n14924), .Z(n15114) );
  XOR U9190 ( .A(n15115), .B(n15114), .Z(n15116) );
  XOR U9191 ( .A(n14926), .B(n15116), .Z(n15121) );
  NANDN U9192 ( .A(n14928), .B(n14927), .Z(n14932) );
  NANDN U9193 ( .A(n14930), .B(n14929), .Z(n14931) );
  NAND U9194 ( .A(n14932), .B(n14931), .Z(n15120) );
  XOR U9195 ( .A(n15138), .B(n15139), .Z(n15140) );
  NAND U9196 ( .A(n14934), .B(n14933), .Z(n14938) );
  NANDN U9197 ( .A(n14936), .B(n14935), .Z(n14937) );
  AND U9198 ( .A(n14938), .B(n14937), .Z(n14999) );
  XOR U9199 ( .A(n15000), .B(n14999), .Z(n15001) );
  XOR U9200 ( .A(n15002), .B(n15001), .Z(n14982) );
  NAND U9201 ( .A(n14940), .B(n14939), .Z(n14944) );
  NAND U9202 ( .A(n14942), .B(n14941), .Z(n14943) );
  AND U9203 ( .A(n14944), .B(n14943), .Z(n14981) );
  NANDN U9204 ( .A(n14946), .B(n14945), .Z(n14950) );
  NANDN U9205 ( .A(n14948), .B(n14947), .Z(n14949) );
  AND U9206 ( .A(n14950), .B(n14949), .Z(n14983) );
  XOR U9207 ( .A(n14984), .B(n14983), .Z(n14972) );
  NANDN U9208 ( .A(n14952), .B(n14951), .Z(n14956) );
  NANDN U9209 ( .A(n14954), .B(n14953), .Z(n14955) );
  AND U9210 ( .A(n14956), .B(n14955), .Z(n14969) );
  NANDN U9211 ( .A(n14958), .B(n14957), .Z(n14962) );
  NAND U9212 ( .A(n14960), .B(n14959), .Z(n14961) );
  NAND U9213 ( .A(n14962), .B(n14961), .Z(n14970) );
  XNOR U9214 ( .A(n14969), .B(n14970), .Z(n14971) );
  XNOR U9215 ( .A(n14972), .B(n14971), .Z(n14975) );
  XNOR U9216 ( .A(n14976), .B(n14975), .Z(n14978) );
  NANDN U9217 ( .A(n14964), .B(n14963), .Z(n14968) );
  NAND U9218 ( .A(n14966), .B(n14965), .Z(n14967) );
  AND U9219 ( .A(n14968), .B(n14967), .Z(n14977) );
  XOR U9220 ( .A(n14978), .B(n14977), .Z(N62) );
  NANDN U9221 ( .A(n14970), .B(n14969), .Z(n14974) );
  NANDN U9222 ( .A(n14972), .B(n14971), .Z(n14973) );
  AND U9223 ( .A(n14974), .B(n14973), .Z(n15170) );
  NANDN U9224 ( .A(n14976), .B(n14975), .Z(n14980) );
  NAND U9225 ( .A(n14978), .B(n14977), .Z(n14979) );
  NAND U9226 ( .A(n14980), .B(n14979), .Z(n15171) );
  NANDN U9227 ( .A(n14982), .B(n14981), .Z(n14986) );
  NAND U9228 ( .A(n14984), .B(n14983), .Z(n14985) );
  NAND U9229 ( .A(n14986), .B(n14985), .Z(n15457) );
  NAND U9230 ( .A(n14988), .B(n14987), .Z(n14992) );
  NAND U9231 ( .A(n14990), .B(n14989), .Z(n14991) );
  AND U9232 ( .A(n14992), .B(n14991), .Z(n15175) );
  NAND U9233 ( .A(n14994), .B(n14993), .Z(n14998) );
  NAND U9234 ( .A(n14996), .B(n14995), .Z(n14997) );
  AND U9235 ( .A(n14998), .B(n14997), .Z(n15177) );
  NAND U9236 ( .A(n15000), .B(n14999), .Z(n15004) );
  NAND U9237 ( .A(n15002), .B(n15001), .Z(n15003) );
  AND U9238 ( .A(n15004), .B(n15003), .Z(n15176) );
  XOR U9239 ( .A(n15177), .B(n15176), .Z(n15174) );
  XOR U9240 ( .A(n15175), .B(n15174), .Z(n15456) );
  NAND U9241 ( .A(n15006), .B(n15005), .Z(n15010) );
  NAND U9242 ( .A(n15008), .B(n15007), .Z(n15009) );
  AND U9243 ( .A(n15010), .B(n15009), .Z(n15194) );
  NAND U9244 ( .A(n15012), .B(n15011), .Z(n15016) );
  NANDN U9245 ( .A(n15014), .B(n15013), .Z(n15015) );
  NAND U9246 ( .A(n15016), .B(n15015), .Z(n15195) );
  XNOR U9247 ( .A(n15194), .B(n15195), .Z(n15193) );
  NAND U9248 ( .A(n15018), .B(n15017), .Z(n15022) );
  NAND U9249 ( .A(n15020), .B(n15019), .Z(n15021) );
  AND U9250 ( .A(n15022), .B(n15021), .Z(n15192) );
  XOR U9251 ( .A(n15193), .B(n15192), .Z(n15425) );
  NAND U9252 ( .A(n15024), .B(n15023), .Z(n15028) );
  NAND U9253 ( .A(n15026), .B(n15025), .Z(n15027) );
  NAND U9254 ( .A(n15028), .B(n15027), .Z(n15200) );
  AND U9255 ( .A(x[1]), .B(y[29]), .Z(n15243) );
  AND U9256 ( .A(x[15]), .B(y[15]), .Z(n15242) );
  XOR U9257 ( .A(n15243), .B(n15242), .Z(n15241) );
  AND U9258 ( .A(x[27]), .B(y[3]), .Z(n15240) );
  XOR U9259 ( .A(n15241), .B(n15240), .Z(n15203) );
  AND U9260 ( .A(x[12]), .B(y[18]), .Z(n15283) );
  XOR U9261 ( .A(n15284), .B(n15283), .Z(n15298) );
  AND U9262 ( .A(x[9]), .B(y[21]), .Z(n15030) );
  NAND U9263 ( .A(y[20]), .B(x[10]), .Z(n15029) );
  XNOR U9264 ( .A(n15030), .B(n15029), .Z(n15297) );
  XOR U9265 ( .A(n15298), .B(n15297), .Z(n15202) );
  XOR U9266 ( .A(n15203), .B(n15202), .Z(n15201) );
  XOR U9267 ( .A(n15200), .B(n15201), .Z(n15183) );
  NAND U9268 ( .A(n15032), .B(n15031), .Z(n15035) );
  NAND U9269 ( .A(n15300), .B(n15033), .Z(n15034) );
  AND U9270 ( .A(n15035), .B(n15034), .Z(n15182) );
  NAND U9271 ( .A(n15037), .B(n15036), .Z(n15041) );
  NANDN U9272 ( .A(n15039), .B(n15038), .Z(n15040) );
  AND U9273 ( .A(n15041), .B(n15040), .Z(n15180) );
  XNOR U9274 ( .A(n15181), .B(n15180), .Z(n15426) );
  NANDN U9275 ( .A(n15043), .B(n15042), .Z(n15047) );
  NAND U9276 ( .A(n15045), .B(n15044), .Z(n15046) );
  AND U9277 ( .A(n15047), .B(n15046), .Z(n15427) );
  XNOR U9278 ( .A(n15428), .B(n15427), .Z(n15463) );
  NAND U9279 ( .A(n15049), .B(n15048), .Z(n15053) );
  NAND U9280 ( .A(n15051), .B(n15050), .Z(n15052) );
  NAND U9281 ( .A(n15053), .B(n15052), .Z(n15419) );
  AND U9282 ( .A(y[7]), .B(x[23]), .Z(n15055) );
  NAND U9283 ( .A(x[24]), .B(y[6]), .Z(n15054) );
  XNOR U9284 ( .A(n15055), .B(n15054), .Z(n15368) );
  AND U9285 ( .A(y[5]), .B(x[25]), .Z(n15367) );
  XOR U9286 ( .A(n15368), .B(n15367), .Z(n15280) );
  NANDN U9287 ( .A(n15057), .B(n15056), .Z(n15061) );
  NAND U9288 ( .A(n15059), .B(n15058), .Z(n15060) );
  AND U9289 ( .A(n15061), .B(n15060), .Z(n15279) );
  AND U9290 ( .A(n15062), .B(o[29]), .Z(n15318) );
  AND U9291 ( .A(x[16]), .B(y[14]), .Z(n15317) );
  XOR U9292 ( .A(n15318), .B(n15317), .Z(n15316) );
  AND U9293 ( .A(y[2]), .B(x[28]), .Z(n15315) );
  XOR U9294 ( .A(n15316), .B(n15315), .Z(n15278) );
  NAND U9295 ( .A(n15064), .B(n15063), .Z(n15068) );
  NAND U9296 ( .A(n15066), .B(n15065), .Z(n15067) );
  NAND U9297 ( .A(n15068), .B(n15067), .Z(n15409) );
  AND U9298 ( .A(y[4]), .B(x[26]), .Z(n15376) );
  NAND U9299 ( .A(n15069), .B(n15376), .Z(n15073) );
  NAND U9300 ( .A(n15071), .B(n15070), .Z(n15072) );
  NAND U9301 ( .A(n15073), .B(n15072), .Z(n15407) );
  XOR U9302 ( .A(n15408), .B(n15407), .Z(n15421) );
  AND U9303 ( .A(x[0]), .B(y[30]), .Z(n15336) );
  AND U9304 ( .A(y[1]), .B(x[29]), .Z(n15289) );
  XOR U9305 ( .A(o[30]), .B(n15289), .Z(n15338) );
  AND U9306 ( .A(y[0]), .B(x[30]), .Z(n15337) );
  XOR U9307 ( .A(n15338), .B(n15337), .Z(n15335) );
  XOR U9308 ( .A(n15336), .B(n15335), .Z(n15223) );
  AND U9309 ( .A(y[10]), .B(x[20]), .Z(n15389) );
  AND U9310 ( .A(y[22]), .B(x[8]), .Z(n15387) );
  XNOR U9311 ( .A(n15388), .B(n15387), .Z(n15222) );
  NAND U9312 ( .A(n15075), .B(n15074), .Z(n15079) );
  NAND U9313 ( .A(n15077), .B(n15076), .Z(n15078) );
  AND U9314 ( .A(n15079), .B(n15078), .Z(n15220) );
  XOR U9315 ( .A(n15221), .B(n15220), .Z(n15212) );
  AND U9316 ( .A(x[22]), .B(y[8]), .Z(n15254) );
  AND U9317 ( .A(x[7]), .B(y[23]), .Z(n15252) );
  AND U9318 ( .A(y[9]), .B(x[21]), .Z(n15251) );
  XOR U9319 ( .A(n15252), .B(n15251), .Z(n15253) );
  XOR U9320 ( .A(n15254), .B(n15253), .Z(n15233) );
  AND U9321 ( .A(x[2]), .B(y[28]), .Z(n15374) );
  AND U9322 ( .A(x[17]), .B(y[13]), .Z(n15373) );
  XOR U9323 ( .A(n15374), .B(n15373), .Z(n15375) );
  XOR U9324 ( .A(n15376), .B(n15375), .Z(n15235) );
  NAND U9325 ( .A(n15080), .B(n15252), .Z(n15084) );
  NAND U9326 ( .A(n15082), .B(n15081), .Z(n15083) );
  NAND U9327 ( .A(n15084), .B(n15083), .Z(n15234) );
  XOR U9328 ( .A(n15235), .B(n15234), .Z(n15232) );
  XOR U9329 ( .A(n15233), .B(n15232), .Z(n15215) );
  NAND U9330 ( .A(n15086), .B(n15085), .Z(n15089) );
  NAND U9331 ( .A(n15087), .B(n15369), .Z(n15088) );
  AND U9332 ( .A(n15089), .B(n15088), .Z(n15214) );
  XNOR U9333 ( .A(n15212), .B(n15213), .Z(n15422) );
  XOR U9334 ( .A(n15419), .B(n15420), .Z(n15444) );
  NAND U9335 ( .A(n15091), .B(n15090), .Z(n15095) );
  NAND U9336 ( .A(n15092), .B(x[27]), .Z(n15093) );
  NANDN U9337 ( .A(n15093), .B(y[2]), .Z(n15094) );
  AND U9338 ( .A(n15095), .B(n15094), .Z(n15207) );
  NAND U9339 ( .A(n15097), .B(n15096), .Z(n15100) );
  NAND U9340 ( .A(n15098), .B(n15248), .Z(n15099) );
  NAND U9341 ( .A(n15100), .B(n15099), .Z(n15208) );
  AND U9342 ( .A(y[11]), .B(x[19]), .Z(n15247) );
  NAND U9343 ( .A(n15101), .B(n15247), .Z(n15105) );
  NAND U9344 ( .A(n15103), .B(n15102), .Z(n15104) );
  NAND U9345 ( .A(n15105), .B(n15104), .Z(n15226) );
  AND U9346 ( .A(x[18]), .B(y[12]), .Z(n15384) );
  AND U9347 ( .A(x[4]), .B(y[26]), .Z(n15383) );
  XOR U9348 ( .A(n15384), .B(n15383), .Z(n15382) );
  AND U9349 ( .A(x[3]), .B(y[27]), .Z(n15381) );
  XOR U9350 ( .A(n15382), .B(n15381), .Z(n15229) );
  AND U9351 ( .A(x[5]), .B(y[25]), .Z(n15107) );
  NAND U9352 ( .A(x[6]), .B(y[24]), .Z(n15106) );
  XNOR U9353 ( .A(n15107), .B(n15106), .Z(n15246) );
  XOR U9354 ( .A(n15247), .B(n15246), .Z(n15228) );
  XOR U9355 ( .A(n15229), .B(n15228), .Z(n15227) );
  XOR U9356 ( .A(n15226), .B(n15227), .Z(n15209) );
  XOR U9357 ( .A(n15208), .B(n15209), .Z(n15206) );
  XNOR U9358 ( .A(n15207), .B(n15206), .Z(n15186) );
  NAND U9359 ( .A(n15109), .B(n15108), .Z(n15113) );
  NAND U9360 ( .A(n15111), .B(n15110), .Z(n15112) );
  NAND U9361 ( .A(n15113), .B(n15112), .Z(n15188) );
  NAND U9362 ( .A(n15115), .B(n15114), .Z(n15119) );
  NANDN U9363 ( .A(n15117), .B(n15116), .Z(n15118) );
  AND U9364 ( .A(n15119), .B(n15118), .Z(n15189) );
  XNOR U9365 ( .A(n15188), .B(n15189), .Z(n15187) );
  NANDN U9366 ( .A(n15121), .B(n15120), .Z(n15125) );
  NANDN U9367 ( .A(n15123), .B(n15122), .Z(n15124) );
  AND U9368 ( .A(n15125), .B(n15124), .Z(n15445) );
  NAND U9369 ( .A(n15127), .B(n15126), .Z(n15131) );
  NAND U9370 ( .A(n15129), .B(n15128), .Z(n15130) );
  NAND U9371 ( .A(n15131), .B(n15130), .Z(n15439) );
  NANDN U9372 ( .A(n15133), .B(n15132), .Z(n15137) );
  NANDN U9373 ( .A(n15135), .B(n15134), .Z(n15136) );
  AND U9374 ( .A(n15137), .B(n15136), .Z(n15437) );
  XOR U9375 ( .A(n15438), .B(n15437), .Z(n15462) );
  NAND U9376 ( .A(n15139), .B(n15138), .Z(n15143) );
  NANDN U9377 ( .A(n15141), .B(n15140), .Z(n15142) );
  AND U9378 ( .A(n15143), .B(n15142), .Z(n15461) );
  XOR U9379 ( .A(n15463), .B(n15464), .Z(n15455) );
  XNOR U9380 ( .A(n15456), .B(n15455), .Z(n15458) );
  XOR U9381 ( .A(n15457), .B(n15458), .Z(n15168) );
  XNOR U9382 ( .A(n15169), .B(n15168), .Z(N63) );
  XOR U9383 ( .A(n15145), .B(n15144), .Z(n6253) );
  XNOR U9384 ( .A(n15147), .B(n15146), .Z(n6254) );
  XNOR U9385 ( .A(n15149), .B(n15148), .Z(n6255) );
  XNOR U9386 ( .A(n15151), .B(n15150), .Z(n6256) );
  XOR U9387 ( .A(n15153), .B(n15152), .Z(n15154) );
  XNOR U9388 ( .A(n15155), .B(n15154), .Z(n6257) );
  XOR U9389 ( .A(n15157), .B(n15156), .Z(n6258) );
  XOR U9390 ( .A(n15159), .B(n15158), .Z(n15160) );
  XNOR U9391 ( .A(n15161), .B(n15160), .Z(n6259) );
  XOR U9392 ( .A(n15163), .B(n15162), .Z(n12497) );
  XNOR U9393 ( .A(n15165), .B(n15164), .Z(n12496) );
  XOR U9394 ( .A(n15167), .B(n15166), .Z(n12495) );
  NAND U9395 ( .A(n15169), .B(n15168), .Z(n15173) );
  NANDN U9396 ( .A(n15171), .B(n15170), .Z(n15172) );
  AND U9397 ( .A(n15173), .B(n15172), .Z(n15454) );
  NAND U9398 ( .A(n15175), .B(n15174), .Z(n15179) );
  NAND U9399 ( .A(n15177), .B(n15176), .Z(n15178) );
  AND U9400 ( .A(n15179), .B(n15178), .Z(n15436) );
  NAND U9401 ( .A(n15181), .B(n15180), .Z(n15185) );
  NANDN U9402 ( .A(n15183), .B(n15182), .Z(n15184) );
  AND U9403 ( .A(n15185), .B(n15184), .Z(n15418) );
  NANDN U9404 ( .A(n15187), .B(n15186), .Z(n15191) );
  NAND U9405 ( .A(n15189), .B(n15188), .Z(n15190) );
  AND U9406 ( .A(n15191), .B(n15190), .Z(n15199) );
  NAND U9407 ( .A(n15193), .B(n15192), .Z(n15197) );
  NANDN U9408 ( .A(n15195), .B(n15194), .Z(n15196) );
  NAND U9409 ( .A(n15197), .B(n15196), .Z(n15198) );
  XNOR U9410 ( .A(n15199), .B(n15198), .Z(n15416) );
  NAND U9411 ( .A(n15201), .B(n15200), .Z(n15205) );
  NAND U9412 ( .A(n15203), .B(n15202), .Z(n15204) );
  AND U9413 ( .A(n15205), .B(n15204), .Z(n15406) );
  NANDN U9414 ( .A(n15207), .B(n15206), .Z(n15211) );
  NAND U9415 ( .A(n15209), .B(n15208), .Z(n15210) );
  AND U9416 ( .A(n15211), .B(n15210), .Z(n15219) );
  NANDN U9417 ( .A(n15213), .B(n15212), .Z(n15217) );
  NANDN U9418 ( .A(n15215), .B(n15214), .Z(n15216) );
  NAND U9419 ( .A(n15217), .B(n15216), .Z(n15218) );
  XNOR U9420 ( .A(n15219), .B(n15218), .Z(n15404) );
  NAND U9421 ( .A(n15221), .B(n15220), .Z(n15225) );
  NANDN U9422 ( .A(n15223), .B(n15222), .Z(n15224) );
  AND U9423 ( .A(n15225), .B(n15224), .Z(n15402) );
  NAND U9424 ( .A(n15227), .B(n15226), .Z(n15231) );
  NAND U9425 ( .A(n15229), .B(n15228), .Z(n15230) );
  AND U9426 ( .A(n15231), .B(n15230), .Z(n15239) );
  NAND U9427 ( .A(n15233), .B(n15232), .Z(n15237) );
  NAND U9428 ( .A(n15235), .B(n15234), .Z(n15236) );
  NAND U9429 ( .A(n15237), .B(n15236), .Z(n15238) );
  XNOR U9430 ( .A(n15239), .B(n15238), .Z(n15400) );
  NAND U9431 ( .A(n15241), .B(n15240), .Z(n15245) );
  NAND U9432 ( .A(n15243), .B(n15242), .Z(n15244) );
  AND U9433 ( .A(n15245), .B(n15244), .Z(n15276) );
  NAND U9434 ( .A(n15247), .B(n15246), .Z(n15250) );
  AND U9435 ( .A(x[6]), .B(y[25]), .Z(n15290) );
  AND U9436 ( .A(n15248), .B(n15290), .Z(n15249) );
  ANDN U9437 ( .B(n15250), .A(n15249), .Z(n15258) );
  AND U9438 ( .A(n15252), .B(n15251), .Z(n15256) );
  AND U9439 ( .A(n15254), .B(n15253), .Z(n15255) );
  OR U9440 ( .A(n15256), .B(n15255), .Z(n15257) );
  XNOR U9441 ( .A(n15258), .B(n15257), .Z(n15274) );
  AND U9442 ( .A(y[15]), .B(x[16]), .Z(n15260) );
  NAND U9443 ( .A(y[8]), .B(x[23]), .Z(n15259) );
  XNOR U9444 ( .A(n15260), .B(n15259), .Z(n15264) );
  AND U9445 ( .A(x[31]), .B(y[0]), .Z(n15262) );
  NAND U9446 ( .A(y[23]), .B(x[8]), .Z(n15261) );
  XNOR U9447 ( .A(n15262), .B(n15261), .Z(n15263) );
  XOR U9448 ( .A(n15264), .B(n15263), .Z(n15272) );
  AND U9449 ( .A(y[3]), .B(x[28]), .Z(n15266) );
  NAND U9450 ( .A(x[12]), .B(y[19]), .Z(n15265) );
  XNOR U9451 ( .A(n15266), .B(n15265), .Z(n15270) );
  AND U9452 ( .A(x[5]), .B(y[26]), .Z(n15268) );
  NAND U9453 ( .A(y[29]), .B(x[2]), .Z(n15267) );
  XNOR U9454 ( .A(n15268), .B(n15267), .Z(n15269) );
  XNOR U9455 ( .A(n15270), .B(n15269), .Z(n15271) );
  XNOR U9456 ( .A(n15272), .B(n15271), .Z(n15273) );
  XNOR U9457 ( .A(n15274), .B(n15273), .Z(n15275) );
  XNOR U9458 ( .A(n15276), .B(n15275), .Z(n15366) );
  NANDN U9459 ( .A(n15278), .B(n15277), .Z(n15282) );
  NANDN U9460 ( .A(n15280), .B(n15279), .Z(n15281) );
  AND U9461 ( .A(n15282), .B(n15281), .Z(n15364) );
  NAND U9462 ( .A(n15284), .B(n15283), .Z(n15288) );
  ANDN U9463 ( .B(n15286), .A(n15285), .Z(n15287) );
  ANDN U9464 ( .B(n15288), .A(n15287), .Z(n15314) );
  AND U9465 ( .A(y[14]), .B(x[17]), .Z(n15296) );
  AND U9466 ( .A(n15289), .B(o[30]), .Z(n15294) );
  XOR U9467 ( .A(n15290), .B(o[31]), .Z(n15292) );
  AND U9468 ( .A(x[10]), .B(y[21]), .Z(n15299) );
  XNOR U9469 ( .A(n15370), .B(n15299), .Z(n15291) );
  XNOR U9470 ( .A(n15292), .B(n15291), .Z(n15293) );
  XNOR U9471 ( .A(n15294), .B(n15293), .Z(n15295) );
  XNOR U9472 ( .A(n15296), .B(n15295), .Z(n15312) );
  NAND U9473 ( .A(n15298), .B(n15297), .Z(n15302) );
  NAND U9474 ( .A(n15300), .B(n15299), .Z(n15301) );
  AND U9475 ( .A(n15302), .B(n15301), .Z(n15310) );
  AND U9476 ( .A(x[20]), .B(y[11]), .Z(n15304) );
  NAND U9477 ( .A(x[7]), .B(y[24]), .Z(n15303) );
  XNOR U9478 ( .A(n15304), .B(n15303), .Z(n15308) );
  AND U9479 ( .A(y[31]), .B(x[0]), .Z(n15306) );
  NAND U9480 ( .A(x[29]), .B(y[2]), .Z(n15305) );
  XNOR U9481 ( .A(n15306), .B(n15305), .Z(n15307) );
  XNOR U9482 ( .A(n15308), .B(n15307), .Z(n15309) );
  XNOR U9483 ( .A(n15310), .B(n15309), .Z(n15311) );
  XNOR U9484 ( .A(n15312), .B(n15311), .Z(n15313) );
  XNOR U9485 ( .A(n15314), .B(n15313), .Z(n15362) );
  NAND U9486 ( .A(n15316), .B(n15315), .Z(n15320) );
  NAND U9487 ( .A(n15318), .B(n15317), .Z(n15319) );
  AND U9488 ( .A(n15320), .B(n15319), .Z(n15360) );
  AND U9489 ( .A(x[26]), .B(y[5]), .Z(n15322) );
  NAND U9490 ( .A(y[27]), .B(x[4]), .Z(n15321) );
  XNOR U9491 ( .A(n15322), .B(n15321), .Z(n15326) );
  AND U9492 ( .A(x[14]), .B(y[17]), .Z(n15324) );
  NAND U9493 ( .A(x[9]), .B(y[22]), .Z(n15323) );
  XNOR U9494 ( .A(n15324), .B(n15323), .Z(n15325) );
  XOR U9495 ( .A(n15326), .B(n15325), .Z(n15334) );
  AND U9496 ( .A(y[13]), .B(x[18]), .Z(n15328) );
  NAND U9497 ( .A(x[21]), .B(y[10]), .Z(n15327) );
  XNOR U9498 ( .A(n15328), .B(n15327), .Z(n15332) );
  AND U9499 ( .A(y[12]), .B(x[19]), .Z(n15330) );
  NAND U9500 ( .A(x[25]), .B(y[6]), .Z(n15329) );
  XNOR U9501 ( .A(n15330), .B(n15329), .Z(n15331) );
  XNOR U9502 ( .A(n15332), .B(n15331), .Z(n15333) );
  XNOR U9503 ( .A(n15334), .B(n15333), .Z(n15358) );
  NAND U9504 ( .A(n15336), .B(n15335), .Z(n15340) );
  NAND U9505 ( .A(n15338), .B(n15337), .Z(n15339) );
  AND U9506 ( .A(n15340), .B(n15339), .Z(n15356) );
  AND U9507 ( .A(y[28]), .B(x[3]), .Z(n15342) );
  NAND U9508 ( .A(y[20]), .B(x[11]), .Z(n15341) );
  XNOR U9509 ( .A(n15342), .B(n15341), .Z(n15354) );
  AND U9510 ( .A(y[30]), .B(x[1]), .Z(n15344) );
  NAND U9511 ( .A(x[27]), .B(y[4]), .Z(n15343) );
  XNOR U9512 ( .A(n15344), .B(n15343), .Z(n15348) );
  AND U9513 ( .A(x[30]), .B(y[1]), .Z(n15346) );
  NAND U9514 ( .A(y[9]), .B(x[22]), .Z(n15345) );
  XNOR U9515 ( .A(n15346), .B(n15345), .Z(n15347) );
  XOR U9516 ( .A(n15348), .B(n15347), .Z(n15352) );
  XNOR U9517 ( .A(n15350), .B(n15349), .Z(n15351) );
  XNOR U9518 ( .A(n15352), .B(n15351), .Z(n15353) );
  XNOR U9519 ( .A(n15354), .B(n15353), .Z(n15355) );
  XNOR U9520 ( .A(n15356), .B(n15355), .Z(n15357) );
  XNOR U9521 ( .A(n15358), .B(n15357), .Z(n15359) );
  XNOR U9522 ( .A(n15360), .B(n15359), .Z(n15361) );
  XNOR U9523 ( .A(n15362), .B(n15361), .Z(n15363) );
  XNOR U9524 ( .A(n15364), .B(n15363), .Z(n15365) );
  XOR U9525 ( .A(n15366), .B(n15365), .Z(n15398) );
  NAND U9526 ( .A(n15368), .B(n15367), .Z(n15372) );
  NAND U9527 ( .A(n15370), .B(n15369), .Z(n15371) );
  AND U9528 ( .A(n15372), .B(n15371), .Z(n15380) );
  NAND U9529 ( .A(n15374), .B(n15373), .Z(n15378) );
  NAND U9530 ( .A(n15376), .B(n15375), .Z(n15377) );
  AND U9531 ( .A(n15378), .B(n15377), .Z(n15379) );
  XNOR U9532 ( .A(n15380), .B(n15379), .Z(n15396) );
  NAND U9533 ( .A(n15382), .B(n15381), .Z(n15386) );
  NAND U9534 ( .A(n15384), .B(n15383), .Z(n15385) );
  AND U9535 ( .A(n15386), .B(n15385), .Z(n15394) );
  NAND U9536 ( .A(n15388), .B(n15387), .Z(n15392) );
  NANDN U9537 ( .A(n15390), .B(n15389), .Z(n15391) );
  NAND U9538 ( .A(n15392), .B(n15391), .Z(n15393) );
  XNOR U9539 ( .A(n15394), .B(n15393), .Z(n15395) );
  XOR U9540 ( .A(n15396), .B(n15395), .Z(n15397) );
  XNOR U9541 ( .A(n15398), .B(n15397), .Z(n15399) );
  XNOR U9542 ( .A(n15400), .B(n15399), .Z(n15401) );
  XNOR U9543 ( .A(n15402), .B(n15401), .Z(n15403) );
  XNOR U9544 ( .A(n15404), .B(n15403), .Z(n15405) );
  XNOR U9545 ( .A(n15406), .B(n15405), .Z(n15414) );
  NAND U9546 ( .A(n15408), .B(n15407), .Z(n15412) );
  NANDN U9547 ( .A(n15410), .B(n15409), .Z(n15411) );
  NAND U9548 ( .A(n15412), .B(n15411), .Z(n15413) );
  XNOR U9549 ( .A(n15414), .B(n15413), .Z(n15415) );
  XNOR U9550 ( .A(n15416), .B(n15415), .Z(n15417) );
  XNOR U9551 ( .A(n15418), .B(n15417), .Z(n15434) );
  NAND U9552 ( .A(n15420), .B(n15419), .Z(n15424) );
  NANDN U9553 ( .A(n15422), .B(n15421), .Z(n15423) );
  AND U9554 ( .A(n15424), .B(n15423), .Z(n15432) );
  ANDN U9555 ( .B(n15426), .A(n15425), .Z(n15430) );
  AND U9556 ( .A(n15428), .B(n15427), .Z(n15429) );
  OR U9557 ( .A(n15430), .B(n15429), .Z(n15431) );
  XNOR U9558 ( .A(n15432), .B(n15431), .Z(n15433) );
  XNOR U9559 ( .A(n15434), .B(n15433), .Z(n15435) );
  XNOR U9560 ( .A(n15436), .B(n15435), .Z(n15452) );
  NAND U9561 ( .A(n15438), .B(n15437), .Z(n15442) );
  NANDN U9562 ( .A(n15440), .B(n15439), .Z(n15441) );
  AND U9563 ( .A(n15442), .B(n15441), .Z(n15450) );
  NANDN U9564 ( .A(n15444), .B(n15443), .Z(n15448) );
  NANDN U9565 ( .A(n15446), .B(n15445), .Z(n15447) );
  NAND U9566 ( .A(n15448), .B(n15447), .Z(n15449) );
  XNOR U9567 ( .A(n15450), .B(n15449), .Z(n15451) );
  XNOR U9568 ( .A(n15452), .B(n15451), .Z(n15453) );
  XNOR U9569 ( .A(n15454), .B(n15453), .Z(n15470) );
  ANDN U9570 ( .B(n15456), .A(n15455), .Z(n15460) );
  AND U9571 ( .A(n15458), .B(n15457), .Z(n15459) );
  NOR U9572 ( .A(n15460), .B(n15459), .Z(n15468) );
  NANDN U9573 ( .A(n15462), .B(n15461), .Z(n15466) );
  NANDN U9574 ( .A(n15464), .B(n15463), .Z(n15465) );
  AND U9575 ( .A(n15466), .B(n15465), .Z(n15467) );
  XNOR U9576 ( .A(n15468), .B(n15467), .Z(n15469) );
  XNOR U9577 ( .A(n15470), .B(n15469), .Z(n12494) );
endmodule

