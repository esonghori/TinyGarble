
module sum_N256_CC2 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[1]), .B(n507), .Z(n93) );
  XOR U4 ( .A(a[4]), .B(n498), .Z(n60) );
  XOR U5 ( .A(a[7]), .B(n489), .Z(n27) );
  XOR U6 ( .A(a[10]), .B(n480), .Z(n175) );
  XOR U7 ( .A(a[13]), .B(n471), .Z(n100) );
  XOR U8 ( .A(a[16]), .B(n462), .Z(n97) );
  XOR U9 ( .A(a[19]), .B(n453), .Z(n94) );
  XOR U10 ( .A(a[22]), .B(n444), .Z(n90) );
  XOR U11 ( .A(a[25]), .B(n435), .Z(n87) );
  XOR U12 ( .A(a[28]), .B(n426), .Z(n84) );
  XOR U13 ( .A(a[31]), .B(n417), .Z(n80) );
  XOR U14 ( .A(a[34]), .B(n408), .Z(n77) );
  XOR U15 ( .A(a[37]), .B(n399), .Z(n74) );
  XOR U16 ( .A(a[40]), .B(n390), .Z(n70) );
  XOR U17 ( .A(a[43]), .B(n381), .Z(n67) );
  XOR U18 ( .A(a[46]), .B(n372), .Z(n64) );
  XOR U19 ( .A(a[49]), .B(n363), .Z(n61) );
  XOR U20 ( .A(a[52]), .B(n354), .Z(n57) );
  XOR U21 ( .A(a[55]), .B(n345), .Z(n54) );
  XOR U22 ( .A(a[58]), .B(n336), .Z(n51) );
  XOR U23 ( .A(a[61]), .B(n327), .Z(n47) );
  XOR U24 ( .A(a[64]), .B(n318), .Z(n44) );
  XOR U25 ( .A(a[67]), .B(n309), .Z(n41) );
  XOR U26 ( .A(a[70]), .B(n300), .Z(n37) );
  XOR U27 ( .A(a[73]), .B(n291), .Z(n34) );
  XOR U28 ( .A(a[76]), .B(n282), .Z(n31) );
  XOR U29 ( .A(a[79]), .B(n273), .Z(n28) );
  XOR U30 ( .A(a[82]), .B(n264), .Z(n24) );
  XOR U31 ( .A(a[85]), .B(n255), .Z(n21) );
  XOR U32 ( .A(a[88]), .B(n246), .Z(n18) );
  XOR U33 ( .A(a[91]), .B(n237), .Z(n14) );
  XOR U34 ( .A(a[94]), .B(n228), .Z(n11) );
  XOR U35 ( .A(a[97]), .B(n219), .Z(n8) );
  XOR U36 ( .A(a[100]), .B(n209), .Z(n211) );
  XOR U37 ( .A(a[103]), .B(n197), .Z(n199) );
  XOR U38 ( .A(a[106]), .B(n185), .Z(n187) );
  XOR U39 ( .A(a[109]), .B(n172), .Z(n174) );
  XOR U40 ( .A(a[112]), .B(n160), .Z(n162) );
  XOR U41 ( .A(a[115]), .B(n148), .Z(n150) );
  XOR U42 ( .A(a[118]), .B(n136), .Z(n138) );
  XOR U43 ( .A(a[121]), .B(n123), .Z(n125) );
  XOR U44 ( .A(a[124]), .B(n111), .Z(n113) );
  XOR U45 ( .A(a[2]), .B(n504), .Z(n82) );
  XOR U46 ( .A(a[5]), .B(n495), .Z(n49) );
  XOR U47 ( .A(a[8]), .B(n486), .Z(n16) );
  XOR U48 ( .A(a[11]), .B(n477), .Z(n134) );
  XOR U49 ( .A(a[14]), .B(n468), .Z(n99) );
  XOR U50 ( .A(a[17]), .B(n459), .Z(n96) );
  XOR U51 ( .A(a[20]), .B(n450), .Z(n92) );
  XOR U52 ( .A(a[23]), .B(n441), .Z(n89) );
  XOR U53 ( .A(a[26]), .B(n432), .Z(n86) );
  XOR U54 ( .A(a[29]), .B(n423), .Z(n83) );
  XOR U55 ( .A(a[32]), .B(n414), .Z(n79) );
  XOR U56 ( .A(a[35]), .B(n405), .Z(n76) );
  XOR U57 ( .A(a[38]), .B(n396), .Z(n73) );
  XOR U58 ( .A(a[41]), .B(n387), .Z(n69) );
  XOR U59 ( .A(a[44]), .B(n378), .Z(n66) );
  XOR U60 ( .A(a[47]), .B(n369), .Z(n63) );
  XOR U61 ( .A(a[50]), .B(n360), .Z(n59) );
  XOR U62 ( .A(a[53]), .B(n351), .Z(n56) );
  XOR U63 ( .A(a[56]), .B(n342), .Z(n53) );
  XOR U64 ( .A(a[59]), .B(n333), .Z(n50) );
  XOR U65 ( .A(a[62]), .B(n324), .Z(n46) );
  XOR U66 ( .A(a[65]), .B(n315), .Z(n43) );
  XOR U67 ( .A(a[68]), .B(n306), .Z(n40) );
  XOR U68 ( .A(a[71]), .B(n297), .Z(n36) );
  XOR U69 ( .A(a[74]), .B(n288), .Z(n33) );
  XOR U70 ( .A(a[77]), .B(n279), .Z(n30) );
  XOR U71 ( .A(a[80]), .B(n270), .Z(n26) );
  XOR U72 ( .A(a[83]), .B(n261), .Z(n23) );
  XOR U73 ( .A(a[86]), .B(n252), .Z(n20) );
  XOR U74 ( .A(a[89]), .B(n243), .Z(n17) );
  XOR U75 ( .A(a[92]), .B(n234), .Z(n13) );
  XOR U76 ( .A(a[95]), .B(n225), .Z(n10) );
  XOR U77 ( .A(a[98]), .B(n216), .Z(n7) );
  XOR U78 ( .A(a[101]), .B(n205), .Z(n207) );
  XOR U79 ( .A(a[104]), .B(n193), .Z(n195) );
  XOR U80 ( .A(a[107]), .B(n181), .Z(n183) );
  XOR U81 ( .A(a[110]), .B(n168), .Z(n170) );
  XOR U82 ( .A(a[113]), .B(n156), .Z(n158) );
  XOR U83 ( .A(a[116]), .B(n144), .Z(n146) );
  XOR U84 ( .A(a[119]), .B(n131), .Z(n133) );
  XOR U85 ( .A(a[122]), .B(n119), .Z(n121) );
  XOR U86 ( .A(a[125]), .B(n107), .Z(n109) );
  XOR U87 ( .A(a[3]), .B(n501), .Z(n71) );
  XOR U88 ( .A(a[6]), .B(n492), .Z(n38) );
  XOR U89 ( .A(a[9]), .B(n483), .Z(n5) );
  XOR U90 ( .A(a[12]), .B(n474), .Z(n101) );
  XOR U91 ( .A(a[15]), .B(n465), .Z(n98) );
  XOR U92 ( .A(a[18]), .B(n456), .Z(n95) );
  XOR U93 ( .A(a[21]), .B(n447), .Z(n91) );
  XOR U94 ( .A(a[24]), .B(n438), .Z(n88) );
  XOR U95 ( .A(a[27]), .B(n429), .Z(n85) );
  XOR U96 ( .A(a[30]), .B(n420), .Z(n81) );
  XOR U97 ( .A(a[33]), .B(n411), .Z(n78) );
  XOR U98 ( .A(a[36]), .B(n402), .Z(n75) );
  XOR U99 ( .A(a[39]), .B(n393), .Z(n72) );
  XOR U100 ( .A(a[42]), .B(n384), .Z(n68) );
  XOR U101 ( .A(a[45]), .B(n375), .Z(n65) );
  XOR U102 ( .A(a[48]), .B(n366), .Z(n62) );
  XOR U103 ( .A(a[51]), .B(n357), .Z(n58) );
  XOR U104 ( .A(a[54]), .B(n348), .Z(n55) );
  XOR U105 ( .A(a[57]), .B(n339), .Z(n52) );
  XOR U106 ( .A(a[60]), .B(n330), .Z(n48) );
  XOR U107 ( .A(a[63]), .B(n321), .Z(n45) );
  XOR U108 ( .A(a[66]), .B(n312), .Z(n42) );
  XOR U109 ( .A(a[69]), .B(n303), .Z(n39) );
  XOR U110 ( .A(a[72]), .B(n294), .Z(n35) );
  XOR U111 ( .A(a[75]), .B(n285), .Z(n32) );
  XOR U112 ( .A(a[78]), .B(n276), .Z(n29) );
  XOR U113 ( .A(a[81]), .B(n267), .Z(n25) );
  XOR U114 ( .A(a[84]), .B(n258), .Z(n22) );
  XOR U115 ( .A(a[87]), .B(n249), .Z(n19) );
  XOR U116 ( .A(a[90]), .B(n240), .Z(n15) );
  XOR U117 ( .A(a[93]), .B(n231), .Z(n12) );
  XOR U118 ( .A(a[96]), .B(n222), .Z(n9) );
  XOR U119 ( .A(a[99]), .B(n213), .Z(n6) );
  XOR U120 ( .A(a[102]), .B(n201), .Z(n203) );
  XOR U121 ( .A(a[105]), .B(n189), .Z(n191) );
  XOR U122 ( .A(a[108]), .B(n177), .Z(n179) );
  XOR U123 ( .A(a[111]), .B(n164), .Z(n166) );
  XOR U124 ( .A(a[114]), .B(n152), .Z(n154) );
  XOR U125 ( .A(a[117]), .B(n140), .Z(n142) );
  XOR U126 ( .A(a[120]), .B(n127), .Z(n129) );
  XOR U127 ( .A(a[123]), .B(n115), .Z(n117) );
  XOR U128 ( .A(a[126]), .B(n103), .Z(n105) );
  XOR U129 ( .A(n1), .B(n2), .Z(carry_on_d) );
  ANDN U130 ( .B(n3), .A(n4), .Z(n1) );
  XOR U131 ( .A(b[127]), .B(n2), .Z(n3) );
  XNOR U132 ( .A(b[9]), .B(n5), .Z(c[9]) );
  XNOR U133 ( .A(b[99]), .B(n6), .Z(c[99]) );
  XNOR U134 ( .A(b[98]), .B(n7), .Z(c[98]) );
  XNOR U135 ( .A(b[97]), .B(n8), .Z(c[97]) );
  XNOR U136 ( .A(b[96]), .B(n9), .Z(c[96]) );
  XNOR U137 ( .A(b[95]), .B(n10), .Z(c[95]) );
  XNOR U138 ( .A(b[94]), .B(n11), .Z(c[94]) );
  XNOR U139 ( .A(b[93]), .B(n12), .Z(c[93]) );
  XNOR U140 ( .A(b[92]), .B(n13), .Z(c[92]) );
  XNOR U141 ( .A(b[91]), .B(n14), .Z(c[91]) );
  XNOR U142 ( .A(b[90]), .B(n15), .Z(c[90]) );
  XNOR U143 ( .A(b[8]), .B(n16), .Z(c[8]) );
  XNOR U144 ( .A(b[89]), .B(n17), .Z(c[89]) );
  XNOR U145 ( .A(b[88]), .B(n18), .Z(c[88]) );
  XNOR U146 ( .A(b[87]), .B(n19), .Z(c[87]) );
  XNOR U147 ( .A(b[86]), .B(n20), .Z(c[86]) );
  XNOR U148 ( .A(b[85]), .B(n21), .Z(c[85]) );
  XNOR U149 ( .A(b[84]), .B(n22), .Z(c[84]) );
  XNOR U150 ( .A(b[83]), .B(n23), .Z(c[83]) );
  XNOR U151 ( .A(b[82]), .B(n24), .Z(c[82]) );
  XNOR U152 ( .A(b[81]), .B(n25), .Z(c[81]) );
  XNOR U153 ( .A(b[80]), .B(n26), .Z(c[80]) );
  XNOR U154 ( .A(b[7]), .B(n27), .Z(c[7]) );
  XNOR U155 ( .A(b[79]), .B(n28), .Z(c[79]) );
  XNOR U156 ( .A(b[78]), .B(n29), .Z(c[78]) );
  XNOR U157 ( .A(b[77]), .B(n30), .Z(c[77]) );
  XNOR U158 ( .A(b[76]), .B(n31), .Z(c[76]) );
  XNOR U159 ( .A(b[75]), .B(n32), .Z(c[75]) );
  XNOR U160 ( .A(b[74]), .B(n33), .Z(c[74]) );
  XNOR U161 ( .A(b[73]), .B(n34), .Z(c[73]) );
  XNOR U162 ( .A(b[72]), .B(n35), .Z(c[72]) );
  XNOR U163 ( .A(b[71]), .B(n36), .Z(c[71]) );
  XNOR U164 ( .A(b[70]), .B(n37), .Z(c[70]) );
  XNOR U165 ( .A(b[6]), .B(n38), .Z(c[6]) );
  XNOR U166 ( .A(b[69]), .B(n39), .Z(c[69]) );
  XNOR U167 ( .A(b[68]), .B(n40), .Z(c[68]) );
  XNOR U168 ( .A(b[67]), .B(n41), .Z(c[67]) );
  XNOR U169 ( .A(b[66]), .B(n42), .Z(c[66]) );
  XNOR U170 ( .A(b[65]), .B(n43), .Z(c[65]) );
  XNOR U171 ( .A(b[64]), .B(n44), .Z(c[64]) );
  XNOR U172 ( .A(b[63]), .B(n45), .Z(c[63]) );
  XNOR U173 ( .A(b[62]), .B(n46), .Z(c[62]) );
  XNOR U174 ( .A(b[61]), .B(n47), .Z(c[61]) );
  XNOR U175 ( .A(b[60]), .B(n48), .Z(c[60]) );
  XNOR U176 ( .A(b[5]), .B(n49), .Z(c[5]) );
  XNOR U177 ( .A(b[59]), .B(n50), .Z(c[59]) );
  XNOR U178 ( .A(b[58]), .B(n51), .Z(c[58]) );
  XNOR U179 ( .A(b[57]), .B(n52), .Z(c[57]) );
  XNOR U180 ( .A(b[56]), .B(n53), .Z(c[56]) );
  XNOR U181 ( .A(b[55]), .B(n54), .Z(c[55]) );
  XNOR U182 ( .A(b[54]), .B(n55), .Z(c[54]) );
  XNOR U183 ( .A(b[53]), .B(n56), .Z(c[53]) );
  XNOR U184 ( .A(b[52]), .B(n57), .Z(c[52]) );
  XNOR U185 ( .A(b[51]), .B(n58), .Z(c[51]) );
  XNOR U186 ( .A(b[50]), .B(n59), .Z(c[50]) );
  XNOR U187 ( .A(b[4]), .B(n60), .Z(c[4]) );
  XNOR U188 ( .A(b[49]), .B(n61), .Z(c[49]) );
  XNOR U189 ( .A(b[48]), .B(n62), .Z(c[48]) );
  XNOR U190 ( .A(b[47]), .B(n63), .Z(c[47]) );
  XNOR U191 ( .A(b[46]), .B(n64), .Z(c[46]) );
  XNOR U192 ( .A(b[45]), .B(n65), .Z(c[45]) );
  XNOR U193 ( .A(b[44]), .B(n66), .Z(c[44]) );
  XNOR U194 ( .A(b[43]), .B(n67), .Z(c[43]) );
  XNOR U195 ( .A(b[42]), .B(n68), .Z(c[42]) );
  XNOR U196 ( .A(b[41]), .B(n69), .Z(c[41]) );
  XNOR U197 ( .A(b[40]), .B(n70), .Z(c[40]) );
  XNOR U198 ( .A(b[3]), .B(n71), .Z(c[3]) );
  XNOR U199 ( .A(b[39]), .B(n72), .Z(c[39]) );
  XNOR U200 ( .A(b[38]), .B(n73), .Z(c[38]) );
  XNOR U201 ( .A(b[37]), .B(n74), .Z(c[37]) );
  XNOR U202 ( .A(b[36]), .B(n75), .Z(c[36]) );
  XNOR U203 ( .A(b[35]), .B(n76), .Z(c[35]) );
  XNOR U204 ( .A(b[34]), .B(n77), .Z(c[34]) );
  XNOR U205 ( .A(b[33]), .B(n78), .Z(c[33]) );
  XNOR U206 ( .A(b[32]), .B(n79), .Z(c[32]) );
  XNOR U207 ( .A(b[31]), .B(n80), .Z(c[31]) );
  XNOR U208 ( .A(b[30]), .B(n81), .Z(c[30]) );
  XNOR U209 ( .A(b[2]), .B(n82), .Z(c[2]) );
  XNOR U210 ( .A(b[29]), .B(n83), .Z(c[29]) );
  XNOR U211 ( .A(b[28]), .B(n84), .Z(c[28]) );
  XNOR U212 ( .A(b[27]), .B(n85), .Z(c[27]) );
  XNOR U213 ( .A(b[26]), .B(n86), .Z(c[26]) );
  XNOR U214 ( .A(b[25]), .B(n87), .Z(c[25]) );
  XNOR U215 ( .A(b[24]), .B(n88), .Z(c[24]) );
  XNOR U216 ( .A(b[23]), .B(n89), .Z(c[23]) );
  XNOR U217 ( .A(b[22]), .B(n90), .Z(c[22]) );
  XNOR U218 ( .A(b[21]), .B(n91), .Z(c[21]) );
  XNOR U219 ( .A(b[20]), .B(n92), .Z(c[20]) );
  XNOR U220 ( .A(b[1]), .B(n93), .Z(c[1]) );
  XNOR U221 ( .A(b[19]), .B(n94), .Z(c[19]) );
  XNOR U222 ( .A(b[18]), .B(n95), .Z(c[18]) );
  XNOR U223 ( .A(b[17]), .B(n96), .Z(c[17]) );
  XNOR U224 ( .A(b[16]), .B(n97), .Z(c[16]) );
  XNOR U225 ( .A(b[15]), .B(n98), .Z(c[15]) );
  XNOR U226 ( .A(b[14]), .B(n99), .Z(c[14]) );
  XNOR U227 ( .A(b[13]), .B(n100), .Z(c[13]) );
  XNOR U228 ( .A(b[12]), .B(n101), .Z(c[12]) );
  XNOR U229 ( .A(b[127]), .B(n4), .Z(c[127]) );
  XNOR U230 ( .A(a[127]), .B(n2), .Z(n4) );
  XNOR U231 ( .A(n102), .B(n103), .Z(n2) );
  ANDN U232 ( .B(n104), .A(n105), .Z(n102) );
  XNOR U233 ( .A(b[126]), .B(n103), .Z(n104) );
  XNOR U234 ( .A(b[126]), .B(n105), .Z(c[126]) );
  XOR U235 ( .A(n106), .B(n107), .Z(n103) );
  ANDN U236 ( .B(n108), .A(n109), .Z(n106) );
  XNOR U237 ( .A(b[125]), .B(n107), .Z(n108) );
  XNOR U238 ( .A(b[125]), .B(n109), .Z(c[125]) );
  XOR U239 ( .A(n110), .B(n111), .Z(n107) );
  ANDN U240 ( .B(n112), .A(n113), .Z(n110) );
  XNOR U241 ( .A(b[124]), .B(n111), .Z(n112) );
  XNOR U242 ( .A(b[124]), .B(n113), .Z(c[124]) );
  XOR U243 ( .A(n114), .B(n115), .Z(n111) );
  ANDN U244 ( .B(n116), .A(n117), .Z(n114) );
  XNOR U245 ( .A(b[123]), .B(n115), .Z(n116) );
  XNOR U246 ( .A(b[123]), .B(n117), .Z(c[123]) );
  XOR U247 ( .A(n118), .B(n119), .Z(n115) );
  ANDN U248 ( .B(n120), .A(n121), .Z(n118) );
  XNOR U249 ( .A(b[122]), .B(n119), .Z(n120) );
  XNOR U250 ( .A(b[122]), .B(n121), .Z(c[122]) );
  XOR U251 ( .A(n122), .B(n123), .Z(n119) );
  ANDN U252 ( .B(n124), .A(n125), .Z(n122) );
  XNOR U253 ( .A(b[121]), .B(n123), .Z(n124) );
  XNOR U254 ( .A(b[121]), .B(n125), .Z(c[121]) );
  XOR U255 ( .A(n126), .B(n127), .Z(n123) );
  ANDN U256 ( .B(n128), .A(n129), .Z(n126) );
  XNOR U257 ( .A(b[120]), .B(n127), .Z(n128) );
  XNOR U258 ( .A(b[120]), .B(n129), .Z(c[120]) );
  XOR U259 ( .A(n130), .B(n131), .Z(n127) );
  ANDN U260 ( .B(n132), .A(n133), .Z(n130) );
  XNOR U261 ( .A(b[119]), .B(n131), .Z(n132) );
  XNOR U262 ( .A(b[11]), .B(n134), .Z(c[11]) );
  XNOR U263 ( .A(b[119]), .B(n133), .Z(c[119]) );
  XOR U264 ( .A(n135), .B(n136), .Z(n131) );
  ANDN U265 ( .B(n137), .A(n138), .Z(n135) );
  XNOR U266 ( .A(b[118]), .B(n136), .Z(n137) );
  XNOR U267 ( .A(b[118]), .B(n138), .Z(c[118]) );
  XOR U268 ( .A(n139), .B(n140), .Z(n136) );
  ANDN U269 ( .B(n141), .A(n142), .Z(n139) );
  XNOR U270 ( .A(b[117]), .B(n140), .Z(n141) );
  XNOR U271 ( .A(b[117]), .B(n142), .Z(c[117]) );
  XOR U272 ( .A(n143), .B(n144), .Z(n140) );
  ANDN U273 ( .B(n145), .A(n146), .Z(n143) );
  XNOR U274 ( .A(b[116]), .B(n144), .Z(n145) );
  XNOR U275 ( .A(b[116]), .B(n146), .Z(c[116]) );
  XOR U276 ( .A(n147), .B(n148), .Z(n144) );
  ANDN U277 ( .B(n149), .A(n150), .Z(n147) );
  XNOR U278 ( .A(b[115]), .B(n148), .Z(n149) );
  XNOR U279 ( .A(b[115]), .B(n150), .Z(c[115]) );
  XOR U280 ( .A(n151), .B(n152), .Z(n148) );
  ANDN U281 ( .B(n153), .A(n154), .Z(n151) );
  XNOR U282 ( .A(b[114]), .B(n152), .Z(n153) );
  XNOR U283 ( .A(b[114]), .B(n154), .Z(c[114]) );
  XOR U284 ( .A(n155), .B(n156), .Z(n152) );
  ANDN U285 ( .B(n157), .A(n158), .Z(n155) );
  XNOR U286 ( .A(b[113]), .B(n156), .Z(n157) );
  XNOR U287 ( .A(b[113]), .B(n158), .Z(c[113]) );
  XOR U288 ( .A(n159), .B(n160), .Z(n156) );
  ANDN U289 ( .B(n161), .A(n162), .Z(n159) );
  XNOR U290 ( .A(b[112]), .B(n160), .Z(n161) );
  XNOR U291 ( .A(b[112]), .B(n162), .Z(c[112]) );
  XOR U292 ( .A(n163), .B(n164), .Z(n160) );
  ANDN U293 ( .B(n165), .A(n166), .Z(n163) );
  XNOR U294 ( .A(b[111]), .B(n164), .Z(n165) );
  XNOR U295 ( .A(b[111]), .B(n166), .Z(c[111]) );
  XOR U296 ( .A(n167), .B(n168), .Z(n164) );
  ANDN U297 ( .B(n169), .A(n170), .Z(n167) );
  XNOR U298 ( .A(b[110]), .B(n168), .Z(n169) );
  XNOR U299 ( .A(b[110]), .B(n170), .Z(c[110]) );
  XOR U300 ( .A(n171), .B(n172), .Z(n168) );
  ANDN U301 ( .B(n173), .A(n174), .Z(n171) );
  XNOR U302 ( .A(b[109]), .B(n172), .Z(n173) );
  XNOR U303 ( .A(b[10]), .B(n175), .Z(c[10]) );
  XNOR U304 ( .A(b[109]), .B(n174), .Z(c[109]) );
  XOR U305 ( .A(n176), .B(n177), .Z(n172) );
  ANDN U306 ( .B(n178), .A(n179), .Z(n176) );
  XNOR U307 ( .A(b[108]), .B(n177), .Z(n178) );
  XNOR U308 ( .A(b[108]), .B(n179), .Z(c[108]) );
  XOR U309 ( .A(n180), .B(n181), .Z(n177) );
  ANDN U310 ( .B(n182), .A(n183), .Z(n180) );
  XNOR U311 ( .A(b[107]), .B(n181), .Z(n182) );
  XNOR U312 ( .A(b[107]), .B(n183), .Z(c[107]) );
  XOR U313 ( .A(n184), .B(n185), .Z(n181) );
  ANDN U314 ( .B(n186), .A(n187), .Z(n184) );
  XNOR U315 ( .A(b[106]), .B(n185), .Z(n186) );
  XNOR U316 ( .A(b[106]), .B(n187), .Z(c[106]) );
  XOR U317 ( .A(n188), .B(n189), .Z(n185) );
  ANDN U318 ( .B(n190), .A(n191), .Z(n188) );
  XNOR U319 ( .A(b[105]), .B(n189), .Z(n190) );
  XNOR U320 ( .A(b[105]), .B(n191), .Z(c[105]) );
  XOR U321 ( .A(n192), .B(n193), .Z(n189) );
  ANDN U322 ( .B(n194), .A(n195), .Z(n192) );
  XNOR U323 ( .A(b[104]), .B(n193), .Z(n194) );
  XNOR U324 ( .A(b[104]), .B(n195), .Z(c[104]) );
  XOR U325 ( .A(n196), .B(n197), .Z(n193) );
  ANDN U326 ( .B(n198), .A(n199), .Z(n196) );
  XNOR U327 ( .A(b[103]), .B(n197), .Z(n198) );
  XNOR U328 ( .A(b[103]), .B(n199), .Z(c[103]) );
  XOR U329 ( .A(n200), .B(n201), .Z(n197) );
  ANDN U330 ( .B(n202), .A(n203), .Z(n200) );
  XNOR U331 ( .A(b[102]), .B(n201), .Z(n202) );
  XNOR U332 ( .A(b[102]), .B(n203), .Z(c[102]) );
  XOR U333 ( .A(n204), .B(n205), .Z(n201) );
  ANDN U334 ( .B(n206), .A(n207), .Z(n204) );
  XNOR U335 ( .A(b[101]), .B(n205), .Z(n206) );
  XNOR U336 ( .A(b[101]), .B(n207), .Z(c[101]) );
  XOR U337 ( .A(n208), .B(n209), .Z(n205) );
  ANDN U338 ( .B(n210), .A(n211), .Z(n208) );
  XNOR U339 ( .A(b[100]), .B(n209), .Z(n210) );
  XNOR U340 ( .A(b[100]), .B(n211), .Z(c[100]) );
  XOR U341 ( .A(n212), .B(n213), .Z(n209) );
  ANDN U342 ( .B(n214), .A(n6), .Z(n212) );
  XNOR U343 ( .A(b[99]), .B(n213), .Z(n214) );
  XOR U344 ( .A(n215), .B(n216), .Z(n213) );
  ANDN U345 ( .B(n217), .A(n7), .Z(n215) );
  XNOR U346 ( .A(b[98]), .B(n216), .Z(n217) );
  XOR U347 ( .A(n218), .B(n219), .Z(n216) );
  ANDN U348 ( .B(n220), .A(n8), .Z(n218) );
  XNOR U349 ( .A(b[97]), .B(n219), .Z(n220) );
  XOR U350 ( .A(n221), .B(n222), .Z(n219) );
  ANDN U351 ( .B(n223), .A(n9), .Z(n221) );
  XNOR U352 ( .A(b[96]), .B(n222), .Z(n223) );
  XOR U353 ( .A(n224), .B(n225), .Z(n222) );
  ANDN U354 ( .B(n226), .A(n10), .Z(n224) );
  XNOR U355 ( .A(b[95]), .B(n225), .Z(n226) );
  XOR U356 ( .A(n227), .B(n228), .Z(n225) );
  ANDN U357 ( .B(n229), .A(n11), .Z(n227) );
  XNOR U358 ( .A(b[94]), .B(n228), .Z(n229) );
  XOR U359 ( .A(n230), .B(n231), .Z(n228) );
  ANDN U360 ( .B(n232), .A(n12), .Z(n230) );
  XNOR U361 ( .A(b[93]), .B(n231), .Z(n232) );
  XOR U362 ( .A(n233), .B(n234), .Z(n231) );
  ANDN U363 ( .B(n235), .A(n13), .Z(n233) );
  XNOR U364 ( .A(b[92]), .B(n234), .Z(n235) );
  XOR U365 ( .A(n236), .B(n237), .Z(n234) );
  ANDN U366 ( .B(n238), .A(n14), .Z(n236) );
  XNOR U367 ( .A(b[91]), .B(n237), .Z(n238) );
  XOR U368 ( .A(n239), .B(n240), .Z(n237) );
  ANDN U369 ( .B(n241), .A(n15), .Z(n239) );
  XNOR U370 ( .A(b[90]), .B(n240), .Z(n241) );
  XOR U371 ( .A(n242), .B(n243), .Z(n240) );
  ANDN U372 ( .B(n244), .A(n17), .Z(n242) );
  XNOR U373 ( .A(b[89]), .B(n243), .Z(n244) );
  XOR U374 ( .A(n245), .B(n246), .Z(n243) );
  ANDN U375 ( .B(n247), .A(n18), .Z(n245) );
  XNOR U376 ( .A(b[88]), .B(n246), .Z(n247) );
  XOR U377 ( .A(n248), .B(n249), .Z(n246) );
  ANDN U378 ( .B(n250), .A(n19), .Z(n248) );
  XNOR U379 ( .A(b[87]), .B(n249), .Z(n250) );
  XOR U380 ( .A(n251), .B(n252), .Z(n249) );
  ANDN U381 ( .B(n253), .A(n20), .Z(n251) );
  XNOR U382 ( .A(b[86]), .B(n252), .Z(n253) );
  XOR U383 ( .A(n254), .B(n255), .Z(n252) );
  ANDN U384 ( .B(n256), .A(n21), .Z(n254) );
  XNOR U385 ( .A(b[85]), .B(n255), .Z(n256) );
  XOR U386 ( .A(n257), .B(n258), .Z(n255) );
  ANDN U387 ( .B(n259), .A(n22), .Z(n257) );
  XNOR U388 ( .A(b[84]), .B(n258), .Z(n259) );
  XOR U389 ( .A(n260), .B(n261), .Z(n258) );
  ANDN U390 ( .B(n262), .A(n23), .Z(n260) );
  XNOR U391 ( .A(b[83]), .B(n261), .Z(n262) );
  XOR U392 ( .A(n263), .B(n264), .Z(n261) );
  ANDN U393 ( .B(n265), .A(n24), .Z(n263) );
  XNOR U394 ( .A(b[82]), .B(n264), .Z(n265) );
  XOR U395 ( .A(n266), .B(n267), .Z(n264) );
  ANDN U396 ( .B(n268), .A(n25), .Z(n266) );
  XNOR U397 ( .A(b[81]), .B(n267), .Z(n268) );
  XOR U398 ( .A(n269), .B(n270), .Z(n267) );
  ANDN U399 ( .B(n271), .A(n26), .Z(n269) );
  XNOR U400 ( .A(b[80]), .B(n270), .Z(n271) );
  XOR U401 ( .A(n272), .B(n273), .Z(n270) );
  ANDN U402 ( .B(n274), .A(n28), .Z(n272) );
  XNOR U403 ( .A(b[79]), .B(n273), .Z(n274) );
  XOR U404 ( .A(n275), .B(n276), .Z(n273) );
  ANDN U405 ( .B(n277), .A(n29), .Z(n275) );
  XNOR U406 ( .A(b[78]), .B(n276), .Z(n277) );
  XOR U407 ( .A(n278), .B(n279), .Z(n276) );
  ANDN U408 ( .B(n280), .A(n30), .Z(n278) );
  XNOR U409 ( .A(b[77]), .B(n279), .Z(n280) );
  XOR U410 ( .A(n281), .B(n282), .Z(n279) );
  ANDN U411 ( .B(n283), .A(n31), .Z(n281) );
  XNOR U412 ( .A(b[76]), .B(n282), .Z(n283) );
  XOR U413 ( .A(n284), .B(n285), .Z(n282) );
  ANDN U414 ( .B(n286), .A(n32), .Z(n284) );
  XNOR U415 ( .A(b[75]), .B(n285), .Z(n286) );
  XOR U416 ( .A(n287), .B(n288), .Z(n285) );
  ANDN U417 ( .B(n289), .A(n33), .Z(n287) );
  XNOR U418 ( .A(b[74]), .B(n288), .Z(n289) );
  XOR U419 ( .A(n290), .B(n291), .Z(n288) );
  ANDN U420 ( .B(n292), .A(n34), .Z(n290) );
  XNOR U421 ( .A(b[73]), .B(n291), .Z(n292) );
  XOR U422 ( .A(n293), .B(n294), .Z(n291) );
  ANDN U423 ( .B(n295), .A(n35), .Z(n293) );
  XNOR U424 ( .A(b[72]), .B(n294), .Z(n295) );
  XOR U425 ( .A(n296), .B(n297), .Z(n294) );
  ANDN U426 ( .B(n298), .A(n36), .Z(n296) );
  XNOR U427 ( .A(b[71]), .B(n297), .Z(n298) );
  XOR U428 ( .A(n299), .B(n300), .Z(n297) );
  ANDN U429 ( .B(n301), .A(n37), .Z(n299) );
  XNOR U430 ( .A(b[70]), .B(n300), .Z(n301) );
  XOR U431 ( .A(n302), .B(n303), .Z(n300) );
  ANDN U432 ( .B(n304), .A(n39), .Z(n302) );
  XNOR U433 ( .A(b[69]), .B(n303), .Z(n304) );
  XOR U434 ( .A(n305), .B(n306), .Z(n303) );
  ANDN U435 ( .B(n307), .A(n40), .Z(n305) );
  XNOR U436 ( .A(b[68]), .B(n306), .Z(n307) );
  XOR U437 ( .A(n308), .B(n309), .Z(n306) );
  ANDN U438 ( .B(n310), .A(n41), .Z(n308) );
  XNOR U439 ( .A(b[67]), .B(n309), .Z(n310) );
  XOR U440 ( .A(n311), .B(n312), .Z(n309) );
  ANDN U441 ( .B(n313), .A(n42), .Z(n311) );
  XNOR U442 ( .A(b[66]), .B(n312), .Z(n313) );
  XOR U443 ( .A(n314), .B(n315), .Z(n312) );
  ANDN U444 ( .B(n316), .A(n43), .Z(n314) );
  XNOR U445 ( .A(b[65]), .B(n315), .Z(n316) );
  XOR U446 ( .A(n317), .B(n318), .Z(n315) );
  ANDN U447 ( .B(n319), .A(n44), .Z(n317) );
  XNOR U448 ( .A(b[64]), .B(n318), .Z(n319) );
  XOR U449 ( .A(n320), .B(n321), .Z(n318) );
  ANDN U450 ( .B(n322), .A(n45), .Z(n320) );
  XNOR U451 ( .A(b[63]), .B(n321), .Z(n322) );
  XOR U452 ( .A(n323), .B(n324), .Z(n321) );
  ANDN U453 ( .B(n325), .A(n46), .Z(n323) );
  XNOR U454 ( .A(b[62]), .B(n324), .Z(n325) );
  XOR U455 ( .A(n326), .B(n327), .Z(n324) );
  ANDN U456 ( .B(n328), .A(n47), .Z(n326) );
  XNOR U457 ( .A(b[61]), .B(n327), .Z(n328) );
  XOR U458 ( .A(n329), .B(n330), .Z(n327) );
  ANDN U459 ( .B(n331), .A(n48), .Z(n329) );
  XNOR U460 ( .A(b[60]), .B(n330), .Z(n331) );
  XOR U461 ( .A(n332), .B(n333), .Z(n330) );
  ANDN U462 ( .B(n334), .A(n50), .Z(n332) );
  XNOR U463 ( .A(b[59]), .B(n333), .Z(n334) );
  XOR U464 ( .A(n335), .B(n336), .Z(n333) );
  ANDN U465 ( .B(n337), .A(n51), .Z(n335) );
  XNOR U466 ( .A(b[58]), .B(n336), .Z(n337) );
  XOR U467 ( .A(n338), .B(n339), .Z(n336) );
  ANDN U468 ( .B(n340), .A(n52), .Z(n338) );
  XNOR U469 ( .A(b[57]), .B(n339), .Z(n340) );
  XOR U470 ( .A(n341), .B(n342), .Z(n339) );
  ANDN U471 ( .B(n343), .A(n53), .Z(n341) );
  XNOR U472 ( .A(b[56]), .B(n342), .Z(n343) );
  XOR U473 ( .A(n344), .B(n345), .Z(n342) );
  ANDN U474 ( .B(n346), .A(n54), .Z(n344) );
  XNOR U475 ( .A(b[55]), .B(n345), .Z(n346) );
  XOR U476 ( .A(n347), .B(n348), .Z(n345) );
  ANDN U477 ( .B(n349), .A(n55), .Z(n347) );
  XNOR U478 ( .A(b[54]), .B(n348), .Z(n349) );
  XOR U479 ( .A(n350), .B(n351), .Z(n348) );
  ANDN U480 ( .B(n352), .A(n56), .Z(n350) );
  XNOR U481 ( .A(b[53]), .B(n351), .Z(n352) );
  XOR U482 ( .A(n353), .B(n354), .Z(n351) );
  ANDN U483 ( .B(n355), .A(n57), .Z(n353) );
  XNOR U484 ( .A(b[52]), .B(n354), .Z(n355) );
  XOR U485 ( .A(n356), .B(n357), .Z(n354) );
  ANDN U486 ( .B(n358), .A(n58), .Z(n356) );
  XNOR U487 ( .A(b[51]), .B(n357), .Z(n358) );
  XOR U488 ( .A(n359), .B(n360), .Z(n357) );
  ANDN U489 ( .B(n361), .A(n59), .Z(n359) );
  XNOR U490 ( .A(b[50]), .B(n360), .Z(n361) );
  XOR U491 ( .A(n362), .B(n363), .Z(n360) );
  ANDN U492 ( .B(n364), .A(n61), .Z(n362) );
  XNOR U493 ( .A(b[49]), .B(n363), .Z(n364) );
  XOR U494 ( .A(n365), .B(n366), .Z(n363) );
  ANDN U495 ( .B(n367), .A(n62), .Z(n365) );
  XNOR U496 ( .A(b[48]), .B(n366), .Z(n367) );
  XOR U497 ( .A(n368), .B(n369), .Z(n366) );
  ANDN U498 ( .B(n370), .A(n63), .Z(n368) );
  XNOR U499 ( .A(b[47]), .B(n369), .Z(n370) );
  XOR U500 ( .A(n371), .B(n372), .Z(n369) );
  ANDN U501 ( .B(n373), .A(n64), .Z(n371) );
  XNOR U502 ( .A(b[46]), .B(n372), .Z(n373) );
  XOR U503 ( .A(n374), .B(n375), .Z(n372) );
  ANDN U504 ( .B(n376), .A(n65), .Z(n374) );
  XNOR U505 ( .A(b[45]), .B(n375), .Z(n376) );
  XOR U506 ( .A(n377), .B(n378), .Z(n375) );
  ANDN U507 ( .B(n379), .A(n66), .Z(n377) );
  XNOR U508 ( .A(b[44]), .B(n378), .Z(n379) );
  XOR U509 ( .A(n380), .B(n381), .Z(n378) );
  ANDN U510 ( .B(n382), .A(n67), .Z(n380) );
  XNOR U511 ( .A(b[43]), .B(n381), .Z(n382) );
  XOR U512 ( .A(n383), .B(n384), .Z(n381) );
  ANDN U513 ( .B(n385), .A(n68), .Z(n383) );
  XNOR U514 ( .A(b[42]), .B(n384), .Z(n385) );
  XOR U515 ( .A(n386), .B(n387), .Z(n384) );
  ANDN U516 ( .B(n388), .A(n69), .Z(n386) );
  XNOR U517 ( .A(b[41]), .B(n387), .Z(n388) );
  XOR U518 ( .A(n389), .B(n390), .Z(n387) );
  ANDN U519 ( .B(n391), .A(n70), .Z(n389) );
  XNOR U520 ( .A(b[40]), .B(n390), .Z(n391) );
  XOR U521 ( .A(n392), .B(n393), .Z(n390) );
  ANDN U522 ( .B(n394), .A(n72), .Z(n392) );
  XNOR U523 ( .A(b[39]), .B(n393), .Z(n394) );
  XOR U524 ( .A(n395), .B(n396), .Z(n393) );
  ANDN U525 ( .B(n397), .A(n73), .Z(n395) );
  XNOR U526 ( .A(b[38]), .B(n396), .Z(n397) );
  XOR U527 ( .A(n398), .B(n399), .Z(n396) );
  ANDN U528 ( .B(n400), .A(n74), .Z(n398) );
  XNOR U529 ( .A(b[37]), .B(n399), .Z(n400) );
  XOR U530 ( .A(n401), .B(n402), .Z(n399) );
  ANDN U531 ( .B(n403), .A(n75), .Z(n401) );
  XNOR U532 ( .A(b[36]), .B(n402), .Z(n403) );
  XOR U533 ( .A(n404), .B(n405), .Z(n402) );
  ANDN U534 ( .B(n406), .A(n76), .Z(n404) );
  XNOR U535 ( .A(b[35]), .B(n405), .Z(n406) );
  XOR U536 ( .A(n407), .B(n408), .Z(n405) );
  ANDN U537 ( .B(n409), .A(n77), .Z(n407) );
  XNOR U538 ( .A(b[34]), .B(n408), .Z(n409) );
  XOR U539 ( .A(n410), .B(n411), .Z(n408) );
  ANDN U540 ( .B(n412), .A(n78), .Z(n410) );
  XNOR U541 ( .A(b[33]), .B(n411), .Z(n412) );
  XOR U542 ( .A(n413), .B(n414), .Z(n411) );
  ANDN U543 ( .B(n415), .A(n79), .Z(n413) );
  XNOR U544 ( .A(b[32]), .B(n414), .Z(n415) );
  XOR U545 ( .A(n416), .B(n417), .Z(n414) );
  ANDN U546 ( .B(n418), .A(n80), .Z(n416) );
  XNOR U547 ( .A(b[31]), .B(n417), .Z(n418) );
  XOR U548 ( .A(n419), .B(n420), .Z(n417) );
  ANDN U549 ( .B(n421), .A(n81), .Z(n419) );
  XNOR U550 ( .A(b[30]), .B(n420), .Z(n421) );
  XOR U551 ( .A(n422), .B(n423), .Z(n420) );
  ANDN U552 ( .B(n424), .A(n83), .Z(n422) );
  XNOR U553 ( .A(b[29]), .B(n423), .Z(n424) );
  XOR U554 ( .A(n425), .B(n426), .Z(n423) );
  ANDN U555 ( .B(n427), .A(n84), .Z(n425) );
  XNOR U556 ( .A(b[28]), .B(n426), .Z(n427) );
  XOR U557 ( .A(n428), .B(n429), .Z(n426) );
  ANDN U558 ( .B(n430), .A(n85), .Z(n428) );
  XNOR U559 ( .A(b[27]), .B(n429), .Z(n430) );
  XOR U560 ( .A(n431), .B(n432), .Z(n429) );
  ANDN U561 ( .B(n433), .A(n86), .Z(n431) );
  XNOR U562 ( .A(b[26]), .B(n432), .Z(n433) );
  XOR U563 ( .A(n434), .B(n435), .Z(n432) );
  ANDN U564 ( .B(n436), .A(n87), .Z(n434) );
  XNOR U565 ( .A(b[25]), .B(n435), .Z(n436) );
  XOR U566 ( .A(n437), .B(n438), .Z(n435) );
  ANDN U567 ( .B(n439), .A(n88), .Z(n437) );
  XNOR U568 ( .A(b[24]), .B(n438), .Z(n439) );
  XOR U569 ( .A(n440), .B(n441), .Z(n438) );
  ANDN U570 ( .B(n442), .A(n89), .Z(n440) );
  XNOR U571 ( .A(b[23]), .B(n441), .Z(n442) );
  XOR U572 ( .A(n443), .B(n444), .Z(n441) );
  ANDN U573 ( .B(n445), .A(n90), .Z(n443) );
  XNOR U574 ( .A(b[22]), .B(n444), .Z(n445) );
  XOR U575 ( .A(n446), .B(n447), .Z(n444) );
  ANDN U576 ( .B(n448), .A(n91), .Z(n446) );
  XNOR U577 ( .A(b[21]), .B(n447), .Z(n448) );
  XOR U578 ( .A(n449), .B(n450), .Z(n447) );
  ANDN U579 ( .B(n451), .A(n92), .Z(n449) );
  XNOR U580 ( .A(b[20]), .B(n450), .Z(n451) );
  XOR U581 ( .A(n452), .B(n453), .Z(n450) );
  ANDN U582 ( .B(n454), .A(n94), .Z(n452) );
  XNOR U583 ( .A(b[19]), .B(n453), .Z(n454) );
  XOR U584 ( .A(n455), .B(n456), .Z(n453) );
  ANDN U585 ( .B(n457), .A(n95), .Z(n455) );
  XNOR U586 ( .A(b[18]), .B(n456), .Z(n457) );
  XOR U587 ( .A(n458), .B(n459), .Z(n456) );
  ANDN U588 ( .B(n460), .A(n96), .Z(n458) );
  XNOR U589 ( .A(b[17]), .B(n459), .Z(n460) );
  XOR U590 ( .A(n461), .B(n462), .Z(n459) );
  ANDN U591 ( .B(n463), .A(n97), .Z(n461) );
  XNOR U592 ( .A(b[16]), .B(n462), .Z(n463) );
  XOR U593 ( .A(n464), .B(n465), .Z(n462) );
  ANDN U594 ( .B(n466), .A(n98), .Z(n464) );
  XNOR U595 ( .A(b[15]), .B(n465), .Z(n466) );
  XOR U596 ( .A(n467), .B(n468), .Z(n465) );
  ANDN U597 ( .B(n469), .A(n99), .Z(n467) );
  XNOR U598 ( .A(b[14]), .B(n468), .Z(n469) );
  XOR U599 ( .A(n470), .B(n471), .Z(n468) );
  ANDN U600 ( .B(n472), .A(n100), .Z(n470) );
  XNOR U601 ( .A(b[13]), .B(n471), .Z(n472) );
  XOR U602 ( .A(n473), .B(n474), .Z(n471) );
  ANDN U603 ( .B(n475), .A(n101), .Z(n473) );
  XNOR U604 ( .A(b[12]), .B(n474), .Z(n475) );
  XOR U605 ( .A(n476), .B(n477), .Z(n474) );
  ANDN U606 ( .B(n478), .A(n134), .Z(n476) );
  XNOR U607 ( .A(b[11]), .B(n477), .Z(n478) );
  XOR U608 ( .A(n479), .B(n480), .Z(n477) );
  ANDN U609 ( .B(n481), .A(n175), .Z(n479) );
  XNOR U610 ( .A(b[10]), .B(n480), .Z(n481) );
  XOR U611 ( .A(n482), .B(n483), .Z(n480) );
  ANDN U612 ( .B(n484), .A(n5), .Z(n482) );
  XNOR U613 ( .A(b[9]), .B(n483), .Z(n484) );
  XOR U614 ( .A(n485), .B(n486), .Z(n483) );
  ANDN U615 ( .B(n487), .A(n16), .Z(n485) );
  XNOR U616 ( .A(b[8]), .B(n486), .Z(n487) );
  XOR U617 ( .A(n488), .B(n489), .Z(n486) );
  ANDN U618 ( .B(n490), .A(n27), .Z(n488) );
  XNOR U619 ( .A(b[7]), .B(n489), .Z(n490) );
  XOR U620 ( .A(n491), .B(n492), .Z(n489) );
  ANDN U621 ( .B(n493), .A(n38), .Z(n491) );
  XNOR U622 ( .A(b[6]), .B(n492), .Z(n493) );
  XOR U623 ( .A(n494), .B(n495), .Z(n492) );
  ANDN U624 ( .B(n496), .A(n49), .Z(n494) );
  XNOR U625 ( .A(b[5]), .B(n495), .Z(n496) );
  XOR U626 ( .A(n497), .B(n498), .Z(n495) );
  ANDN U627 ( .B(n499), .A(n60), .Z(n497) );
  XNOR U628 ( .A(b[4]), .B(n498), .Z(n499) );
  XOR U629 ( .A(n500), .B(n501), .Z(n498) );
  ANDN U630 ( .B(n502), .A(n71), .Z(n500) );
  XNOR U631 ( .A(b[3]), .B(n501), .Z(n502) );
  XOR U632 ( .A(n503), .B(n504), .Z(n501) );
  ANDN U633 ( .B(n505), .A(n82), .Z(n503) );
  XNOR U634 ( .A(b[2]), .B(n504), .Z(n505) );
  XOR U635 ( .A(n506), .B(n507), .Z(n504) );
  ANDN U636 ( .B(n508), .A(n93), .Z(n506) );
  XNOR U637 ( .A(b[1]), .B(n507), .Z(n508) );
  XOR U638 ( .A(carry_on), .B(n509), .Z(n507) );
  NANDN U639 ( .A(n510), .B(n511), .Z(n509) );
  XOR U640 ( .A(carry_on), .B(b[0]), .Z(n511) );
  XNOR U641 ( .A(b[0]), .B(n510), .Z(c[0]) );
  XNOR U642 ( .A(a[0]), .B(carry_on), .Z(n510) );
endmodule

