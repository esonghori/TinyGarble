
module hamming_N16000_CC64 ( clk, rst, x, y, o );
  input [249:0] x;
  input [249:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U253 ( .A(n1065), .B(n1064), .Z(n1) );
  NAND U254 ( .A(n1062), .B(n1063), .Z(n2) );
  AND U255 ( .A(n1), .B(n2), .Z(n1084) );
  NAND U256 ( .A(n540), .B(n539), .Z(n3) );
  NAND U257 ( .A(n537), .B(n538), .Z(n4) );
  AND U258 ( .A(n3), .B(n4), .Z(n1198) );
  XNOR U259 ( .A(n1150), .B(n1149), .Z(n1121) );
  NAND U260 ( .A(n958), .B(n959), .Z(n5) );
  XOR U261 ( .A(n958), .B(n959), .Z(n6) );
  NANDN U262 ( .A(n957), .B(n6), .Z(n7) );
  NAND U263 ( .A(n5), .B(n7), .Z(n1342) );
  NAND U264 ( .A(n971), .B(n972), .Z(n8) );
  XOR U265 ( .A(n971), .B(n972), .Z(n9) );
  NANDN U266 ( .A(n970), .B(n9), .Z(n10) );
  NAND U267 ( .A(n8), .B(n10), .Z(n1116) );
  NAND U268 ( .A(n744), .B(n746), .Z(n11) );
  XOR U269 ( .A(n744), .B(n746), .Z(n12) );
  NAND U270 ( .A(n12), .B(n745), .Z(n13) );
  NAND U271 ( .A(n11), .B(n13), .Z(n1291) );
  NAND U272 ( .A(n1118), .B(n1120), .Z(n14) );
  XOR U273 ( .A(n1118), .B(n1120), .Z(n15) );
  NAND U274 ( .A(n15), .B(n1119), .Z(n16) );
  NAND U275 ( .A(n14), .B(n16), .Z(n1502) );
  NAND U276 ( .A(n1088), .B(n1089), .Z(n17) );
  XOR U277 ( .A(n1088), .B(n1089), .Z(n18) );
  NANDN U278 ( .A(n1087), .B(n18), .Z(n19) );
  NAND U279 ( .A(n17), .B(n19), .Z(n1424) );
  NAND U280 ( .A(n1249), .B(n1250), .Z(n20) );
  XOR U281 ( .A(n1249), .B(n1250), .Z(n21) );
  NANDN U282 ( .A(n1248), .B(n21), .Z(n22) );
  NAND U283 ( .A(n20), .B(n22), .Z(n1414) );
  NAND U284 ( .A(n1226), .B(n1227), .Z(n23) );
  XOR U285 ( .A(n1226), .B(n1227), .Z(n24) );
  NANDN U286 ( .A(n1225), .B(n24), .Z(n25) );
  NAND U287 ( .A(n23), .B(n25), .Z(n1476) );
  NAND U288 ( .A(n1239), .B(n1240), .Z(n26) );
  XOR U289 ( .A(n1239), .B(n1240), .Z(n27) );
  NANDN U290 ( .A(n1238), .B(n27), .Z(n28) );
  NAND U291 ( .A(n26), .B(n28), .Z(n1473) );
  NAND U292 ( .A(n865), .B(n866), .Z(n29) );
  XOR U293 ( .A(n865), .B(n866), .Z(n30) );
  NANDN U294 ( .A(n864), .B(n30), .Z(n31) );
  NAND U295 ( .A(n29), .B(n31), .Z(n1330) );
  NAND U296 ( .A(n899), .B(n900), .Z(n32) );
  XOR U297 ( .A(n899), .B(n900), .Z(n33) );
  NANDN U298 ( .A(n898), .B(n33), .Z(n34) );
  NAND U299 ( .A(n32), .B(n34), .Z(n1377) );
  XOR U300 ( .A(n1143), .B(n1144), .Z(n35) );
  XNOR U301 ( .A(n1142), .B(n35), .Z(n1359) );
  NAND U302 ( .A(n1399), .B(n1398), .Z(n36) );
  XOR U303 ( .A(n1399), .B(n1398), .Z(n37) );
  NANDN U304 ( .A(n1400), .B(n37), .Z(n38) );
  NAND U305 ( .A(n36), .B(n38), .Z(n1566) );
  NAND U306 ( .A(n1504), .B(n1505), .Z(n39) );
  XOR U307 ( .A(n1504), .B(n1505), .Z(n40) );
  NAND U308 ( .A(n40), .B(n1503), .Z(n41) );
  NAND U309 ( .A(n39), .B(n41), .Z(n1569) );
  NAND U310 ( .A(n1412), .B(n1411), .Z(n42) );
  XOR U311 ( .A(n1412), .B(n1411), .Z(n43) );
  NANDN U312 ( .A(n1413), .B(n43), .Z(n44) );
  NAND U313 ( .A(n42), .B(n44), .Z(n1573) );
  XNOR U314 ( .A(n1506), .B(n1508), .Z(n45) );
  XNOR U315 ( .A(n1507), .B(n45), .Z(n1458) );
  XNOR U316 ( .A(n1624), .B(n1623), .Z(n1618) );
  NAND U317 ( .A(n1575), .B(n1576), .Z(n46) );
  XOR U318 ( .A(n1575), .B(n1576), .Z(n47) );
  NANDN U319 ( .A(n1574), .B(n47), .Z(n48) );
  NAND U320 ( .A(n46), .B(n48), .Z(n1615) );
  XOR U321 ( .A(n1318), .B(n1316), .Z(n49) );
  NANDN U322 ( .A(n1317), .B(n49), .Z(n50) );
  NAND U323 ( .A(n1318), .B(n1316), .Z(n51) );
  AND U324 ( .A(n50), .B(n51), .Z(n1521) );
  NAND U325 ( .A(n1278), .B(n1279), .Z(n52) );
  XOR U326 ( .A(n1278), .B(n1279), .Z(n53) );
  NANDN U327 ( .A(n1277), .B(n53), .Z(n54) );
  NAND U328 ( .A(n52), .B(n54), .Z(n1429) );
  NAND U329 ( .A(n1587), .B(n1589), .Z(n55) );
  XOR U330 ( .A(n1587), .B(n1589), .Z(n56) );
  NAND U331 ( .A(n56), .B(n1588), .Z(n57) );
  NAND U332 ( .A(n55), .B(n57), .Z(n1613) );
  NAND U333 ( .A(n868), .B(n869), .Z(n58) );
  XOR U334 ( .A(n868), .B(n869), .Z(n59) );
  NANDN U335 ( .A(n867), .B(n59), .Z(n60) );
  NAND U336 ( .A(n58), .B(n60), .Z(n1340) );
  NAND U337 ( .A(n942), .B(n943), .Z(n61) );
  XOR U338 ( .A(n942), .B(n943), .Z(n62) );
  NANDN U339 ( .A(n941), .B(n62), .Z(n63) );
  NAND U340 ( .A(n61), .B(n63), .Z(n1118) );
  NAND U341 ( .A(n917), .B(n916), .Z(n64) );
  NAND U342 ( .A(n914), .B(n915), .Z(n65) );
  NAND U343 ( .A(n64), .B(n65), .Z(n1088) );
  NAND U344 ( .A(n1055), .B(n1054), .Z(n66) );
  NAND U345 ( .A(n1052), .B(n1053), .Z(n67) );
  NAND U346 ( .A(n66), .B(n67), .Z(n1086) );
  XNOR U347 ( .A(n1199), .B(n1198), .Z(n1200) );
  NAND U348 ( .A(n955), .B(n956), .Z(n68) );
  XOR U349 ( .A(n955), .B(n956), .Z(n69) );
  NANDN U350 ( .A(n954), .B(n69), .Z(n70) );
  NAND U351 ( .A(n68), .B(n70), .Z(n1343) );
  NAND U352 ( .A(n987), .B(n989), .Z(n71) );
  XOR U353 ( .A(n987), .B(n989), .Z(n72) );
  NAND U354 ( .A(n72), .B(n988), .Z(n73) );
  NAND U355 ( .A(n71), .B(n73), .Z(n1300) );
  NAND U356 ( .A(n962), .B(n963), .Z(n74) );
  XOR U357 ( .A(n962), .B(n963), .Z(n75) );
  NANDN U358 ( .A(n961), .B(n75), .Z(n76) );
  NAND U359 ( .A(n74), .B(n76), .Z(n1115) );
  NAND U360 ( .A(n505), .B(n506), .Z(n77) );
  XOR U361 ( .A(n505), .B(n506), .Z(n78) );
  NANDN U362 ( .A(n504), .B(n78), .Z(n79) );
  NAND U363 ( .A(n77), .B(n79), .Z(n1220) );
  NAND U364 ( .A(n477), .B(n478), .Z(n80) );
  XOR U365 ( .A(n477), .B(n478), .Z(n81) );
  NANDN U366 ( .A(n476), .B(n81), .Z(n82) );
  NAND U367 ( .A(n80), .B(n82), .Z(n1174) );
  NAND U368 ( .A(n1067), .B(n1069), .Z(n83) );
  XOR U369 ( .A(n1067), .B(n1069), .Z(n84) );
  NAND U370 ( .A(n84), .B(n1068), .Z(n85) );
  NAND U371 ( .A(n83), .B(n85), .Z(n1293) );
  NAND U372 ( .A(n1236), .B(n1237), .Z(n86) );
  XOR U373 ( .A(n1236), .B(n1237), .Z(n87) );
  NANDN U374 ( .A(n1235), .B(n87), .Z(n88) );
  NAND U375 ( .A(n86), .B(n88), .Z(n1471) );
  NAND U376 ( .A(n1352), .B(n1353), .Z(n89) );
  XOR U377 ( .A(n1352), .B(n1353), .Z(n90) );
  NANDN U378 ( .A(n1351), .B(n90), .Z(n91) );
  NAND U379 ( .A(n89), .B(n91), .Z(n1489) );
  NAND U380 ( .A(n1209), .B(n1210), .Z(n92) );
  XOR U381 ( .A(n1209), .B(n1210), .Z(n93) );
  NANDN U382 ( .A(n1208), .B(n93), .Z(n94) );
  NAND U383 ( .A(n92), .B(n94), .Z(n1484) );
  XOR U384 ( .A(n1121), .B(n1123), .Z(n95) );
  XNOR U385 ( .A(n1122), .B(n95), .Z(n1332) );
  XNOR U386 ( .A(n1550), .B(n1551), .Z(n1571) );
  NAND U387 ( .A(n1474), .B(n1476), .Z(n96) );
  XOR U388 ( .A(n1474), .B(n1476), .Z(n97) );
  NAND U389 ( .A(n97), .B(n1475), .Z(n98) );
  NAND U390 ( .A(n96), .B(n98), .Z(n1558) );
  NAND U391 ( .A(n1274), .B(n1275), .Z(n99) );
  XOR U392 ( .A(n1274), .B(n1275), .Z(n100) );
  NANDN U393 ( .A(n1273), .B(n100), .Z(n101) );
  NAND U394 ( .A(n99), .B(n101), .Z(n1444) );
  XOR U395 ( .A(n1359), .B(n1357), .Z(n102) );
  NANDN U396 ( .A(n1358), .B(n102), .Z(n103) );
  NAND U397 ( .A(n1359), .B(n1357), .Z(n104) );
  AND U398 ( .A(n103), .B(n104), .Z(n1516) );
  NAND U399 ( .A(n1564), .B(n1566), .Z(n105) );
  XOR U400 ( .A(n1564), .B(n1566), .Z(n106) );
  NAND U401 ( .A(n106), .B(n1565), .Z(n107) );
  NAND U402 ( .A(n105), .B(n107), .Z(n1620) );
  XNOR U403 ( .A(n1497), .B(n1496), .Z(n1522) );
  XOR U404 ( .A(n1456), .B(n1458), .Z(n108) );
  XNOR U405 ( .A(n1457), .B(n108), .Z(n1453) );
  NAND U406 ( .A(n1579), .B(n1580), .Z(n109) );
  XOR U407 ( .A(n1579), .B(n1580), .Z(n110) );
  NANDN U408 ( .A(n1578), .B(n110), .Z(n111) );
  NAND U409 ( .A(n109), .B(n111), .Z(n1612) );
  NAND U410 ( .A(n1537), .B(n1538), .Z(n112) );
  XOR U411 ( .A(n1537), .B(n1538), .Z(n113) );
  NANDN U412 ( .A(n1536), .B(n113), .Z(n114) );
  NAND U413 ( .A(n112), .B(n114), .Z(n1609) );
  NAND U414 ( .A(oglobal[4]), .B(n1628), .Z(n115) );
  XOR U415 ( .A(oglobal[4]), .B(n1628), .Z(n116) );
  NANDN U416 ( .A(n1627), .B(n116), .Z(n117) );
  NAND U417 ( .A(n115), .B(n117), .Z(n1631) );
  XNOR U418 ( .A(n898), .B(n899), .Z(n118) );
  XNOR U419 ( .A(n900), .B(n118), .Z(n402) );
  XOR U420 ( .A(n396), .B(n394), .Z(n119) );
  NANDN U421 ( .A(n395), .B(n119), .Z(n120) );
  NAND U422 ( .A(n396), .B(n394), .Z(n121) );
  AND U423 ( .A(n120), .B(n121), .Z(n1318) );
  NAND U424 ( .A(n951), .B(n952), .Z(n122) );
  XOR U425 ( .A(n951), .B(n952), .Z(n123) );
  NANDN U426 ( .A(n950), .B(n123), .Z(n124) );
  NAND U427 ( .A(n122), .B(n124), .Z(n1119) );
  NAND U428 ( .A(n1044), .B(n1043), .Z(n125) );
  NAND U429 ( .A(n1041), .B(n1042), .Z(n126) );
  NAND U430 ( .A(n125), .B(n126), .Z(n1079) );
  NAND U431 ( .A(n913), .B(n912), .Z(n127) );
  NAND U432 ( .A(n910), .B(n911), .Z(n128) );
  NAND U433 ( .A(n127), .B(n128), .Z(n1089) );
  NAND U434 ( .A(n995), .B(n994), .Z(n129) );
  NAND U435 ( .A(n992), .B(n993), .Z(n130) );
  NAND U436 ( .A(n129), .B(n130), .Z(n1159) );
  XNOR U437 ( .A(n1154), .B(n1153), .Z(n1155) );
  XNOR U438 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U439 ( .A(n937), .B(n938), .Z(n131) );
  XOR U440 ( .A(n937), .B(n938), .Z(n132) );
  NANDN U441 ( .A(n936), .B(n132), .Z(n133) );
  NAND U442 ( .A(n131), .B(n133), .Z(n1309) );
  NAND U443 ( .A(n1028), .B(n1030), .Z(n134) );
  XOR U444 ( .A(n1028), .B(n1030), .Z(n135) );
  NAND U445 ( .A(n135), .B(n1029), .Z(n136) );
  NAND U446 ( .A(n134), .B(n136), .Z(n1303) );
  XNOR U447 ( .A(n1229), .B(n1228), .Z(n137) );
  XNOR U448 ( .A(n1231), .B(n137), .Z(n1298) );
  NAND U449 ( .A(n606), .B(n607), .Z(n138) );
  XOR U450 ( .A(n606), .B(n607), .Z(n139) );
  NANDN U451 ( .A(n605), .B(n139), .Z(n140) );
  NAND U452 ( .A(n138), .B(n140), .Z(n1137) );
  NAND U453 ( .A(n441), .B(n442), .Z(n141) );
  XOR U454 ( .A(n441), .B(n442), .Z(n142) );
  NANDN U455 ( .A(n440), .B(n142), .Z(n143) );
  NAND U456 ( .A(n141), .B(n143), .Z(n1111) );
  NAND U457 ( .A(n723), .B(n724), .Z(n144) );
  XOR U458 ( .A(n723), .B(n724), .Z(n145) );
  NANDN U459 ( .A(n722), .B(n145), .Z(n146) );
  NAND U460 ( .A(n144), .B(n146), .Z(n1143) );
  NAND U461 ( .A(n805), .B(n806), .Z(n147) );
  XOR U462 ( .A(n805), .B(n806), .Z(n148) );
  NANDN U463 ( .A(n804), .B(n148), .Z(n149) );
  NAND U464 ( .A(n147), .B(n149), .Z(n1129) );
  NAND U465 ( .A(n1299), .B(n1301), .Z(n150) );
  XOR U466 ( .A(n1299), .B(n1301), .Z(n151) );
  NAND U467 ( .A(n151), .B(n1300), .Z(n152) );
  NAND U468 ( .A(n150), .B(n152), .Z(n1398) );
  NAND U469 ( .A(n1339), .B(n1341), .Z(n153) );
  XOR U470 ( .A(n1339), .B(n1341), .Z(n154) );
  NAND U471 ( .A(n154), .B(n1340), .Z(n155) );
  NAND U472 ( .A(n153), .B(n155), .Z(n1396) );
  NAND U473 ( .A(n1115), .B(n1117), .Z(n156) );
  XOR U474 ( .A(n1115), .B(n1117), .Z(n157) );
  NAND U475 ( .A(n157), .B(n1116), .Z(n158) );
  NAND U476 ( .A(n156), .B(n158), .Z(n1500) );
  NAND U477 ( .A(n1092), .B(n1093), .Z(n159) );
  XOR U478 ( .A(n1092), .B(n1093), .Z(n160) );
  NANDN U479 ( .A(n1091), .B(n160), .Z(n161) );
  NAND U480 ( .A(n159), .B(n161), .Z(n1465) );
  NAND U481 ( .A(n1085), .B(n1086), .Z(n162) );
  XOR U482 ( .A(n1085), .B(n1086), .Z(n163) );
  NANDN U483 ( .A(n1084), .B(n163), .Z(n164) );
  NAND U484 ( .A(n162), .B(n164), .Z(n1425) );
  NAND U485 ( .A(n1164), .B(n1165), .Z(n165) );
  XOR U486 ( .A(n1164), .B(n1165), .Z(n166) );
  NANDN U487 ( .A(n1163), .B(n166), .Z(n167) );
  NAND U488 ( .A(n165), .B(n167), .Z(n1418) );
  NAND U489 ( .A(n1349), .B(n1350), .Z(n168) );
  XOR U490 ( .A(n1349), .B(n1350), .Z(n169) );
  NANDN U491 ( .A(n1348), .B(n169), .Z(n170) );
  NAND U492 ( .A(n168), .B(n170), .Z(n1487) );
  NAND U493 ( .A(n1206), .B(n1207), .Z(n171) );
  XOR U494 ( .A(n1206), .B(n1207), .Z(n172) );
  NANDN U495 ( .A(n1205), .B(n172), .Z(n173) );
  NAND U496 ( .A(n171), .B(n173), .Z(n1482) );
  XNOR U497 ( .A(n456), .B(n455), .Z(n457) );
  NAND U498 ( .A(n902), .B(n903), .Z(n174) );
  XOR U499 ( .A(n902), .B(n903), .Z(n175) );
  NANDN U500 ( .A(n901), .B(n175), .Z(n176) );
  NAND U501 ( .A(n174), .B(n176), .Z(n1375) );
  NAND U502 ( .A(n404), .B(n406), .Z(n177) );
  XOR U503 ( .A(n404), .B(n406), .Z(n178) );
  NAND U504 ( .A(n178), .B(n405), .Z(n179) );
  NAND U505 ( .A(n177), .B(n179), .Z(n1370) );
  NAND U506 ( .A(n1218), .B(n1220), .Z(n180) );
  XOR U507 ( .A(n1218), .B(n1220), .Z(n181) );
  NAND U508 ( .A(n181), .B(n1219), .Z(n182) );
  NAND U509 ( .A(n180), .B(n182), .Z(n1503) );
  XOR U510 ( .A(n1292), .B(n1290), .Z(n183) );
  NANDN U511 ( .A(n1291), .B(n183), .Z(n184) );
  NAND U512 ( .A(n1292), .B(n1290), .Z(n185) );
  AND U513 ( .A(n184), .B(n185), .Z(n1495) );
  NAND U514 ( .A(n1479), .B(n1480), .Z(n186) );
  XOR U515 ( .A(n1479), .B(n1480), .Z(n187) );
  NANDN U516 ( .A(n1478), .B(n187), .Z(n188) );
  NAND U517 ( .A(n186), .B(n188), .Z(n1546) );
  XOR U518 ( .A(n1362), .B(n1363), .Z(n189) );
  XNOR U519 ( .A(n1360), .B(n189), .Z(n1278) );
  NAND U520 ( .A(n1406), .B(n1407), .Z(n190) );
  XOR U521 ( .A(n1406), .B(n1407), .Z(n191) );
  NANDN U522 ( .A(n1405), .B(n191), .Z(n192) );
  NAND U523 ( .A(n190), .B(n192), .Z(n1540) );
  NAND U524 ( .A(n1571), .B(n1573), .Z(n193) );
  XOR U525 ( .A(n1571), .B(n1573), .Z(n194) );
  NAND U526 ( .A(n194), .B(n1572), .Z(n195) );
  NAND U527 ( .A(n193), .B(n195), .Z(n1616) );
  XOR U528 ( .A(n1280), .B(n1282), .Z(n196) );
  XNOR U529 ( .A(n1281), .B(n196), .Z(n1328) );
  NAND U530 ( .A(n1619), .B(n1620), .Z(n197) );
  XOR U531 ( .A(n1619), .B(n1620), .Z(n198) );
  NANDN U532 ( .A(n1618), .B(n198), .Z(n199) );
  NAND U533 ( .A(n197), .B(n199), .Z(n1633) );
  XOR U534 ( .A(n1032), .B(n1034), .Z(n200) );
  XNOR U535 ( .A(n1033), .B(n200), .Z(n401) );
  NAND U536 ( .A(n398), .B(n399), .Z(n201) );
  XOR U537 ( .A(n398), .B(n399), .Z(n202) );
  NANDN U538 ( .A(n397), .B(n202), .Z(n203) );
  NAND U539 ( .A(n201), .B(n203), .Z(n1316) );
  XNOR U540 ( .A(n1453), .B(n1454), .Z(n204) );
  XNOR U541 ( .A(n1452), .B(n204), .Z(n1431) );
  NAND U542 ( .A(n1591), .B(n1593), .Z(n205) );
  XOR U543 ( .A(n1591), .B(n1593), .Z(n206) );
  NAND U544 ( .A(n206), .B(n1592), .Z(n207) );
  NAND U545 ( .A(n205), .B(n207), .Z(n1604) );
  NAND U546 ( .A(n1612), .B(n1614), .Z(n208) );
  XOR U547 ( .A(n1612), .B(n1614), .Z(n209) );
  NAND U548 ( .A(n209), .B(n1613), .Z(n210) );
  NAND U549 ( .A(n208), .B(n210), .Z(n1641) );
  XOR U550 ( .A(oglobal[5]), .B(n1632), .Z(n211) );
  NAND U551 ( .A(n211), .B(n1631), .Z(n212) );
  NAND U552 ( .A(oglobal[5]), .B(n1632), .Z(n213) );
  AND U553 ( .A(n212), .B(n213), .Z(n1655) );
  XNOR U554 ( .A(n799), .B(n798), .Z(n800) );
  XNOR U555 ( .A(n450), .B(n449), .Z(n451) );
  XNOR U556 ( .A(n420), .B(n419), .Z(n421) );
  XNOR U557 ( .A(n1169), .B(n1168), .Z(n1312) );
  NAND U558 ( .A(n411), .B(n412), .Z(n214) );
  XOR U559 ( .A(n411), .B(n412), .Z(n215) );
  NANDN U560 ( .A(n410), .B(n215), .Z(n216) );
  NAND U561 ( .A(n214), .B(n216), .Z(n1183) );
  XNOR U562 ( .A(n1236), .B(n1235), .Z(n217) );
  XNOR U563 ( .A(n1237), .B(n217), .Z(n1173) );
  NAND U564 ( .A(n438), .B(n439), .Z(n218) );
  XOR U565 ( .A(n438), .B(n439), .Z(n219) );
  NANDN U566 ( .A(n437), .B(n219), .Z(n220) );
  NAND U567 ( .A(n218), .B(n220), .Z(n1109) );
  NAND U568 ( .A(n1297), .B(n1298), .Z(n221) );
  XOR U569 ( .A(n1297), .B(n1298), .Z(n222) );
  NANDN U570 ( .A(n1296), .B(n222), .Z(n223) );
  NAND U571 ( .A(n221), .B(n223), .Z(n1399) );
  NAND U572 ( .A(n1252), .B(n1253), .Z(n224) );
  XOR U573 ( .A(n1252), .B(n1253), .Z(n225) );
  NANDN U574 ( .A(n1251), .B(n225), .Z(n226) );
  NAND U575 ( .A(n224), .B(n226), .Z(n1416) );
  NAND U576 ( .A(n1223), .B(n1224), .Z(n227) );
  XOR U577 ( .A(n1223), .B(n1224), .Z(n228) );
  NANDN U578 ( .A(n1222), .B(n228), .Z(n229) );
  NAND U579 ( .A(n227), .B(n229), .Z(n1474) );
  NAND U580 ( .A(n1160), .B(n1161), .Z(n230) );
  XOR U581 ( .A(n1160), .B(n1161), .Z(n231) );
  NANDN U582 ( .A(n1159), .B(n231), .Z(n232) );
  NAND U583 ( .A(n230), .B(n232), .Z(n1469) );
  XNOR U584 ( .A(n686), .B(n685), .Z(n687) );
  XNOR U585 ( .A(n815), .B(n814), .Z(n816) );
  XNOR U586 ( .A(n847), .B(n846), .Z(n848) );
  XNOR U587 ( .A(n520), .B(n519), .Z(n521) );
  XNOR U588 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U589 ( .A(n615), .B(n614), .Z(n616) );
  NAND U590 ( .A(n1307), .B(n1308), .Z(n233) );
  XOR U591 ( .A(n1307), .B(n1308), .Z(n234) );
  NANDN U592 ( .A(n1306), .B(n234), .Z(n235) );
  NAND U593 ( .A(n233), .B(n235), .Z(n1412) );
  NAND U594 ( .A(n434), .B(n435), .Z(n236) );
  XOR U595 ( .A(n434), .B(n435), .Z(n237) );
  NANDN U596 ( .A(n433), .B(n237), .Z(n238) );
  NAND U597 ( .A(n236), .B(n238), .Z(n1369) );
  NAND U598 ( .A(n529), .B(n530), .Z(n239) );
  XOR U599 ( .A(n529), .B(n530), .Z(n240) );
  NANDN U600 ( .A(n528), .B(n240), .Z(n241) );
  NAND U601 ( .A(n239), .B(n241), .Z(n1362) );
  NAND U602 ( .A(n1337), .B(n1338), .Z(n242) );
  XOR U603 ( .A(n1337), .B(n1338), .Z(n243) );
  NANDN U604 ( .A(n1336), .B(n243), .Z(n244) );
  NAND U605 ( .A(n242), .B(n244), .Z(n1460) );
  NAND U606 ( .A(n1396), .B(n1397), .Z(n245) );
  XOR U607 ( .A(n1396), .B(n1397), .Z(n246) );
  NANDN U608 ( .A(n1395), .B(n246), .Z(n247) );
  NAND U609 ( .A(n245), .B(n247), .Z(n1564) );
  NAND U610 ( .A(n1465), .B(n1467), .Z(n248) );
  XOR U611 ( .A(n1465), .B(n1467), .Z(n249) );
  NAND U612 ( .A(n249), .B(n1466), .Z(n250) );
  NAND U613 ( .A(n248), .B(n250), .Z(n1575) );
  NAND U614 ( .A(n1409), .B(n1408), .Z(n251) );
  XOR U615 ( .A(n1409), .B(n1408), .Z(n252) );
  NANDN U616 ( .A(n1410), .B(n252), .Z(n253) );
  NAND U617 ( .A(n251), .B(n253), .Z(n1572) );
  NAND U618 ( .A(n1423), .B(n1425), .Z(n254) );
  XOR U619 ( .A(n1423), .B(n1425), .Z(n255) );
  NAND U620 ( .A(n255), .B(n1424), .Z(n256) );
  NAND U621 ( .A(n254), .B(n256), .Z(n1549) );
  NAND U622 ( .A(n1471), .B(n1473), .Z(n257) );
  XOR U623 ( .A(n1471), .B(n1473), .Z(n258) );
  NAND U624 ( .A(n258), .B(n1472), .Z(n259) );
  NAND U625 ( .A(n257), .B(n259), .Z(n1559) );
  NAND U626 ( .A(n1482), .B(n1484), .Z(n260) );
  XOR U627 ( .A(n1482), .B(n1484), .Z(n261) );
  NAND U628 ( .A(n261), .B(n1483), .Z(n262) );
  NAND U629 ( .A(n260), .B(n262), .Z(n1556) );
  NAND U630 ( .A(n1567), .B(n1569), .Z(n263) );
  XOR U631 ( .A(n1567), .B(n1569), .Z(n264) );
  NAND U632 ( .A(n264), .B(n1568), .Z(n265) );
  NAND U633 ( .A(n263), .B(n265), .Z(n1619) );
  NAND U634 ( .A(n1547), .B(oglobal[3]), .Z(n266) );
  XOR U635 ( .A(n1547), .B(oglobal[3]), .Z(n267) );
  NANDN U636 ( .A(n1546), .B(n267), .Z(n268) );
  NAND U637 ( .A(n266), .B(n268), .Z(n1628) );
  XOR U638 ( .A(n955), .B(n954), .Z(n269) );
  XNOR U639 ( .A(n956), .B(n269), .Z(n1033) );
  XOR U640 ( .A(n1282), .B(n1280), .Z(n270) );
  NANDN U641 ( .A(n1281), .B(n270), .Z(n271) );
  NAND U642 ( .A(n1282), .B(n1280), .Z(n272) );
  AND U643 ( .A(n271), .B(n272), .Z(n1428) );
  NAND U644 ( .A(n1521), .B(n1522), .Z(n273) );
  XOR U645 ( .A(n1521), .B(n1522), .Z(n274) );
  NANDN U646 ( .A(n1523), .B(n274), .Z(n275) );
  NAND U647 ( .A(n273), .B(n275), .Z(n1591) );
  NAND U648 ( .A(n1327), .B(n1328), .Z(n276) );
  XOR U649 ( .A(n1327), .B(n1328), .Z(n277) );
  NANDN U650 ( .A(n1326), .B(n277), .Z(n278) );
  NAND U651 ( .A(n276), .B(n278), .Z(n1390) );
  NAND U652 ( .A(n1453), .B(n1454), .Z(n279) );
  XOR U653 ( .A(n1453), .B(n1454), .Z(n280) );
  NANDN U654 ( .A(n1452), .B(n280), .Z(n281) );
  NAND U655 ( .A(n279), .B(n281), .Z(n1534) );
  XNOR U656 ( .A(n1608), .B(n1609), .Z(n1605) );
  XNOR U657 ( .A(n1643), .B(n1642), .Z(n1647) );
  NAND U658 ( .A(n1075), .B(n1076), .Z(n282) );
  XOR U659 ( .A(n1075), .B(n1076), .Z(n283) );
  NANDN U660 ( .A(n1074), .B(n283), .Z(n284) );
  NAND U661 ( .A(n282), .B(n284), .Z(n1284) );
  XOR U662 ( .A(n1655), .B(n1654), .Z(n285) );
  NANDN U663 ( .A(oglobal[6]), .B(n285), .Z(n286) );
  NAND U664 ( .A(n1655), .B(n1654), .Z(n287) );
  AND U665 ( .A(n286), .B(n287), .Z(n1664) );
  XNOR U666 ( .A(n1167), .B(n1166), .Z(n1168) );
  XNOR U667 ( .A(n1187), .B(n1186), .Z(n1188) );
  XOR U668 ( .A(n1088), .B(n1087), .Z(n288) );
  XNOR U669 ( .A(n1089), .B(n288), .Z(n1310) );
  NAND U670 ( .A(n502), .B(n503), .Z(n289) );
  XOR U671 ( .A(n502), .B(n503), .Z(n290) );
  NANDN U672 ( .A(n501), .B(n290), .Z(n291) );
  NAND U673 ( .A(n289), .B(n291), .Z(n1219) );
  NAND U674 ( .A(n408), .B(n409), .Z(n292) );
  XOR U675 ( .A(n408), .B(n409), .Z(n293) );
  NANDN U676 ( .A(n407), .B(n293), .Z(n294) );
  NAND U677 ( .A(n292), .B(n294), .Z(n1181) );
  NAND U678 ( .A(n479), .B(n481), .Z(n295) );
  XOR U679 ( .A(n479), .B(n481), .Z(n296) );
  NAND U680 ( .A(n296), .B(n480), .Z(n297) );
  NAND U681 ( .A(n295), .B(n297), .Z(n1176) );
  XNOR U682 ( .A(n1349), .B(n1348), .Z(n298) );
  XNOR U683 ( .A(n1350), .B(n298), .Z(n1128) );
  NAND U684 ( .A(n1294), .B(n1295), .Z(n299) );
  XOR U685 ( .A(n1294), .B(n1295), .Z(n300) );
  NANDN U686 ( .A(n1293), .B(n300), .Z(n301) );
  NAND U687 ( .A(n299), .B(n301), .Z(n1400) );
  XNOR U688 ( .A(n768), .B(n767), .Z(n769) );
  XNOR U689 ( .A(n774), .B(n773), .Z(n775) );
  XNOR U690 ( .A(n697), .B(n696), .Z(n698) );
  XNOR U691 ( .A(n809), .B(n808), .Z(n810) );
  XNOR U692 ( .A(n828), .B(n827), .Z(n829) );
  XNOR U693 ( .A(n483), .B(n482), .Z(n484) );
  XNOR U694 ( .A(n877), .B(n876), .Z(n878) );
  XNOR U695 ( .A(n889), .B(n888), .Z(n890) );
  XNOR U696 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U697 ( .A(n834), .B(n833), .Z(n835) );
  XNOR U698 ( .A(n691), .B(oglobal[0]), .Z(n692) );
  XNOR U699 ( .A(n508), .B(n507), .Z(n509) );
  XNOR U700 ( .A(n489), .B(n488), .Z(n490) );
  XNOR U701 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U702 ( .A(n821), .B(n820), .Z(n822) );
  XNOR U703 ( .A(n859), .B(n858), .Z(n860) );
  XNOR U704 ( .A(n426), .B(n425), .Z(n427) );
  XNOR U705 ( .A(n414), .B(n413), .Z(n415) );
  XNOR U706 ( .A(n514), .B(n513), .Z(n515) );
  XNOR U707 ( .A(n495), .B(n494), .Z(n496) );
  XNOR U708 ( .A(n853), .B(n852), .Z(n854) );
  XNOR U709 ( .A(n444), .B(n443), .Z(n445) );
  XNOR U710 ( .A(n754), .B(n753), .Z(n755) );
  XNOR U711 ( .A(n760), .B(n759), .Z(n761) );
  NAND U712 ( .A(n1304), .B(n1305), .Z(n302) );
  XOR U713 ( .A(n1304), .B(n1305), .Z(n303) );
  NANDN U714 ( .A(n1303), .B(n303), .Z(n304) );
  NAND U715 ( .A(n302), .B(n304), .Z(n1413) );
  XOR U716 ( .A(n1034), .B(n1032), .Z(n305) );
  NANDN U717 ( .A(n1033), .B(n305), .Z(n306) );
  NAND U718 ( .A(n1034), .B(n1032), .Z(n307) );
  AND U719 ( .A(n306), .B(n307), .Z(n1267) );
  NAND U720 ( .A(n1143), .B(n1142), .Z(n308) );
  XOR U721 ( .A(n1143), .B(n1142), .Z(n309) );
  NANDN U722 ( .A(n1144), .B(n309), .Z(n310) );
  NAND U723 ( .A(n308), .B(n310), .Z(n1408) );
  NAND U724 ( .A(n1402), .B(n1403), .Z(n311) );
  XOR U725 ( .A(n1402), .B(n1403), .Z(n312) );
  NAND U726 ( .A(n312), .B(n1401), .Z(n313) );
  NAND U727 ( .A(n311), .B(n313), .Z(n1565) );
  NAND U728 ( .A(n1500), .B(n1502), .Z(n314) );
  XOR U729 ( .A(n1500), .B(n1502), .Z(n315) );
  NAND U730 ( .A(n315), .B(n1501), .Z(n316) );
  NAND U731 ( .A(n314), .B(n316), .Z(n1567) );
  NAND U732 ( .A(n1414), .B(n1416), .Z(n317) );
  XOR U733 ( .A(n1414), .B(n1416), .Z(n318) );
  NAND U734 ( .A(n318), .B(n1415), .Z(n319) );
  NAND U735 ( .A(n317), .B(n319), .Z(n1551) );
  NAND U736 ( .A(n1469), .B(n1470), .Z(n320) );
  XOR U737 ( .A(n1469), .B(n1470), .Z(n321) );
  NANDN U738 ( .A(n1468), .B(n321), .Z(n322) );
  NAND U739 ( .A(n320), .B(n322), .Z(n1561) );
  XOR U740 ( .A(n723), .B(n722), .Z(n323) );
  XNOR U741 ( .A(n724), .B(n323), .Z(n873) );
  XOR U742 ( .A(n1358), .B(n1359), .Z(n324) );
  XNOR U743 ( .A(n1357), .B(n324), .Z(n1281) );
  NAND U744 ( .A(n1264), .B(n1265), .Z(n325) );
  XOR U745 ( .A(n1264), .B(n1265), .Z(n326) );
  NANDN U746 ( .A(n1263), .B(n326), .Z(n327) );
  NAND U747 ( .A(n325), .B(n327), .Z(n1446) );
  XNOR U748 ( .A(n1461), .B(n1462), .Z(n1514) );
  NAND U749 ( .A(n1457), .B(n1458), .Z(n328) );
  XOR U750 ( .A(n1457), .B(n1458), .Z(n329) );
  NANDN U751 ( .A(n1456), .B(n329), .Z(n330) );
  NAND U752 ( .A(n328), .B(n330), .Z(n1582) );
  NAND U753 ( .A(n1434), .B(n1436), .Z(n331) );
  XOR U754 ( .A(n1434), .B(n1436), .Z(n332) );
  NAND U755 ( .A(n332), .B(n1435), .Z(n333) );
  NAND U756 ( .A(n331), .B(n333), .Z(n1589) );
  NAND U757 ( .A(n1555), .B(n1557), .Z(n334) );
  XOR U758 ( .A(n1555), .B(n1557), .Z(n335) );
  NAND U759 ( .A(n335), .B(n1556), .Z(n336) );
  NAND U760 ( .A(n334), .B(n336), .Z(n1622) );
  XNOR U761 ( .A(n958), .B(n957), .Z(n337) );
  XNOR U762 ( .A(n959), .B(n337), .Z(n901) );
  XNOR U763 ( .A(n505), .B(n504), .Z(n338) );
  XNOR U764 ( .A(n506), .B(n338), .Z(n434) );
  XNOR U765 ( .A(n477), .B(n476), .Z(n339) );
  XNOR U766 ( .A(n478), .B(n339), .Z(n465) );
  XNOR U767 ( .A(n411), .B(n410), .Z(n340) );
  XNOR U768 ( .A(n412), .B(n340), .Z(n864) );
  XNOR U769 ( .A(n868), .B(n867), .Z(n341) );
  XNOR U770 ( .A(n869), .B(n341), .Z(n471) );
  XOR U771 ( .A(n1278), .B(n1277), .Z(n342) );
  XNOR U772 ( .A(n1279), .B(n342), .Z(n1327) );
  NAND U773 ( .A(n1615), .B(n1617), .Z(n343) );
  XOR U774 ( .A(n1615), .B(n1617), .Z(n344) );
  NAND U775 ( .A(n344), .B(n1616), .Z(n345) );
  NAND U776 ( .A(n343), .B(n345), .Z(n1634) );
  NAND U777 ( .A(n401), .B(n402), .Z(n346) );
  XOR U778 ( .A(n401), .B(n402), .Z(n347) );
  NANDN U779 ( .A(n400), .B(n347), .Z(n348) );
  NAND U780 ( .A(n346), .B(n348), .Z(n1317) );
  XOR U781 ( .A(n1385), .B(n1386), .Z(n349) );
  NANDN U782 ( .A(n1387), .B(n349), .Z(n350) );
  NAND U783 ( .A(n1385), .B(n1386), .Z(n351) );
  AND U784 ( .A(n350), .B(n351), .Z(n1528) );
  NAND U785 ( .A(n1533), .B(n1535), .Z(n352) );
  XOR U786 ( .A(n1533), .B(n1535), .Z(n353) );
  NAND U787 ( .A(n353), .B(n1534), .Z(n354) );
  NAND U788 ( .A(n352), .B(n354), .Z(n1600) );
  NAND U789 ( .A(n1604), .B(n1605), .Z(n355) );
  XOR U790 ( .A(n1604), .B(n1605), .Z(n356) );
  NANDN U791 ( .A(n1603), .B(n356), .Z(n357) );
  NAND U792 ( .A(n355), .B(n357), .Z(n1650) );
  XOR U793 ( .A(oglobal[7]), .B(n1664), .Z(n358) );
  NANDN U794 ( .A(n1665), .B(n358), .Z(n359) );
  NAND U795 ( .A(oglobal[7]), .B(n1664), .Z(n360) );
  AND U796 ( .A(n359), .B(n360), .Z(n1666) );
  NAND U797 ( .A(n1670), .B(oglobal[12]), .Z(n361) );
  XNOR U798 ( .A(oglobal[13]), .B(n361), .Z(o[13]) );
  XOR U799 ( .A(x[34]), .B(y[34]), .Z(n770) );
  XOR U800 ( .A(x[38]), .B(y[38]), .Z(n767) );
  XNOR U801 ( .A(x[36]), .B(y[36]), .Z(n768) );
  XOR U802 ( .A(n770), .B(n769), .Z(n989) );
  XOR U803 ( .A(x[28]), .B(y[28]), .Z(n1018) );
  XOR U804 ( .A(x[32]), .B(y[32]), .Z(n1016) );
  XOR U805 ( .A(x[30]), .B(y[30]), .Z(n1015) );
  XOR U806 ( .A(n1016), .B(n1015), .Z(n1017) );
  XOR U807 ( .A(n1018), .B(n1017), .Z(n988) );
  XOR U808 ( .A(x[40]), .B(y[40]), .Z(n776) );
  XOR U809 ( .A(x[44]), .B(y[44]), .Z(n773) );
  XNOR U810 ( .A(x[42]), .B(y[42]), .Z(n774) );
  XOR U811 ( .A(n776), .B(n775), .Z(n987) );
  XNOR U812 ( .A(n988), .B(n987), .Z(n362) );
  XNOR U813 ( .A(n989), .B(n362), .Z(n406) );
  XOR U814 ( .A(x[16]), .B(y[16]), .Z(n688) );
  XOR U815 ( .A(x[20]), .B(y[20]), .Z(n685) );
  XNOR U816 ( .A(x[18]), .B(y[18]), .Z(n686) );
  XOR U817 ( .A(n688), .B(n687), .Z(n1067) );
  XOR U818 ( .A(x[22]), .B(y[22]), .Z(n1012) );
  XOR U819 ( .A(x[26]), .B(y[26]), .Z(n1010) );
  XOR U820 ( .A(x[24]), .B(y[24]), .Z(n1009) );
  XOR U821 ( .A(n1010), .B(n1009), .Z(n1011) );
  XOR U822 ( .A(n1012), .B(n1011), .Z(n1069) );
  XOR U823 ( .A(x[10]), .B(y[10]), .Z(n699) );
  XOR U824 ( .A(x[14]), .B(y[14]), .Z(n696) );
  XNOR U825 ( .A(x[12]), .B(y[12]), .Z(n697) );
  XOR U826 ( .A(n699), .B(n698), .Z(n1068) );
  XNOR U827 ( .A(n1069), .B(n1068), .Z(n363) );
  XNOR U828 ( .A(n1067), .B(n363), .Z(n405) );
  XOR U829 ( .A(x[58]), .B(y[58]), .Z(n641) );
  XOR U830 ( .A(x[62]), .B(y[62]), .Z(n639) );
  XNOR U831 ( .A(x[60]), .B(y[60]), .Z(n640) );
  XOR U832 ( .A(n639), .B(n640), .Z(n642) );
  XNOR U833 ( .A(n641), .B(n642), .Z(n943) );
  XOR U834 ( .A(x[46]), .B(y[46]), .Z(n789) );
  XOR U835 ( .A(x[50]), .B(y[50]), .Z(n787) );
  XOR U836 ( .A(x[48]), .B(y[48]), .Z(n786) );
  XOR U837 ( .A(n787), .B(n786), .Z(n788) );
  XNOR U838 ( .A(n789), .B(n788), .Z(n941) );
  XOR U839 ( .A(x[52]), .B(y[52]), .Z(n795) );
  XOR U840 ( .A(x[56]), .B(y[56]), .Z(n793) );
  XOR U841 ( .A(x[54]), .B(y[54]), .Z(n792) );
  XOR U842 ( .A(n793), .B(n792), .Z(n794) );
  XOR U843 ( .A(n795), .B(n794), .Z(n942) );
  XOR U844 ( .A(n941), .B(n942), .Z(n364) );
  XNOR U845 ( .A(n943), .B(n364), .Z(n404) );
  XNOR U846 ( .A(n405), .B(n404), .Z(n365) );
  XOR U847 ( .A(n406), .B(n365), .Z(n396) );
  XOR U848 ( .A(x[157]), .B(y[157]), .Z(n595) );
  XOR U849 ( .A(x[205]), .B(y[205]), .Z(n593) );
  XOR U850 ( .A(x[155]), .B(y[155]), .Z(n592) );
  XOR U851 ( .A(n593), .B(n592), .Z(n594) );
  XOR U852 ( .A(n595), .B(n594), .Z(n408) );
  XOR U853 ( .A(x[153]), .B(y[153]), .Z(n568) );
  XOR U854 ( .A(x[207]), .B(y[207]), .Z(n566) );
  XNOR U855 ( .A(x[151]), .B(y[151]), .Z(n567) );
  XOR U856 ( .A(n566), .B(n567), .Z(n569) );
  XNOR U857 ( .A(n568), .B(n569), .Z(n409) );
  XOR U858 ( .A(x[161]), .B(y[161]), .Z(n601) );
  XOR U859 ( .A(x[203]), .B(y[203]), .Z(n599) );
  XOR U860 ( .A(x[159]), .B(y[159]), .Z(n598) );
  XOR U861 ( .A(n599), .B(n598), .Z(n600) );
  XNOR U862 ( .A(n601), .B(n600), .Z(n407) );
  XOR U863 ( .A(n409), .B(n407), .Z(n366) );
  XOR U864 ( .A(n408), .B(n366), .Z(n435) );
  XOR U865 ( .A(x[145]), .B(y[145]), .Z(n574) );
  XOR U866 ( .A(x[211]), .B(y[211]), .Z(n572) );
  XNOR U867 ( .A(x[143]), .B(y[143]), .Z(n573) );
  XOR U868 ( .A(n572), .B(n573), .Z(n575) );
  XOR U869 ( .A(n574), .B(n575), .Z(n504) );
  XOR U870 ( .A(x[141]), .B(y[141]), .Z(n540) );
  XOR U871 ( .A(x[213]), .B(y[213]), .Z(n538) );
  XOR U872 ( .A(x[139]), .B(y[139]), .Z(n537) );
  XOR U873 ( .A(n538), .B(n537), .Z(n539) );
  XOR U874 ( .A(n540), .B(n539), .Z(n506) );
  XOR U875 ( .A(x[149]), .B(y[149]), .Z(n580) );
  XOR U876 ( .A(x[209]), .B(y[209]), .Z(n578) );
  XNOR U877 ( .A(x[147]), .B(y[147]), .Z(n579) );
  XOR U878 ( .A(n578), .B(n579), .Z(n581) );
  XNOR U879 ( .A(n580), .B(n581), .Z(n505) );
  XOR U880 ( .A(x[165]), .B(y[165]), .Z(n589) );
  XOR U881 ( .A(x[201]), .B(y[201]), .Z(n587) );
  XOR U882 ( .A(x[163]), .B(y[163]), .Z(n586) );
  XOR U883 ( .A(n587), .B(n586), .Z(n588) );
  XOR U884 ( .A(n589), .B(n588), .Z(n1028) );
  XOR U885 ( .A(x[177]), .B(y[177]), .Z(n749) );
  XOR U886 ( .A(x[191]), .B(y[191]), .Z(n747) );
  XNOR U887 ( .A(x[183]), .B(y[183]), .Z(n748) );
  XOR U888 ( .A(n747), .B(n748), .Z(n750) );
  XNOR U889 ( .A(n749), .B(n750), .Z(n712) );
  XOR U890 ( .A(x[185]), .B(y[185]), .Z(n710) );
  XOR U891 ( .A(x[181]), .B(y[181]), .Z(n709) );
  XOR U892 ( .A(n710), .B(n709), .Z(n711) );
  XOR U893 ( .A(n712), .B(n711), .Z(n1030) );
  XOR U894 ( .A(x[173]), .B(y[173]), .Z(n706) );
  XOR U895 ( .A(x[197]), .B(y[197]), .Z(n704) );
  XOR U896 ( .A(x[171]), .B(y[171]), .Z(n703) );
  XOR U897 ( .A(n704), .B(n703), .Z(n705) );
  XOR U898 ( .A(n706), .B(n705), .Z(n1029) );
  XNOR U899 ( .A(n1030), .B(n1029), .Z(n367) );
  XNOR U900 ( .A(n1028), .B(n367), .Z(n433) );
  XOR U901 ( .A(n434), .B(n433), .Z(n368) );
  XOR U902 ( .A(n435), .B(n368), .Z(n395) );
  XOR U903 ( .A(x[88]), .B(y[88]), .Z(n666) );
  XOR U904 ( .A(x[92]), .B(y[92]), .Z(n664) );
  XNOR U905 ( .A(x[90]), .B(y[90]), .Z(n665) );
  XOR U906 ( .A(n664), .B(n665), .Z(n667) );
  XOR U907 ( .A(n666), .B(n667), .Z(n964) );
  XOR U908 ( .A(x[94]), .B(y[94]), .Z(n811) );
  XOR U909 ( .A(x[98]), .B(y[98]), .Z(n808) );
  XNOR U910 ( .A(x[96]), .B(y[96]), .Z(n809) );
  XOR U911 ( .A(n811), .B(n810), .Z(n967) );
  XOR U912 ( .A(x[82]), .B(y[82]), .Z(n678) );
  XOR U913 ( .A(x[86]), .B(y[86]), .Z(n676) );
  XNOR U914 ( .A(x[84]), .B(y[84]), .Z(n677) );
  XOR U915 ( .A(n676), .B(n677), .Z(n679) );
  XNOR U916 ( .A(n678), .B(n679), .Z(n965) );
  XNOR U917 ( .A(n967), .B(n965), .Z(n369) );
  XOR U918 ( .A(n964), .B(n369), .Z(n903) );
  XOR U919 ( .A(x[106]), .B(y[106]), .Z(n817) );
  XOR U920 ( .A(x[110]), .B(y[110]), .Z(n814) );
  XNOR U921 ( .A(x[108]), .B(y[108]), .Z(n815) );
  XNOR U922 ( .A(n817), .B(n816), .Z(n957) );
  XOR U923 ( .A(x[112]), .B(y[112]), .Z(n849) );
  XOR U924 ( .A(x[116]), .B(y[116]), .Z(n846) );
  XNOR U925 ( .A(x[114]), .B(y[114]), .Z(n847) );
  XOR U926 ( .A(n849), .B(n848), .Z(n959) );
  XOR U927 ( .A(x[100]), .B(y[100]), .Z(n917) );
  XOR U928 ( .A(x[104]), .B(y[104]), .Z(n915) );
  XOR U929 ( .A(x[102]), .B(y[102]), .Z(n914) );
  XOR U930 ( .A(n915), .B(n914), .Z(n916) );
  XOR U931 ( .A(n917), .B(n916), .Z(n958) );
  XOR U932 ( .A(x[70]), .B(y[70]), .Z(n659) );
  XOR U933 ( .A(x[74]), .B(y[74]), .Z(n657) );
  XNOR U934 ( .A(x[72]), .B(y[72]), .Z(n658) );
  XOR U935 ( .A(n657), .B(n658), .Z(n660) );
  XOR U936 ( .A(n659), .B(n660), .Z(n970) );
  XOR U937 ( .A(x[76]), .B(y[76]), .Z(n647) );
  XOR U938 ( .A(x[80]), .B(y[80]), .Z(n645) );
  XNOR U939 ( .A(x[78]), .B(y[78]), .Z(n646) );
  XOR U940 ( .A(n645), .B(n646), .Z(n648) );
  XNOR U941 ( .A(n647), .B(n648), .Z(n972) );
  XOR U942 ( .A(x[64]), .B(y[64]), .Z(n635) );
  XOR U943 ( .A(x[68]), .B(y[68]), .Z(n633) );
  XNOR U944 ( .A(x[66]), .B(y[66]), .Z(n634) );
  XOR U945 ( .A(n633), .B(n634), .Z(n636) );
  XNOR U946 ( .A(n635), .B(n636), .Z(n971) );
  XNOR U947 ( .A(n972), .B(n971), .Z(n370) );
  XOR U948 ( .A(n970), .B(n370), .Z(n902) );
  XOR U949 ( .A(n901), .B(n902), .Z(n371) );
  XOR U950 ( .A(n903), .B(n371), .Z(n394) );
  XOR U951 ( .A(n395), .B(n394), .Z(n372) );
  XNOR U952 ( .A(n396), .B(n372), .Z(n1076) );
  XOR U953 ( .A(x[172]), .B(y[172]), .Z(n485) );
  XOR U954 ( .A(x[176]), .B(y[176]), .Z(n482) );
  XNOR U955 ( .A(x[174]), .B(y[174]), .Z(n483) );
  XNOR U956 ( .A(n485), .B(n484), .Z(n950) );
  XOR U957 ( .A(x[178]), .B(y[178]), .Z(n830) );
  XOR U958 ( .A(x[182]), .B(y[182]), .Z(n827) );
  XNOR U959 ( .A(x[180]), .B(y[180]), .Z(n828) );
  XOR U960 ( .A(n830), .B(n829), .Z(n952) );
  XOR U961 ( .A(x[247]), .B(y[247]), .Z(n920) );
  XOR U962 ( .A(x[249]), .B(y[249]), .Z(n918) );
  XNOR U963 ( .A(x[2]), .B(y[2]), .Z(n919) );
  XOR U964 ( .A(n918), .B(n919), .Z(n921) );
  XNOR U965 ( .A(n920), .B(n921), .Z(n951) );
  XNOR U966 ( .A(n952), .B(n951), .Z(n373) );
  XOR U967 ( .A(n950), .B(n373), .Z(n900) );
  XOR U968 ( .A(x[228]), .B(y[228]), .Z(n653) );
  XOR U969 ( .A(x[241]), .B(y[241]), .Z(n651) );
  XNOR U970 ( .A(x[230]), .B(y[230]), .Z(n652) );
  XOR U971 ( .A(n651), .B(n652), .Z(n654) );
  XOR U972 ( .A(n653), .B(n654), .Z(n870) );
  XOR U973 ( .A(x[208]), .B(y[208]), .Z(n422) );
  XOR U974 ( .A(x[210]), .B(y[210]), .Z(n419) );
  XNOR U975 ( .A(x[17]), .B(y[17]), .Z(n420) );
  XNOR U976 ( .A(n422), .B(n421), .Z(n722) );
  XOR U977 ( .A(x[212]), .B(y[212]), .Z(n452) );
  XOR U978 ( .A(x[237]), .B(y[237]), .Z(n449) );
  XNOR U979 ( .A(x[214]), .B(y[214]), .Z(n450) );
  XOR U980 ( .A(n452), .B(n451), .Z(n724) );
  XOR U981 ( .A(x[236]), .B(y[236]), .Z(n801) );
  XOR U982 ( .A(x[243]), .B(y[243]), .Z(n798) );
  XNOR U983 ( .A(x[238]), .B(y[238]), .Z(n799) );
  XOR U984 ( .A(n801), .B(n800), .Z(n723) );
  XOR U985 ( .A(x[224]), .B(y[224]), .Z(n672) );
  XOR U986 ( .A(x[226]), .B(y[226]), .Z(n670) );
  XNOR U987 ( .A(x[9]), .B(y[9]), .Z(n671) );
  XOR U988 ( .A(n670), .B(n671), .Z(n673) );
  XNOR U989 ( .A(n672), .B(n673), .Z(n871) );
  XNOR U990 ( .A(n873), .B(n871), .Z(n374) );
  XOR U991 ( .A(n870), .B(n374), .Z(n899) );
  XOR U992 ( .A(x[244]), .B(y[244]), .Z(n1024) );
  XOR U993 ( .A(x[246]), .B(y[246]), .Z(n1022) );
  XOR U994 ( .A(x[245]), .B(y[245]), .Z(n1021) );
  XOR U995 ( .A(n1022), .B(n1021), .Z(n1023) );
  XOR U996 ( .A(n1024), .B(n1023), .Z(n974) );
  XOR U997 ( .A(x[196]), .B(y[196]), .Z(n879) );
  XOR U998 ( .A(x[233]), .B(y[233]), .Z(n876) );
  XNOR U999 ( .A(x[198]), .B(y[198]), .Z(n877) );
  XOR U1000 ( .A(n879), .B(n878), .Z(n977) );
  XOR U1001 ( .A(x[192]), .B(y[192]), .Z(n891) );
  XOR U1002 ( .A(x[194]), .B(y[194]), .Z(n888) );
  XNOR U1003 ( .A(x[25]), .B(y[25]), .Z(n889) );
  XOR U1004 ( .A(n891), .B(n890), .Z(n975) );
  XNOR U1005 ( .A(n977), .B(n975), .Z(n375) );
  XOR U1006 ( .A(n974), .B(n375), .Z(n898) );
  XOR U1007 ( .A(x[148]), .B(y[148]), .Z(n522) );
  XOR U1008 ( .A(x[152]), .B(y[152]), .Z(n519) );
  XNOR U1009 ( .A(x[150]), .B(y[150]), .Z(n520) );
  XOR U1010 ( .A(n522), .B(n521), .Z(n963) );
  XOR U1011 ( .A(x[136]), .B(y[136]), .Z(n428) );
  XOR U1012 ( .A(x[140]), .B(y[140]), .Z(n425) );
  XNOR U1013 ( .A(x[138]), .B(y[138]), .Z(n426) );
  XNOR U1014 ( .A(n428), .B(n427), .Z(n961) );
  XOR U1015 ( .A(x[142]), .B(y[142]), .Z(n416) );
  XOR U1016 ( .A(x[146]), .B(y[146]), .Z(n413) );
  XNOR U1017 ( .A(x[144]), .B(y[144]), .Z(n414) );
  XOR U1018 ( .A(n416), .B(n415), .Z(n962) );
  XOR U1019 ( .A(n961), .B(n962), .Z(n376) );
  XOR U1020 ( .A(n963), .B(n376), .Z(n1034) );
  XOR U1021 ( .A(x[124]), .B(y[124]), .Z(n458) );
  XOR U1022 ( .A(x[128]), .B(y[128]), .Z(n455) );
  XNOR U1023 ( .A(x[126]), .B(y[126]), .Z(n456) );
  XNOR U1024 ( .A(n458), .B(n457), .Z(n954) );
  XOR U1025 ( .A(x[130]), .B(y[130]), .Z(n446) );
  XOR U1026 ( .A(x[134]), .B(y[134]), .Z(n443) );
  XNOR U1027 ( .A(x[132]), .B(y[132]), .Z(n444) );
  XOR U1028 ( .A(n446), .B(n445), .Z(n956) );
  XOR U1029 ( .A(x[118]), .B(y[118]), .Z(n855) );
  XOR U1030 ( .A(x[122]), .B(y[122]), .Z(n852) );
  XNOR U1031 ( .A(x[120]), .B(y[120]), .Z(n853) );
  XOR U1032 ( .A(n855), .B(n854), .Z(n955) );
  XOR U1033 ( .A(x[166]), .B(y[166]), .Z(n885) );
  XOR U1034 ( .A(x[170]), .B(y[170]), .Z(n882) );
  XNOR U1035 ( .A(x[168]), .B(y[168]), .Z(n883) );
  XOR U1036 ( .A(n885), .B(n884), .Z(n946) );
  XOR U1037 ( .A(x[154]), .B(y[154]), .Z(n516) );
  XOR U1038 ( .A(x[158]), .B(y[158]), .Z(n513) );
  XNOR U1039 ( .A(x[156]), .B(y[156]), .Z(n514) );
  XNOR U1040 ( .A(n516), .B(n515), .Z(n944) );
  XOR U1041 ( .A(x[160]), .B(y[160]), .Z(n497) );
  XOR U1042 ( .A(x[164]), .B(y[164]), .Z(n494) );
  XNOR U1043 ( .A(x[162]), .B(y[162]), .Z(n495) );
  XOR U1044 ( .A(n497), .B(n496), .Z(n945) );
  XOR U1045 ( .A(n944), .B(n945), .Z(n377) );
  XOR U1046 ( .A(n946), .B(n377), .Z(n1032) );
  XOR U1047 ( .A(x[184]), .B(y[184]), .Z(n842) );
  XOR U1048 ( .A(x[186]), .B(y[186]), .Z(n839) );
  XNOR U1049 ( .A(x[29]), .B(y[29]), .Z(n840) );
  XOR U1050 ( .A(n842), .B(n841), .Z(n982) );
  XOR U1051 ( .A(x[248]), .B(y[248]), .Z(n693) );
  XNOR U1052 ( .A(x[4]), .B(y[4]), .Z(n691) );
  XOR U1053 ( .A(n693), .B(n692), .Z(n981) );
  XOR U1054 ( .A(x[188]), .B(y[188]), .Z(n836) );
  XOR U1055 ( .A(x[231]), .B(y[231]), .Z(n833) );
  XNOR U1056 ( .A(x[190]), .B(y[190]), .Z(n834) );
  XOR U1057 ( .A(n836), .B(n835), .Z(n980) );
  XNOR U1058 ( .A(n981), .B(n980), .Z(n378) );
  XOR U1059 ( .A(n982), .B(n378), .Z(n530) );
  XOR U1060 ( .A(x[232]), .B(y[232]), .Z(n630) );
  XOR U1061 ( .A(x[234]), .B(y[234]), .Z(n627) );
  XNOR U1062 ( .A(x[5]), .B(y[5]), .Z(n628) );
  XNOR U1063 ( .A(n627), .B(n628), .Z(n629) );
  XOR U1064 ( .A(n630), .B(n629), .Z(n606) );
  XOR U1065 ( .A(x[220]), .B(y[220]), .Z(n823) );
  XOR U1066 ( .A(x[239]), .B(y[239]), .Z(n820) );
  XNOR U1067 ( .A(x[222]), .B(y[222]), .Z(n821) );
  XOR U1068 ( .A(n823), .B(n822), .Z(n607) );
  XOR U1069 ( .A(x[216]), .B(y[216]), .Z(n861) );
  XOR U1070 ( .A(x[218]), .B(y[218]), .Z(n858) );
  XNOR U1071 ( .A(x[13]), .B(y[13]), .Z(n859) );
  XNOR U1072 ( .A(n861), .B(n860), .Z(n605) );
  XOR U1073 ( .A(n607), .B(n605), .Z(n379) );
  XOR U1074 ( .A(n606), .B(n379), .Z(n529) );
  XOR U1075 ( .A(x[240]), .B(y[240]), .Z(n782) );
  XOR U1076 ( .A(x[242]), .B(y[242]), .Z(n779) );
  XNOR U1077 ( .A(x[1]), .B(y[1]), .Z(n780) );
  XOR U1078 ( .A(n782), .B(n781), .Z(n806) );
  XOR U1079 ( .A(x[204]), .B(y[204]), .Z(n510) );
  XOR U1080 ( .A(x[235]), .B(y[235]), .Z(n507) );
  XNOR U1081 ( .A(x[206]), .B(y[206]), .Z(n508) );
  XNOR U1082 ( .A(n510), .B(n509), .Z(n804) );
  XOR U1083 ( .A(x[200]), .B(y[200]), .Z(n491) );
  XOR U1084 ( .A(x[202]), .B(y[202]), .Z(n488) );
  XNOR U1085 ( .A(x[21]), .B(y[21]), .Z(n489) );
  XOR U1086 ( .A(n491), .B(n490), .Z(n805) );
  XOR U1087 ( .A(n804), .B(n805), .Z(n380) );
  XNOR U1088 ( .A(n806), .B(n380), .Z(n528) );
  XOR U1089 ( .A(n529), .B(n528), .Z(n381) );
  XOR U1090 ( .A(n530), .B(n381), .Z(n400) );
  XOR U1091 ( .A(n401), .B(n400), .Z(n382) );
  XOR U1092 ( .A(n402), .B(n382), .Z(n1074) );
  XOR U1093 ( .A(x[133]), .B(y[133]), .Z(n543) );
  XOR U1094 ( .A(x[217]), .B(y[217]), .Z(n541) );
  XNOR U1095 ( .A(x[131]), .B(y[131]), .Z(n542) );
  XOR U1096 ( .A(n541), .B(n542), .Z(n544) );
  XOR U1097 ( .A(n543), .B(n544), .Z(n476) );
  XOR U1098 ( .A(x[129]), .B(y[129]), .Z(n617) );
  XOR U1099 ( .A(x[219]), .B(y[219]), .Z(n614) );
  XNOR U1100 ( .A(x[127]), .B(y[127]), .Z(n615) );
  XOR U1101 ( .A(n617), .B(n616), .Z(n478) );
  XOR U1102 ( .A(x[137]), .B(y[137]), .Z(n533) );
  XOR U1103 ( .A(x[215]), .B(y[215]), .Z(n531) );
  XNOR U1104 ( .A(x[135]), .B(y[135]), .Z(n532) );
  XOR U1105 ( .A(n531), .B(n532), .Z(n534) );
  XNOR U1106 ( .A(n533), .B(n534), .Z(n477) );
  XOR U1107 ( .A(x[121]), .B(y[121]), .Z(n623) );
  XOR U1108 ( .A(x[223]), .B(y[223]), .Z(n621) );
  XOR U1109 ( .A(x[119]), .B(y[119]), .Z(n620) );
  XOR U1110 ( .A(n621), .B(n620), .Z(n622) );
  XOR U1111 ( .A(n623), .B(n622), .Z(n502) );
  XOR U1112 ( .A(x[117]), .B(y[117]), .Z(n549) );
  XOR U1113 ( .A(x[225]), .B(y[225]), .Z(n547) );
  XNOR U1114 ( .A(x[115]), .B(y[115]), .Z(n548) );
  XOR U1115 ( .A(n547), .B(n548), .Z(n550) );
  XNOR U1116 ( .A(n549), .B(n550), .Z(n503) );
  XOR U1117 ( .A(x[125]), .B(y[125]), .Z(n611) );
  XOR U1118 ( .A(x[221]), .B(y[221]), .Z(n609) );
  XOR U1119 ( .A(x[123]), .B(y[123]), .Z(n608) );
  XOR U1120 ( .A(n609), .B(n608), .Z(n610) );
  XNOR U1121 ( .A(n611), .B(n610), .Z(n501) );
  XOR U1122 ( .A(n503), .B(n501), .Z(n383) );
  XOR U1123 ( .A(n502), .B(n383), .Z(n464) );
  XOR U1124 ( .A(x[169]), .B(y[169]), .Z(n718) );
  XOR U1125 ( .A(x[199]), .B(y[199]), .Z(n716) );
  XOR U1126 ( .A(x[167]), .B(y[167]), .Z(n715) );
  XOR U1127 ( .A(n716), .B(n715), .Z(n717) );
  XOR U1128 ( .A(n718), .B(n717), .Z(n746) );
  XOR U1129 ( .A(x[187]), .B(y[187]), .Z(n762) );
  XOR U1130 ( .A(x[189]), .B(y[189]), .Z(n759) );
  XNOR U1131 ( .A(x[179]), .B(y[179]), .Z(n760) );
  XOR U1132 ( .A(n762), .B(n761), .Z(n745) );
  XOR U1133 ( .A(x[193]), .B(y[193]), .Z(n756) );
  XOR U1134 ( .A(x[195]), .B(y[195]), .Z(n753) );
  XNOR U1135 ( .A(x[175]), .B(y[175]), .Z(n754) );
  XOR U1136 ( .A(n756), .B(n755), .Z(n744) );
  XNOR U1137 ( .A(n745), .B(n744), .Z(n384) );
  XNOR U1138 ( .A(n746), .B(n384), .Z(n463) );
  XOR U1139 ( .A(n464), .B(n463), .Z(n385) );
  XOR U1140 ( .A(n465), .B(n385), .Z(n399) );
  XOR U1141 ( .A(x[33]), .B(y[33]), .Z(n932) );
  XOR U1142 ( .A(x[31]), .B(y[31]), .Z(n930) );
  XNOR U1143 ( .A(x[27]), .B(y[27]), .Z(n931) );
  XOR U1144 ( .A(n930), .B(n931), .Z(n933) );
  XNOR U1145 ( .A(n932), .B(n933), .Z(n442) );
  XOR U1146 ( .A(x[45]), .B(y[45]), .Z(n1058) );
  XOR U1147 ( .A(x[43]), .B(y[43]), .Z(n1057) );
  XOR U1148 ( .A(x[41]), .B(y[41]), .Z(n1056) );
  XOR U1149 ( .A(n1057), .B(n1056), .Z(n1059) );
  XNOR U1150 ( .A(n1058), .B(n1059), .Z(n440) );
  XOR U1151 ( .A(x[39]), .B(y[39]), .Z(n1055) );
  XOR U1152 ( .A(x[37]), .B(y[37]), .Z(n1053) );
  XOR U1153 ( .A(x[35]), .B(y[35]), .Z(n1052) );
  XOR U1154 ( .A(n1053), .B(n1052), .Z(n1054) );
  XOR U1155 ( .A(n1055), .B(n1054), .Z(n441) );
  XOR U1156 ( .A(n440), .B(n441), .Z(n386) );
  XNOR U1157 ( .A(n442), .B(n386), .Z(n866) );
  XOR U1158 ( .A(x[57]), .B(y[57]), .Z(n1037) );
  XOR U1159 ( .A(x[55]), .B(y[55]), .Z(n1036) );
  XOR U1160 ( .A(x[53]), .B(y[53]), .Z(n1035) );
  XOR U1161 ( .A(n1036), .B(n1035), .Z(n1038) );
  XNOR U1162 ( .A(n1037), .B(n1038), .Z(n410) );
  XOR U1163 ( .A(x[51]), .B(y[51]), .Z(n1065) );
  XOR U1164 ( .A(x[49]), .B(y[49]), .Z(n1063) );
  XOR U1165 ( .A(x[47]), .B(y[47]), .Z(n1062) );
  XOR U1166 ( .A(n1063), .B(n1062), .Z(n1064) );
  XOR U1167 ( .A(n1065), .B(n1064), .Z(n412) );
  XOR U1168 ( .A(x[63]), .B(y[63]), .Z(n1044) );
  XOR U1169 ( .A(x[61]), .B(y[61]), .Z(n1042) );
  XOR U1170 ( .A(x[59]), .B(y[59]), .Z(n1041) );
  XOR U1171 ( .A(n1042), .B(n1041), .Z(n1043) );
  XOR U1172 ( .A(n1044), .B(n1043), .Z(n411) );
  XOR U1173 ( .A(x[11]), .B(y[11]), .Z(n906) );
  XOR U1174 ( .A(x[7]), .B(y[7]), .Z(n905) );
  XOR U1175 ( .A(x[3]), .B(y[3]), .Z(n904) );
  XOR U1176 ( .A(n905), .B(n904), .Z(n907) );
  XNOR U1177 ( .A(n906), .B(n907), .Z(n437) );
  XOR U1178 ( .A(x[0]), .B(y[0]), .Z(n913) );
  XOR U1179 ( .A(x[8]), .B(y[8]), .Z(n911) );
  XOR U1180 ( .A(x[6]), .B(y[6]), .Z(n910) );
  XOR U1181 ( .A(n911), .B(n910), .Z(n912) );
  XOR U1182 ( .A(n913), .B(n912), .Z(n439) );
  XOR U1183 ( .A(x[23]), .B(y[23]), .Z(n926) );
  XOR U1184 ( .A(x[19]), .B(y[19]), .Z(n924) );
  XNOR U1185 ( .A(x[15]), .B(y[15]), .Z(n925) );
  XOR U1186 ( .A(n924), .B(n925), .Z(n927) );
  XNOR U1187 ( .A(n926), .B(n927), .Z(n438) );
  XNOR U1188 ( .A(n439), .B(n438), .Z(n387) );
  XOR U1189 ( .A(n437), .B(n387), .Z(n865) );
  XOR U1190 ( .A(n864), .B(n865), .Z(n388) );
  XOR U1191 ( .A(n866), .B(n388), .Z(n397) );
  XOR U1192 ( .A(x[109]), .B(y[109]), .Z(n555) );
  XOR U1193 ( .A(x[229]), .B(y[229]), .Z(n553) );
  XNOR U1194 ( .A(x[107]), .B(y[107]), .Z(n554) );
  XOR U1195 ( .A(n553), .B(n554), .Z(n556) );
  XOR U1196 ( .A(n555), .B(n556), .Z(n867) );
  XOR U1197 ( .A(x[105]), .B(y[105]), .Z(n739) );
  XOR U1198 ( .A(x[103]), .B(y[103]), .Z(n737) );
  XNOR U1199 ( .A(x[101]), .B(y[101]), .Z(n738) );
  XOR U1200 ( .A(n737), .B(n738), .Z(n740) );
  XNOR U1201 ( .A(n739), .B(n740), .Z(n869) );
  XOR U1202 ( .A(x[113]), .B(y[113]), .Z(n561) );
  XOR U1203 ( .A(x[227]), .B(y[227]), .Z(n559) );
  XNOR U1204 ( .A(x[111]), .B(y[111]), .Z(n560) );
  XOR U1205 ( .A(n559), .B(n560), .Z(n562) );
  XNOR U1206 ( .A(n561), .B(n562), .Z(n868) );
  XOR U1207 ( .A(x[75]), .B(y[75]), .Z(n999) );
  XOR U1208 ( .A(x[73]), .B(y[73]), .Z(n996) );
  XNOR U1209 ( .A(x[71]), .B(y[71]), .Z(n997) );
  XNOR U1210 ( .A(n996), .B(n997), .Z(n998) );
  XNOR U1211 ( .A(n999), .B(n998), .Z(n938) );
  XOR U1212 ( .A(x[81]), .B(y[81]), .Z(n1005) );
  XOR U1213 ( .A(x[79]), .B(y[79]), .Z(n1002) );
  XNOR U1214 ( .A(x[77]), .B(y[77]), .Z(n1003) );
  XNOR U1215 ( .A(n1002), .B(n1003), .Z(n1004) );
  XNOR U1216 ( .A(n1005), .B(n1004), .Z(n937) );
  XOR U1217 ( .A(x[69]), .B(y[69]), .Z(n1048) );
  XOR U1218 ( .A(x[67]), .B(y[67]), .Z(n1045) );
  XNOR U1219 ( .A(x[65]), .B(y[65]), .Z(n1046) );
  XNOR U1220 ( .A(n1045), .B(n1046), .Z(n1047) );
  XOR U1221 ( .A(n1048), .B(n1047), .Z(n936) );
  XOR U1222 ( .A(n937), .B(n936), .Z(n389) );
  XNOR U1223 ( .A(n938), .B(n389), .Z(n470) );
  XOR U1224 ( .A(x[87]), .B(y[87]), .Z(n995) );
  XOR U1225 ( .A(x[85]), .B(y[85]), .Z(n993) );
  XOR U1226 ( .A(x[83]), .B(y[83]), .Z(n992) );
  XOR U1227 ( .A(n993), .B(n992), .Z(n994) );
  XOR U1228 ( .A(n995), .B(n994), .Z(n481) );
  XOR U1229 ( .A(x[99]), .B(y[99]), .Z(n733) );
  XOR U1230 ( .A(x[97]), .B(y[97]), .Z(n731) );
  XNOR U1231 ( .A(x[95]), .B(y[95]), .Z(n732) );
  XOR U1232 ( .A(n731), .B(n732), .Z(n734) );
  XNOR U1233 ( .A(n733), .B(n734), .Z(n480) );
  XOR U1234 ( .A(x[93]), .B(y[93]), .Z(n727) );
  XOR U1235 ( .A(x[91]), .B(y[91]), .Z(n725) );
  XNOR U1236 ( .A(x[89]), .B(y[89]), .Z(n726) );
  XOR U1237 ( .A(n725), .B(n726), .Z(n728) );
  XNOR U1238 ( .A(n727), .B(n728), .Z(n479) );
  XNOR U1239 ( .A(n480), .B(n479), .Z(n390) );
  XNOR U1240 ( .A(n481), .B(n390), .Z(n469) );
  XOR U1241 ( .A(n470), .B(n469), .Z(n391) );
  XOR U1242 ( .A(n471), .B(n391), .Z(n398) );
  XOR U1243 ( .A(n397), .B(n398), .Z(n392) );
  XOR U1244 ( .A(n399), .B(n392), .Z(n1075) );
  XNOR U1245 ( .A(n1074), .B(n1075), .Z(n393) );
  XNOR U1246 ( .A(n1076), .B(n393), .Z(o[0]) );
  XOR U1247 ( .A(n1316), .B(n1317), .Z(n403) );
  XNOR U1248 ( .A(n1318), .B(n403), .Z(n1286) );
  NANDN U1249 ( .A(n414), .B(n413), .Z(n418) );
  NAND U1250 ( .A(n416), .B(n415), .Z(n417) );
  NAND U1251 ( .A(n418), .B(n417), .Z(n1207) );
  NANDN U1252 ( .A(n420), .B(n419), .Z(n424) );
  NAND U1253 ( .A(n422), .B(n421), .Z(n423) );
  NAND U1254 ( .A(n424), .B(n423), .Z(n1206) );
  NANDN U1255 ( .A(n426), .B(n425), .Z(n430) );
  NAND U1256 ( .A(n428), .B(n427), .Z(n429) );
  AND U1257 ( .A(n430), .B(n429), .Z(n1205) );
  XOR U1258 ( .A(n1206), .B(n1205), .Z(n431) );
  XOR U1259 ( .A(n1207), .B(n431), .Z(n1180) );
  IV U1260 ( .A(n1180), .Z(n1179) );
  XOR U1261 ( .A(n1183), .B(n1179), .Z(n432) );
  XOR U1262 ( .A(n1181), .B(n432), .Z(n1368) );
  IV U1263 ( .A(n1368), .Z(n1367) );
  XOR U1264 ( .A(n1367), .B(n1369), .Z(n436) );
  XOR U1265 ( .A(n1370), .B(n436), .Z(n1277) );
  NANDN U1266 ( .A(n444), .B(n443), .Z(n448) );
  NAND U1267 ( .A(n446), .B(n445), .Z(n447) );
  NAND U1268 ( .A(n448), .B(n447), .Z(n1256) );
  NANDN U1269 ( .A(n450), .B(n449), .Z(n454) );
  NAND U1270 ( .A(n452), .B(n451), .Z(n453) );
  NAND U1271 ( .A(n454), .B(n453), .Z(n1255) );
  NANDN U1272 ( .A(n456), .B(n455), .Z(n460) );
  NAND U1273 ( .A(n458), .B(n457), .Z(n459) );
  AND U1274 ( .A(n460), .B(n459), .Z(n1254) );
  XOR U1275 ( .A(n1255), .B(n1254), .Z(n461) );
  XOR U1276 ( .A(n1256), .B(n461), .Z(n1108) );
  IV U1277 ( .A(n1108), .Z(n1107) );
  XOR U1278 ( .A(n1111), .B(n1107), .Z(n462) );
  XOR U1279 ( .A(n1109), .B(n462), .Z(n1273) );
  NANDN U1280 ( .A(n464), .B(n463), .Z(n468) );
  ANDN U1281 ( .B(n464), .A(n463), .Z(n466) );
  OR U1282 ( .A(n466), .B(n465), .Z(n467) );
  AND U1283 ( .A(n468), .B(n467), .Z(n1275) );
  NANDN U1284 ( .A(n470), .B(n469), .Z(n474) );
  ANDN U1285 ( .B(n470), .A(n469), .Z(n472) );
  OR U1286 ( .A(n472), .B(n471), .Z(n473) );
  AND U1287 ( .A(n474), .B(n473), .Z(n1274) );
  XNOR U1288 ( .A(n1275), .B(n1274), .Z(n475) );
  XOR U1289 ( .A(n1273), .B(n475), .Z(n1279) );
  NANDN U1290 ( .A(n483), .B(n482), .Z(n487) );
  NAND U1291 ( .A(n485), .B(n484), .Z(n486) );
  NAND U1292 ( .A(n487), .B(n486), .Z(n1235) );
  NANDN U1293 ( .A(n489), .B(n488), .Z(n493) );
  NAND U1294 ( .A(n491), .B(n490), .Z(n492) );
  AND U1295 ( .A(n493), .B(n492), .Z(n1237) );
  NANDN U1296 ( .A(n495), .B(n494), .Z(n499) );
  NAND U1297 ( .A(n497), .B(n496), .Z(n498) );
  AND U1298 ( .A(n499), .B(n498), .Z(n1236) );
  XOR U1299 ( .A(n1176), .B(n1173), .Z(n500) );
  XOR U1300 ( .A(n1174), .B(n500), .Z(n1363) );
  NANDN U1301 ( .A(n508), .B(n507), .Z(n512) );
  NAND U1302 ( .A(n510), .B(n509), .Z(n511) );
  NAND U1303 ( .A(n512), .B(n511), .Z(n1238) );
  IV U1304 ( .A(n1238), .Z(n526) );
  NANDN U1305 ( .A(n514), .B(n513), .Z(n518) );
  NAND U1306 ( .A(n516), .B(n515), .Z(n517) );
  AND U1307 ( .A(n518), .B(n517), .Z(n1240) );
  NANDN U1308 ( .A(n520), .B(n519), .Z(n524) );
  NAND U1309 ( .A(n522), .B(n521), .Z(n523) );
  AND U1310 ( .A(n524), .B(n523), .Z(n1239) );
  XNOR U1311 ( .A(n1240), .B(n1239), .Z(n525) );
  XOR U1312 ( .A(n526), .B(n525), .Z(n1218) );
  XOR U1313 ( .A(n1220), .B(n1218), .Z(n527) );
  XOR U1314 ( .A(n1219), .B(n527), .Z(n1361) );
  IV U1315 ( .A(n1361), .Z(n1360) );
  NANDN U1316 ( .A(n532), .B(n531), .Z(n536) );
  NANDN U1317 ( .A(n534), .B(n533), .Z(n535) );
  AND U1318 ( .A(n536), .B(n535), .Z(n1201) );
  NANDN U1319 ( .A(n542), .B(n541), .Z(n546) );
  NANDN U1320 ( .A(n544), .B(n543), .Z(n545) );
  NAND U1321 ( .A(n546), .B(n545), .Z(n1199) );
  XNOR U1322 ( .A(n1201), .B(n1200), .Z(n1308) );
  NANDN U1323 ( .A(n548), .B(n547), .Z(n552) );
  NANDN U1324 ( .A(n550), .B(n549), .Z(n551) );
  AND U1325 ( .A(n552), .B(n551), .Z(n1248) );
  NANDN U1326 ( .A(n554), .B(n553), .Z(n558) );
  NANDN U1327 ( .A(n556), .B(n555), .Z(n557) );
  NAND U1328 ( .A(n558), .B(n557), .Z(n1250) );
  NANDN U1329 ( .A(n560), .B(n559), .Z(n564) );
  NANDN U1330 ( .A(n562), .B(n561), .Z(n563) );
  NAND U1331 ( .A(n564), .B(n563), .Z(n1249) );
  XNOR U1332 ( .A(n1250), .B(n1249), .Z(n565) );
  XOR U1333 ( .A(n1248), .B(n565), .Z(n1307) );
  NANDN U1334 ( .A(n567), .B(n566), .Z(n571) );
  NANDN U1335 ( .A(n569), .B(n568), .Z(n570) );
  AND U1336 ( .A(n571), .B(n570), .Z(n1208) );
  NANDN U1337 ( .A(n573), .B(n572), .Z(n577) );
  NANDN U1338 ( .A(n575), .B(n574), .Z(n576) );
  NAND U1339 ( .A(n577), .B(n576), .Z(n1210) );
  NANDN U1340 ( .A(n579), .B(n578), .Z(n583) );
  NANDN U1341 ( .A(n581), .B(n580), .Z(n582) );
  NAND U1342 ( .A(n583), .B(n582), .Z(n1209) );
  XNOR U1343 ( .A(n1210), .B(n1209), .Z(n584) );
  XNOR U1344 ( .A(n1208), .B(n584), .Z(n1306) );
  XOR U1345 ( .A(n1307), .B(n1306), .Z(n585) );
  XNOR U1346 ( .A(n1308), .B(n585), .Z(n1265) );
  NAND U1347 ( .A(n587), .B(n586), .Z(n591) );
  NAND U1348 ( .A(n589), .B(n588), .Z(n590) );
  AND U1349 ( .A(n591), .B(n590), .Z(n1094) );
  NAND U1350 ( .A(n593), .B(n592), .Z(n597) );
  NAND U1351 ( .A(n595), .B(n594), .Z(n596) );
  NAND U1352 ( .A(n597), .B(n596), .Z(n1096) );
  NAND U1353 ( .A(n599), .B(n598), .Z(n603) );
  NAND U1354 ( .A(n601), .B(n600), .Z(n602) );
  NAND U1355 ( .A(n603), .B(n602), .Z(n1095) );
  XNOR U1356 ( .A(n1096), .B(n1095), .Z(n604) );
  XOR U1357 ( .A(n1094), .B(n604), .Z(n1138) );
  NAND U1358 ( .A(n609), .B(n608), .Z(n613) );
  NAND U1359 ( .A(n611), .B(n610), .Z(n612) );
  AND U1360 ( .A(n613), .B(n612), .Z(n1189) );
  NANDN U1361 ( .A(n615), .B(n614), .Z(n619) );
  NAND U1362 ( .A(n617), .B(n616), .Z(n618) );
  AND U1363 ( .A(n619), .B(n618), .Z(n1186) );
  NAND U1364 ( .A(n621), .B(n620), .Z(n625) );
  NAND U1365 ( .A(n623), .B(n622), .Z(n624) );
  NAND U1366 ( .A(n625), .B(n624), .Z(n1187) );
  XOR U1367 ( .A(n1189), .B(n1188), .Z(n1136) );
  IV U1368 ( .A(n1136), .Z(n1135) );
  XOR U1369 ( .A(n1137), .B(n1135), .Z(n626) );
  XOR U1370 ( .A(n1138), .B(n626), .Z(n1264) );
  NANDN U1371 ( .A(n628), .B(n627), .Z(n632) );
  NAND U1372 ( .A(n630), .B(n629), .Z(n631) );
  NAND U1373 ( .A(n632), .B(n631), .Z(n1228) );
  NANDN U1374 ( .A(n634), .B(n633), .Z(n638) );
  NANDN U1375 ( .A(n636), .B(n635), .Z(n637) );
  AND U1376 ( .A(n638), .B(n637), .Z(n1231) );
  NANDN U1377 ( .A(n640), .B(n639), .Z(n644) );
  NANDN U1378 ( .A(n642), .B(n641), .Z(n643) );
  AND U1379 ( .A(n644), .B(n643), .Z(n1229) );
  NANDN U1380 ( .A(n646), .B(n645), .Z(n650) );
  NANDN U1381 ( .A(n648), .B(n647), .Z(n649) );
  NAND U1382 ( .A(n650), .B(n649), .Z(n1194) );
  NANDN U1383 ( .A(n652), .B(n651), .Z(n656) );
  NANDN U1384 ( .A(n654), .B(n653), .Z(n655) );
  NAND U1385 ( .A(n656), .B(n655), .Z(n1193) );
  NANDN U1386 ( .A(n658), .B(n657), .Z(n662) );
  NANDN U1387 ( .A(n660), .B(n659), .Z(n661) );
  AND U1388 ( .A(n662), .B(n661), .Z(n1192) );
  XOR U1389 ( .A(n1193), .B(n1192), .Z(n663) );
  XNOR U1390 ( .A(n1194), .B(n663), .Z(n1297) );
  NANDN U1391 ( .A(n665), .B(n664), .Z(n669) );
  NANDN U1392 ( .A(n667), .B(n666), .Z(n668) );
  NAND U1393 ( .A(n669), .B(n668), .Z(n1213) );
  NANDN U1394 ( .A(n671), .B(n670), .Z(n675) );
  NANDN U1395 ( .A(n673), .B(n672), .Z(n674) );
  NAND U1396 ( .A(n675), .B(n674), .Z(n1212) );
  NANDN U1397 ( .A(n677), .B(n676), .Z(n681) );
  NANDN U1398 ( .A(n679), .B(n678), .Z(n680) );
  AND U1399 ( .A(n681), .B(n680), .Z(n1211) );
  XOR U1400 ( .A(n1212), .B(n1211), .Z(n682) );
  XOR U1401 ( .A(n1213), .B(n682), .Z(n1296) );
  XOR U1402 ( .A(n1297), .B(n1296), .Z(n683) );
  XOR U1403 ( .A(n1298), .B(n683), .Z(n1263) );
  XOR U1404 ( .A(n1264), .B(n1263), .Z(n684) );
  XOR U1405 ( .A(n1265), .B(n684), .Z(n1282) );
  NANDN U1406 ( .A(n686), .B(n685), .Z(n690) );
  NAND U1407 ( .A(n688), .B(n687), .Z(n689) );
  NAND U1408 ( .A(n690), .B(n689), .Z(n1165) );
  NANDN U1409 ( .A(n691), .B(oglobal[0]), .Z(n695) );
  NAND U1410 ( .A(n693), .B(n692), .Z(n694) );
  NAND U1411 ( .A(n695), .B(n694), .Z(n1164) );
  NANDN U1412 ( .A(n697), .B(n696), .Z(n701) );
  NAND U1413 ( .A(n699), .B(n698), .Z(n700) );
  AND U1414 ( .A(n701), .B(n700), .Z(n1163) );
  XOR U1415 ( .A(n1164), .B(n1163), .Z(n702) );
  XOR U1416 ( .A(n1165), .B(n702), .Z(n1144) );
  NAND U1417 ( .A(n704), .B(n703), .Z(n708) );
  NAND U1418 ( .A(n706), .B(n705), .Z(n707) );
  AND U1419 ( .A(n708), .B(n707), .Z(n1100) );
  NAND U1420 ( .A(n710), .B(n709), .Z(n714) );
  NAND U1421 ( .A(n712), .B(n711), .Z(n713) );
  NAND U1422 ( .A(n714), .B(n713), .Z(n1102) );
  NAND U1423 ( .A(n716), .B(n715), .Z(n720) );
  NAND U1424 ( .A(n718), .B(n717), .Z(n719) );
  NAND U1425 ( .A(n720), .B(n719), .Z(n1101) );
  XNOR U1426 ( .A(n1102), .B(n1101), .Z(n721) );
  XOR U1427 ( .A(n1100), .B(n721), .Z(n1142) );
  NANDN U1428 ( .A(n726), .B(n725), .Z(n730) );
  NANDN U1429 ( .A(n728), .B(n727), .Z(n729) );
  NAND U1430 ( .A(n730), .B(n729), .Z(n1253) );
  NANDN U1431 ( .A(n732), .B(n731), .Z(n736) );
  NANDN U1432 ( .A(n734), .B(n733), .Z(n735) );
  NAND U1433 ( .A(n736), .B(n735), .Z(n1252) );
  NANDN U1434 ( .A(n738), .B(n737), .Z(n742) );
  NANDN U1435 ( .A(n740), .B(n739), .Z(n741) );
  AND U1436 ( .A(n742), .B(n741), .Z(n1251) );
  XOR U1437 ( .A(n1252), .B(n1251), .Z(n743) );
  XOR U1438 ( .A(n1253), .B(n743), .Z(n1292) );
  NANDN U1439 ( .A(n748), .B(n747), .Z(n752) );
  NANDN U1440 ( .A(n750), .B(n749), .Z(n751) );
  NAND U1441 ( .A(n752), .B(n751), .Z(n1354) );
  XOR U1442 ( .A(n1354), .B(oglobal[1]), .Z(n1353) );
  NANDN U1443 ( .A(n754), .B(n753), .Z(n758) );
  NAND U1444 ( .A(n756), .B(n755), .Z(n757) );
  NAND U1445 ( .A(n758), .B(n757), .Z(n1352) );
  NANDN U1446 ( .A(n760), .B(n759), .Z(n764) );
  NAND U1447 ( .A(n762), .B(n761), .Z(n763) );
  AND U1448 ( .A(n764), .B(n763), .Z(n1351) );
  XOR U1449 ( .A(n1352), .B(n1351), .Z(n765) );
  XOR U1450 ( .A(n1353), .B(n765), .Z(n1290) );
  XOR U1451 ( .A(n1291), .B(n1290), .Z(n766) );
  XOR U1452 ( .A(n1292), .B(n766), .Z(n1357) );
  NANDN U1453 ( .A(n768), .B(n767), .Z(n772) );
  NAND U1454 ( .A(n770), .B(n769), .Z(n771) );
  NAND U1455 ( .A(n772), .B(n771), .Z(n1241) );
  NANDN U1456 ( .A(n774), .B(n773), .Z(n778) );
  NAND U1457 ( .A(n776), .B(n775), .Z(n777) );
  AND U1458 ( .A(n778), .B(n777), .Z(n1244) );
  NANDN U1459 ( .A(n780), .B(n779), .Z(n784) );
  NAND U1460 ( .A(n782), .B(n781), .Z(n783) );
  AND U1461 ( .A(n784), .B(n783), .Z(n1242) );
  XNOR U1462 ( .A(n1244), .B(n1242), .Z(n785) );
  XOR U1463 ( .A(n1241), .B(n785), .Z(n1131) );
  NAND U1464 ( .A(n787), .B(n786), .Z(n791) );
  NAND U1465 ( .A(n789), .B(n788), .Z(n790) );
  AND U1466 ( .A(n791), .B(n790), .Z(n1348) );
  NAND U1467 ( .A(n793), .B(n792), .Z(n797) );
  NAND U1468 ( .A(n795), .B(n794), .Z(n796) );
  NAND U1469 ( .A(n797), .B(n796), .Z(n1350) );
  NANDN U1470 ( .A(n799), .B(n798), .Z(n803) );
  NAND U1471 ( .A(n801), .B(n800), .Z(n802) );
  NAND U1472 ( .A(n803), .B(n802), .Z(n1349) );
  IV U1473 ( .A(n1128), .Z(n1130) );
  XOR U1474 ( .A(n1130), .B(n1129), .Z(n807) );
  XOR U1475 ( .A(n1131), .B(n807), .Z(n1358) );
  NANDN U1476 ( .A(n809), .B(n808), .Z(n813) );
  NAND U1477 ( .A(n811), .B(n810), .Z(n812) );
  AND U1478 ( .A(n813), .B(n812), .Z(n1153) );
  NANDN U1479 ( .A(n815), .B(n814), .Z(n819) );
  NAND U1480 ( .A(n817), .B(n816), .Z(n818) );
  NAND U1481 ( .A(n819), .B(n818), .Z(n1154) );
  NANDN U1482 ( .A(n821), .B(n820), .Z(n825) );
  NAND U1483 ( .A(n823), .B(n822), .Z(n824) );
  NAND U1484 ( .A(n825), .B(n824), .Z(n1156) );
  IV U1485 ( .A(n1156), .Z(n826) );
  XOR U1486 ( .A(n1155), .B(n826), .Z(n1123) );
  NANDN U1487 ( .A(n828), .B(n827), .Z(n832) );
  NAND U1488 ( .A(n830), .B(n829), .Z(n831) );
  NAND U1489 ( .A(n832), .B(n831), .Z(n1222) );
  NANDN U1490 ( .A(n834), .B(n833), .Z(n838) );
  NAND U1491 ( .A(n836), .B(n835), .Z(n837) );
  AND U1492 ( .A(n838), .B(n837), .Z(n1224) );
  NANDN U1493 ( .A(n840), .B(n839), .Z(n844) );
  NAND U1494 ( .A(n842), .B(n841), .Z(n843) );
  AND U1495 ( .A(n844), .B(n843), .Z(n1223) );
  XNOR U1496 ( .A(n1224), .B(n1223), .Z(n845) );
  XNOR U1497 ( .A(n1222), .B(n845), .Z(n1122) );
  NANDN U1498 ( .A(n847), .B(n846), .Z(n851) );
  NAND U1499 ( .A(n849), .B(n848), .Z(n850) );
  AND U1500 ( .A(n851), .B(n850), .Z(n1147) );
  NANDN U1501 ( .A(n853), .B(n852), .Z(n857) );
  NAND U1502 ( .A(n855), .B(n854), .Z(n856) );
  NAND U1503 ( .A(n857), .B(n856), .Z(n1148) );
  NANDN U1504 ( .A(n859), .B(n858), .Z(n863) );
  NAND U1505 ( .A(n861), .B(n860), .Z(n862) );
  NAND U1506 ( .A(n863), .B(n862), .Z(n1150) );
  NANDN U1507 ( .A(n871), .B(n870), .Z(n875) );
  ANDN U1508 ( .B(n871), .A(n870), .Z(n872) );
  OR U1509 ( .A(n873), .B(n872), .Z(n874) );
  AND U1510 ( .A(n875), .B(n874), .Z(n1341) );
  NANDN U1511 ( .A(n877), .B(n876), .Z(n881) );
  NAND U1512 ( .A(n879), .B(n878), .Z(n880) );
  NAND U1513 ( .A(n881), .B(n880), .Z(n1225) );
  IV U1514 ( .A(n1225), .Z(n895) );
  NANDN U1515 ( .A(n883), .B(n882), .Z(n887) );
  NAND U1516 ( .A(n885), .B(n884), .Z(n886) );
  AND U1517 ( .A(n887), .B(n886), .Z(n1227) );
  NANDN U1518 ( .A(n889), .B(n888), .Z(n893) );
  NAND U1519 ( .A(n891), .B(n890), .Z(n892) );
  AND U1520 ( .A(n893), .B(n892), .Z(n1226) );
  XNOR U1521 ( .A(n1227), .B(n1226), .Z(n894) );
  XOR U1522 ( .A(n895), .B(n894), .Z(n1339) );
  XOR U1523 ( .A(n1341), .B(n1339), .Z(n896) );
  XOR U1524 ( .A(n1340), .B(n896), .Z(n1331) );
  IV U1525 ( .A(n1331), .Z(n1329) );
  XOR U1526 ( .A(n1330), .B(n1329), .Z(n897) );
  XNOR U1527 ( .A(n1332), .B(n897), .Z(n1280) );
  NAND U1528 ( .A(n905), .B(n904), .Z(n909) );
  NAND U1529 ( .A(n907), .B(n906), .Z(n908) );
  AND U1530 ( .A(n909), .B(n908), .Z(n1087) );
  NANDN U1531 ( .A(n919), .B(n918), .Z(n923) );
  NANDN U1532 ( .A(n921), .B(n920), .Z(n922) );
  AND U1533 ( .A(n923), .B(n922), .Z(n1169) );
  NANDN U1534 ( .A(n925), .B(n924), .Z(n929) );
  NANDN U1535 ( .A(n927), .B(n926), .Z(n928) );
  AND U1536 ( .A(n929), .B(n928), .Z(n1167) );
  NANDN U1537 ( .A(n931), .B(n930), .Z(n935) );
  NANDN U1538 ( .A(n933), .B(n932), .Z(n934) );
  NAND U1539 ( .A(n935), .B(n934), .Z(n1166) );
  XNOR U1540 ( .A(n1312), .B(n1309), .Z(n939) );
  XOR U1541 ( .A(n1310), .B(n939), .Z(n1376) );
  IV U1542 ( .A(n1376), .Z(n1374) );
  XOR U1543 ( .A(n1375), .B(n1374), .Z(n940) );
  XNOR U1544 ( .A(n1377), .B(n940), .Z(n1321) );
  NANDN U1545 ( .A(n945), .B(n944), .Z(n949) );
  ANDN U1546 ( .B(n945), .A(n944), .Z(n947) );
  OR U1547 ( .A(n947), .B(n946), .Z(n948) );
  AND U1548 ( .A(n949), .B(n948), .Z(n1120) );
  XOR U1549 ( .A(n1120), .B(n1119), .Z(n953) );
  XOR U1550 ( .A(n1118), .B(n953), .Z(n1345) );
  XNOR U1551 ( .A(n1343), .B(n1342), .Z(n960) );
  XOR U1552 ( .A(n1345), .B(n960), .Z(n1338) );
  NANDN U1553 ( .A(n965), .B(n964), .Z(n969) );
  ANDN U1554 ( .B(n965), .A(n964), .Z(n966) );
  OR U1555 ( .A(n967), .B(n966), .Z(n968) );
  AND U1556 ( .A(n969), .B(n968), .Z(n1117) );
  XOR U1557 ( .A(n1117), .B(n1116), .Z(n973) );
  XNOR U1558 ( .A(n1115), .B(n973), .Z(n1337) );
  OR U1559 ( .A(n975), .B(n974), .Z(n979) );
  AND U1560 ( .A(n975), .B(n974), .Z(n976) );
  OR U1561 ( .A(n977), .B(n976), .Z(n978) );
  AND U1562 ( .A(n979), .B(n978), .Z(n1299) );
  OR U1563 ( .A(n981), .B(n980), .Z(n986) );
  AND U1564 ( .A(n981), .B(n980), .Z(n984) );
  IV U1565 ( .A(n982), .Z(n983) );
  NANDN U1566 ( .A(n984), .B(n983), .Z(n985) );
  AND U1567 ( .A(n986), .B(n985), .Z(n1301) );
  XOR U1568 ( .A(n1301), .B(n1300), .Z(n990) );
  XOR U1569 ( .A(n1299), .B(n990), .Z(n1336) );
  XOR U1570 ( .A(n1337), .B(n1336), .Z(n991) );
  XOR U1571 ( .A(n1338), .B(n991), .Z(n1320) );
  NANDN U1572 ( .A(n997), .B(n996), .Z(n1001) );
  NAND U1573 ( .A(n999), .B(n998), .Z(n1000) );
  AND U1574 ( .A(n1001), .B(n1000), .Z(n1161) );
  NANDN U1575 ( .A(n1003), .B(n1002), .Z(n1007) );
  NAND U1576 ( .A(n1005), .B(n1004), .Z(n1006) );
  AND U1577 ( .A(n1007), .B(n1006), .Z(n1160) );
  XNOR U1578 ( .A(n1161), .B(n1160), .Z(n1008) );
  XOR U1579 ( .A(n1159), .B(n1008), .Z(n1305) );
  NAND U1580 ( .A(n1010), .B(n1009), .Z(n1014) );
  NAND U1581 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U1582 ( .A(n1014), .B(n1013), .Z(n1092) );
  NAND U1583 ( .A(n1016), .B(n1015), .Z(n1020) );
  NAND U1584 ( .A(n1018), .B(n1017), .Z(n1019) );
  NAND U1585 ( .A(n1020), .B(n1019), .Z(n1093) );
  NAND U1586 ( .A(n1022), .B(n1021), .Z(n1026) );
  NAND U1587 ( .A(n1024), .B(n1023), .Z(n1025) );
  AND U1588 ( .A(n1026), .B(n1025), .Z(n1091) );
  XOR U1589 ( .A(n1093), .B(n1091), .Z(n1027) );
  XOR U1590 ( .A(n1092), .B(n1027), .Z(n1304) );
  XNOR U1591 ( .A(n1304), .B(n1303), .Z(n1031) );
  XOR U1592 ( .A(n1305), .B(n1031), .Z(n1269) );
  NAND U1593 ( .A(n1036), .B(n1035), .Z(n1040) );
  NAND U1594 ( .A(n1038), .B(n1037), .Z(n1039) );
  NAND U1595 ( .A(n1040), .B(n1039), .Z(n1080) );
  NANDN U1596 ( .A(n1046), .B(n1045), .Z(n1050) );
  NAND U1597 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U1598 ( .A(n1050), .B(n1049), .Z(n1078) );
  XOR U1599 ( .A(n1079), .B(n1078), .Z(n1051) );
  XOR U1600 ( .A(n1080), .B(n1051), .Z(n1295) );
  NAND U1601 ( .A(n1057), .B(n1056), .Z(n1061) );
  NAND U1602 ( .A(n1059), .B(n1058), .Z(n1060) );
  NAND U1603 ( .A(n1061), .B(n1060), .Z(n1085) );
  XOR U1604 ( .A(n1085), .B(n1084), .Z(n1066) );
  XOR U1605 ( .A(n1086), .B(n1066), .Z(n1294) );
  XNOR U1606 ( .A(n1294), .B(n1293), .Z(n1070) );
  XOR U1607 ( .A(n1295), .B(n1070), .Z(n1266) );
  IV U1608 ( .A(n1266), .Z(n1268) );
  XOR U1609 ( .A(n1267), .B(n1268), .Z(n1071) );
  XOR U1610 ( .A(n1269), .B(n1071), .Z(n1319) );
  XNOR U1611 ( .A(n1320), .B(n1319), .Z(n1072) );
  XOR U1612 ( .A(n1321), .B(n1072), .Z(n1326) );
  XNOR U1613 ( .A(n1328), .B(n1326), .Z(n1073) );
  XOR U1614 ( .A(n1327), .B(n1073), .Z(n1285) );
  IV U1615 ( .A(n1285), .Z(n1283) );
  XOR U1616 ( .A(n1283), .B(n1284), .Z(n1077) );
  XNOR U1617 ( .A(n1286), .B(n1077), .Z(o[1]) );
  NANDN U1618 ( .A(n1079), .B(n1078), .Z(n1083) );
  ANDN U1619 ( .B(n1079), .A(n1078), .Z(n1081) );
  OR U1620 ( .A(n1081), .B(n1080), .Z(n1082) );
  AND U1621 ( .A(n1083), .B(n1082), .Z(n1423) );
  XOR U1622 ( .A(n1425), .B(n1424), .Z(n1090) );
  XOR U1623 ( .A(n1423), .B(n1090), .Z(n1402) );
  NANDN U1624 ( .A(n1095), .B(n1094), .Z(n1099) );
  ANDN U1625 ( .B(n1095), .A(n1094), .Z(n1097) );
  OR U1626 ( .A(n1097), .B(n1096), .Z(n1098) );
  AND U1627 ( .A(n1099), .B(n1098), .Z(n1467) );
  NANDN U1628 ( .A(n1101), .B(n1100), .Z(n1105) );
  ANDN U1629 ( .B(n1101), .A(n1100), .Z(n1103) );
  OR U1630 ( .A(n1103), .B(n1102), .Z(n1104) );
  AND U1631 ( .A(n1105), .B(n1104), .Z(n1466) );
  XNOR U1632 ( .A(n1467), .B(n1466), .Z(n1106) );
  XNOR U1633 ( .A(n1465), .B(n1106), .Z(n1403) );
  OR U1634 ( .A(n1109), .B(n1107), .Z(n1113) );
  ANDN U1635 ( .B(n1109), .A(n1108), .Z(n1110) );
  OR U1636 ( .A(n1111), .B(n1110), .Z(n1112) );
  AND U1637 ( .A(n1113), .B(n1112), .Z(n1401) );
  XNOR U1638 ( .A(n1403), .B(n1401), .Z(n1114) );
  XOR U1639 ( .A(n1402), .B(n1114), .Z(n1440) );
  NANDN U1640 ( .A(n1122), .B(n1121), .Z(n1126) );
  ANDN U1641 ( .B(n1122), .A(n1121), .Z(n1124) );
  NANDN U1642 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U1643 ( .A(n1126), .B(n1125), .Z(n1501) );
  XOR U1644 ( .A(n1502), .B(n1501), .Z(n1127) );
  XOR U1645 ( .A(n1500), .B(n1127), .Z(n1438) );
  IV U1646 ( .A(n1438), .Z(n1437) );
  NANDN U1647 ( .A(n1128), .B(n1129), .Z(n1134) );
  NOR U1648 ( .A(n1130), .B(n1129), .Z(n1132) );
  OR U1649 ( .A(n1132), .B(n1131), .Z(n1133) );
  AND U1650 ( .A(n1134), .B(n1133), .Z(n1410) );
  OR U1651 ( .A(n1137), .B(n1135), .Z(n1141) );
  ANDN U1652 ( .B(n1137), .A(n1136), .Z(n1139) );
  OR U1653 ( .A(n1139), .B(n1138), .Z(n1140) );
  AND U1654 ( .A(n1141), .B(n1140), .Z(n1409) );
  XNOR U1655 ( .A(n1409), .B(n1408), .Z(n1145) );
  XNOR U1656 ( .A(n1410), .B(n1145), .Z(n1439) );
  XOR U1657 ( .A(n1437), .B(n1439), .Z(n1146) );
  XOR U1658 ( .A(n1440), .B(n1146), .Z(n1454) );
  NANDN U1659 ( .A(n1148), .B(n1147), .Z(n1152) );
  NANDN U1660 ( .A(n1150), .B(n1149), .Z(n1151) );
  AND U1661 ( .A(n1152), .B(n1151), .Z(n1468) );
  NANDN U1662 ( .A(n1154), .B(n1153), .Z(n1158) );
  NANDN U1663 ( .A(n1156), .B(n1155), .Z(n1157) );
  NAND U1664 ( .A(n1158), .B(n1157), .Z(n1470) );
  XOR U1665 ( .A(n1470), .B(n1469), .Z(n1162) );
  XOR U1666 ( .A(n1468), .B(n1162), .Z(n1420) );
  IV U1667 ( .A(n1420), .Z(n1172) );
  NANDN U1668 ( .A(n1167), .B(n1166), .Z(n1171) );
  NANDN U1669 ( .A(n1169), .B(n1168), .Z(n1170) );
  AND U1670 ( .A(n1171), .B(n1170), .Z(n1417) );
  XNOR U1671 ( .A(n1418), .B(n1417), .Z(n1419) );
  XOR U1672 ( .A(n1172), .B(n1419), .Z(n1508) );
  OR U1673 ( .A(n1174), .B(n1173), .Z(n1178) );
  AND U1674 ( .A(n1174), .B(n1173), .Z(n1175) );
  OR U1675 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1676 ( .A(n1178), .B(n1177), .Z(n1507) );
  OR U1677 ( .A(n1181), .B(n1179), .Z(n1185) );
  ANDN U1678 ( .B(n1181), .A(n1180), .Z(n1182) );
  OR U1679 ( .A(n1183), .B(n1182), .Z(n1184) );
  AND U1680 ( .A(n1185), .B(n1184), .Z(n1506) );
  NANDN U1681 ( .A(n1187), .B(n1186), .Z(n1191) );
  NAND U1682 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U1683 ( .A(n1191), .B(n1190), .Z(n1480) );
  NANDN U1684 ( .A(n1193), .B(n1192), .Z(n1197) );
  ANDN U1685 ( .B(n1193), .A(n1192), .Z(n1195) );
  OR U1686 ( .A(n1195), .B(n1194), .Z(n1196) );
  AND U1687 ( .A(n1197), .B(n1196), .Z(n1478) );
  NANDN U1688 ( .A(n1199), .B(n1198), .Z(n1203) );
  NAND U1689 ( .A(n1201), .B(n1200), .Z(n1202) );
  NAND U1690 ( .A(n1203), .B(n1202), .Z(n1479) );
  XOR U1691 ( .A(n1478), .B(n1479), .Z(n1204) );
  XOR U1692 ( .A(n1480), .B(n1204), .Z(n1504) );
  NANDN U1693 ( .A(n1212), .B(n1211), .Z(n1216) );
  ANDN U1694 ( .B(n1212), .A(n1211), .Z(n1214) );
  OR U1695 ( .A(n1214), .B(n1213), .Z(n1215) );
  AND U1696 ( .A(n1216), .B(n1215), .Z(n1483) );
  XNOR U1697 ( .A(n1484), .B(n1483), .Z(n1217) );
  XNOR U1698 ( .A(n1482), .B(n1217), .Z(n1505) );
  XNOR U1699 ( .A(n1505), .B(n1503), .Z(n1221) );
  XOR U1700 ( .A(n1504), .B(n1221), .Z(n1457) );
  NANDN U1701 ( .A(n1229), .B(n1228), .Z(n1233) );
  ANDN U1702 ( .B(n1229), .A(n1228), .Z(n1230) );
  OR U1703 ( .A(n1231), .B(n1230), .Z(n1232) );
  AND U1704 ( .A(n1233), .B(n1232), .Z(n1475) );
  XOR U1705 ( .A(n1476), .B(n1475), .Z(n1234) );
  XNOR U1706 ( .A(n1474), .B(n1234), .Z(n1407) );
  NANDN U1707 ( .A(n1242), .B(n1241), .Z(n1246) );
  ANDN U1708 ( .B(n1242), .A(n1241), .Z(n1243) );
  OR U1709 ( .A(n1244), .B(n1243), .Z(n1245) );
  AND U1710 ( .A(n1246), .B(n1245), .Z(n1472) );
  XNOR U1711 ( .A(n1473), .B(n1472), .Z(n1247) );
  XOR U1712 ( .A(n1471), .B(n1247), .Z(n1406) );
  NANDN U1713 ( .A(n1255), .B(n1254), .Z(n1259) );
  ANDN U1714 ( .B(n1255), .A(n1254), .Z(n1257) );
  OR U1715 ( .A(n1257), .B(n1256), .Z(n1258) );
  AND U1716 ( .A(n1259), .B(n1258), .Z(n1415) );
  XNOR U1717 ( .A(n1416), .B(n1415), .Z(n1260) );
  XOR U1718 ( .A(n1414), .B(n1260), .Z(n1405) );
  IV U1719 ( .A(n1405), .Z(n1261) );
  XOR U1720 ( .A(n1406), .B(n1261), .Z(n1262) );
  XOR U1721 ( .A(n1407), .B(n1262), .Z(n1456) );
  NANDN U1722 ( .A(n1266), .B(n1267), .Z(n1272) );
  NOR U1723 ( .A(n1268), .B(n1267), .Z(n1270) );
  OR U1724 ( .A(n1270), .B(n1269), .Z(n1271) );
  AND U1725 ( .A(n1272), .B(n1271), .Z(n1445) );
  XNOR U1726 ( .A(n1445), .B(n1444), .Z(n1276) );
  XNOR U1727 ( .A(n1446), .B(n1276), .Z(n1452) );
  XNOR U1728 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U1729 ( .A(n1431), .B(n1430), .Z(n1387) );
  NANDN U1730 ( .A(n1283), .B(n1284), .Z(n1289) );
  NOR U1731 ( .A(n1285), .B(n1284), .Z(n1287) );
  OR U1732 ( .A(n1287), .B(n1286), .Z(n1288) );
  AND U1733 ( .A(n1289), .B(n1288), .Z(n1385) );
  XNOR U1734 ( .A(n1399), .B(n1398), .Z(n1302) );
  XNOR U1735 ( .A(n1400), .B(n1302), .Z(n1494) );
  XNOR U1736 ( .A(n1495), .B(n1494), .Z(n1496) );
  NANDN U1737 ( .A(n1310), .B(n1309), .Z(n1314) );
  ANDN U1738 ( .B(n1310), .A(n1309), .Z(n1311) );
  OR U1739 ( .A(n1312), .B(n1311), .Z(n1313) );
  AND U1740 ( .A(n1314), .B(n1313), .Z(n1411) );
  XNOR U1741 ( .A(n1412), .B(n1411), .Z(n1315) );
  XOR U1742 ( .A(n1413), .B(n1315), .Z(n1497) );
  NANDN U1743 ( .A(n1320), .B(n1319), .Z(n1324) );
  ANDN U1744 ( .B(n1320), .A(n1319), .Z(n1322) );
  OR U1745 ( .A(n1322), .B(n1321), .Z(n1323) );
  AND U1746 ( .A(n1324), .B(n1323), .Z(n1523) );
  XNOR U1747 ( .A(n1521), .B(n1523), .Z(n1325) );
  XOR U1748 ( .A(n1522), .B(n1325), .Z(n1391) );
  NANDN U1749 ( .A(n1329), .B(n1330), .Z(n1335) );
  NOR U1750 ( .A(n1331), .B(n1330), .Z(n1333) );
  OR U1751 ( .A(n1333), .B(n1332), .Z(n1334) );
  AND U1752 ( .A(n1335), .B(n1334), .Z(n1462) );
  OR U1753 ( .A(n1343), .B(n1342), .Z(n1347) );
  AND U1754 ( .A(n1343), .B(n1342), .Z(n1344) );
  OR U1755 ( .A(n1345), .B(n1344), .Z(n1346) );
  AND U1756 ( .A(n1347), .B(n1346), .Z(n1397) );
  AND U1757 ( .A(oglobal[1]), .B(n1354), .Z(n1477) );
  XOR U1758 ( .A(oglobal[2]), .B(n1477), .Z(n1485) );
  IV U1759 ( .A(n1485), .Z(n1486) );
  XOR U1760 ( .A(n1489), .B(n1486), .Z(n1355) );
  XOR U1761 ( .A(n1487), .B(n1355), .Z(n1395) );
  XOR U1762 ( .A(n1397), .B(n1395), .Z(n1356) );
  XNOR U1763 ( .A(n1396), .B(n1356), .Z(n1459) );
  XOR U1764 ( .A(n1460), .B(n1459), .Z(n1461) );
  IV U1765 ( .A(n1514), .Z(n1515) );
  OR U1766 ( .A(n1362), .B(n1360), .Z(n1366) );
  ANDN U1767 ( .B(n1362), .A(n1361), .Z(n1364) );
  NANDN U1768 ( .A(n1364), .B(n1363), .Z(n1365) );
  AND U1769 ( .A(n1366), .B(n1365), .Z(n1434) );
  OR U1770 ( .A(n1369), .B(n1367), .Z(n1373) );
  ANDN U1771 ( .B(n1369), .A(n1368), .Z(n1371) );
  NANDN U1772 ( .A(n1371), .B(n1370), .Z(n1372) );
  AND U1773 ( .A(n1373), .B(n1372), .Z(n1436) );
  NANDN U1774 ( .A(n1374), .B(n1375), .Z(n1380) );
  NOR U1775 ( .A(n1376), .B(n1375), .Z(n1378) );
  NANDN U1776 ( .A(n1378), .B(n1377), .Z(n1379) );
  AND U1777 ( .A(n1380), .B(n1379), .Z(n1435) );
  XNOR U1778 ( .A(n1436), .B(n1435), .Z(n1381) );
  XNOR U1779 ( .A(n1434), .B(n1381), .Z(n1517) );
  XNOR U1780 ( .A(n1516), .B(n1517), .Z(n1382) );
  XOR U1781 ( .A(n1515), .B(n1382), .Z(n1388) );
  IV U1782 ( .A(n1388), .Z(n1389) );
  XOR U1783 ( .A(n1390), .B(n1389), .Z(n1383) );
  XOR U1784 ( .A(n1391), .B(n1383), .Z(n1386) );
  XOR U1785 ( .A(n1385), .B(n1386), .Z(n1384) );
  XNOR U1786 ( .A(n1387), .B(n1384), .Z(o[2]) );
  OR U1787 ( .A(n1390), .B(n1388), .Z(n1394) );
  ANDN U1788 ( .B(n1390), .A(n1389), .Z(n1392) );
  OR U1789 ( .A(n1392), .B(n1391), .Z(n1393) );
  AND U1790 ( .A(n1394), .B(n1393), .Z(n1533) );
  XOR U1791 ( .A(n1566), .B(n1565), .Z(n1404) );
  XNOR U1792 ( .A(n1564), .B(n1404), .Z(n1542) );
  NANDN U1793 ( .A(n1418), .B(n1417), .Z(n1422) );
  NANDN U1794 ( .A(n1420), .B(n1419), .Z(n1421) );
  NAND U1795 ( .A(n1422), .B(n1421), .Z(n1548) );
  XOR U1796 ( .A(n1548), .B(n1549), .Z(n1550) );
  XOR U1797 ( .A(n1573), .B(n1571), .Z(n1426) );
  XOR U1798 ( .A(n1572), .B(n1426), .Z(n1541) );
  IV U1799 ( .A(n1541), .Z(n1539) );
  XOR U1800 ( .A(n1540), .B(n1539), .Z(n1427) );
  XNOR U1801 ( .A(n1542), .B(n1427), .Z(n1537) );
  NANDN U1802 ( .A(n1429), .B(n1428), .Z(n1433) );
  NAND U1803 ( .A(n1431), .B(n1430), .Z(n1432) );
  AND U1804 ( .A(n1433), .B(n1432), .Z(n1538) );
  OR U1805 ( .A(n1439), .B(n1437), .Z(n1443) );
  ANDN U1806 ( .B(n1439), .A(n1438), .Z(n1441) );
  OR U1807 ( .A(n1441), .B(n1440), .Z(n1442) );
  AND U1808 ( .A(n1443), .B(n1442), .Z(n1588) );
  OR U1809 ( .A(n1445), .B(n1444), .Z(n1449) );
  AND U1810 ( .A(n1445), .B(n1444), .Z(n1447) );
  NANDN U1811 ( .A(n1447), .B(n1446), .Z(n1448) );
  AND U1812 ( .A(n1449), .B(n1448), .Z(n1587) );
  XNOR U1813 ( .A(n1588), .B(n1587), .Z(n1450) );
  XOR U1814 ( .A(n1589), .B(n1450), .Z(n1536) );
  XOR U1815 ( .A(n1538), .B(n1536), .Z(n1451) );
  XNOR U1816 ( .A(n1537), .B(n1451), .Z(n1535) );
  XNOR U1817 ( .A(n1535), .B(n1534), .Z(n1455) );
  XNOR U1818 ( .A(n1533), .B(n1455), .Z(n1530) );
  NANDN U1819 ( .A(n1460), .B(n1459), .Z(n1464) );
  OR U1820 ( .A(n1462), .B(n1461), .Z(n1463) );
  NAND U1821 ( .A(n1464), .B(n1463), .Z(n1581) );
  XNOR U1822 ( .A(n1582), .B(n1581), .Z(n1584) );
  XOR U1823 ( .A(n1559), .B(n1558), .Z(n1560) );
  XNOR U1824 ( .A(n1561), .B(n1560), .Z(n1576) );
  AND U1825 ( .A(n1477), .B(oglobal[2]), .Z(n1547) );
  XNOR U1826 ( .A(oglobal[3]), .B(n1546), .Z(n1481) );
  XOR U1827 ( .A(n1547), .B(n1481), .Z(n1557) );
  OR U1828 ( .A(n1487), .B(n1485), .Z(n1491) );
  ANDN U1829 ( .B(n1487), .A(n1486), .Z(n1488) );
  OR U1830 ( .A(n1489), .B(n1488), .Z(n1490) );
  AND U1831 ( .A(n1491), .B(n1490), .Z(n1555) );
  XNOR U1832 ( .A(n1556), .B(n1555), .Z(n1492) );
  XOR U1833 ( .A(n1557), .B(n1492), .Z(n1574) );
  XOR U1834 ( .A(n1576), .B(n1574), .Z(n1493) );
  XOR U1835 ( .A(n1575), .B(n1493), .Z(n1579) );
  NANDN U1836 ( .A(n1495), .B(n1494), .Z(n1499) );
  NANDN U1837 ( .A(n1497), .B(n1496), .Z(n1498) );
  NAND U1838 ( .A(n1499), .B(n1498), .Z(n1580) );
  OR U1839 ( .A(n1507), .B(n1506), .Z(n1511) );
  AND U1840 ( .A(n1507), .B(n1506), .Z(n1509) );
  NANDN U1841 ( .A(n1509), .B(n1508), .Z(n1510) );
  AND U1842 ( .A(n1511), .B(n1510), .Z(n1568) );
  XNOR U1843 ( .A(n1569), .B(n1568), .Z(n1512) );
  XNOR U1844 ( .A(n1567), .B(n1512), .Z(n1578) );
  XOR U1845 ( .A(n1580), .B(n1578), .Z(n1513) );
  XOR U1846 ( .A(n1579), .B(n1513), .Z(n1583) );
  XNOR U1847 ( .A(n1584), .B(n1583), .Z(n1593) );
  OR U1848 ( .A(n1516), .B(n1514), .Z(n1520) );
  ANDN U1849 ( .B(n1516), .A(n1515), .Z(n1518) );
  OR U1850 ( .A(n1518), .B(n1517), .Z(n1519) );
  AND U1851 ( .A(n1520), .B(n1519), .Z(n1592) );
  XNOR U1852 ( .A(n1592), .B(n1591), .Z(n1524) );
  XOR U1853 ( .A(n1593), .B(n1524), .Z(n1527) );
  IV U1854 ( .A(n1527), .Z(n1526) );
  XOR U1855 ( .A(n1530), .B(n1526), .Z(n1525) );
  XNOR U1856 ( .A(n1528), .B(n1525), .Z(o[3]) );
  OR U1857 ( .A(n1528), .B(n1526), .Z(n1532) );
  ANDN U1858 ( .B(n1528), .A(n1527), .Z(n1529) );
  OR U1859 ( .A(n1530), .B(n1529), .Z(n1531) );
  AND U1860 ( .A(n1532), .B(n1531), .Z(n1598) );
  NANDN U1861 ( .A(n1539), .B(n1540), .Z(n1545) );
  NOR U1862 ( .A(n1541), .B(n1540), .Z(n1543) );
  OR U1863 ( .A(n1543), .B(n1542), .Z(n1544) );
  AND U1864 ( .A(n1545), .B(n1544), .Z(n1607) );
  NANDN U1865 ( .A(n1549), .B(n1548), .Z(n1553) );
  OR U1866 ( .A(n1551), .B(n1550), .Z(n1552) );
  NAND U1867 ( .A(n1553), .B(n1552), .Z(n1627) );
  XOR U1868 ( .A(n1627), .B(oglobal[4]), .Z(n1554) );
  XOR U1869 ( .A(n1628), .B(n1554), .Z(n1623) );
  OR U1870 ( .A(n1559), .B(n1558), .Z(n1563) );
  NANDN U1871 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1872 ( .A(n1563), .B(n1562), .Z(n1621) );
  XOR U1873 ( .A(n1622), .B(n1621), .Z(n1624) );
  XNOR U1874 ( .A(n1620), .B(n1619), .Z(n1570) );
  XOR U1875 ( .A(n1618), .B(n1570), .Z(n1617) );
  XNOR U1876 ( .A(n1616), .B(n1615), .Z(n1577) );
  XNOR U1877 ( .A(n1617), .B(n1577), .Z(n1606) );
  XOR U1878 ( .A(n1607), .B(n1606), .Z(n1608) );
  NANDN U1879 ( .A(n1582), .B(n1581), .Z(n1586) );
  NAND U1880 ( .A(n1584), .B(n1583), .Z(n1585) );
  AND U1881 ( .A(n1586), .B(n1585), .Z(n1614) );
  XNOR U1882 ( .A(n1614), .B(n1613), .Z(n1590) );
  XOR U1883 ( .A(n1612), .B(n1590), .Z(n1603) );
  XOR U1884 ( .A(n1603), .B(n1604), .Z(n1594) );
  XOR U1885 ( .A(n1605), .B(n1594), .Z(n1597) );
  IV U1886 ( .A(n1597), .Z(n1596) );
  XOR U1887 ( .A(n1600), .B(n1596), .Z(n1595) );
  XNOR U1888 ( .A(n1598), .B(n1595), .Z(o[4]) );
  OR U1889 ( .A(n1598), .B(n1596), .Z(n1602) );
  ANDN U1890 ( .B(n1598), .A(n1597), .Z(n1599) );
  OR U1891 ( .A(n1600), .B(n1599), .Z(n1601) );
  AND U1892 ( .A(n1602), .B(n1601), .Z(n1648) );
  NANDN U1893 ( .A(n1607), .B(n1606), .Z(n1611) );
  OR U1894 ( .A(n1609), .B(n1608), .Z(n1610) );
  NAND U1895 ( .A(n1611), .B(n1610), .Z(n1642) );
  XOR U1896 ( .A(n1634), .B(n1633), .Z(n1636) );
  NANDN U1897 ( .A(n1622), .B(n1621), .Z(n1626) );
  NANDN U1898 ( .A(n1624), .B(n1623), .Z(n1625) );
  AND U1899 ( .A(n1626), .B(n1625), .Z(n1632) );
  XNOR U1900 ( .A(oglobal[5]), .B(n1631), .Z(n1629) );
  XOR U1901 ( .A(n1632), .B(n1629), .Z(n1635) );
  XNOR U1902 ( .A(n1636), .B(n1635), .Z(n1640) );
  XOR U1903 ( .A(n1641), .B(n1640), .Z(n1643) );
  IV U1904 ( .A(n1647), .Z(n1646) );
  XOR U1905 ( .A(n1650), .B(n1646), .Z(n1630) );
  XNOR U1906 ( .A(n1648), .B(n1630), .Z(o[5]) );
  OR U1907 ( .A(n1634), .B(n1633), .Z(n1638) );
  NAND U1908 ( .A(n1636), .B(n1635), .Z(n1637) );
  NAND U1909 ( .A(n1638), .B(n1637), .Z(n1654) );
  XOR U1910 ( .A(oglobal[6]), .B(n1654), .Z(n1639) );
  XOR U1911 ( .A(n1655), .B(n1639), .Z(n1657) );
  IV U1912 ( .A(n1657), .Z(n1656) );
  NANDN U1913 ( .A(n1641), .B(n1640), .Z(n1645) );
  NANDN U1914 ( .A(n1643), .B(n1642), .Z(n1644) );
  AND U1915 ( .A(n1645), .B(n1644), .Z(n1660) );
  OR U1916 ( .A(n1648), .B(n1646), .Z(n1652) );
  ANDN U1917 ( .B(n1648), .A(n1647), .Z(n1649) );
  OR U1918 ( .A(n1650), .B(n1649), .Z(n1651) );
  AND U1919 ( .A(n1652), .B(n1651), .Z(n1658) );
  XNOR U1920 ( .A(n1660), .B(n1658), .Z(n1653) );
  XOR U1921 ( .A(n1656), .B(n1653), .Z(o[6]) );
  OR U1922 ( .A(n1658), .B(n1656), .Z(n1662) );
  ANDN U1923 ( .B(n1658), .A(n1657), .Z(n1659) );
  OR U1924 ( .A(n1660), .B(n1659), .Z(n1661) );
  AND U1925 ( .A(n1662), .B(n1661), .Z(n1665) );
  XOR U1926 ( .A(n1664), .B(n1665), .Z(n1663) );
  XNOR U1927 ( .A(oglobal[7]), .B(n1663), .Z(o[7]) );
  XNOR U1928 ( .A(n1666), .B(oglobal[8]), .Z(o[8]) );
  ANDN U1929 ( .B(oglobal[8]), .A(n1666), .Z(n1667) );
  XOR U1930 ( .A(n1667), .B(oglobal[9]), .Z(o[9]) );
  AND U1931 ( .A(n1667), .B(oglobal[9]), .Z(n1668) );
  XOR U1932 ( .A(n1668), .B(oglobal[10]), .Z(o[10]) );
  AND U1933 ( .A(n1668), .B(oglobal[10]), .Z(n1669) );
  XOR U1934 ( .A(n1669), .B(oglobal[11]), .Z(o[11]) );
  AND U1935 ( .A(n1669), .B(oglobal[11]), .Z(n1670) );
  XOR U1936 ( .A(oglobal[12]), .B(n1670), .Z(o[12]) );
endmodule

