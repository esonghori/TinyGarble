
module Lite_MIPS ( clk, rst, inst_mem_in_wire, data_mem_in_wire, 
        data_mem_out_wire );
  input [2047:0] inst_mem_in_wire;
  input [2047:0] data_mem_in_wire;
  output [2047:0] data_mem_out_wire;
  input clk, rst;
  wire   N24, N25, N26, N27, N28, N29, \PC_Next/n311 , \PC_Next/n310 ,
         \PC_Next/n309 , \PC_Next/n308 , \PC_Next/N45 , \PC_Next/N44 ,
         \PC_Next/N43 , \PC_Next/N42 , \PC_Next/N41 , \PC_Next/N40 ,
         \PC_Next/N39 , \PC_Next/N38 , \PC_Next/N37 , \PC_Next/N36 ,
         \PC_Next/N35 , \PC_Next/N34 , \PC_Next/N33 , \PC_Next/N32 ,
         \PC_Next/N31 , \PC_Next/N30 , \PC_Next/N29 , \PC_Next/N28 ,
         \PC_Next/N27 , \PC_Next/N26 , \PC_Next/N25 , \PC_Next/N24 ,
         \PC_Next/N23 , \PC_Next/N22 , \PC_Next/N21 , \PC_Next/N20 ,
         \PC_Next/N19 , \PC_Next/N18 , \PC_Next/N17 , \PC_Next/N16 ,
         \PC_Next/pc_future[27] , \PC_Next/pc_future[26] ,
         \PC_Next/pc_future[25] , \PC_Next/pc_future[24] ,
         \PC_Next/pc_future[23] , \PC_Next/pc_future[22] ,
         \PC_Next/pc_future[21] , \PC_Next/pc_future[20] ,
         \PC_Next/pc_future[19] , \PC_Next/pc_future[18] ,
         \PC_Next/pc_future[17] , \PC_Next/pc_future[16] ,
         \PC_Next/pc_future[15] , \PC_Next/pc_future[14] ,
         \PC_Next/pc_future[13] , \PC_Next/pc_future[12] ,
         \PC_Next/pc_future[11] , \PC_Next/pc_future[10] ,
         \PC_Next/pc_future[9] , \PC_Next/pc_future[8] ,
         \PC_Next/pc_future[7] , \PC_Next/pc_future[6] ,
         \PC_Next/pc_future[5] , \PC_Next/pc_future[4] ,
         \PC_Next/pc_future[3] , \PC_Next/pc_future[2] , \Inst_Mem/n1984 ,
         \Inst_Mem/n1983 , \Inst_Mem/n1982 , \Inst_Mem/n1981 ,
         \Inst_Mem/n1980 , \Inst_Mem/n1979 , \Inst_Mem/n1978 ,
         \Inst_Mem/n1977 , \Inst_Mem/n1976 , \Inst_Mem/n1975 ,
         \Inst_Mem/n1974 , \Inst_Mem/n1973 , \Inst_Mem/n1972 ,
         \Inst_Mem/n1971 , \Inst_Mem/n1970 , \Inst_Mem/n1969 ,
         \Inst_Mem/n1968 , \Inst_Mem/n1967 , \Inst_Mem/n1966 ,
         \Inst_Mem/n1965 , \Inst_Mem/n1964 , \Inst_Mem/n1963 ,
         \Inst_Mem/n1962 , \Inst_Mem/n1961 , \Inst_Mem/n1960 ,
         \Inst_Mem/n1959 , \Inst_Mem/n1958 , \Inst_Mem/n1957 ,
         \Inst_Mem/n1956 , \Inst_Mem/n1955 , \Inst_Mem/n1954 ,
         \Inst_Mem/n1953 , \Inst_Mem/n1952 , \Inst_Mem/n1951 ,
         \Inst_Mem/n1950 , \Inst_Mem/n1949 , \Inst_Mem/n1948 ,
         \Inst_Mem/n1947 , \Inst_Mem/n1946 , \Inst_Mem/n1945 ,
         \Inst_Mem/n1944 , \Inst_Mem/n1943 , \Inst_Mem/n1942 ,
         \Inst_Mem/n1941 , \Inst_Mem/n1940 , \Inst_Mem/n1939 ,
         \Inst_Mem/n1938 , \Inst_Mem/n1937 , \Inst_Mem/n1936 ,
         \Inst_Mem/n1935 , \Inst_Mem/n1934 , \Inst_Mem/n1933 ,
         \Inst_Mem/n1932 , \Inst_Mem/n1931 , \Inst_Mem/n1930 ,
         \Inst_Mem/n1929 , \Inst_Mem/n1928 , \Inst_Mem/n1927 ,
         \Inst_Mem/n1926 , \Inst_Mem/n1925 , \Inst_Mem/n1924 ,
         \Inst_Mem/n1923 , \Inst_Mem/n1922 , \Inst_Mem/n1921 ,
         \Inst_Mem/n1920 , \Inst_Mem/n1919 , \Inst_Mem/n1918 ,
         \Inst_Mem/n1917 , \Inst_Mem/n1916 , \Inst_Mem/n1915 ,
         \Inst_Mem/n1914 , \Inst_Mem/n1913 , \Inst_Mem/n1912 ,
         \Inst_Mem/n1911 , \Inst_Mem/n1910 , \Inst_Mem/n1909 ,
         \Inst_Mem/n1908 , \Inst_Mem/n1907 , \Inst_Mem/n1906 ,
         \Inst_Mem/n1905 , \Inst_Mem/n1904 , \Inst_Mem/n1903 ,
         \Inst_Mem/n1902 , \Inst_Mem/n1901 , \Inst_Mem/n1900 ,
         \Inst_Mem/n1899 , \Inst_Mem/n1898 , \Inst_Mem/n1897 ,
         \Inst_Mem/n1896 , \Inst_Mem/n1895 , \Inst_Mem/n1894 ,
         \Inst_Mem/n1893 , \Inst_Mem/n1892 , \Inst_Mem/n1891 ,
         \Inst_Mem/n1890 , \Inst_Mem/n1889 , \Inst_Mem/n1888 ,
         \Inst_Mem/n1887 , \Inst_Mem/n1886 , \Inst_Mem/n1885 ,
         \Inst_Mem/n1884 , \Inst_Mem/n1883 , \Inst_Mem/n1882 ,
         \Inst_Mem/n1881 , \Inst_Mem/n1880 , \Inst_Mem/n1879 ,
         \Inst_Mem/n1878 , \Inst_Mem/n1877 , \Inst_Mem/n1876 ,
         \Inst_Mem/n1875 , \Inst_Mem/n1874 , \Inst_Mem/n1873 ,
         \Inst_Mem/n1872 , \Inst_Mem/n1871 , \Inst_Mem/n1870 ,
         \Inst_Mem/n1869 , \Inst_Mem/n1868 , \Inst_Mem/n1867 ,
         \Inst_Mem/n1866 , \Inst_Mem/n1865 , \Inst_Mem/n1864 ,
         \Inst_Mem/n1863 , \Inst_Mem/n1862 , \Inst_Mem/n1861 ,
         \Inst_Mem/n1860 , \Inst_Mem/n1859 , \Inst_Mem/n1858 ,
         \Inst_Mem/n1857 , \Inst_Mem/n1856 , \Inst_Mem/n1855 ,
         \Inst_Mem/n1854 , \Inst_Mem/n1853 , \Inst_Mem/n1852 ,
         \Inst_Mem/n1851 , \Inst_Mem/n1850 , \Inst_Mem/n1849 ,
         \Inst_Mem/n1848 , \Inst_Mem/n1847 , \Inst_Mem/n1846 ,
         \Inst_Mem/n1845 , \Inst_Mem/n1844 , \Inst_Mem/n1843 ,
         \Inst_Mem/n1842 , \Inst_Mem/n1841 , \Inst_Mem/n1840 ,
         \Inst_Mem/n1839 , \Inst_Mem/n1838 , \Inst_Mem/n1837 ,
         \Inst_Mem/n1836 , \Inst_Mem/n1835 , \Inst_Mem/n1834 ,
         \Inst_Mem/n1833 , \Inst_Mem/n1832 , \Inst_Mem/n1831 ,
         \Inst_Mem/n1830 , \Inst_Mem/n1829 , \Inst_Mem/n1828 ,
         \Inst_Mem/n1827 , \Inst_Mem/n1826 , \Inst_Mem/n1825 ,
         \Inst_Mem/n1824 , \Inst_Mem/n1823 , \Inst_Mem/n1822 ,
         \Inst_Mem/n1821 , \Inst_Mem/n1820 , \Inst_Mem/n1819 ,
         \Inst_Mem/n1818 , \Inst_Mem/n1817 , \Inst_Mem/n1816 ,
         \Inst_Mem/n1815 , \Inst_Mem/n1814 , \Inst_Mem/n1813 ,
         \Inst_Mem/n1812 , \Inst_Mem/n1811 , \Inst_Mem/n1810 ,
         \Inst_Mem/n1809 , \Inst_Mem/n1808 , \Inst_Mem/n1807 ,
         \Inst_Mem/n1806 , \Inst_Mem/n1805 , \Inst_Mem/n1804 ,
         \Inst_Mem/n1803 , \Inst_Mem/n1802 , \Inst_Mem/n1801 ,
         \Inst_Mem/n1800 , \Inst_Mem/n1799 , \Inst_Mem/n1798 ,
         \Inst_Mem/n1797 , \Inst_Mem/n1796 , \Inst_Mem/n1795 ,
         \Inst_Mem/n1794 , \Inst_Mem/n1793 , \Inst_Mem/n1792 ,
         \Inst_Mem/n1791 , \Inst_Mem/n1790 , \Inst_Mem/n1789 ,
         \Inst_Mem/n1788 , \Inst_Mem/n1787 , \Inst_Mem/n1786 ,
         \Inst_Mem/n1785 , \Inst_Mem/n1784 , \Inst_Mem/n1783 ,
         \Inst_Mem/n1782 , \Inst_Mem/n1781 , \Inst_Mem/n1780 ,
         \Inst_Mem/n1779 , \Inst_Mem/n1778 , \Inst_Mem/n1777 ,
         \Inst_Mem/n1776 , \Inst_Mem/n1775 , \Inst_Mem/n1774 ,
         \Inst_Mem/n1773 , \Inst_Mem/n1772 , \Inst_Mem/n1771 ,
         \Inst_Mem/n1770 , \Inst_Mem/n1769 , \Inst_Mem/n1768 ,
         \Inst_Mem/n1767 , \Inst_Mem/n1766 , \Inst_Mem/n1765 ,
         \Inst_Mem/n1764 , \Inst_Mem/n1763 , \Inst_Mem/n1762 ,
         \Inst_Mem/n1761 , \Inst_Mem/n1760 , \Inst_Mem/n1759 ,
         \Inst_Mem/n1758 , \Inst_Mem/n1757 , \Inst_Mem/n1756 ,
         \Inst_Mem/n1755 , \Inst_Mem/n1754 , \Inst_Mem/n1753 ,
         \Inst_Mem/n1752 , \Inst_Mem/n1751 , \Inst_Mem/n1750 ,
         \Inst_Mem/n1749 , \Inst_Mem/n1748 , \Inst_Mem/n1747 ,
         \Inst_Mem/n1746 , \Inst_Mem/n1745 , \Inst_Mem/n1744 ,
         \Inst_Mem/n1743 , \Inst_Mem/n1742 , \Inst_Mem/n1741 ,
         \Inst_Mem/n1740 , \Inst_Mem/n1739 , \Inst_Mem/n1738 ,
         \Inst_Mem/n1737 , \Inst_Mem/n1736 , \Inst_Mem/n1735 ,
         \Inst_Mem/n1734 , \Inst_Mem/n1733 , \Inst_Mem/n1732 ,
         \Inst_Mem/n1731 , \Inst_Mem/n1730 , \Inst_Mem/n1729 ,
         \Inst_Mem/n1728 , \Inst_Mem/n1727 , \Inst_Mem/n1726 ,
         \Inst_Mem/n1725 , \Inst_Mem/n1724 , \Inst_Mem/n1723 ,
         \Inst_Mem/n1722 , \Inst_Mem/n1721 , \Inst_Mem/n1720 ,
         \Inst_Mem/n1719 , \Inst_Mem/n1718 , \Inst_Mem/n1717 ,
         \Inst_Mem/n1716 , \Inst_Mem/n1715 , \Inst_Mem/n1714 ,
         \Inst_Mem/n1713 , \Inst_Mem/n1712 , \Inst_Mem/n1711 ,
         \Inst_Mem/n1710 , \Inst_Mem/n1709 , \Inst_Mem/n1708 ,
         \Inst_Mem/n1707 , \Inst_Mem/n1706 , \Inst_Mem/n1705 ,
         \Inst_Mem/n1704 , \Inst_Mem/n1703 , \Inst_Mem/n1702 ,
         \Inst_Mem/n1701 , \Inst_Mem/n1700 , \Inst_Mem/n1699 ,
         \Inst_Mem/n1698 , \Inst_Mem/n1697 , \Inst_Mem/n1696 ,
         \Inst_Mem/n1695 , \Inst_Mem/n1694 , \Inst_Mem/n1693 ,
         \Inst_Mem/n1692 , \Inst_Mem/n1691 , \Inst_Mem/n1690 ,
         \Inst_Mem/n1689 , \Inst_Mem/n1688 , \Inst_Mem/n1687 ,
         \Inst_Mem/n1686 , \Inst_Mem/n1685 , \Inst_Mem/n1684 ,
         \Inst_Mem/n1683 , \Inst_Mem/n1682 , \Inst_Mem/n1681 ,
         \Inst_Mem/n1680 , \Inst_Mem/n1679 , \Inst_Mem/n1678 ,
         \Inst_Mem/n1677 , \Inst_Mem/n1676 , \Inst_Mem/n1675 ,
         \Inst_Mem/n1674 , \Inst_Mem/n1673 , \Inst_Mem/n1672 ,
         \Inst_Mem/n1671 , \Inst_Mem/n1670 , \Inst_Mem/n1669 ,
         \Inst_Mem/n1668 , \Inst_Mem/n1667 , \Inst_Mem/n1666 ,
         \Inst_Mem/n1665 , \Inst_Mem/n1664 , \Inst_Mem/n1663 ,
         \Inst_Mem/n1662 , \Inst_Mem/n1661 , \Inst_Mem/n1660 ,
         \Inst_Mem/n1659 , \Inst_Mem/n1658 , \Inst_Mem/n1657 ,
         \Inst_Mem/n1656 , \Inst_Mem/n1655 , \Inst_Mem/n1654 ,
         \Inst_Mem/n1653 , \Inst_Mem/n1652 , \Inst_Mem/n1651 ,
         \Inst_Mem/n1650 , \Inst_Mem/n1649 , \Inst_Mem/n1648 ,
         \Inst_Mem/n1647 , \Inst_Mem/n1646 , \Inst_Mem/n1645 ,
         \Inst_Mem/n1644 , \Inst_Mem/n1643 , \Inst_Mem/n1642 ,
         \Inst_Mem/n1641 , \Inst_Mem/n1640 , \Inst_Mem/n1639 ,
         \Inst_Mem/n1638 , \Inst_Mem/n1637 , \Inst_Mem/n1636 ,
         \Inst_Mem/n1635 , \Inst_Mem/n1634 , \Inst_Mem/n1633 ,
         \Inst_Mem/n1632 , \Inst_Mem/n1631 , \Inst_Mem/n1630 ,
         \Inst_Mem/n1629 , \Inst_Mem/n1628 , \Inst_Mem/n1627 ,
         \Inst_Mem/n1626 , \Inst_Mem/n1625 , \Inst_Mem/n1624 ,
         \Inst_Mem/n1623 , \Inst_Mem/n1622 , \Inst_Mem/n1621 ,
         \Inst_Mem/n1620 , \Inst_Mem/n1619 , \Inst_Mem/n1618 ,
         \Inst_Mem/n1617 , \Inst_Mem/n1616 , \Inst_Mem/n1615 ,
         \Inst_Mem/n1614 , \Inst_Mem/n1613 , \Inst_Mem/n1612 ,
         \Inst_Mem/n1611 , \Inst_Mem/n1610 , \Inst_Mem/n1609 ,
         \Inst_Mem/n1608 , \Inst_Mem/n1607 , \Inst_Mem/n1606 ,
         \Inst_Mem/n1605 , \Inst_Mem/n1604 , \Inst_Mem/n1603 ,
         \Inst_Mem/n1602 , \Inst_Mem/n1601 , \Inst_Mem/n1600 ,
         \Inst_Mem/n1599 , \Inst_Mem/n1598 , \Inst_Mem/n1597 ,
         \Inst_Mem/n1596 , \Inst_Mem/n1595 , \Inst_Mem/n1594 ,
         \Inst_Mem/n1593 , \Inst_Mem/n1592 , \Inst_Mem/n1591 ,
         \Inst_Mem/n1590 , \Inst_Mem/n1589 , \Inst_Mem/n1588 ,
         \Inst_Mem/n1587 , \Inst_Mem/n1586 , \Inst_Mem/n1585 ,
         \Inst_Mem/n1584 , \Inst_Mem/n1583 , \Inst_Mem/n1582 ,
         \Inst_Mem/n1581 , \Inst_Mem/n1580 , \Inst_Mem/n1579 ,
         \Inst_Mem/n1578 , \Inst_Mem/n1577 , \Inst_Mem/n1576 ,
         \Inst_Mem/n1575 , \Inst_Mem/n1574 , \Inst_Mem/n1573 ,
         \Inst_Mem/n1572 , \Inst_Mem/n1571 , \Inst_Mem/n1570 ,
         \Inst_Mem/n1569 , \Inst_Mem/n1568 , \Inst_Mem/n1567 ,
         \Inst_Mem/n1566 , \Inst_Mem/n1565 , \Inst_Mem/n1564 ,
         \Inst_Mem/n1563 , \Inst_Mem/n1562 , \Inst_Mem/n1561 ,
         \Inst_Mem/n1560 , \Inst_Mem/n1559 , \Inst_Mem/n1558 ,
         \Inst_Mem/n1557 , \Inst_Mem/n1556 , \Inst_Mem/n1555 ,
         \Inst_Mem/n1554 , \Inst_Mem/n1553 , \Inst_Mem/n1552 ,
         \Inst_Mem/n1551 , \Inst_Mem/n1550 , \Inst_Mem/n1549 ,
         \Inst_Mem/n1548 , \Inst_Mem/n1547 , \Inst_Mem/n1546 ,
         \Inst_Mem/n1545 , \Inst_Mem/n1544 , \Inst_Mem/n1543 ,
         \Inst_Mem/n1542 , \Inst_Mem/n1541 , \Inst_Mem/n1540 ,
         \Inst_Mem/n1539 , \Inst_Mem/n1538 , \Inst_Mem/n1537 ,
         \Inst_Mem/n1536 , \Inst_Mem/n1535 , \Inst_Mem/n1534 ,
         \Inst_Mem/n1533 , \Inst_Mem/n1532 , \Inst_Mem/n1531 ,
         \Inst_Mem/n1530 , \Inst_Mem/n1529 , \Inst_Mem/n1528 ,
         \Inst_Mem/n1527 , \Inst_Mem/n1526 , \Inst_Mem/n1525 ,
         \Inst_Mem/n1524 , \Inst_Mem/n1523 , \Inst_Mem/n1522 ,
         \Inst_Mem/n1521 , \Inst_Mem/n1520 , \Inst_Mem/n1519 ,
         \Inst_Mem/n1518 , \Inst_Mem/n1517 , \Inst_Mem/n1516 ,
         \Inst_Mem/n1515 , \Inst_Mem/n1514 , \Inst_Mem/n1513 ,
         \Inst_Mem/n1512 , \Inst_Mem/n1511 , \Inst_Mem/n1510 ,
         \Inst_Mem/n1509 , \Inst_Mem/n1508 , \Inst_Mem/n1507 ,
         \Inst_Mem/n1506 , \Inst_Mem/n1505 , \Inst_Mem/n1504 ,
         \Inst_Mem/n1503 , \Inst_Mem/n1502 , \Inst_Mem/n1501 ,
         \Inst_Mem/n1500 , \Inst_Mem/n1499 , \Inst_Mem/n1498 ,
         \Inst_Mem/n1497 , \Inst_Mem/n1496 , \Inst_Mem/n1495 ,
         \Inst_Mem/n1494 , \Inst_Mem/n1493 , \Inst_Mem/n1492 ,
         \Inst_Mem/n1491 , \Inst_Mem/n1490 , \Inst_Mem/n1489 ,
         \Inst_Mem/n1488 , \Inst_Mem/n1487 , \Inst_Mem/n1486 ,
         \Inst_Mem/n1485 , \Inst_Mem/n1484 , \Inst_Mem/n1483 ,
         \Inst_Mem/n1482 , \Inst_Mem/n1481 , \Inst_Mem/n1480 ,
         \Inst_Mem/n1479 , \Inst_Mem/n1478 , \Inst_Mem/n1477 ,
         \Inst_Mem/n1476 , \Inst_Mem/n1475 , \Inst_Mem/n1474 ,
         \Inst_Mem/n1473 , \Inst_Mem/n1472 , \Inst_Mem/n1471 ,
         \Inst_Mem/n1470 , \Inst_Mem/n1469 , \Inst_Mem/n1468 ,
         \Inst_Mem/n1467 , \Inst_Mem/n1466 , \Inst_Mem/n1465 ,
         \Inst_Mem/n1464 , \Inst_Mem/n1463 , \Inst_Mem/n1462 ,
         \Inst_Mem/n1461 , \Inst_Mem/n1460 , \Inst_Mem/n1459 ,
         \Inst_Mem/n1458 , \Inst_Mem/n1457 , \Inst_Mem/n1456 ,
         \Inst_Mem/n1455 , \Inst_Mem/n1454 , \Inst_Mem/n1453 ,
         \Inst_Mem/n1452 , \Inst_Mem/n1451 , \Inst_Mem/n1450 ,
         \Inst_Mem/n1449 , \Inst_Mem/n1448 , \Inst_Mem/n1447 ,
         \Inst_Mem/n1446 , \Inst_Mem/n1445 , \Inst_Mem/n1444 ,
         \Inst_Mem/n1443 , \Inst_Mem/n1442 , \Inst_Mem/n1441 ,
         \Inst_Mem/n1440 , \Inst_Mem/n1439 , \Inst_Mem/n1438 ,
         \Inst_Mem/n1437 , \Inst_Mem/n1436 , \Inst_Mem/n1435 ,
         \Inst_Mem/n1434 , \Inst_Mem/n1433 , \Inst_Mem/n1432 ,
         \Inst_Mem/n1431 , \Inst_Mem/n1430 , \Inst_Mem/n1429 ,
         \Inst_Mem/n1428 , \Inst_Mem/n1427 , \Inst_Mem/n1426 ,
         \Inst_Mem/n1425 , \Inst_Mem/n1424 , \Inst_Mem/n1423 ,
         \Inst_Mem/n1422 , \Inst_Mem/n1421 , \Inst_Mem/n1420 ,
         \Inst_Mem/n1419 , \Inst_Mem/n1418 , \Inst_Mem/n1417 ,
         \Inst_Mem/n1416 , \Inst_Mem/n1415 , \Inst_Mem/n1414 ,
         \Inst_Mem/n1413 , \Inst_Mem/n1412 , \Inst_Mem/n1411 ,
         \Inst_Mem/n1410 , \Inst_Mem/n1409 , \Inst_Mem/n1408 ,
         \Inst_Mem/n1407 , \Inst_Mem/n1406 , \Inst_Mem/n1405 ,
         \Inst_Mem/n1404 , \Inst_Mem/n1403 , \Inst_Mem/n1402 ,
         \Inst_Mem/n1401 , \Inst_Mem/n1400 , \Inst_Mem/n1399 ,
         \Inst_Mem/n1398 , \Inst_Mem/n1397 , \Inst_Mem/n1396 ,
         \Inst_Mem/n1395 , \Inst_Mem/n1394 , \Inst_Mem/n1393 ,
         \Inst_Mem/n1392 , \Inst_Mem/n1391 , \Inst_Mem/n1390 ,
         \Inst_Mem/n1389 , \Inst_Mem/n1388 , \Inst_Mem/n1387 ,
         \Inst_Mem/n1386 , \Inst_Mem/n1385 , \Inst_Mem/n1384 ,
         \Inst_Mem/n1383 , \Inst_Mem/n1382 , \Inst_Mem/n1381 ,
         \Inst_Mem/n1380 , \Inst_Mem/n1379 , \Inst_Mem/n1378 ,
         \Inst_Mem/n1377 , \Inst_Mem/n1376 , \Inst_Mem/n1375 ,
         \Inst_Mem/n1374 , \Inst_Mem/n1373 , \Inst_Mem/n1372 ,
         \Inst_Mem/n1371 , \Inst_Mem/n1370 , \Inst_Mem/n1369 ,
         \Inst_Mem/n1368 , \Inst_Mem/n1367 , \Inst_Mem/n1366 ,
         \Inst_Mem/n1365 , \Inst_Mem/n1364 , \Inst_Mem/n1363 ,
         \Inst_Mem/n1362 , \Inst_Mem/n1361 , \Inst_Mem/n1360 ,
         \Inst_Mem/n1359 , \Inst_Mem/n1358 , \Inst_Mem/n1357 ,
         \Inst_Mem/n1356 , \Inst_Mem/n1355 , \Inst_Mem/n1354 ,
         \Inst_Mem/n1353 , \Inst_Mem/n1352 , \Inst_Mem/n1351 ,
         \Inst_Mem/n1350 , \Inst_Mem/n1349 , \Inst_Mem/n1348 ,
         \Inst_Mem/n1347 , \Inst_Mem/n1346 , \Inst_Mem/n1345 ,
         \Inst_Mem/n1344 , \Inst_Mem/n1343 , \Inst_Mem/n1342 ,
         \Inst_Mem/n1341 , \Inst_Mem/n1340 , \Inst_Mem/n1339 ,
         \Inst_Mem/n1338 , \Inst_Mem/n1337 , \Inst_Mem/n1336 ,
         \Inst_Mem/n1335 , \Inst_Mem/n1334 , \Inst_Mem/n1333 ,
         \Inst_Mem/n1332 , \Inst_Mem/n1331 , \Inst_Mem/n1330 ,
         \Inst_Mem/n1329 , \Inst_Mem/n1328 , \Inst_Mem/n1327 ,
         \Inst_Mem/n1326 , \Inst_Mem/n1325 , \Inst_Mem/n1324 ,
         \Inst_Mem/n1323 , \Inst_Mem/n1322 , \Inst_Mem/n1321 ,
         \Inst_Mem/n1320 , \Inst_Mem/n1319 , \Inst_Mem/n1318 ,
         \Inst_Mem/n1317 , \Inst_Mem/n1316 , \Inst_Mem/n1315 ,
         \Inst_Mem/n1314 , \Inst_Mem/n1313 , \Inst_Mem/n1312 ,
         \Inst_Mem/n1311 , \Inst_Mem/n1310 , \Inst_Mem/n1309 ,
         \Inst_Mem/n1308 , \Inst_Mem/n1307 , \Inst_Mem/n1306 ,
         \Inst_Mem/n1305 , \Inst_Mem/n1304 , \Inst_Mem/n1303 ,
         \Inst_Mem/n1302 , \Inst_Mem/n1301 , \Inst_Mem/n1300 ,
         \Inst_Mem/n1299 , \Inst_Mem/n1298 , \Inst_Mem/n1297 ,
         \Inst_Mem/n1296 , \Inst_Mem/n1295 , \Inst_Mem/n1294 ,
         \Inst_Mem/n1293 , \Inst_Mem/n1292 , \Inst_Mem/n1291 ,
         \Inst_Mem/n1290 , \Inst_Mem/n1289 , \Inst_Mem/n1288 ,
         \Inst_Mem/n1287 , \Inst_Mem/n1286 , \Inst_Mem/n1285 ,
         \Inst_Mem/n1284 , \Inst_Mem/n1283 , \Inst_Mem/n1282 ,
         \Inst_Mem/n1281 , \Inst_Mem/n1280 , \Inst_Mem/n1279 ,
         \Inst_Mem/n1278 , \Inst_Mem/n1277 , \Inst_Mem/n1276 ,
         \Inst_Mem/n1275 , \Inst_Mem/n1274 , \Inst_Mem/n1273 ,
         \Inst_Mem/n1272 , \Inst_Mem/n1271 , \Inst_Mem/n1270 ,
         \Inst_Mem/n1269 , \Inst_Mem/n1268 , \Inst_Mem/n1267 ,
         \Inst_Mem/n1266 , \Inst_Mem/n1265 , \Inst_Mem/n1264 ,
         \Inst_Mem/n1263 , \Inst_Mem/n1262 , \Inst_Mem/n1261 ,
         \Inst_Mem/n1260 , \Inst_Mem/n1259 , \Inst_Mem/n1258 ,
         \Inst_Mem/n1257 , \Inst_Mem/n1256 , \Inst_Mem/n1255 ,
         \Inst_Mem/n1254 , \Inst_Mem/n1253 , \Inst_Mem/n1252 ,
         \Inst_Mem/n1251 , \Inst_Mem/n1250 , \Inst_Mem/n1249 ,
         \Inst_Mem/n1248 , \Inst_Mem/n1247 , \Inst_Mem/n1246 ,
         \Inst_Mem/n1245 , \Inst_Mem/n1244 , \Inst_Mem/n1243 ,
         \Inst_Mem/n1242 , \Inst_Mem/n1241 , \Inst_Mem/n1240 ,
         \Inst_Mem/n1239 , \Inst_Mem/n1238 , \Inst_Mem/n1237 ,
         \Inst_Mem/n1236 , \Inst_Mem/n1235 , \Inst_Mem/n1234 ,
         \Inst_Mem/n1233 , \Inst_Mem/n1232 , \Inst_Mem/n1231 ,
         \Inst_Mem/n1230 , \Inst_Mem/n1229 , \Inst_Mem/n1228 ,
         \Inst_Mem/n1227 , \Inst_Mem/n1226 , \Inst_Mem/n1225 ,
         \Inst_Mem/n1224 , \Inst_Mem/n1223 , \Inst_Mem/n1222 ,
         \Inst_Mem/n1221 , \Inst_Mem/n1220 , \Inst_Mem/n1219 ,
         \Inst_Mem/n1218 , \Inst_Mem/n1217 , \Inst_Mem/n1216 ,
         \Inst_Mem/n1215 , \Inst_Mem/n1214 , \Inst_Mem/n1213 ,
         \Inst_Mem/n1212 , \Inst_Mem/n1211 , \Inst_Mem/n1210 ,
         \Inst_Mem/n1209 , \Inst_Mem/n1208 , \Inst_Mem/n1207 ,
         \Inst_Mem/n1206 , \Inst_Mem/n1205 , \Inst_Mem/n1204 ,
         \Inst_Mem/n1203 , \Inst_Mem/n1202 , \Inst_Mem/n1201 ,
         \Inst_Mem/n1200 , \Inst_Mem/n1199 , \Inst_Mem/n1198 ,
         \Inst_Mem/n1197 , \Inst_Mem/n1196 , \Inst_Mem/n1195 ,
         \Inst_Mem/n1194 , \Inst_Mem/n1193 , \Inst_Mem/n1192 ,
         \Inst_Mem/n1191 , \Inst_Mem/n1190 , \Inst_Mem/n1189 ,
         \Inst_Mem/n1188 , \Inst_Mem/n1187 , \Inst_Mem/n1186 ,
         \Inst_Mem/n1185 , \Inst_Mem/n1184 , \Inst_Mem/n1183 ,
         \Inst_Mem/n1182 , \Inst_Mem/n1181 , \Inst_Mem/n1180 ,
         \Inst_Mem/n1179 , \Inst_Mem/n1178 , \Inst_Mem/n1177 ,
         \Inst_Mem/n1176 , \Inst_Mem/n1175 , \Inst_Mem/n1174 ,
         \Inst_Mem/n1173 , \Inst_Mem/n1172 , \Inst_Mem/n1171 ,
         \Inst_Mem/n1170 , \Inst_Mem/n1169 , \Inst_Mem/n1168 ,
         \Inst_Mem/n1167 , \Inst_Mem/n1166 , \Inst_Mem/n1165 ,
         \Inst_Mem/n1164 , \Inst_Mem/n1163 , \Inst_Mem/n1162 ,
         \Inst_Mem/n1161 , \Inst_Mem/n1160 , \Inst_Mem/n1159 ,
         \Inst_Mem/n1158 , \Inst_Mem/n1157 , \Inst_Mem/n1156 ,
         \Inst_Mem/n1155 , \Inst_Mem/n1154 , \Inst_Mem/n1153 ,
         \Inst_Mem/n1152 , \Inst_Mem/n1151 , \Inst_Mem/n1150 ,
         \Inst_Mem/n1149 , \Inst_Mem/n1148 , \Inst_Mem/n1147 ,
         \Inst_Mem/n1146 , \Inst_Mem/n1145 , \Inst_Mem/n1144 ,
         \Inst_Mem/n1143 , \Inst_Mem/n1142 , \Inst_Mem/n1141 ,
         \Inst_Mem/n1140 , \Inst_Mem/n1139 , \Inst_Mem/n1138 ,
         \Inst_Mem/n1137 , \Inst_Mem/n1136 , \Inst_Mem/n1135 ,
         \Inst_Mem/n1134 , \Inst_Mem/n1133 , \Inst_Mem/n1132 ,
         \Inst_Mem/n1131 , \Inst_Mem/n1130 , \Inst_Mem/n1129 ,
         \Inst_Mem/n1128 , \Inst_Mem/n1127 , \Inst_Mem/n1126 ,
         \Inst_Mem/n1125 , \Inst_Mem/n1124 , \Inst_Mem/n1123 ,
         \Inst_Mem/n1122 , \Inst_Mem/n1121 , \Inst_Mem/n1120 ,
         \Inst_Mem/n1119 , \Inst_Mem/n1118 , \Inst_Mem/n1117 ,
         \Inst_Mem/n1116 , \Inst_Mem/n1115 , \Inst_Mem/n1114 ,
         \Inst_Mem/n1113 , \Inst_Mem/n1112 , \Inst_Mem/n1111 ,
         \Inst_Mem/n1110 , \Inst_Mem/n1109 , \Inst_Mem/n1108 ,
         \Inst_Mem/n1107 , \Inst_Mem/n1106 , \Inst_Mem/n1105 ,
         \Inst_Mem/n1104 , \Inst_Mem/n1103 , \Inst_Mem/n1102 ,
         \Inst_Mem/n1101 , \Inst_Mem/n1100 , \Inst_Mem/n1099 ,
         \Inst_Mem/n1098 , \Inst_Mem/n1097 , \Inst_Mem/n1096 ,
         \Inst_Mem/n1095 , \Inst_Mem/n1094 , \Inst_Mem/n1093 ,
         \Inst_Mem/n1092 , \Inst_Mem/n1091 , \Inst_Mem/n1090 ,
         \Inst_Mem/n1089 , \Inst_Mem/n1088 , \Inst_Mem/n1087 ,
         \Inst_Mem/n1086 , \Inst_Mem/n1085 , \Inst_Mem/n1084 ,
         \Inst_Mem/n1083 , \Inst_Mem/n1082 , \Inst_Mem/n1081 ,
         \Inst_Mem/n1080 , \Inst_Mem/n1079 , \Inst_Mem/n1078 ,
         \Inst_Mem/n1077 , \Inst_Mem/n1076 , \Inst_Mem/n1075 ,
         \Inst_Mem/n1074 , \Inst_Mem/n1073 , \Inst_Mem/n1072 ,
         \Inst_Mem/n1071 , \Inst_Mem/n1070 , \Inst_Mem/n1069 ,
         \Inst_Mem/n1068 , \Inst_Mem/n1067 , \Inst_Mem/n1066 ,
         \Inst_Mem/n1065 , \Inst_Mem/n1064 , \Inst_Mem/n1063 ,
         \Inst_Mem/n1062 , \Inst_Mem/n1061 , \Inst_Mem/n1060 ,
         \Inst_Mem/n1059 , \Inst_Mem/n1058 , \Inst_Mem/n1057 ,
         \Inst_Mem/n1056 , \Inst_Mem/n1055 , \Inst_Mem/n1054 ,
         \Inst_Mem/n1053 , \Inst_Mem/n1052 , \Inst_Mem/n1051 ,
         \Inst_Mem/n1050 , \Inst_Mem/n1049 , \Inst_Mem/n1048 ,
         \Inst_Mem/n1047 , \Inst_Mem/n1046 , \Inst_Mem/n1045 ,
         \Inst_Mem/n1044 , \Inst_Mem/n1043 , \Inst_Mem/n1042 ,
         \Inst_Mem/n1041 , \Inst_Mem/n1040 , \Inst_Mem/n1039 ,
         \Inst_Mem/n1038 , \Inst_Mem/n1037 , \Inst_Mem/n1036 ,
         \Inst_Mem/n1035 , \Inst_Mem/n1034 , \Inst_Mem/n1033 ,
         \Inst_Mem/n1032 , \Inst_Mem/n1031 , \Inst_Mem/n1030 ,
         \Inst_Mem/n1029 , \Inst_Mem/n1028 , \Inst_Mem/n1027 ,
         \Inst_Mem/n1026 , \Inst_Mem/n1025 , \Inst_Mem/n1024 ,
         \Inst_Mem/n1023 , \Inst_Mem/n1022 , \Inst_Mem/n1021 ,
         \Inst_Mem/n1020 , \Inst_Mem/n1019 , \Inst_Mem/n1018 ,
         \Inst_Mem/n1017 , \Inst_Mem/n1016 , \Inst_Mem/n1015 ,
         \Inst_Mem/n1014 , \Inst_Mem/n1013 , \Inst_Mem/n1012 ,
         \Inst_Mem/n1011 , \Inst_Mem/n1010 , \Inst_Mem/n1009 ,
         \Inst_Mem/n1008 , \Inst_Mem/n1007 , \Inst_Mem/n1006 ,
         \Inst_Mem/n1005 , \Inst_Mem/n1004 , \Inst_Mem/n1003 ,
         \Inst_Mem/n1002 , \Inst_Mem/n1001 , \Inst_Mem/n1000 , \Inst_Mem/n999 ,
         \Inst_Mem/n998 , \Inst_Mem/n997 , \Inst_Mem/n996 , \Inst_Mem/n995 ,
         \Inst_Mem/n994 , \Inst_Mem/n993 , \Inst_Mem/n992 , \Inst_Mem/n991 ,
         \Inst_Mem/n990 , \Inst_Mem/n989 , \Inst_Mem/n988 , \Inst_Mem/n987 ,
         \Inst_Mem/n986 , \Inst_Mem/n985 , \Inst_Mem/n984 , \Inst_Mem/n983 ,
         \Inst_Mem/n982 , \Inst_Mem/n981 , \Inst_Mem/n980 , \Inst_Mem/n979 ,
         \Inst_Mem/n978 , \Inst_Mem/n977 , \Inst_Mem/n976 , \Inst_Mem/n975 ,
         \Inst_Mem/n974 , \Inst_Mem/n973 , \Inst_Mem/n972 , \Inst_Mem/n971 ,
         \Inst_Mem/n970 , \Inst_Mem/n969 , \Inst_Mem/n968 , \Inst_Mem/n967 ,
         \Inst_Mem/n966 , \Inst_Mem/n965 , \Inst_Mem/n964 , \Inst_Mem/n963 ,
         \Inst_Mem/n962 , \Inst_Mem/n961 , \Inst_Mem/n960 , \Inst_Mem/n959 ,
         \Inst_Mem/n958 , \Inst_Mem/n957 , \Inst_Mem/n956 , \Inst_Mem/n955 ,
         \Inst_Mem/n954 , \Inst_Mem/n953 , \Inst_Mem/n952 , \Inst_Mem/n951 ,
         \Inst_Mem/n950 , \Inst_Mem/n949 , \Inst_Mem/n948 , \Inst_Mem/n947 ,
         \Inst_Mem/n946 , \Inst_Mem/n945 , \Inst_Mem/n944 , \Inst_Mem/n943 ,
         \Inst_Mem/n942 , \Inst_Mem/n941 , \Inst_Mem/n940 , \Inst_Mem/n939 ,
         \Inst_Mem/n938 , \Inst_Mem/n937 , \Inst_Mem/n936 , \Inst_Mem/n935 ,
         \Inst_Mem/n934 , \Inst_Mem/n933 , \Inst_Mem/n932 , \Inst_Mem/n931 ,
         \Inst_Mem/n930 , \Inst_Mem/n929 , \Inst_Mem/n928 , \Inst_Mem/n927 ,
         \Inst_Mem/n926 , \Inst_Mem/n925 , \Inst_Mem/n924 , \Inst_Mem/n923 ,
         \Inst_Mem/n922 , \Inst_Mem/n921 , \Inst_Mem/n920 , \Inst_Mem/n919 ,
         \Inst_Mem/n918 , \Inst_Mem/n917 , \Inst_Mem/n916 , \Inst_Mem/n915 ,
         \Inst_Mem/n914 , \Inst_Mem/n913 , \Inst_Mem/n912 , \Inst_Mem/n911 ,
         \Inst_Mem/n910 , \Inst_Mem/n909 , \Inst_Mem/n908 , \Inst_Mem/n907 ,
         \Inst_Mem/n906 , \Inst_Mem/n905 , \Inst_Mem/n904 , \Inst_Mem/n903 ,
         \Inst_Mem/n902 , \Inst_Mem/n901 , \Inst_Mem/n900 , \Inst_Mem/n899 ,
         \Inst_Mem/n898 , \Inst_Mem/n897 , \Inst_Mem/n896 , \Inst_Mem/n895 ,
         \Inst_Mem/n894 , \Inst_Mem/n893 , \Inst_Mem/n892 , \Inst_Mem/n891 ,
         \Inst_Mem/n890 , \Inst_Mem/n889 , \Inst_Mem/n888 , \Inst_Mem/n887 ,
         \Inst_Mem/n886 , \Inst_Mem/n885 , \Inst_Mem/n884 , \Inst_Mem/n883 ,
         \Inst_Mem/n882 , \Inst_Mem/n881 , \Inst_Mem/n880 , \Inst_Mem/n879 ,
         \Inst_Mem/n878 , \Inst_Mem/n877 , \Inst_Mem/n876 , \Inst_Mem/n875 ,
         \Inst_Mem/n874 , \Inst_Mem/n873 , \Inst_Mem/n872 , \Inst_Mem/n871 ,
         \Inst_Mem/n870 , \Inst_Mem/n869 , \Inst_Mem/n868 , \Inst_Mem/n867 ,
         \Inst_Mem/n866 , \Inst_Mem/n865 , \Inst_Mem/n864 , \Inst_Mem/n863 ,
         \Inst_Mem/n862 , \Inst_Mem/n861 , \Inst_Mem/n860 , \Inst_Mem/n859 ,
         \Inst_Mem/n858 , \Inst_Mem/n857 , \Inst_Mem/n856 , \Inst_Mem/n855 ,
         \Inst_Mem/n854 , \Inst_Mem/n853 , \Inst_Mem/n852 , \Inst_Mem/n851 ,
         \Inst_Mem/n850 , \Inst_Mem/n849 , \Inst_Mem/n848 , \Inst_Mem/n847 ,
         \Inst_Mem/n846 , \Inst_Mem/n845 , \Inst_Mem/n844 , \Inst_Mem/n843 ,
         \Inst_Mem/n842 , \Inst_Mem/n841 , \Inst_Mem/n840 , \Inst_Mem/n839 ,
         \Inst_Mem/n838 , \Inst_Mem/n837 , \Inst_Mem/n836 , \Inst_Mem/n835 ,
         \Inst_Mem/n834 , \Inst_Mem/n833 , \Inst_Mem/n832 , \Inst_Mem/n831 ,
         \Inst_Mem/n830 , \Inst_Mem/n829 , \Inst_Mem/n828 , \Inst_Mem/n827 ,
         \Inst_Mem/n826 , \Inst_Mem/n825 , \Inst_Mem/n824 , \Inst_Mem/n823 ,
         \Inst_Mem/n822 , \Inst_Mem/n821 , \Inst_Mem/n820 , \Inst_Mem/n819 ,
         \Inst_Mem/n818 , \Inst_Mem/n817 , \Inst_Mem/n816 , \Inst_Mem/n815 ,
         \Inst_Mem/n814 , \Inst_Mem/n813 , \Inst_Mem/n812 , \Inst_Mem/n811 ,
         \Inst_Mem/n810 , \Inst_Mem/n809 , \Inst_Mem/n808 , \Inst_Mem/n807 ,
         \Inst_Mem/n806 , \Inst_Mem/n805 , \Inst_Mem/n804 , \Inst_Mem/n803 ,
         \Inst_Mem/n802 , \Inst_Mem/n801 , \Inst_Mem/n800 , \Inst_Mem/n799 ,
         \Inst_Mem/n798 , \Inst_Mem/n797 , \Inst_Mem/n796 , \Inst_Mem/n795 ,
         \Inst_Mem/n794 , \Inst_Mem/n793 , \Inst_Mem/n792 , \Inst_Mem/n791 ,
         \Inst_Mem/n790 , \Inst_Mem/n789 , \Inst_Mem/n788 , \Inst_Mem/n787 ,
         \Inst_Mem/n786 , \Inst_Mem/n785 , \Inst_Mem/n784 , \Inst_Mem/n783 ,
         \Inst_Mem/n782 , \Inst_Mem/n781 , \Inst_Mem/n780 , \Inst_Mem/n779 ,
         \Inst_Mem/n778 , \Inst_Mem/n777 , \Inst_Mem/n776 , \Inst_Mem/n775 ,
         \Inst_Mem/n774 , \Inst_Mem/n773 , \Inst_Mem/n772 , \Inst_Mem/n771 ,
         \Inst_Mem/n770 , \Inst_Mem/n769 , \Inst_Mem/n768 , \Inst_Mem/n767 ,
         \Inst_Mem/n766 , \Inst_Mem/n765 , \Inst_Mem/n764 , \Inst_Mem/n763 ,
         \Inst_Mem/n762 , \Inst_Mem/n761 , \Inst_Mem/n760 , \Inst_Mem/n759 ,
         \Inst_Mem/n758 , \Inst_Mem/n757 , \Inst_Mem/n756 , \Inst_Mem/n755 ,
         \Inst_Mem/n754 , \Inst_Mem/n753 , \Inst_Mem/n752 , \Inst_Mem/n751 ,
         \Inst_Mem/n750 , \Inst_Mem/n749 , \Inst_Mem/n748 , \Inst_Mem/n747 ,
         \Inst_Mem/n746 , \Inst_Mem/n745 , \Inst_Mem/n744 , \Inst_Mem/n743 ,
         \Inst_Mem/n742 , \Inst_Mem/n741 , \Inst_Mem/n740 , \Inst_Mem/n739 ,
         \Inst_Mem/n738 , \Inst_Mem/n737 , \Inst_Mem/n736 , \Inst_Mem/n735 ,
         \Inst_Mem/n734 , \Inst_Mem/n733 , \Inst_Mem/n732 , \Inst_Mem/n731 ,
         \Inst_Mem/n730 , \Inst_Mem/n729 , \Inst_Mem/n728 , \Inst_Mem/n727 ,
         \Inst_Mem/n726 , \Inst_Mem/n725 , \Inst_Mem/n724 , \Inst_Mem/n723 ,
         \Inst_Mem/n722 , \Inst_Mem/n721 , \Inst_Mem/n720 , \Inst_Mem/n719 ,
         \Inst_Mem/n718 , \Inst_Mem/n717 , \Inst_Mem/n716 , \Inst_Mem/n715 ,
         \Inst_Mem/n714 , \Inst_Mem/n713 , \Inst_Mem/n712 , \Inst_Mem/n711 ,
         \Inst_Mem/n710 , \Inst_Mem/n709 , \Inst_Mem/n708 , \Inst_Mem/n707 ,
         \Inst_Mem/n706 , \Inst_Mem/n705 , \Inst_Mem/n704 , \Inst_Mem/n703 ,
         \Inst_Mem/n702 , \Inst_Mem/n701 , \Inst_Mem/n700 , \Inst_Mem/n699 ,
         \Inst_Mem/n698 , \Inst_Mem/n697 , \Inst_Mem/n696 , \Inst_Mem/n695 ,
         \Inst_Mem/n694 , \Inst_Mem/n693 , \Inst_Mem/n692 , \Inst_Mem/n691 ,
         \Inst_Mem/n690 , \Inst_Mem/n689 , \Inst_Mem/n688 , \Inst_Mem/n687 ,
         \Inst_Mem/n686 , \Inst_Mem/n685 , \Inst_Mem/n684 , \Inst_Mem/n683 ,
         \Inst_Mem/n682 , \Inst_Mem/n681 , \Inst_Mem/n680 , \Inst_Mem/n679 ,
         \Inst_Mem/n678 , \Inst_Mem/n677 , \Inst_Mem/n676 , \Inst_Mem/n675 ,
         \Inst_Mem/n674 , \Inst_Mem/n673 , \Inst_Mem/n672 , \Inst_Mem/n671 ,
         \Inst_Mem/n670 , \Inst_Mem/n669 , \Inst_Mem/n668 , \Inst_Mem/n667 ,
         \Inst_Mem/n666 , \Inst_Mem/n665 , \Inst_Mem/n664 , \Inst_Mem/n663 ,
         \Inst_Mem/n662 , \Inst_Mem/n661 , \Inst_Mem/n660 , \Inst_Mem/n659 ,
         \Inst_Mem/n658 , \Inst_Mem/n657 , \Inst_Mem/n656 , \Inst_Mem/n655 ,
         \Inst_Mem/n654 , \Inst_Mem/n653 , \Inst_Mem/n652 , \Inst_Mem/n651 ,
         \Inst_Mem/n650 , \Inst_Mem/n649 , \Inst_Mem/n648 , \Inst_Mem/n647 ,
         \Inst_Mem/n646 , \Inst_Mem/n645 , \Inst_Mem/n644 , \Inst_Mem/n643 ,
         \Inst_Mem/n642 , \Inst_Mem/n641 , \Inst_Mem/n640 , \Inst_Mem/n639 ,
         \Inst_Mem/n638 , \Inst_Mem/n637 , \Inst_Mem/n636 , \Inst_Mem/n635 ,
         \Inst_Mem/n634 , \Inst_Mem/n633 , \Inst_Mem/n632 , \Inst_Mem/n631 ,
         \Inst_Mem/n630 , \Inst_Mem/n629 , \Inst_Mem/n628 , \Inst_Mem/n627 ,
         \Inst_Mem/n626 , \Inst_Mem/n625 , \Inst_Mem/n624 , \Inst_Mem/n623 ,
         \Inst_Mem/n622 , \Inst_Mem/n621 , \Inst_Mem/n620 , \Inst_Mem/n619 ,
         \Inst_Mem/n618 , \Inst_Mem/n617 , \Inst_Mem/n616 , \Inst_Mem/n615 ,
         \Inst_Mem/n614 , \Inst_Mem/n613 , \Inst_Mem/n612 , \Inst_Mem/n611 ,
         \Inst_Mem/n610 , \Inst_Mem/n609 , \Inst_Mem/n608 , \Inst_Mem/n607 ,
         \Inst_Mem/n606 , \Inst_Mem/n605 , \Inst_Mem/n604 , \Inst_Mem/n603 ,
         \Inst_Mem/n602 , \Inst_Mem/n601 , \Inst_Mem/n600 , \Inst_Mem/n599 ,
         \Inst_Mem/n598 , \Inst_Mem/n597 , \Inst_Mem/n596 , \Inst_Mem/n595 ,
         \Inst_Mem/n594 , \Inst_Mem/n593 , \Inst_Mem/n592 , \Inst_Mem/n591 ,
         \Inst_Mem/n590 , \Inst_Mem/n589 , \Inst_Mem/n588 , \Inst_Mem/n587 ,
         \Inst_Mem/n586 , \Inst_Mem/n585 , \Inst_Mem/n584 , \Inst_Mem/n583 ,
         \Inst_Mem/n582 , \Inst_Mem/n581 , \Inst_Mem/n580 , \Inst_Mem/n579 ,
         \Inst_Mem/n578 , \Inst_Mem/n577 , \Inst_Mem/n576 , \Inst_Mem/n575 ,
         \Inst_Mem/n574 , \Inst_Mem/n573 , \Inst_Mem/n572 , \Inst_Mem/n571 ,
         \Inst_Mem/n570 , \Inst_Mem/n569 , \Inst_Mem/n568 , \Inst_Mem/n567 ,
         \Inst_Mem/n566 , \Inst_Mem/n565 , \Inst_Mem/n564 , \Inst_Mem/n563 ,
         \Inst_Mem/n562 , \Inst_Mem/n561 , \Inst_Mem/n560 , \Inst_Mem/n559 ,
         \Inst_Mem/n558 , \Inst_Mem/n557 , \Inst_Mem/n556 , \Inst_Mem/n555 ,
         \Inst_Mem/n554 , \Inst_Mem/n553 , \Inst_Mem/n552 , \Inst_Mem/n551 ,
         \Inst_Mem/n550 , \Inst_Mem/n549 , \Inst_Mem/n548 , \Inst_Mem/n547 ,
         \Inst_Mem/n546 , \Inst_Mem/n545 , \Inst_Mem/n544 , \Inst_Mem/n543 ,
         \Inst_Mem/n542 , \Inst_Mem/n541 , \Inst_Mem/n540 , \Inst_Mem/n539 ,
         \Inst_Mem/n538 , \Inst_Mem/n537 , \Inst_Mem/n536 , \Inst_Mem/n535 ,
         \Inst_Mem/n534 , \Inst_Mem/n533 , \Inst_Mem/n532 , \Inst_Mem/n531 ,
         \Inst_Mem/n530 , \Inst_Mem/n529 , \Inst_Mem/n528 , \Inst_Mem/n527 ,
         \Inst_Mem/n526 , \Inst_Mem/n525 , \Inst_Mem/n524 , \Inst_Mem/n523 ,
         \Inst_Mem/n522 , \Inst_Mem/n521 , \Inst_Mem/n520 , \Inst_Mem/n519 ,
         \Inst_Mem/n518 , \Inst_Mem/n517 , \Inst_Mem/n516 , \Inst_Mem/n515 ,
         \Inst_Mem/n514 , \Inst_Mem/n513 , \Inst_Mem/n512 , \Inst_Mem/n511 ,
         \Inst_Mem/n510 , \Inst_Mem/n509 , \Inst_Mem/n508 , \Inst_Mem/n507 ,
         \Inst_Mem/n506 , \Inst_Mem/n505 , \Inst_Mem/n504 , \Inst_Mem/n503 ,
         \Inst_Mem/n502 , \Inst_Mem/n501 , \Inst_Mem/n500 , \Inst_Mem/n499 ,
         \Inst_Mem/n498 , \Inst_Mem/n497 , \Inst_Mem/n496 , \Inst_Mem/n495 ,
         \Inst_Mem/n494 , \Inst_Mem/n493 , \Inst_Mem/n492 , \Inst_Mem/n491 ,
         \Inst_Mem/n490 , \Inst_Mem/n489 , \Inst_Mem/n488 , \Inst_Mem/n487 ,
         \Inst_Mem/n486 , \Inst_Mem/n485 , \Inst_Mem/n484 , \Inst_Mem/n483 ,
         \Inst_Mem/n482 , \Inst_Mem/n481 , \Inst_Mem/n480 , \Inst_Mem/n479 ,
         \Inst_Mem/n478 , \Inst_Mem/n477 , \Inst_Mem/n476 , \Inst_Mem/n475 ,
         \Inst_Mem/n474 , \Inst_Mem/n473 , \Inst_Mem/n472 , \Inst_Mem/n471 ,
         \Inst_Mem/n470 , \Inst_Mem/n469 , \Inst_Mem/n468 , \Inst_Mem/n467 ,
         \Inst_Mem/n466 , \Inst_Mem/n465 , \Inst_Mem/n464 , \Inst_Mem/n463 ,
         \Inst_Mem/n462 , \Inst_Mem/n461 , \Inst_Mem/n460 , \Inst_Mem/n459 ,
         \Inst_Mem/n458 , \Inst_Mem/n457 , \Inst_Mem/n456 , \Inst_Mem/n455 ,
         \Inst_Mem/n454 , \Inst_Mem/n453 , \Inst_Mem/n452 , \Inst_Mem/n451 ,
         \Inst_Mem/n450 , \Inst_Mem/n449 , \Inst_Mem/n448 , \Inst_Mem/n447 ,
         \Inst_Mem/n446 , \Inst_Mem/n445 , \Inst_Mem/n444 , \Inst_Mem/n443 ,
         \Inst_Mem/n442 , \Inst_Mem/n441 , \Inst_Mem/n440 , \Inst_Mem/n439 ,
         \Inst_Mem/n438 , \Inst_Mem/n437 , \Inst_Mem/n436 , \Inst_Mem/n435 ,
         \Inst_Mem/n434 , \Inst_Mem/n433 , \Inst_Mem/n432 , \Inst_Mem/n431 ,
         \Inst_Mem/n430 , \Inst_Mem/n429 , \Inst_Mem/n428 , \Inst_Mem/n427 ,
         \Inst_Mem/n426 , \Inst_Mem/n425 , \Inst_Mem/n424 , \Inst_Mem/n423 ,
         \Inst_Mem/n422 , \Inst_Mem/n421 , \Inst_Mem/n420 , \Inst_Mem/n419 ,
         \Inst_Mem/n418 , \Inst_Mem/n417 , \Inst_Mem/n416 , \Inst_Mem/n415 ,
         \Inst_Mem/n414 , \Inst_Mem/n413 , \Inst_Mem/n412 , \Inst_Mem/n411 ,
         \Inst_Mem/n410 , \Inst_Mem/n409 , \Inst_Mem/n408 , \Inst_Mem/n407 ,
         \Inst_Mem/n406 , \Inst_Mem/n405 , \Inst_Mem/n404 , \Inst_Mem/n403 ,
         \Inst_Mem/n402 , \Inst_Mem/n401 , \Inst_Mem/n400 , \Inst_Mem/n399 ,
         \Inst_Mem/n398 , \Inst_Mem/n397 , \Inst_Mem/n396 , \Inst_Mem/n395 ,
         \Inst_Mem/n394 , \Inst_Mem/n393 , \Inst_Mem/n392 , \Inst_Mem/n391 ,
         \Inst_Mem/n390 , \Inst_Mem/n389 , \Inst_Mem/n388 , \Inst_Mem/n387 ,
         \Inst_Mem/n386 , \Inst_Mem/n385 , \Inst_Mem/n384 , \Inst_Mem/n383 ,
         \Inst_Mem/n382 , \Inst_Mem/n381 , \Inst_Mem/n380 , \Inst_Mem/n379 ,
         \Inst_Mem/n378 , \Inst_Mem/n377 , \Inst_Mem/n376 , \Inst_Mem/n375 ,
         \Inst_Mem/n374 , \Inst_Mem/n373 , \Inst_Mem/n372 , \Inst_Mem/n371 ,
         \Inst_Mem/n370 , \Inst_Mem/n369 , \Inst_Mem/n368 , \Inst_Mem/n367 ,
         \Inst_Mem/n366 , \Inst_Mem/n365 , \Inst_Mem/n364 , \Inst_Mem/n363 ,
         \Inst_Mem/n362 , \Inst_Mem/n361 , \Inst_Mem/n360 , \Inst_Mem/n359 ,
         \Inst_Mem/n358 , \Inst_Mem/n357 , \Inst_Mem/n356 , \Inst_Mem/n355 ,
         \Inst_Mem/n354 , \Inst_Mem/n353 , \Inst_Mem/n352 , \Inst_Mem/n351 ,
         \Inst_Mem/n350 , \Inst_Mem/n349 , \Inst_Mem/n348 , \Inst_Mem/n347 ,
         \Inst_Mem/n346 , \Inst_Mem/n345 , \Inst_Mem/n344 , \Inst_Mem/n343 ,
         \Inst_Mem/n342 , \Inst_Mem/n341 , \Inst_Mem/n340 , \Inst_Mem/n339 ,
         \Inst_Mem/n338 , \Inst_Mem/n337 , \Inst_Mem/n336 , \Inst_Mem/n335 ,
         \Inst_Mem/n334 , \Inst_Mem/n333 , \Inst_Mem/n332 , \Inst_Mem/n331 ,
         \Inst_Mem/n330 , \Inst_Mem/n329 , \Inst_Mem/n328 , \Inst_Mem/n327 ,
         \Inst_Mem/n326 , \Inst_Mem/n325 , \Inst_Mem/n324 , \Inst_Mem/n323 ,
         \Inst_Mem/n322 , \Inst_Mem/n321 , \Inst_Mem/n320 , \Inst_Mem/n319 ,
         \Inst_Mem/n318 , \Inst_Mem/n317 , \Inst_Mem/n316 , \Inst_Mem/n315 ,
         \Inst_Mem/n314 , \Inst_Mem/n313 , \Inst_Mem/n312 , \Inst_Mem/n311 ,
         \Inst_Mem/n310 , \Inst_Mem/n309 , \Inst_Mem/n308 , \Inst_Mem/n307 ,
         \Inst_Mem/n306 , \Inst_Mem/n305 , \Inst_Mem/n304 , \Inst_Mem/n303 ,
         \Inst_Mem/n302 , \Inst_Mem/n301 , \Inst_Mem/n300 , \Inst_Mem/n299 ,
         \Inst_Mem/n298 , \Inst_Mem/n297 , \Inst_Mem/n296 , \Inst_Mem/n295 ,
         \Inst_Mem/n294 , \Inst_Mem/n293 , \Inst_Mem/n292 , \Inst_Mem/n291 ,
         \Inst_Mem/n290 , \Inst_Mem/n289 , \Inst_Mem/n288 , \Inst_Mem/n287 ,
         \Inst_Mem/n286 , \Inst_Mem/n285 , \Inst_Mem/n284 , \Inst_Mem/n283 ,
         \Inst_Mem/n282 , \Inst_Mem/n281 , \Inst_Mem/n280 , \Inst_Mem/n279 ,
         \Inst_Mem/n278 , \Inst_Mem/n277 , \Inst_Mem/n276 , \Inst_Mem/n275 ,
         \Inst_Mem/n274 , \Inst_Mem/n273 , \Inst_Mem/n272 , \Inst_Mem/n271 ,
         \Inst_Mem/n270 , \Inst_Mem/n269 , \Inst_Mem/n268 , \Inst_Mem/n267 ,
         \Inst_Mem/n266 , \Inst_Mem/n265 , \Inst_Mem/n264 , \Inst_Mem/n263 ,
         \Inst_Mem/n262 , \Inst_Mem/n261 , \Inst_Mem/n260 , \Inst_Mem/n259 ,
         \Inst_Mem/n258 , \Inst_Mem/n257 , \Inst_Mem/n256 , \Inst_Mem/n255 ,
         \Inst_Mem/n254 , \Inst_Mem/n253 , \Inst_Mem/n252 , \Inst_Mem/n251 ,
         \Inst_Mem/n250 , \Inst_Mem/n249 , \Inst_Mem/n248 , \Inst_Mem/n247 ,
         \Inst_Mem/n246 , \Inst_Mem/n245 , \Inst_Mem/n244 , \Inst_Mem/n243 ,
         \Inst_Mem/n242 , \Inst_Mem/n241 , \Inst_Mem/n240 , \Inst_Mem/n239 ,
         \Inst_Mem/n238 , \Inst_Mem/n237 , \Inst_Mem/n236 , \Inst_Mem/n235 ,
         \Inst_Mem/n234 , \Inst_Mem/n233 , \Inst_Mem/n232 , \Inst_Mem/n231 ,
         \Inst_Mem/n230 , \Inst_Mem/n229 , \Inst_Mem/n228 , \Inst_Mem/n227 ,
         \Inst_Mem/n226 , \Inst_Mem/n225 , \Inst_Mem/n224 , \Inst_Mem/n223 ,
         \Inst_Mem/n222 , \Inst_Mem/n221 , \Inst_Mem/n220 , \Inst_Mem/n219 ,
         \Inst_Mem/n218 , \Inst_Mem/n217 , \Inst_Mem/n216 , \Inst_Mem/n215 ,
         \Inst_Mem/n214 , \Inst_Mem/n213 , \Inst_Mem/n212 , \Inst_Mem/n211 ,
         \Inst_Mem/n210 , \Inst_Mem/n209 , \Inst_Mem/n208 , \Inst_Mem/n207 ,
         \Inst_Mem/n206 , \Inst_Mem/n205 , \Inst_Mem/n204 , \Inst_Mem/n203 ,
         \Inst_Mem/n202 , \Inst_Mem/n201 , \Inst_Mem/n200 , \Inst_Mem/n199 ,
         \Inst_Mem/n198 , \Inst_Mem/n197 , \Inst_Mem/n196 , \Inst_Mem/n195 ,
         \Inst_Mem/n194 , \Inst_Mem/n193 , \Inst_Mem/n192 , \Inst_Mem/n191 ,
         \Inst_Mem/n190 , \Inst_Mem/n189 , \Inst_Mem/n188 , \Inst_Mem/n187 ,
         \Inst_Mem/n186 , \Inst_Mem/n185 , \Inst_Mem/n184 , \Inst_Mem/n183 ,
         \Inst_Mem/n182 , \Inst_Mem/n181 , \Inst_Mem/n180 , \Inst_Mem/n179 ,
         \Inst_Mem/n178 , \Inst_Mem/n177 , \Inst_Mem/n176 , \Inst_Mem/n175 ,
         \Inst_Mem/n174 , \Inst_Mem/n173 , \Inst_Mem/n172 , \Inst_Mem/n171 ,
         \Inst_Mem/n170 , \Inst_Mem/n169 , \Inst_Mem/n168 , \Inst_Mem/n167 ,
         \Inst_Mem/n166 , \Inst_Mem/n165 , \Inst_Mem/n164 , \Inst_Mem/n163 ,
         \Inst_Mem/n162 , \Inst_Mem/n161 , \Inst_Mem/n160 , \Inst_Mem/n159 ,
         \Inst_Mem/n158 , \Inst_Mem/n157 , \Inst_Mem/n156 , \Inst_Mem/n155 ,
         \Inst_Mem/n154 , \Inst_Mem/n153 , \Inst_Mem/n152 , \Inst_Mem/n151 ,
         \Inst_Mem/n150 , \Inst_Mem/n149 , \Inst_Mem/n148 , \Inst_Mem/n147 ,
         \Inst_Mem/n146 , \Inst_Mem/n145 , \Inst_Mem/n144 , \Inst_Mem/n143 ,
         \Inst_Mem/n142 , \Inst_Mem/n141 , \Inst_Mem/n140 , \Inst_Mem/n139 ,
         \Inst_Mem/n138 , \Inst_Mem/n137 , \Inst_Mem/n136 , \Inst_Mem/n135 ,
         \Inst_Mem/n134 , \Inst_Mem/n133 , \Inst_Mem/n132 , \Inst_Mem/n131 ,
         \Inst_Mem/n130 , \Inst_Mem/n129 , \Inst_Mem/n128 , \Inst_Mem/n127 ,
         \Inst_Mem/n126 , \Inst_Mem/n125 , \Inst_Mem/n124 , \Inst_Mem/n123 ,
         \Inst_Mem/n122 , \Inst_Mem/n121 , \Inst_Mem/n120 , \Inst_Mem/n119 ,
         \Inst_Mem/n118 , \Inst_Mem/n117 , \Inst_Mem/n116 , \Inst_Mem/n115 ,
         \Inst_Mem/n114 , \Inst_Mem/n113 , \Inst_Mem/n112 , \Inst_Mem/n111 ,
         \Inst_Mem/n110 , \Inst_Mem/n109 , \Inst_Mem/n108 , \Inst_Mem/n107 ,
         \Inst_Mem/n106 , \Inst_Mem/n105 , \Inst_Mem/n104 , \Inst_Mem/n103 ,
         \Inst_Mem/n102 , \Inst_Mem/n101 , \Inst_Mem/n100 , \Inst_Mem/n99 ,
         \Inst_Mem/n98 , \Inst_Mem/n97 , \Inst_Mem/n96 , \Inst_Mem/n95 ,
         \Inst_Mem/n94 , \Inst_Mem/n93 , \Inst_Mem/n92 , \Inst_Mem/n91 ,
         \Inst_Mem/n90 , \Inst_Mem/n89 , \Inst_Mem/n88 , \Inst_Mem/n87 ,
         \Inst_Mem/n86 , \Inst_Mem/n85 , \Inst_Mem/n84 , \Inst_Mem/n83 ,
         \Inst_Mem/n82 , \Inst_Mem/n81 , \Inst_Mem/n80 , \Inst_Mem/n79 ,
         \Inst_Mem/n78 , \Inst_Mem/n77 , \Inst_Mem/n76 , \Inst_Mem/n75 ,
         \Inst_Mem/n74 , \Inst_Mem/n73 , \Inst_Mem/n72 , \Inst_Mem/n71 ,
         \Inst_Mem/n70 , \Inst_Mem/n69 , \Inst_Mem/n68 , \Inst_Mem/n67 ,
         \Inst_Mem/n66 , \Inst_Mem/n65 , \Inst_Mem/n64 , \Inst_Mem/n63 ,
         \Inst_Mem/n62 , \Inst_Mem/n61 , \Inst_Mem/n60 , \Inst_Mem/n59 ,
         \Inst_Mem/n58 , \Inst_Mem/n57 , \Inst_Mem/n56 , \Inst_Mem/n55 ,
         \Inst_Mem/n54 , \Inst_Mem/n53 , \Inst_Mem/n52 , \Inst_Mem/n51 ,
         \Inst_Mem/n50 , \Inst_Mem/n49 , \Inst_Mem/n48 , \Inst_Mem/n47 ,
         \Inst_Mem/n46 , \Inst_Mem/n45 , \Inst_Mem/n44 , \Inst_Mem/n43 ,
         \Inst_Mem/n42 , \Inst_Mem/n41 , \Inst_Mem/n40 , \Inst_Mem/n39 ,
         \Inst_Mem/n38 , \Inst_Mem/n37 , \Inst_Mem/n36 , \Inst_Mem/n35 ,
         \Inst_Mem/n34 , \Inst_Mem/n33 , \Inst_Mem/n32 , \Inst_Mem/n31 ,
         \Inst_Mem/n30 , \Inst_Mem/n29 , \Inst_Mem/n28 , \Inst_Mem/n27 ,
         \Inst_Mem/n26 , \Inst_Mem/n25 , \Inst_Mem/n24 , \Inst_Mem/n23 ,
         \Inst_Mem/n22 , \Inst_Mem/n21 , \Inst_Mem/n20 , \Inst_Mem/n19 ,
         \Inst_Mem/n18 , \Inst_Mem/n17 , \Inst_Mem/n16 , \Inst_Mem/n15 ,
         \Inst_Mem/n14 , \Inst_Mem/n13 , \Inst_Mem/n12 , \Inst_Mem/n11 ,
         \Inst_Mem/n10 , \Inst_Mem/n9 , \Inst_Mem/n8 , \Inst_Mem/n7 ,
         \Inst_Mem/n6 , \Inst_Mem/n5 , \Inst_Mem/n4 , \Inst_Mem/n3 ,
         \Inst_Mem/n2 , \Inst_Mem/n1 , \Data_Mem/n8247 , \Data_Mem/n8246 ,
         \Data_Mem/n8245 , \Data_Mem/n8244 , \Data_Mem/n8243 ,
         \Data_Mem/n8242 , \Data_Mem/n8241 , \Data_Mem/n8240 ,
         \Data_Mem/n8239 , \Data_Mem/n8238 , \Data_Mem/n8237 ,
         \Data_Mem/n8236 , \Data_Mem/n8235 , \Data_Mem/n8234 ,
         \Data_Mem/n8233 , \Data_Mem/n8232 , \Data_Mem/n8231 ,
         \Data_Mem/n8230 , \Data_Mem/n8229 , \Data_Mem/n8228 ,
         \Data_Mem/n8227 , \Data_Mem/n8226 , \Data_Mem/n8225 ,
         \Data_Mem/n8224 , \Data_Mem/n8223 , \Data_Mem/n8222 ,
         \Data_Mem/n8221 , \Data_Mem/n8220 , \Data_Mem/n8219 ,
         \Data_Mem/n8218 , \Data_Mem/n8217 , \Data_Mem/n8216 ,
         \Data_Mem/n8215 , \Data_Mem/n8214 , \Data_Mem/n8213 ,
         \Data_Mem/n8212 , \Data_Mem/n8211 , \Data_Mem/n8210 ,
         \Data_Mem/n8209 , \Data_Mem/n8208 , \Data_Mem/n8207 ,
         \Data_Mem/n8206 , \Data_Mem/n8205 , \Data_Mem/n8204 ,
         \Data_Mem/n8203 , \Data_Mem/n8202 , \Data_Mem/n8201 ,
         \Data_Mem/n8200 , \Data_Mem/n8199 , \Data_Mem/n8198 ,
         \Data_Mem/n8197 , \Data_Mem/n8196 , \Data_Mem/n8195 ,
         \Data_Mem/n8194 , \Data_Mem/n8193 , \Data_Mem/n8192 ,
         \Data_Mem/n8191 , \Data_Mem/n8190 , \Data_Mem/n8189 ,
         \Data_Mem/n8188 , \Data_Mem/n8187 , \Data_Mem/n8186 ,
         \Data_Mem/n8185 , \Data_Mem/n8184 , \Data_Mem/n8183 ,
         \Data_Mem/n8182 , \Data_Mem/n8181 , \Data_Mem/n8180 ,
         \Data_Mem/n8179 , \Data_Mem/n8178 , \Data_Mem/n8177 ,
         \Data_Mem/n8176 , \Data_Mem/n8175 , \Data_Mem/n8174 ,
         \Data_Mem/n8173 , \Data_Mem/n8172 , \Data_Mem/n8171 ,
         \Data_Mem/n8170 , \Data_Mem/n8169 , \Data_Mem/n8168 ,
         \Data_Mem/n8167 , \Data_Mem/n8166 , \Data_Mem/n8165 ,
         \Data_Mem/n8164 , \Data_Mem/n8163 , \Data_Mem/n8162 ,
         \Data_Mem/n8161 , \Data_Mem/n8160 , \Data_Mem/n8159 ,
         \Data_Mem/n8158 , \Data_Mem/n8157 , \Data_Mem/n8156 ,
         \Data_Mem/n8155 , \Data_Mem/n8154 , \Data_Mem/n8153 ,
         \Data_Mem/n8152 , \Data_Mem/n8151 , \Data_Mem/n8150 ,
         \Data_Mem/n8149 , \Data_Mem/n8148 , \Data_Mem/n8147 ,
         \Data_Mem/n8146 , \Data_Mem/n8145 , \Data_Mem/n8144 ,
         \Data_Mem/n8143 , \Data_Mem/n8142 , \Data_Mem/n8141 ,
         \Data_Mem/n8140 , \Data_Mem/n8139 , \Data_Mem/n8138 ,
         \Data_Mem/n8137 , \Data_Mem/n8136 , \Data_Mem/n8135 ,
         \Data_Mem/n8134 , \Data_Mem/n8133 , \Data_Mem/n8132 ,
         \Data_Mem/n8131 , \Data_Mem/n8130 , \Data_Mem/n8129 ,
         \Data_Mem/n8128 , \Data_Mem/n8127 , \Data_Mem/n8126 ,
         \Data_Mem/n8125 , \Data_Mem/n8124 , \Data_Mem/n8123 ,
         \Data_Mem/n8122 , \Data_Mem/n8121 , \Data_Mem/n8120 ,
         \Data_Mem/n8119 , \Data_Mem/n8118 , \Data_Mem/n8117 ,
         \Data_Mem/n8116 , \Data_Mem/n8115 , \Data_Mem/n8114 ,
         \Data_Mem/n8113 , \Data_Mem/n8112 , \Data_Mem/n8111 ,
         \Data_Mem/n8110 , \Data_Mem/n8109 , \Data_Mem/n8108 ,
         \Data_Mem/n8107 , \Data_Mem/n8106 , \Data_Mem/n8105 ,
         \Data_Mem/n8104 , \Data_Mem/n8103 , \Data_Mem/n8102 ,
         \Data_Mem/n8101 , \Data_Mem/n8100 , \Data_Mem/n8099 ,
         \Data_Mem/n8098 , \Data_Mem/n8097 , \Data_Mem/n8096 ,
         \Data_Mem/n8095 , \Data_Mem/n8094 , \Data_Mem/n8093 ,
         \Data_Mem/n8092 , \Data_Mem/n8091 , \Data_Mem/n8090 ,
         \Data_Mem/n8089 , \Data_Mem/n8088 , \Data_Mem/n8087 ,
         \Data_Mem/n8086 , \Data_Mem/n8085 , \Data_Mem/n8084 ,
         \Data_Mem/n8083 , \Data_Mem/n8082 , \Data_Mem/n8081 ,
         \Data_Mem/n8080 , \Data_Mem/n8079 , \Data_Mem/n8078 ,
         \Data_Mem/n8077 , \Data_Mem/n8076 , \Data_Mem/n8075 ,
         \Data_Mem/n8074 , \Data_Mem/n8073 , \Data_Mem/n8072 ,
         \Data_Mem/n8071 , \Data_Mem/n8070 , \Data_Mem/n8069 ,
         \Data_Mem/n8068 , \Data_Mem/n8067 , \Data_Mem/n8066 ,
         \Data_Mem/n8065 , \Data_Mem/n8064 , \Data_Mem/n8063 ,
         \Data_Mem/n8062 , \Data_Mem/n8061 , \Data_Mem/n8060 ,
         \Data_Mem/n8059 , \Data_Mem/n8058 , \Data_Mem/n8057 ,
         \Data_Mem/n8056 , \Data_Mem/n8055 , \Data_Mem/n8054 ,
         \Data_Mem/n8053 , \Data_Mem/n8052 , \Data_Mem/n8051 ,
         \Data_Mem/n8050 , \Data_Mem/n8049 , \Data_Mem/n8048 ,
         \Data_Mem/n8047 , \Data_Mem/n8046 , \Data_Mem/n8045 ,
         \Data_Mem/n8044 , \Data_Mem/n8043 , \Data_Mem/n8042 ,
         \Data_Mem/n8041 , \Data_Mem/n8040 , \Data_Mem/n8039 ,
         \Data_Mem/n8038 , \Data_Mem/n8037 , \Data_Mem/n8036 ,
         \Data_Mem/n8035 , \Data_Mem/n8034 , \Data_Mem/n8033 ,
         \Data_Mem/n8032 , \Data_Mem/n8031 , \Data_Mem/n8030 ,
         \Data_Mem/n8029 , \Data_Mem/n8028 , \Data_Mem/n8027 ,
         \Data_Mem/n8026 , \Data_Mem/n8025 , \Data_Mem/n8024 ,
         \Data_Mem/n8023 , \Data_Mem/n8022 , \Data_Mem/n8021 ,
         \Data_Mem/n8020 , \Data_Mem/n8019 , \Data_Mem/n8018 ,
         \Data_Mem/n8017 , \Data_Mem/n8016 , \Data_Mem/n8015 ,
         \Data_Mem/n8014 , \Data_Mem/n8013 , \Data_Mem/n8012 ,
         \Data_Mem/n8011 , \Data_Mem/n8010 , \Data_Mem/n8009 ,
         \Data_Mem/n8008 , \Data_Mem/n8007 , \Data_Mem/n8006 ,
         \Data_Mem/n8005 , \Data_Mem/n8004 , \Data_Mem/n8003 ,
         \Data_Mem/n8002 , \Data_Mem/n8001 , \Data_Mem/n8000 ,
         \Data_Mem/n7999 , \Data_Mem/n7998 , \Data_Mem/n7997 ,
         \Data_Mem/n7996 , \Data_Mem/n7995 , \Data_Mem/n7994 ,
         \Data_Mem/n7993 , \Data_Mem/n7992 , \Data_Mem/n7991 ,
         \Data_Mem/n7990 , \Data_Mem/n7989 , \Data_Mem/n7988 ,
         \Data_Mem/n7987 , \Data_Mem/n7986 , \Data_Mem/n7985 ,
         \Data_Mem/n7984 , \Data_Mem/n7983 , \Data_Mem/n7982 ,
         \Data_Mem/n7981 , \Data_Mem/n7980 , \Data_Mem/n7979 ,
         \Data_Mem/n7978 , \Data_Mem/n7977 , \Data_Mem/n7976 ,
         \Data_Mem/n7975 , \Data_Mem/n7974 , \Data_Mem/n7973 ,
         \Data_Mem/n7972 , \Data_Mem/n7971 , \Data_Mem/n7970 ,
         \Data_Mem/n7969 , \Data_Mem/n7968 , \Data_Mem/n7967 ,
         \Data_Mem/n7966 , \Data_Mem/n7965 , \Data_Mem/n7964 ,
         \Data_Mem/n7963 , \Data_Mem/n7962 , \Data_Mem/n7961 ,
         \Data_Mem/n7960 , \Data_Mem/n7959 , \Data_Mem/n7958 ,
         \Data_Mem/n7957 , \Data_Mem/n7956 , \Data_Mem/n7955 ,
         \Data_Mem/n7954 , \Data_Mem/n7953 , \Data_Mem/n7952 ,
         \Data_Mem/n7951 , \Data_Mem/n7950 , \Data_Mem/n7949 ,
         \Data_Mem/n7948 , \Data_Mem/n7947 , \Data_Mem/n7946 ,
         \Data_Mem/n7945 , \Data_Mem/n7944 , \Data_Mem/n7943 ,
         \Data_Mem/n7942 , \Data_Mem/n7941 , \Data_Mem/n7940 ,
         \Data_Mem/n7939 , \Data_Mem/n7938 , \Data_Mem/n7937 ,
         \Data_Mem/n7936 , \Data_Mem/n7935 , \Data_Mem/n7934 ,
         \Data_Mem/n7933 , \Data_Mem/n7932 , \Data_Mem/n7931 ,
         \Data_Mem/n7930 , \Data_Mem/n7929 , \Data_Mem/n7928 ,
         \Data_Mem/n7927 , \Data_Mem/n7926 , \Data_Mem/n7925 ,
         \Data_Mem/n7924 , \Data_Mem/n7923 , \Data_Mem/n7922 ,
         \Data_Mem/n7921 , \Data_Mem/n7920 , \Data_Mem/n7919 ,
         \Data_Mem/n7918 , \Data_Mem/n7917 , \Data_Mem/n7916 ,
         \Data_Mem/n7915 , \Data_Mem/n7914 , \Data_Mem/n7913 ,
         \Data_Mem/n7912 , \Data_Mem/n7911 , \Data_Mem/n7910 ,
         \Data_Mem/n7909 , \Data_Mem/n7908 , \Data_Mem/n7907 ,
         \Data_Mem/n7906 , \Data_Mem/n7905 , \Data_Mem/n7904 ,
         \Data_Mem/n7903 , \Data_Mem/n7902 , \Data_Mem/n7901 ,
         \Data_Mem/n7900 , \Data_Mem/n7899 , \Data_Mem/n7898 ,
         \Data_Mem/n7897 , \Data_Mem/n7896 , \Data_Mem/n7895 ,
         \Data_Mem/n7894 , \Data_Mem/n7893 , \Data_Mem/n7892 ,
         \Data_Mem/n7891 , \Data_Mem/n7890 , \Data_Mem/n7889 ,
         \Data_Mem/n7888 , \Data_Mem/n7887 , \Data_Mem/n7886 ,
         \Data_Mem/n7885 , \Data_Mem/n7884 , \Data_Mem/n7883 ,
         \Data_Mem/n7882 , \Data_Mem/n7881 , \Data_Mem/n7880 ,
         \Data_Mem/n7879 , \Data_Mem/n7878 , \Data_Mem/n7877 ,
         \Data_Mem/n7876 , \Data_Mem/n7875 , \Data_Mem/n7874 ,
         \Data_Mem/n7873 , \Data_Mem/n7872 , \Data_Mem/n7871 ,
         \Data_Mem/n7870 , \Data_Mem/n7869 , \Data_Mem/n7868 ,
         \Data_Mem/n7867 , \Data_Mem/n7866 , \Data_Mem/n7865 ,
         \Data_Mem/n7864 , \Data_Mem/n7863 , \Data_Mem/n7862 ,
         \Data_Mem/n7861 , \Data_Mem/n7860 , \Data_Mem/n7859 ,
         \Data_Mem/n7858 , \Data_Mem/n7857 , \Data_Mem/n7856 ,
         \Data_Mem/n7855 , \Data_Mem/n7854 , \Data_Mem/n7853 ,
         \Data_Mem/n7852 , \Data_Mem/n7851 , \Data_Mem/n7850 ,
         \Data_Mem/n7849 , \Data_Mem/n7848 , \Data_Mem/n7847 ,
         \Data_Mem/n7846 , \Data_Mem/n7845 , \Data_Mem/n7844 ,
         \Data_Mem/n7843 , \Data_Mem/n7842 , \Data_Mem/n7841 ,
         \Data_Mem/n7840 , \Data_Mem/n7839 , \Data_Mem/n7838 ,
         \Data_Mem/n7837 , \Data_Mem/n7836 , \Data_Mem/n7835 ,
         \Data_Mem/n7834 , \Data_Mem/n7833 , \Data_Mem/n7832 ,
         \Data_Mem/n7831 , \Data_Mem/n7830 , \Data_Mem/n7829 ,
         \Data_Mem/n7828 , \Data_Mem/n7827 , \Data_Mem/n7826 ,
         \Data_Mem/n7825 , \Data_Mem/n7824 , \Data_Mem/n7823 ,
         \Data_Mem/n7822 , \Data_Mem/n7821 , \Data_Mem/n7820 ,
         \Data_Mem/n7819 , \Data_Mem/n7818 , \Data_Mem/n7817 ,
         \Data_Mem/n7816 , \Data_Mem/n7815 , \Data_Mem/n7814 ,
         \Data_Mem/n7813 , \Data_Mem/n7812 , \Data_Mem/n7811 ,
         \Data_Mem/n7810 , \Data_Mem/n7809 , \Data_Mem/n7808 ,
         \Data_Mem/n7807 , \Data_Mem/n7806 , \Data_Mem/n7805 ,
         \Data_Mem/n7804 , \Data_Mem/n7803 , \Data_Mem/n7802 ,
         \Data_Mem/n7801 , \Data_Mem/n7800 , \Data_Mem/n7799 ,
         \Data_Mem/n7798 , \Data_Mem/n7797 , \Data_Mem/n7796 ,
         \Data_Mem/n7795 , \Data_Mem/n7794 , \Data_Mem/n7793 ,
         \Data_Mem/n7792 , \Data_Mem/n7791 , \Data_Mem/n7790 ,
         \Data_Mem/n7789 , \Data_Mem/n7788 , \Data_Mem/n7787 ,
         \Data_Mem/n7786 , \Data_Mem/n7785 , \Data_Mem/n7784 ,
         \Data_Mem/n7783 , \Data_Mem/n7782 , \Data_Mem/n7781 ,
         \Data_Mem/n7780 , \Data_Mem/n7779 , \Data_Mem/n7778 ,
         \Data_Mem/n7777 , \Data_Mem/n7776 , \Data_Mem/n7775 ,
         \Data_Mem/n7774 , \Data_Mem/n7773 , \Data_Mem/n7772 ,
         \Data_Mem/n7771 , \Data_Mem/n7770 , \Data_Mem/n7769 ,
         \Data_Mem/n7768 , \Data_Mem/n7767 , \Data_Mem/n7766 ,
         \Data_Mem/n7765 , \Data_Mem/n7764 , \Data_Mem/n7763 ,
         \Data_Mem/n7762 , \Data_Mem/n7761 , \Data_Mem/n7760 ,
         \Data_Mem/n7759 , \Data_Mem/n7758 , \Data_Mem/n7757 ,
         \Data_Mem/n7756 , \Data_Mem/n7755 , \Data_Mem/n7754 ,
         \Data_Mem/n7753 , \Data_Mem/n7752 , \Data_Mem/n7751 ,
         \Data_Mem/n7750 , \Data_Mem/n7749 , \Data_Mem/n7748 ,
         \Data_Mem/n7747 , \Data_Mem/n7746 , \Data_Mem/n7745 ,
         \Data_Mem/n7744 , \Data_Mem/n7743 , \Data_Mem/n7742 ,
         \Data_Mem/n7741 , \Data_Mem/n7740 , \Data_Mem/n7739 ,
         \Data_Mem/n7738 , \Data_Mem/n7737 , \Data_Mem/n7736 ,
         \Data_Mem/n7735 , \Data_Mem/n7734 , \Data_Mem/n7733 ,
         \Data_Mem/n7732 , \Data_Mem/n7731 , \Data_Mem/n7730 ,
         \Data_Mem/n7729 , \Data_Mem/n7728 , \Data_Mem/n7727 ,
         \Data_Mem/n7726 , \Data_Mem/n7725 , \Data_Mem/n7724 ,
         \Data_Mem/n7723 , \Data_Mem/n7722 , \Data_Mem/n7721 ,
         \Data_Mem/n7720 , \Data_Mem/n7719 , \Data_Mem/n7718 ,
         \Data_Mem/n7717 , \Data_Mem/n7716 , \Data_Mem/n7715 ,
         \Data_Mem/n7714 , \Data_Mem/n7713 , \Data_Mem/n7712 ,
         \Data_Mem/n7711 , \Data_Mem/n7710 , \Data_Mem/n7709 ,
         \Data_Mem/n7708 , \Data_Mem/n7707 , \Data_Mem/n7706 ,
         \Data_Mem/n7705 , \Data_Mem/n7704 , \Data_Mem/n7703 ,
         \Data_Mem/n7702 , \Data_Mem/n7701 , \Data_Mem/n7700 ,
         \Data_Mem/n7699 , \Data_Mem/n7698 , \Data_Mem/n7697 ,
         \Data_Mem/n7696 , \Data_Mem/n7695 , \Data_Mem/n7694 ,
         \Data_Mem/n7693 , \Data_Mem/n7692 , \Data_Mem/n7691 ,
         \Data_Mem/n7690 , \Data_Mem/n7689 , \Data_Mem/n7688 ,
         \Data_Mem/n7687 , \Data_Mem/n7686 , \Data_Mem/n7685 ,
         \Data_Mem/n7684 , \Data_Mem/n7683 , \Data_Mem/n7682 ,
         \Data_Mem/n7681 , \Data_Mem/n7680 , \Data_Mem/n7679 ,
         \Data_Mem/n7678 , \Data_Mem/n7677 , \Data_Mem/n7676 ,
         \Data_Mem/n7675 , \Data_Mem/n7674 , \Data_Mem/n7673 ,
         \Data_Mem/n7672 , \Data_Mem/n7671 , \Data_Mem/n7670 ,
         \Data_Mem/n7669 , \Data_Mem/n7668 , \Data_Mem/n7667 ,
         \Data_Mem/n7666 , \Data_Mem/n7665 , \Data_Mem/n7664 ,
         \Data_Mem/n7663 , \Data_Mem/n7662 , \Data_Mem/n7661 ,
         \Data_Mem/n7660 , \Data_Mem/n7659 , \Data_Mem/n7658 ,
         \Data_Mem/n7657 , \Data_Mem/n7656 , \Data_Mem/n7655 ,
         \Data_Mem/n7654 , \Data_Mem/n7653 , \Data_Mem/n7652 ,
         \Data_Mem/n7651 , \Data_Mem/n7650 , \Data_Mem/n7649 ,
         \Data_Mem/n7648 , \Data_Mem/n7647 , \Data_Mem/n7646 ,
         \Data_Mem/n7645 , \Data_Mem/n7644 , \Data_Mem/n7643 ,
         \Data_Mem/n7642 , \Data_Mem/n7641 , \Data_Mem/n7640 ,
         \Data_Mem/n7639 , \Data_Mem/n7638 , \Data_Mem/n7637 ,
         \Data_Mem/n7636 , \Data_Mem/n7635 , \Data_Mem/n7634 ,
         \Data_Mem/n7633 , \Data_Mem/n7632 , \Data_Mem/n7631 ,
         \Data_Mem/n7630 , \Data_Mem/n7629 , \Data_Mem/n7628 ,
         \Data_Mem/n7627 , \Data_Mem/n7626 , \Data_Mem/n7625 ,
         \Data_Mem/n7624 , \Data_Mem/n7623 , \Data_Mem/n7622 ,
         \Data_Mem/n7621 , \Data_Mem/n7620 , \Data_Mem/n7619 ,
         \Data_Mem/n7618 , \Data_Mem/n7617 , \Data_Mem/n7616 ,
         \Data_Mem/n7615 , \Data_Mem/n7614 , \Data_Mem/n7613 ,
         \Data_Mem/n7612 , \Data_Mem/n7611 , \Data_Mem/n7610 ,
         \Data_Mem/n7609 , \Data_Mem/n7608 , \Data_Mem/n7607 ,
         \Data_Mem/n7606 , \Data_Mem/n7605 , \Data_Mem/n7604 ,
         \Data_Mem/n7603 , \Data_Mem/n7602 , \Data_Mem/n7601 ,
         \Data_Mem/n7600 , \Data_Mem/n7599 , \Data_Mem/n7598 ,
         \Data_Mem/n7597 , \Data_Mem/n7596 , \Data_Mem/n7595 ,
         \Data_Mem/n7594 , \Data_Mem/n7593 , \Data_Mem/n7592 ,
         \Data_Mem/n7591 , \Data_Mem/n7590 , \Data_Mem/n7589 ,
         \Data_Mem/n7588 , \Data_Mem/n7587 , \Data_Mem/n7586 ,
         \Data_Mem/n7585 , \Data_Mem/n7584 , \Data_Mem/n7583 ,
         \Data_Mem/n7582 , \Data_Mem/n7581 , \Data_Mem/n7580 ,
         \Data_Mem/n7579 , \Data_Mem/n7578 , \Data_Mem/n7577 ,
         \Data_Mem/n7576 , \Data_Mem/n7575 , \Data_Mem/n7574 ,
         \Data_Mem/n7573 , \Data_Mem/n7572 , \Data_Mem/n7571 ,
         \Data_Mem/n7570 , \Data_Mem/n7569 , \Data_Mem/n7568 ,
         \Data_Mem/n7567 , \Data_Mem/n7566 , \Data_Mem/n7565 ,
         \Data_Mem/n7564 , \Data_Mem/n7563 , \Data_Mem/n7562 ,
         \Data_Mem/n7561 , \Data_Mem/n7560 , \Data_Mem/n7559 ,
         \Data_Mem/n7558 , \Data_Mem/n7557 , \Data_Mem/n7556 ,
         \Data_Mem/n7555 , \Data_Mem/n7554 , \Data_Mem/n7553 ,
         \Data_Mem/n7552 , \Data_Mem/n7551 , \Data_Mem/n7550 ,
         \Data_Mem/n7549 , \Data_Mem/n7548 , \Data_Mem/n7547 ,
         \Data_Mem/n7546 , \Data_Mem/n7545 , \Data_Mem/n7544 ,
         \Data_Mem/n7543 , \Data_Mem/n7542 , \Data_Mem/n7541 ,
         \Data_Mem/n7540 , \Data_Mem/n7539 , \Data_Mem/n7538 ,
         \Data_Mem/n7537 , \Data_Mem/n7536 , \Data_Mem/n7535 ,
         \Data_Mem/n7534 , \Data_Mem/n7533 , \Data_Mem/n7532 ,
         \Data_Mem/n7531 , \Data_Mem/n7530 , \Data_Mem/n7529 ,
         \Data_Mem/n7528 , \Data_Mem/n7527 , \Data_Mem/n7526 ,
         \Data_Mem/n7525 , \Data_Mem/n7524 , \Data_Mem/n7523 ,
         \Data_Mem/n7522 , \Data_Mem/n7521 , \Data_Mem/n7520 ,
         \Data_Mem/n7519 , \Data_Mem/n7518 , \Data_Mem/n7517 ,
         \Data_Mem/n7516 , \Data_Mem/n7515 , \Data_Mem/n7514 ,
         \Data_Mem/n7513 , \Data_Mem/n7512 , \Data_Mem/n7511 ,
         \Data_Mem/n7510 , \Data_Mem/n7509 , \Data_Mem/n7508 ,
         \Data_Mem/n7507 , \Data_Mem/n7506 , \Data_Mem/n7505 ,
         \Data_Mem/n7504 , \Data_Mem/n7503 , \Data_Mem/n7502 ,
         \Data_Mem/n7501 , \Data_Mem/n7500 , \Data_Mem/n7499 ,
         \Data_Mem/n7498 , \Data_Mem/n7497 , \Data_Mem/n7496 ,
         \Data_Mem/n7495 , \Data_Mem/n7494 , \Data_Mem/n7493 ,
         \Data_Mem/n7492 , \Data_Mem/n7491 , \Data_Mem/n7490 ,
         \Data_Mem/n7489 , \Data_Mem/n7488 , \Data_Mem/n7487 ,
         \Data_Mem/n7486 , \Data_Mem/n7485 , \Data_Mem/n7484 ,
         \Data_Mem/n7483 , \Data_Mem/n7482 , \Data_Mem/n7481 ,
         \Data_Mem/n7480 , \Data_Mem/n7479 , \Data_Mem/n7478 ,
         \Data_Mem/n7477 , \Data_Mem/n7476 , \Data_Mem/n7475 ,
         \Data_Mem/n7474 , \Data_Mem/n7473 , \Data_Mem/n7472 ,
         \Data_Mem/n7471 , \Data_Mem/n7470 , \Data_Mem/n7469 ,
         \Data_Mem/n7468 , \Data_Mem/n7467 , \Data_Mem/n7466 ,
         \Data_Mem/n7465 , \Data_Mem/n7464 , \Data_Mem/n7463 ,
         \Data_Mem/n7462 , \Data_Mem/n7461 , \Data_Mem/n7460 ,
         \Data_Mem/n7459 , \Data_Mem/n7458 , \Data_Mem/n7457 ,
         \Data_Mem/n7456 , \Data_Mem/n7455 , \Data_Mem/n7454 ,
         \Data_Mem/n7453 , \Data_Mem/n7452 , \Data_Mem/n7451 ,
         \Data_Mem/n7450 , \Data_Mem/n7449 , \Data_Mem/n7448 ,
         \Data_Mem/n7447 , \Data_Mem/n7446 , \Data_Mem/n7445 ,
         \Data_Mem/n7444 , \Data_Mem/n7443 , \Data_Mem/n7442 ,
         \Data_Mem/n7441 , \Data_Mem/n7440 , \Data_Mem/n7439 ,
         \Data_Mem/n7438 , \Data_Mem/n7437 , \Data_Mem/n7436 ,
         \Data_Mem/n7435 , \Data_Mem/n7434 , \Data_Mem/n7433 ,
         \Data_Mem/n7432 , \Data_Mem/n7431 , \Data_Mem/n7430 ,
         \Data_Mem/n7429 , \Data_Mem/n7428 , \Data_Mem/n7427 ,
         \Data_Mem/n7426 , \Data_Mem/n7425 , \Data_Mem/n7424 ,
         \Data_Mem/n7423 , \Data_Mem/n7422 , \Data_Mem/n7421 ,
         \Data_Mem/n7420 , \Data_Mem/n7419 , \Data_Mem/n7418 ,
         \Data_Mem/n7417 , \Data_Mem/n7416 , \Data_Mem/n7415 ,
         \Data_Mem/n7414 , \Data_Mem/n7413 , \Data_Mem/n7412 ,
         \Data_Mem/n7411 , \Data_Mem/n7410 , \Data_Mem/n7409 ,
         \Data_Mem/n7408 , \Data_Mem/n7407 , \Data_Mem/n7406 ,
         \Data_Mem/n7405 , \Data_Mem/n7404 , \Data_Mem/n7403 ,
         \Data_Mem/n7402 , \Data_Mem/n7401 , \Data_Mem/n7400 ,
         \Data_Mem/n7399 , \Data_Mem/n7398 , \Data_Mem/n7397 ,
         \Data_Mem/n7396 , \Data_Mem/n7395 , \Data_Mem/n7394 ,
         \Data_Mem/n7393 , \Data_Mem/n7392 , \Data_Mem/n7391 ,
         \Data_Mem/n7390 , \Data_Mem/n7389 , \Data_Mem/n7388 ,
         \Data_Mem/n7387 , \Data_Mem/n7386 , \Data_Mem/n7385 ,
         \Data_Mem/n7384 , \Data_Mem/n7383 , \Data_Mem/n7382 ,
         \Data_Mem/n7381 , \Data_Mem/n7380 , \Data_Mem/n7379 ,
         \Data_Mem/n7378 , \Data_Mem/n7377 , \Data_Mem/n7376 ,
         \Data_Mem/n7375 , \Data_Mem/n7374 , \Data_Mem/n7373 ,
         \Data_Mem/n7372 , \Data_Mem/n7371 , \Data_Mem/n7370 ,
         \Data_Mem/n7369 , \Data_Mem/n7368 , \Data_Mem/n7367 ,
         \Data_Mem/n7366 , \Data_Mem/n7365 , \Data_Mem/n7364 ,
         \Data_Mem/n7363 , \Data_Mem/n7362 , \Data_Mem/n7361 ,
         \Data_Mem/n7360 , \Data_Mem/n7359 , \Data_Mem/n7358 ,
         \Data_Mem/n7357 , \Data_Mem/n7356 , \Data_Mem/n7355 ,
         \Data_Mem/n7354 , \Data_Mem/n7353 , \Data_Mem/n7352 ,
         \Data_Mem/n7351 , \Data_Mem/n7350 , \Data_Mem/n7349 ,
         \Data_Mem/n7348 , \Data_Mem/n7347 , \Data_Mem/n7346 ,
         \Data_Mem/n7345 , \Data_Mem/n7344 , \Data_Mem/n7343 ,
         \Data_Mem/n7342 , \Data_Mem/n7341 , \Data_Mem/n7340 ,
         \Data_Mem/n7339 , \Data_Mem/n7338 , \Data_Mem/n7337 ,
         \Data_Mem/n7336 , \Data_Mem/n7335 , \Data_Mem/n7334 ,
         \Data_Mem/n7333 , \Data_Mem/n7332 , \Data_Mem/n7331 ,
         \Data_Mem/n7330 , \Data_Mem/n7329 , \Data_Mem/n7328 ,
         \Data_Mem/n7327 , \Data_Mem/n7326 , \Data_Mem/n7325 ,
         \Data_Mem/n7324 , \Data_Mem/n7323 , \Data_Mem/n7322 ,
         \Data_Mem/n7321 , \Data_Mem/n7320 , \Data_Mem/n7319 ,
         \Data_Mem/n7318 , \Data_Mem/n7317 , \Data_Mem/n7316 ,
         \Data_Mem/n7315 , \Data_Mem/n7314 , \Data_Mem/n7313 ,
         \Data_Mem/n7312 , \Data_Mem/n7311 , \Data_Mem/n7310 ,
         \Data_Mem/n7309 , \Data_Mem/n7308 , \Data_Mem/n7307 ,
         \Data_Mem/n7306 , \Data_Mem/n7305 , \Data_Mem/n7304 ,
         \Data_Mem/n7303 , \Data_Mem/n7302 , \Data_Mem/n7301 ,
         \Data_Mem/n7300 , \Data_Mem/n7299 , \Data_Mem/n7298 ,
         \Data_Mem/n7297 , \Data_Mem/n7296 , \Data_Mem/n7295 ,
         \Data_Mem/n7294 , \Data_Mem/n7293 , \Data_Mem/n7292 ,
         \Data_Mem/n7291 , \Data_Mem/n7290 , \Data_Mem/n7289 ,
         \Data_Mem/n7288 , \Data_Mem/n7287 , \Data_Mem/n7286 ,
         \Data_Mem/n7285 , \Data_Mem/n7284 , \Data_Mem/n7283 ,
         \Data_Mem/n7282 , \Data_Mem/n7281 , \Data_Mem/n7280 ,
         \Data_Mem/n7279 , \Data_Mem/n7278 , \Data_Mem/n7277 ,
         \Data_Mem/n7276 , \Data_Mem/n7275 , \Data_Mem/n7274 ,
         \Data_Mem/n7273 , \Data_Mem/n7272 , \Data_Mem/n7271 ,
         \Data_Mem/n7270 , \Data_Mem/n7269 , \Data_Mem/n7268 ,
         \Data_Mem/n7267 , \Data_Mem/n7266 , \Data_Mem/n7265 ,
         \Data_Mem/n7264 , \Data_Mem/n7263 , \Data_Mem/n7262 ,
         \Data_Mem/n7261 , \Data_Mem/n7260 , \Data_Mem/n7259 ,
         \Data_Mem/n7258 , \Data_Mem/n7257 , \Data_Mem/n7256 ,
         \Data_Mem/n7255 , \Data_Mem/n7254 , \Data_Mem/n7253 ,
         \Data_Mem/n7252 , \Data_Mem/n7251 , \Data_Mem/n7250 ,
         \Data_Mem/n7249 , \Data_Mem/n7248 , \Data_Mem/n7247 ,
         \Data_Mem/n7246 , \Data_Mem/n7245 , \Data_Mem/n7244 ,
         \Data_Mem/n7243 , \Data_Mem/n7242 , \Data_Mem/n7241 ,
         \Data_Mem/n7240 , \Data_Mem/n7239 , \Data_Mem/n7238 ,
         \Data_Mem/n7237 , \Data_Mem/n7236 , \Data_Mem/n7235 ,
         \Data_Mem/n7234 , \Data_Mem/n7233 , \Data_Mem/n7232 ,
         \Data_Mem/n7231 , \Data_Mem/n7230 , \Data_Mem/n7229 ,
         \Data_Mem/n7228 , \Data_Mem/n7227 , \Data_Mem/n7226 ,
         \Data_Mem/n7225 , \Data_Mem/n7224 , \Data_Mem/n7223 ,
         \Data_Mem/n7222 , \Data_Mem/n7221 , \Data_Mem/n7220 ,
         \Data_Mem/n7219 , \Data_Mem/n7218 , \Data_Mem/n7217 ,
         \Data_Mem/n7216 , \Data_Mem/n7215 , \Data_Mem/n7214 ,
         \Data_Mem/n7213 , \Data_Mem/n7212 , \Data_Mem/n7211 ,
         \Data_Mem/n7210 , \Data_Mem/n7209 , \Data_Mem/n7208 ,
         \Data_Mem/n7207 , \Data_Mem/n7206 , \Data_Mem/n7205 ,
         \Data_Mem/n7204 , \Data_Mem/n7203 , \Data_Mem/n7202 ,
         \Data_Mem/n7201 , \Data_Mem/n7200 , \Data_Mem/n7199 ,
         \Data_Mem/n7198 , \Data_Mem/n7197 , \Data_Mem/n7196 ,
         \Data_Mem/n7195 , \Data_Mem/n7194 , \Data_Mem/n7193 ,
         \Data_Mem/n7192 , \Data_Mem/n7191 , \Data_Mem/n7190 ,
         \Data_Mem/n7189 , \Data_Mem/n7188 , \Data_Mem/n7187 ,
         \Data_Mem/n7186 , \Data_Mem/n7185 , \Data_Mem/n7184 ,
         \Data_Mem/n7183 , \Data_Mem/n7182 , \Data_Mem/n7181 ,
         \Data_Mem/n7180 , \Data_Mem/n7179 , \Data_Mem/n7178 ,
         \Data_Mem/n7177 , \Data_Mem/n7176 , \Data_Mem/n7175 ,
         \Data_Mem/n7174 , \Data_Mem/n7173 , \Data_Mem/n7172 ,
         \Data_Mem/n7171 , \Data_Mem/n7170 , \Data_Mem/n7169 ,
         \Data_Mem/n7168 , \Data_Mem/n7167 , \Data_Mem/n7166 ,
         \Data_Mem/n7165 , \Data_Mem/n7164 , \Data_Mem/n7163 ,
         \Data_Mem/n7162 , \Data_Mem/n7161 , \Data_Mem/n7160 ,
         \Data_Mem/n7159 , \Data_Mem/n7158 , \Data_Mem/n7157 ,
         \Data_Mem/n7156 , \Data_Mem/n7155 , \Data_Mem/n7154 ,
         \Data_Mem/n7153 , \Data_Mem/n7152 , \Data_Mem/n7151 ,
         \Data_Mem/n7150 , \Data_Mem/n7149 , \Data_Mem/n7148 ,
         \Data_Mem/n7147 , \Data_Mem/n7146 , \Data_Mem/n7145 ,
         \Data_Mem/n7144 , \Data_Mem/n7143 , \Data_Mem/n7142 ,
         \Data_Mem/n7141 , \Data_Mem/n7140 , \Data_Mem/n7139 ,
         \Data_Mem/n7138 , \Data_Mem/n7137 , \Data_Mem/n7136 ,
         \Data_Mem/n7135 , \Data_Mem/n7134 , \Data_Mem/n7133 ,
         \Data_Mem/n7132 , \Data_Mem/n7131 , \Data_Mem/n7130 ,
         \Data_Mem/n7129 , \Data_Mem/n7128 , \Data_Mem/n7127 ,
         \Data_Mem/n7126 , \Data_Mem/n7125 , \Data_Mem/n7124 ,
         \Data_Mem/n7123 , \Data_Mem/n7122 , \Data_Mem/n7121 ,
         \Data_Mem/n7120 , \Data_Mem/n7119 , \Data_Mem/n7118 ,
         \Data_Mem/n7117 , \Data_Mem/n7116 , \Data_Mem/n7115 ,
         \Data_Mem/n7114 , \Data_Mem/n7113 , \Data_Mem/n7112 ,
         \Data_Mem/n7111 , \Data_Mem/n7110 , \Data_Mem/n7109 ,
         \Data_Mem/n7108 , \Data_Mem/n7107 , \Data_Mem/n7106 ,
         \Data_Mem/n7105 , \Data_Mem/n7104 , \Data_Mem/n7103 ,
         \Data_Mem/n7102 , \Data_Mem/n7101 , \Data_Mem/n7100 ,
         \Data_Mem/n7099 , \Data_Mem/n7098 , \Data_Mem/n7097 ,
         \Data_Mem/n7096 , \Data_Mem/n7095 , \Data_Mem/n7094 ,
         \Data_Mem/n7093 , \Data_Mem/n7092 , \Data_Mem/n7091 ,
         \Data_Mem/n7090 , \Data_Mem/n7089 , \Data_Mem/n7088 ,
         \Data_Mem/n7087 , \Data_Mem/n7086 , \Data_Mem/n7085 ,
         \Data_Mem/n7084 , \Data_Mem/n7083 , \Data_Mem/n7082 ,
         \Data_Mem/n7081 , \Data_Mem/n7080 , \Data_Mem/n7079 ,
         \Data_Mem/n7078 , \Data_Mem/n7077 , \Data_Mem/n7076 ,
         \Data_Mem/n7075 , \Data_Mem/n7074 , \Data_Mem/n7073 ,
         \Data_Mem/n7072 , \Data_Mem/n7071 , \Data_Mem/n7070 ,
         \Data_Mem/n7069 , \Data_Mem/n7068 , \Data_Mem/n7067 ,
         \Data_Mem/n7066 , \Data_Mem/n7065 , \Data_Mem/n7064 ,
         \Data_Mem/n7063 , \Data_Mem/n7062 , \Data_Mem/n7061 ,
         \Data_Mem/n7060 , \Data_Mem/n7059 , \Data_Mem/n7058 ,
         \Data_Mem/n7057 , \Data_Mem/n7056 , \Data_Mem/n7055 ,
         \Data_Mem/n7054 , \Data_Mem/n7053 , \Data_Mem/n7052 ,
         \Data_Mem/n7051 , \Data_Mem/n7050 , \Data_Mem/n7049 ,
         \Data_Mem/n7048 , \Data_Mem/n7047 , \Data_Mem/n7046 ,
         \Data_Mem/n7045 , \Data_Mem/n7044 , \Data_Mem/n7043 ,
         \Data_Mem/n7042 , \Data_Mem/n7041 , \Data_Mem/n7040 ,
         \Data_Mem/n7039 , \Data_Mem/n7038 , \Data_Mem/n7037 ,
         \Data_Mem/n7036 , \Data_Mem/n7035 , \Data_Mem/n7034 ,
         \Data_Mem/n7033 , \Data_Mem/n7032 , \Data_Mem/n7031 ,
         \Data_Mem/n7030 , \Data_Mem/n7029 , \Data_Mem/n7028 ,
         \Data_Mem/n7027 , \Data_Mem/n7026 , \Data_Mem/n7025 ,
         \Data_Mem/n7024 , \Data_Mem/n7023 , \Data_Mem/n7022 ,
         \Data_Mem/n7021 , \Data_Mem/n7020 , \Data_Mem/n7019 ,
         \Data_Mem/n7018 , \Data_Mem/n7017 , \Data_Mem/n7016 ,
         \Data_Mem/n7015 , \Data_Mem/n7014 , \Data_Mem/n7013 ,
         \Data_Mem/n7012 , \Data_Mem/n7011 , \Data_Mem/n7010 ,
         \Data_Mem/n7009 , \Data_Mem/n7008 , \Data_Mem/n7007 ,
         \Data_Mem/n7006 , \Data_Mem/n7005 , \Data_Mem/n7004 ,
         \Data_Mem/n7003 , \Data_Mem/n7002 , \Data_Mem/n7001 ,
         \Data_Mem/n7000 , \Data_Mem/n6999 , \Data_Mem/n6998 ,
         \Data_Mem/n6997 , \Data_Mem/n6996 , \Data_Mem/n6995 ,
         \Data_Mem/n6994 , \Data_Mem/n6993 , \Data_Mem/n6992 ,
         \Data_Mem/n6991 , \Data_Mem/n6990 , \Data_Mem/n6989 ,
         \Data_Mem/n6988 , \Data_Mem/n6987 , \Data_Mem/n6986 ,
         \Data_Mem/n6985 , \Data_Mem/n6984 , \Data_Mem/n6983 ,
         \Data_Mem/n6982 , \Data_Mem/n6981 , \Data_Mem/n6980 ,
         \Data_Mem/n6979 , \Data_Mem/n6978 , \Data_Mem/n6977 ,
         \Data_Mem/n6976 , \Data_Mem/n6975 , \Data_Mem/n6974 ,
         \Data_Mem/n6973 , \Data_Mem/n6972 , \Data_Mem/n6971 ,
         \Data_Mem/n6970 , \Data_Mem/n6969 , \Data_Mem/n6968 ,
         \Data_Mem/n6967 , \Data_Mem/n6966 , \Data_Mem/n6965 ,
         \Data_Mem/n6964 , \Data_Mem/n6963 , \Data_Mem/n6962 ,
         \Data_Mem/n6961 , \Data_Mem/n6960 , \Data_Mem/n6959 ,
         \Data_Mem/n6958 , \Data_Mem/n6957 , \Data_Mem/n6956 ,
         \Data_Mem/n6955 , \Data_Mem/n6954 , \Data_Mem/n6953 ,
         \Data_Mem/n6952 , \Data_Mem/n6951 , \Data_Mem/n6950 ,
         \Data_Mem/n6949 , \Data_Mem/n6948 , \Data_Mem/n6947 ,
         \Data_Mem/n6946 , \Data_Mem/n6945 , \Data_Mem/n6944 ,
         \Data_Mem/n6943 , \Data_Mem/n6942 , \Data_Mem/n6941 ,
         \Data_Mem/n6940 , \Data_Mem/n6939 , \Data_Mem/n6938 ,
         \Data_Mem/n6937 , \Data_Mem/n6936 , \Data_Mem/n6935 ,
         \Data_Mem/n6934 , \Data_Mem/n6933 , \Data_Mem/n6932 ,
         \Data_Mem/n6931 , \Data_Mem/n6930 , \Data_Mem/n6929 ,
         \Data_Mem/n6928 , \Data_Mem/n6927 , \Data_Mem/n6926 ,
         \Data_Mem/n6925 , \Data_Mem/n6924 , \Data_Mem/n6923 ,
         \Data_Mem/n6922 , \Data_Mem/n6921 , \Data_Mem/n6920 ,
         \Data_Mem/n6919 , \Data_Mem/n6918 , \Data_Mem/n6917 ,
         \Data_Mem/n6916 , \Data_Mem/n6915 , \Data_Mem/n6914 ,
         \Data_Mem/n6913 , \Data_Mem/n6912 , \Data_Mem/n6911 ,
         \Data_Mem/n6910 , \Data_Mem/n6909 , \Data_Mem/n6908 ,
         \Data_Mem/n6907 , \Data_Mem/n6906 , \Data_Mem/n6905 ,
         \Data_Mem/n6904 , \Data_Mem/n6903 , \Data_Mem/n6902 ,
         \Data_Mem/n6901 , \Data_Mem/n6900 , \Data_Mem/n6899 ,
         \Data_Mem/n6898 , \Data_Mem/n6897 , \Data_Mem/n6896 ,
         \Data_Mem/n6895 , \Data_Mem/n6894 , \Data_Mem/n6893 ,
         \Data_Mem/n6892 , \Data_Mem/n6891 , \Data_Mem/n6890 ,
         \Data_Mem/n6889 , \Data_Mem/n6888 , \Data_Mem/n6887 ,
         \Data_Mem/n6886 , \Data_Mem/n6885 , \Data_Mem/n6884 ,
         \Data_Mem/n6883 , \Data_Mem/n6882 , \Data_Mem/n6881 ,
         \Data_Mem/n6880 , \Data_Mem/n6879 , \Data_Mem/n6878 ,
         \Data_Mem/n6877 , \Data_Mem/n6876 , \Data_Mem/n6875 ,
         \Data_Mem/n6874 , \Data_Mem/n6873 , \Data_Mem/n6872 ,
         \Data_Mem/n6871 , \Data_Mem/n6870 , \Data_Mem/n6869 ,
         \Data_Mem/n6868 , \Data_Mem/n6867 , \Data_Mem/n6866 ,
         \Data_Mem/n6865 , \Data_Mem/n6864 , \Data_Mem/n6863 ,
         \Data_Mem/n6862 , \Data_Mem/n6861 , \Data_Mem/n6860 ,
         \Data_Mem/n6859 , \Data_Mem/n6858 , \Data_Mem/n6857 ,
         \Data_Mem/n6856 , \Data_Mem/n6855 , \Data_Mem/n6854 ,
         \Data_Mem/n6853 , \Data_Mem/n6852 , \Data_Mem/n6851 ,
         \Data_Mem/n6850 , \Data_Mem/n6849 , \Data_Mem/n6848 ,
         \Data_Mem/n6847 , \Data_Mem/n6846 , \Data_Mem/n6845 ,
         \Data_Mem/n6844 , \Data_Mem/n6843 , \Data_Mem/n6842 ,
         \Data_Mem/n6841 , \Data_Mem/n6840 , \Data_Mem/n6839 ,
         \Data_Mem/n6838 , \Data_Mem/n6837 , \Data_Mem/n6836 ,
         \Data_Mem/n6835 , \Data_Mem/n6834 , \Data_Mem/n6833 ,
         \Data_Mem/n6832 , \Data_Mem/n6831 , \Data_Mem/n6830 ,
         \Data_Mem/n6829 , \Data_Mem/n6828 , \Data_Mem/n6827 ,
         \Data_Mem/n6826 , \Data_Mem/n6825 , \Data_Mem/n6824 ,
         \Data_Mem/n6823 , \Data_Mem/n6822 , \Data_Mem/n6821 ,
         \Data_Mem/n6820 , \Data_Mem/n6819 , \Data_Mem/n6818 ,
         \Data_Mem/n6817 , \Data_Mem/n6816 , \Data_Mem/n6815 ,
         \Data_Mem/n6814 , \Data_Mem/n6813 , \Data_Mem/n6812 ,
         \Data_Mem/n6811 , \Data_Mem/n6810 , \Data_Mem/n6809 ,
         \Data_Mem/n6808 , \Data_Mem/n6807 , \Data_Mem/n6806 ,
         \Data_Mem/n6805 , \Data_Mem/n6804 , \Data_Mem/n6803 ,
         \Data_Mem/n6802 , \Data_Mem/n6801 , \Data_Mem/n6800 ,
         \Data_Mem/n6799 , \Data_Mem/n6798 , \Data_Mem/n6797 ,
         \Data_Mem/n6796 , \Data_Mem/n6795 , \Data_Mem/n6794 ,
         \Data_Mem/n6793 , \Data_Mem/n6792 , \Data_Mem/n6791 ,
         \Data_Mem/n6790 , \Data_Mem/n6789 , \Data_Mem/n6788 ,
         \Data_Mem/n6787 , \Data_Mem/n6786 , \Data_Mem/n6785 ,
         \Data_Mem/n6784 , \Data_Mem/n6783 , \Data_Mem/n6782 ,
         \Data_Mem/n6781 , \Data_Mem/n6780 , \Data_Mem/n6779 ,
         \Data_Mem/n6778 , \Data_Mem/n6777 , \Data_Mem/n6776 ,
         \Data_Mem/n6775 , \Data_Mem/n6774 , \Data_Mem/n6773 ,
         \Data_Mem/n6772 , \Data_Mem/n6771 , \Data_Mem/n6770 ,
         \Data_Mem/n6769 , \Data_Mem/n6768 , \Data_Mem/n6767 ,
         \Data_Mem/n6766 , \Data_Mem/n6765 , \Data_Mem/n6764 ,
         \Data_Mem/n6763 , \Data_Mem/n6762 , \Data_Mem/n6761 ,
         \Data_Mem/n6760 , \Data_Mem/n6759 , \Data_Mem/n6758 ,
         \Data_Mem/n6757 , \Data_Mem/n6756 , \Data_Mem/n6755 ,
         \Data_Mem/n6754 , \Data_Mem/n6753 , \Data_Mem/n6752 ,
         \Data_Mem/n6751 , \Data_Mem/n6750 , \Data_Mem/n6749 ,
         \Data_Mem/n6748 , \Data_Mem/n6747 , \Data_Mem/n6746 ,
         \Data_Mem/n6745 , \Data_Mem/n6744 , \Data_Mem/n6743 ,
         \Data_Mem/n6742 , \Data_Mem/n6741 , \Data_Mem/n6740 ,
         \Data_Mem/n6739 , \Data_Mem/n6738 , \Data_Mem/n6737 ,
         \Data_Mem/n6736 , \Data_Mem/n6735 , \Data_Mem/n6734 ,
         \Data_Mem/n6733 , \Data_Mem/n6732 , \Data_Mem/n6731 ,
         \Data_Mem/n6730 , \Data_Mem/n6729 , \Data_Mem/n6728 ,
         \Data_Mem/n6727 , \Data_Mem/n6726 , \Data_Mem/n6725 ,
         \Data_Mem/n6724 , \Data_Mem/n6723 , \Data_Mem/n6722 ,
         \Data_Mem/n6721 , \Data_Mem/n6720 , \Data_Mem/n6719 ,
         \Data_Mem/n6718 , \Data_Mem/n6717 , \Data_Mem/n6716 ,
         \Data_Mem/n6715 , \Data_Mem/n6714 , \Data_Mem/n6713 ,
         \Data_Mem/n6712 , \Data_Mem/n6711 , \Data_Mem/n6710 ,
         \Data_Mem/n6709 , \Data_Mem/n6708 , \Data_Mem/n6707 ,
         \Data_Mem/n6706 , \Data_Mem/n6705 , \Data_Mem/n6704 ,
         \Data_Mem/n6703 , \Data_Mem/n6702 , \Data_Mem/n6701 ,
         \Data_Mem/n6700 , \Data_Mem/n6699 , \Data_Mem/n6698 ,
         \Data_Mem/n6697 , \Data_Mem/n6696 , \Data_Mem/n6695 ,
         \Data_Mem/n6694 , \Data_Mem/n6693 , \Data_Mem/n6692 ,
         \Data_Mem/n6691 , \Data_Mem/n6690 , \Data_Mem/n6689 ,
         \Data_Mem/n6688 , \Data_Mem/n6687 , \Data_Mem/n6686 ,
         \Data_Mem/n6685 , \Data_Mem/n6684 , \Data_Mem/n6683 ,
         \Data_Mem/n6682 , \Data_Mem/n6681 , \Data_Mem/n6680 ,
         \Data_Mem/n6679 , \Data_Mem/n6678 , \Data_Mem/n6677 ,
         \Data_Mem/n6676 , \Data_Mem/n6675 , \Data_Mem/n6674 ,
         \Data_Mem/n6673 , \Data_Mem/n6672 , \Data_Mem/n6671 ,
         \Data_Mem/n6670 , \Data_Mem/n6669 , \Data_Mem/n6668 ,
         \Data_Mem/n6667 , \Data_Mem/n6666 , \Data_Mem/n6665 ,
         \Data_Mem/n6664 , \Data_Mem/n6663 , \Data_Mem/n6662 ,
         \Data_Mem/n6661 , \Data_Mem/n6660 , \Data_Mem/n6659 ,
         \Data_Mem/n6658 , \Data_Mem/n6657 , \Data_Mem/n6656 ,
         \Data_Mem/n6655 , \Data_Mem/n6654 , \Data_Mem/n6653 ,
         \Data_Mem/n6652 , \Data_Mem/n6651 , \Data_Mem/n6650 ,
         \Data_Mem/n6649 , \Data_Mem/n6648 , \Data_Mem/n6647 ,
         \Data_Mem/n6646 , \Data_Mem/n6645 , \Data_Mem/n6644 ,
         \Data_Mem/n6643 , \Data_Mem/n6642 , \Data_Mem/n6641 ,
         \Data_Mem/n6640 , \Data_Mem/n6639 , \Data_Mem/n6638 ,
         \Data_Mem/n6637 , \Data_Mem/n6636 , \Data_Mem/n6635 ,
         \Data_Mem/n6634 , \Data_Mem/n6633 , \Data_Mem/n6632 ,
         \Data_Mem/n6631 , \Data_Mem/n6630 , \Data_Mem/n6629 ,
         \Data_Mem/n6628 , \Data_Mem/n6627 , \Data_Mem/n6626 ,
         \Data_Mem/n6625 , \Data_Mem/n6624 , \Data_Mem/n6623 ,
         \Data_Mem/n6622 , \Data_Mem/n6621 , \Data_Mem/n6620 ,
         \Data_Mem/n6619 , \Data_Mem/n6618 , \Data_Mem/n6617 ,
         \Data_Mem/n6616 , \Data_Mem/n6615 , \Data_Mem/n6614 ,
         \Data_Mem/n6613 , \Data_Mem/n6612 , \Data_Mem/n6611 ,
         \Data_Mem/n6610 , \Data_Mem/n6609 , \Data_Mem/n6608 ,
         \Data_Mem/n6607 , \Data_Mem/n6606 , \Data_Mem/n6605 ,
         \Data_Mem/n6604 , \Data_Mem/n6603 , \Data_Mem/n6602 ,
         \Data_Mem/n6601 , \Data_Mem/n6600 , \Data_Mem/n6599 ,
         \Data_Mem/n6598 , \Data_Mem/n6597 , \Data_Mem/n6596 ,
         \Data_Mem/n6595 , \Data_Mem/n6594 , \Data_Mem/n6593 ,
         \Data_Mem/n6592 , \Data_Mem/n6591 , \Data_Mem/n6590 ,
         \Data_Mem/n6589 , \Data_Mem/n6588 , \Data_Mem/n6587 ,
         \Data_Mem/n6586 , \Data_Mem/n6585 , \Data_Mem/n6584 ,
         \Data_Mem/n6583 , \Data_Mem/n6582 , \Data_Mem/n6581 ,
         \Data_Mem/n6580 , \Data_Mem/n6579 , \Data_Mem/n6578 ,
         \Data_Mem/n6577 , \Data_Mem/n6576 , \Data_Mem/n6575 ,
         \Data_Mem/n6574 , \Data_Mem/n6573 , \Data_Mem/n6572 ,
         \Data_Mem/n6571 , \Data_Mem/n6570 , \Data_Mem/n6569 ,
         \Data_Mem/n6568 , \Data_Mem/n6567 , \Data_Mem/n6566 ,
         \Data_Mem/n6565 , \Data_Mem/n6564 , \Data_Mem/n6563 ,
         \Data_Mem/n6562 , \Data_Mem/n6561 , \Data_Mem/n6560 ,
         \Data_Mem/n6559 , \Data_Mem/n6558 , \Data_Mem/n6557 ,
         \Data_Mem/n6556 , \Data_Mem/n6555 , \Data_Mem/n6554 ,
         \Data_Mem/n6553 , \Data_Mem/n6552 , \Data_Mem/n6551 ,
         \Data_Mem/n6550 , \Data_Mem/n6549 , \Data_Mem/n6548 ,
         \Data_Mem/n6547 , \Data_Mem/n6546 , \Data_Mem/n6545 ,
         \Data_Mem/n6544 , \Data_Mem/n6543 , \Data_Mem/n6542 ,
         \Data_Mem/n6541 , \Data_Mem/n6540 , \Data_Mem/n6539 ,
         \Data_Mem/n6538 , \Data_Mem/n6537 , \Data_Mem/n6536 ,
         \Data_Mem/n6535 , \Data_Mem/n6534 , \Data_Mem/n6533 ,
         \Data_Mem/n6532 , \Data_Mem/n6531 , \Data_Mem/n6530 ,
         \Data_Mem/n6529 , \Data_Mem/n6528 , \Data_Mem/n6527 ,
         \Data_Mem/n6526 , \Data_Mem/n6525 , \Data_Mem/n6524 ,
         \Data_Mem/n6523 , \Data_Mem/n6522 , \Data_Mem/n6521 ,
         \Data_Mem/n6520 , \Data_Mem/n6519 , \Data_Mem/n6518 ,
         \Data_Mem/n6517 , \Data_Mem/n6516 , \Data_Mem/n6515 ,
         \Data_Mem/n6514 , \Data_Mem/n6513 , \Data_Mem/n6512 ,
         \Data_Mem/n6511 , \Data_Mem/n6510 , \Data_Mem/n6509 ,
         \Data_Mem/n6508 , \Data_Mem/n6507 , \Data_Mem/n6506 ,
         \Data_Mem/n6505 , \Data_Mem/n6504 , \Data_Mem/n6503 ,
         \Data_Mem/n6502 , \Data_Mem/n6501 , \Data_Mem/n6500 ,
         \Data_Mem/n6499 , \Data_Mem/n6498 , \Data_Mem/n6497 ,
         \Data_Mem/n6496 , \Data_Mem/n6495 , \Data_Mem/n6494 ,
         \Data_Mem/n6493 , \Data_Mem/n6492 , \Data_Mem/n6491 ,
         \Data_Mem/n6490 , \Data_Mem/n6489 , \Data_Mem/n6488 ,
         \Data_Mem/n6487 , \Data_Mem/n6486 , \Data_Mem/n6485 ,
         \Data_Mem/n6484 , \Data_Mem/n6483 , \Data_Mem/n6482 ,
         \Data_Mem/n6481 , \Data_Mem/n6480 , \Data_Mem/n6479 ,
         \Data_Mem/n6478 , \Data_Mem/n6477 , \Data_Mem/n6476 ,
         \Data_Mem/n6475 , \Data_Mem/n6474 , \Data_Mem/n6473 ,
         \Data_Mem/n6472 , \Data_Mem/n6471 , \Data_Mem/n6470 ,
         \Data_Mem/n6469 , \Data_Mem/n6468 , \Data_Mem/n6467 ,
         \Data_Mem/n6466 , \Data_Mem/n6465 , \Data_Mem/n6464 ,
         \Data_Mem/n6463 , \Data_Mem/n6462 , \Data_Mem/n6461 ,
         \Data_Mem/n6460 , \Data_Mem/n6459 , \Data_Mem/n6458 ,
         \Data_Mem/n6457 , \Data_Mem/n6456 , \Data_Mem/n6455 ,
         \Data_Mem/n6454 , \Data_Mem/n6453 , \Data_Mem/n6452 ,
         \Data_Mem/n6451 , \Data_Mem/n6450 , \Data_Mem/n6449 ,
         \Data_Mem/n6448 , \Data_Mem/n6447 , \Data_Mem/n6446 ,
         \Data_Mem/n6445 , \Data_Mem/n6444 , \Data_Mem/n6443 ,
         \Data_Mem/n6442 , \Data_Mem/n6441 , \Data_Mem/n6440 ,
         \Data_Mem/n6439 , \Data_Mem/n6438 , \Data_Mem/n6437 ,
         \Data_Mem/n6436 , \Data_Mem/n6435 , \Data_Mem/n6434 ,
         \Data_Mem/n6433 , \Data_Mem/n6432 , \Data_Mem/n6431 ,
         \Data_Mem/n6430 , \Data_Mem/n6429 , \Data_Mem/n6428 ,
         \Data_Mem/n6427 , \Data_Mem/n6426 , \Data_Mem/n6425 ,
         \Data_Mem/n6424 , \Data_Mem/n6423 , \Data_Mem/n6422 ,
         \Data_Mem/n6421 , \Data_Mem/n6420 , \Data_Mem/n6419 ,
         \Data_Mem/n6418 , \Data_Mem/n6417 , \Data_Mem/n6416 ,
         \Data_Mem/n6415 , \Data_Mem/n6414 , \Data_Mem/n6413 ,
         \Data_Mem/n6412 , \Data_Mem/n6411 , \Data_Mem/n6410 ,
         \Data_Mem/n6409 , \Data_Mem/n6408 , \Data_Mem/n6407 ,
         \Data_Mem/n6406 , \Data_Mem/n6405 , \Data_Mem/n6404 ,
         \Data_Mem/n6403 , \Data_Mem/n6402 , \Data_Mem/n6401 ,
         \Data_Mem/n6400 , \Data_Mem/n6399 , \Data_Mem/n6398 ,
         \Data_Mem/n6397 , \Data_Mem/n6396 , \Data_Mem/n6395 ,
         \Data_Mem/n6394 , \Data_Mem/n6393 , \Data_Mem/n6392 ,
         \Data_Mem/n6391 , \Data_Mem/n6390 , \Data_Mem/n6389 ,
         \Data_Mem/n6388 , \Data_Mem/n6387 , \Data_Mem/n6386 ,
         \Data_Mem/n6385 , \Data_Mem/n6384 , \Data_Mem/n6383 ,
         \Data_Mem/n6382 , \Data_Mem/n6381 , \Data_Mem/n6380 ,
         \Data_Mem/n6379 , \Data_Mem/n6378 , \Data_Mem/n6377 ,
         \Data_Mem/n6376 , \Data_Mem/n6375 , \Data_Mem/n6374 ,
         \Data_Mem/n6373 , \Data_Mem/n6372 , \Data_Mem/n6371 ,
         \Data_Mem/n6370 , \Data_Mem/n6369 , \Data_Mem/n6368 ,
         \Data_Mem/n6367 , \Data_Mem/n6366 , \Data_Mem/n6365 ,
         \Data_Mem/n6364 , \Data_Mem/n6363 , \Data_Mem/n6362 ,
         \Data_Mem/n6361 , \Data_Mem/n6360 , \Data_Mem/n6359 ,
         \Data_Mem/n6358 , \Data_Mem/n6357 , \Data_Mem/n6356 ,
         \Data_Mem/n6355 , \Data_Mem/n6354 , \Data_Mem/n6353 ,
         \Data_Mem/n6352 , \Data_Mem/n6351 , \Data_Mem/n6350 ,
         \Data_Mem/n6349 , \Data_Mem/n6348 , \Data_Mem/n6347 ,
         \Data_Mem/n6346 , \Data_Mem/n6345 , \Data_Mem/n6344 ,
         \Data_Mem/n6343 , \Data_Mem/n6342 , \Data_Mem/n6341 ,
         \Data_Mem/n6340 , \Data_Mem/n6339 , \Data_Mem/n6338 ,
         \Data_Mem/n6337 , \Data_Mem/n6336 , \Data_Mem/n6335 ,
         \Data_Mem/n6334 , \Data_Mem/n6333 , \Data_Mem/n6332 ,
         \Data_Mem/n6331 , \Data_Mem/n6330 , \Data_Mem/n6329 ,
         \Data_Mem/n6328 , \Data_Mem/n6327 , \Data_Mem/n6326 ,
         \Data_Mem/n6325 , \Data_Mem/n6324 , \Data_Mem/n6323 ,
         \Data_Mem/n6322 , \Data_Mem/n6321 , \Data_Mem/n6320 ,
         \Data_Mem/n6319 , \Data_Mem/n6318 , \Data_Mem/n6317 ,
         \Data_Mem/n6316 , \Data_Mem/n6315 , \Data_Mem/n6314 ,
         \Data_Mem/n6313 , \Data_Mem/n6312 , \Data_Mem/n6311 ,
         \Data_Mem/n6310 , \Data_Mem/n6309 , \Data_Mem/n6308 ,
         \Data_Mem/n6307 , \Data_Mem/n6306 , \Data_Mem/n6305 ,
         \Data_Mem/n6304 , \Data_Mem/n6303 , \Data_Mem/n6302 ,
         \Data_Mem/n6301 , \Data_Mem/n6300 , \Data_Mem/n6299 ,
         \Data_Mem/n6298 , \Data_Mem/n6297 , \Data_Mem/n6296 ,
         \Data_Mem/n6295 , \Data_Mem/n6294 , \Data_Mem/n6293 ,
         \Data_Mem/n6292 , \Data_Mem/n6291 , \Data_Mem/n6290 ,
         \Data_Mem/n6289 , \Data_Mem/n6288 , \Data_Mem/n6287 ,
         \Data_Mem/n6286 , \Data_Mem/n6285 , \Data_Mem/n6284 ,
         \Data_Mem/n6283 , \Data_Mem/n6282 , \Data_Mem/n6281 ,
         \Data_Mem/n6280 , \Data_Mem/n6279 , \Data_Mem/n6278 ,
         \Data_Mem/n6277 , \Data_Mem/n6276 , \Data_Mem/n6275 ,
         \Data_Mem/n6274 , \Data_Mem/n6273 , \Data_Mem/n6272 ,
         \Data_Mem/n6271 , \Data_Mem/n6270 , \Data_Mem/n6269 ,
         \Data_Mem/n6268 , \Data_Mem/n6267 , \Data_Mem/n6266 ,
         \Data_Mem/n6265 , \Data_Mem/n6264 , \Data_Mem/n6263 ,
         \Data_Mem/n6262 , \Data_Mem/n6261 , \Data_Mem/n6260 ,
         \Data_Mem/n6259 , \Data_Mem/n6258 , \Data_Mem/n6257 ,
         \Data_Mem/n6256 , \Data_Mem/n6255 , \Data_Mem/n6254 ,
         \Data_Mem/n6253 , \Data_Mem/n6252 , \Data_Mem/n6251 ,
         \Data_Mem/n6250 , \Data_Mem/n6249 , \Data_Mem/n6248 ,
         \Data_Mem/n6247 , \Data_Mem/n6246 , \Data_Mem/n6245 ,
         \Data_Mem/n6244 , \Data_Mem/n6243 , \Data_Mem/n6242 ,
         \Data_Mem/n6241 , \Data_Mem/n6240 , \Data_Mem/n6239 ,
         \Data_Mem/n6238 , \Data_Mem/n6237 , \Data_Mem/n6236 ,
         \Data_Mem/n6235 , \Data_Mem/n6234 , \Data_Mem/n6233 ,
         \Data_Mem/n6232 , \Data_Mem/n6231 , \Data_Mem/n6230 ,
         \Data_Mem/n6229 , \Data_Mem/n6228 , \Data_Mem/n6227 ,
         \Data_Mem/n6226 , \Data_Mem/n6225 , \Data_Mem/n6224 ,
         \Data_Mem/n6223 , \Data_Mem/n6222 , \Data_Mem/n6221 ,
         \Data_Mem/n6220 , \Data_Mem/n6219 , \Data_Mem/n6218 ,
         \Data_Mem/n6217 , \Data_Mem/n6216 , \Data_Mem/n6215 ,
         \Data_Mem/n6214 , \Data_Mem/n6213 , \Data_Mem/n6212 ,
         \Data_Mem/n6211 , \Data_Mem/n6210 , \Data_Mem/n6209 ,
         \Data_Mem/n6208 , \Data_Mem/n6207 , \Data_Mem/n6206 ,
         \Data_Mem/n6205 , \Data_Mem/n6204 , \Data_Mem/n6203 ,
         \Data_Mem/n6202 , \Data_Mem/n6201 , \Data_Mem/n6200 ,
         \Data_Mem/n6199 , \Data_Mem/n6198 , \Data_Mem/n6197 ,
         \Data_Mem/n6196 , \Data_Mem/n6195 , \Data_Mem/n6194 ,
         \Data_Mem/n6193 , \Data_Mem/n6192 , \Data_Mem/n6191 ,
         \Data_Mem/n6190 , \Data_Mem/n6189 , \Data_Mem/n6188 ,
         \Data_Mem/n6187 , \Data_Mem/n6186 , \Data_Mem/n6185 ,
         \Data_Mem/n6184 , \Data_Mem/n6183 , \Data_Mem/n6182 ,
         \Data_Mem/n6181 , \Data_Mem/n6180 , \Data_Mem/n6179 ,
         \Data_Mem/n6178 , \Data_Mem/n6177 , \Data_Mem/n6176 ,
         \Data_Mem/n6175 , \Data_Mem/n6174 , \Data_Mem/n6173 ,
         \Data_Mem/n6172 , \Data_Mem/n6171 , \Data_Mem/n6170 ,
         \Data_Mem/n6169 , \Data_Mem/n6168 , \Data_Mem/n6167 ,
         \Data_Mem/n6166 , \Data_Mem/n6165 , \Data_Mem/n6164 ,
         \Data_Mem/n6163 , \Data_Mem/n6162 , \Data_Mem/n6161 ,
         \Data_Mem/n6160 , \Data_Mem/n6159 , \Data_Mem/n6158 ,
         \Data_Mem/n6157 , \Data_Mem/n6156 , \Data_Mem/n6155 ,
         \Data_Mem/n6154 , \Data_Mem/n6153 , \Data_Mem/n6152 ,
         \Data_Mem/n6151 , \Data_Mem/n6150 , \Data_Mem/n6149 ,
         \Data_Mem/n6148 , \Data_Mem/n6147 , \Data_Mem/n6146 ,
         \Data_Mem/n6145 , \Data_Mem/n6144 , \Data_Mem/n6143 ,
         \Data_Mem/n6142 , \Data_Mem/n6141 , \Data_Mem/n6140 ,
         \Data_Mem/n6139 , \Data_Mem/n6138 , \Data_Mem/n6137 ,
         \Data_Mem/n6136 , \Data_Mem/n6135 , \Data_Mem/n6134 ,
         \Data_Mem/n6133 , \Data_Mem/n6132 , \Data_Mem/n6131 ,
         \Data_Mem/n6130 , \Data_Mem/n6129 , \Data_Mem/n6128 ,
         \Data_Mem/n6127 , \Data_Mem/n6126 , \Data_Mem/n6125 ,
         \Data_Mem/n6124 , \Data_Mem/n6123 , \Data_Mem/n6122 ,
         \Data_Mem/n6121 , \Data_Mem/n6120 , \Data_Mem/n6119 ,
         \Data_Mem/n6118 , \Data_Mem/n6117 , \Data_Mem/n6116 ,
         \Data_Mem/n6115 , \Data_Mem/n6114 , \Data_Mem/n6113 ,
         \Data_Mem/n6112 , \Data_Mem/n6111 , \Data_Mem/n6110 ,
         \Data_Mem/n6109 , \Data_Mem/n6108 , \Data_Mem/n6107 ,
         \Data_Mem/n6106 , \Data_Mem/n6105 , \Data_Mem/n6104 ,
         \Data_Mem/n6103 , \Data_Mem/n6102 , \Data_Mem/n6101 ,
         \Data_Mem/n6100 , \Data_Mem/n6099 , \Data_Mem/n6098 ,
         \Data_Mem/n6097 , \Data_Mem/n6096 , \Data_Mem/n6095 ,
         \Data_Mem/n6094 , \Data_Mem/n6093 , \Data_Mem/n6092 ,
         \Data_Mem/n6091 , \Data_Mem/n6090 , \Data_Mem/n6089 ,
         \Data_Mem/n6088 , \Data_Mem/n6087 , \Data_Mem/n6086 ,
         \Data_Mem/n6085 , \Data_Mem/n6084 , \Data_Mem/n6083 ,
         \Data_Mem/n6082 , \Data_Mem/n6081 , \Data_Mem/n6080 ,
         \Data_Mem/n6079 , \Data_Mem/n6078 , \Data_Mem/n6077 ,
         \Data_Mem/n6076 , \Data_Mem/n6075 , \Data_Mem/n6074 ,
         \Data_Mem/n6073 , \Data_Mem/n6072 , \Data_Mem/n6071 ,
         \Data_Mem/n6070 , \Data_Mem/n6069 , \Data_Mem/n6068 ,
         \Data_Mem/n6067 , \Data_Mem/n6066 , \Data_Mem/n6065 ,
         \Data_Mem/n6064 , \Data_Mem/n6063 , \Data_Mem/n6062 ,
         \Data_Mem/n6061 , \Data_Mem/n6060 , \Data_Mem/n6059 ,
         \Data_Mem/n6058 , \Data_Mem/n6057 , \Data_Mem/n6056 ,
         \Data_Mem/n6055 , \Data_Mem/n6054 , \Data_Mem/n6053 ,
         \Data_Mem/n6052 , \Data_Mem/n6051 , \Data_Mem/n6050 ,
         \Data_Mem/n6049 , \Data_Mem/n6048 , \Data_Mem/n6047 ,
         \Data_Mem/n6046 , \Data_Mem/n6045 , \Data_Mem/n6044 ,
         \Data_Mem/n6043 , \Data_Mem/n6042 , \Data_Mem/n6041 ,
         \Data_Mem/n6040 , \Data_Mem/n6039 , \Data_Mem/n6038 ,
         \Data_Mem/n6037 , \Data_Mem/n6036 , \Data_Mem/n6035 ,
         \Data_Mem/n6034 , \Data_Mem/n6033 , \Data_Mem/n6032 ,
         \Data_Mem/n6031 , \Data_Mem/n6030 , \Data_Mem/n6029 ,
         \Data_Mem/n6028 , \Data_Mem/n6027 , \Data_Mem/n6026 ,
         \Data_Mem/n6025 , \Data_Mem/n6024 , \Data_Mem/n6023 ,
         \Data_Mem/n6022 , \Data_Mem/n6021 , \Data_Mem/n6020 ,
         \Data_Mem/n6019 , \Data_Mem/n6018 , \Data_Mem/n6017 ,
         \Data_Mem/n6016 , \Data_Mem/n6015 , \Data_Mem/n6014 ,
         \Data_Mem/n6013 , \Data_Mem/n6012 , \Data_Mem/n6011 ,
         \Data_Mem/n6010 , \Data_Mem/n6009 , \Data_Mem/n6008 ,
         \Data_Mem/n6007 , \Data_Mem/n6006 , \Data_Mem/n6005 ,
         \Data_Mem/n6004 , \Data_Mem/n6003 , \Data_Mem/n6002 ,
         \Data_Mem/n6001 , \Data_Mem/n6000 , \Data_Mem/n5999 ,
         \Data_Mem/n5998 , \Data_Mem/n5997 , \Data_Mem/n5996 ,
         \Data_Mem/n5995 , \Data_Mem/n5994 , \Data_Mem/n5993 ,
         \Data_Mem/n5992 , \Data_Mem/n5991 , \Data_Mem/n5990 ,
         \Data_Mem/n5989 , \Data_Mem/n5988 , \Data_Mem/n5987 ,
         \Data_Mem/n5986 , \Data_Mem/n5985 , \Data_Mem/n5984 ,
         \Data_Mem/n5983 , \Data_Mem/n5982 , \Data_Mem/n5981 ,
         \Data_Mem/n5980 , \Data_Mem/n5979 , \Data_Mem/n5978 ,
         \Data_Mem/n5977 , \Data_Mem/n5976 , \Data_Mem/n5975 ,
         \Data_Mem/n5974 , \Data_Mem/n5973 , \Data_Mem/n5972 ,
         \Data_Mem/n5971 , \Data_Mem/n5970 , \Data_Mem/n5969 ,
         \Data_Mem/n5968 , \Data_Mem/n5967 , \Data_Mem/n5966 ,
         \Data_Mem/n5965 , \Data_Mem/n5964 , \Data_Mem/n5963 ,
         \Data_Mem/n5962 , \Data_Mem/n5961 , \Data_Mem/n5960 ,
         \Data_Mem/n5959 , \Data_Mem/n5958 , \Data_Mem/n5957 ,
         \Data_Mem/n5956 , \Data_Mem/n5955 , \Data_Mem/n5954 ,
         \Data_Mem/n5953 , \Data_Mem/n5952 , \Data_Mem/n5951 ,
         \Data_Mem/n5950 , \Data_Mem/n5949 , \Data_Mem/n5948 ,
         \Data_Mem/n5947 , \Data_Mem/n5946 , \Data_Mem/n5945 ,
         \Data_Mem/n5944 , \Data_Mem/n5943 , \Data_Mem/n5942 ,
         \Data_Mem/n5941 , \Data_Mem/n5940 , \Data_Mem/n5939 ,
         \Data_Mem/n5938 , \Data_Mem/n5937 , \Data_Mem/n5936 ,
         \Data_Mem/n5935 , \Data_Mem/n5934 , \Data_Mem/n5933 ,
         \Data_Mem/n5932 , \Data_Mem/n5931 , \Data_Mem/n5930 ,
         \Data_Mem/n5929 , \Data_Mem/n5928 , \Data_Mem/n5927 ,
         \Data_Mem/n5926 , \Data_Mem/n5925 , \Data_Mem/n5924 ,
         \Data_Mem/n5923 , \Data_Mem/n5922 , \Data_Mem/n5921 ,
         \Data_Mem/n5920 , \Data_Mem/n5919 , \Data_Mem/n5918 ,
         \Data_Mem/n5917 , \Data_Mem/n5916 , \Data_Mem/n5915 ,
         \Data_Mem/n5914 , \Data_Mem/n5913 , \Data_Mem/n5912 ,
         \Data_Mem/n5911 , \Data_Mem/n5910 , \Data_Mem/n5909 ,
         \Data_Mem/n5908 , \Data_Mem/n5907 , \Data_Mem/n5906 ,
         \Data_Mem/n5905 , \Data_Mem/n5904 , \Data_Mem/n5903 ,
         \Data_Mem/n5902 , \Data_Mem/n5901 , \Data_Mem/n5900 ,
         \Data_Mem/n5899 , \Data_Mem/n5898 , \Data_Mem/n5897 ,
         \Data_Mem/n5896 , \Data_Mem/n5895 , \Data_Mem/n5894 ,
         \Data_Mem/n5893 , \Data_Mem/n5892 , \Data_Mem/n5891 ,
         \Data_Mem/n5890 , \Data_Mem/n5889 , \Data_Mem/n5888 ,
         \Data_Mem/n5887 , \Data_Mem/n5886 , \Data_Mem/n5885 ,
         \Data_Mem/n5884 , \Data_Mem/n5883 , \Data_Mem/n5882 ,
         \Data_Mem/n5881 , \Data_Mem/n5880 , \Data_Mem/n5879 ,
         \Data_Mem/n5878 , \Data_Mem/n5877 , \Data_Mem/n5876 ,
         \Data_Mem/n5875 , \Data_Mem/n5874 , \Data_Mem/n5873 ,
         \Data_Mem/n5872 , \Data_Mem/n5871 , \Data_Mem/n5870 ,
         \Data_Mem/n5869 , \Data_Mem/n5868 , \Data_Mem/n5867 ,
         \Data_Mem/n5866 , \Data_Mem/n5865 , \Data_Mem/n5864 ,
         \Data_Mem/n5863 , \Data_Mem/n5862 , \Data_Mem/n5861 ,
         \Data_Mem/n5860 , \Data_Mem/n5859 , \Data_Mem/n5858 ,
         \Data_Mem/n5857 , \Data_Mem/n5856 , \Data_Mem/n5855 ,
         \Data_Mem/n5854 , \Data_Mem/n5853 , \Data_Mem/n5852 ,
         \Data_Mem/n5851 , \Data_Mem/n5850 , \Data_Mem/n5849 ,
         \Data_Mem/n5848 , \Data_Mem/n5847 , \Data_Mem/n5846 ,
         \Data_Mem/n5845 , \Data_Mem/n5844 , \Data_Mem/n5843 ,
         \Data_Mem/n5842 , \Data_Mem/n5841 , \Data_Mem/n5840 ,
         \Data_Mem/n5839 , \Data_Mem/n5838 , \Data_Mem/n5837 ,
         \Data_Mem/n5836 , \Data_Mem/n5835 , \Data_Mem/n5834 ,
         \Data_Mem/n5833 , \Data_Mem/n5832 , \Data_Mem/n5831 ,
         \Data_Mem/n5830 , \Data_Mem/n5829 , \Data_Mem/n5828 ,
         \Data_Mem/n5827 , \Data_Mem/n5826 , \Data_Mem/n5825 ,
         \Data_Mem/n5824 , \Data_Mem/n5823 , \Data_Mem/n5822 ,
         \Data_Mem/n5821 , \Data_Mem/n5820 , \Data_Mem/n5819 ,
         \Data_Mem/n5818 , \Data_Mem/n5817 , \Data_Mem/n5816 ,
         \Data_Mem/n5815 , \Data_Mem/n5814 , \Data_Mem/n5813 ,
         \Data_Mem/n5812 , \Data_Mem/n5811 , \Data_Mem/n5810 ,
         \Data_Mem/n5809 , \Data_Mem/n5808 , \Data_Mem/n5807 ,
         \Data_Mem/n5806 , \Data_Mem/n5805 , \Data_Mem/n5804 ,
         \Data_Mem/n5803 , \Data_Mem/n5802 , \Data_Mem/n5801 ,
         \Data_Mem/n5800 , \Data_Mem/n5799 , \Data_Mem/n5798 ,
         \Data_Mem/n5797 , \Data_Mem/n5796 , \Data_Mem/n5795 ,
         \Data_Mem/n5794 , \Data_Mem/n5793 , \Data_Mem/n5792 ,
         \Data_Mem/n5791 , \Data_Mem/n5790 , \Data_Mem/n5789 ,
         \Data_Mem/n5788 , \Data_Mem/n5787 , \Data_Mem/n5786 ,
         \Data_Mem/n5785 , \Data_Mem/n5784 , \Data_Mem/n5783 ,
         \Data_Mem/n5782 , \Data_Mem/n5781 , \Data_Mem/n5780 ,
         \Data_Mem/n5779 , \Data_Mem/n5778 , \Data_Mem/n5777 ,
         \Data_Mem/n5776 , \Data_Mem/n5775 , \Data_Mem/n5774 ,
         \Data_Mem/n5773 , \Data_Mem/n5772 , \Data_Mem/n5771 ,
         \Data_Mem/n5770 , \Data_Mem/n5769 , \Data_Mem/n5768 ,
         \Data_Mem/n5767 , \Data_Mem/n5766 , \Data_Mem/n5765 ,
         \Data_Mem/n5764 , \Data_Mem/n5763 , \Data_Mem/n5762 ,
         \Data_Mem/n5761 , \Data_Mem/n5760 , \Data_Mem/n5759 ,
         \Data_Mem/n5758 , \Data_Mem/n5757 , \Data_Mem/n5756 ,
         \Data_Mem/n5755 , \Data_Mem/n5754 , \Data_Mem/n5753 ,
         \Data_Mem/n5752 , \Data_Mem/n5751 , \Data_Mem/n5750 ,
         \Data_Mem/n5749 , \Data_Mem/n5748 , \Data_Mem/n5747 ,
         \Data_Mem/n5746 , \Data_Mem/n5745 , \Data_Mem/n5744 ,
         \Data_Mem/n5743 , \Data_Mem/n5742 , \Data_Mem/n5741 ,
         \Data_Mem/n5740 , \Data_Mem/n5739 , \Data_Mem/n5738 ,
         \Data_Mem/n5737 , \Data_Mem/n5736 , \Data_Mem/n5735 ,
         \Data_Mem/n5734 , \Data_Mem/n5733 , \Data_Mem/n5732 ,
         \Data_Mem/n5731 , \Data_Mem/n5730 , \Data_Mem/n5729 ,
         \Data_Mem/n5728 , \Data_Mem/n5727 , \Data_Mem/n5726 ,
         \Data_Mem/n5725 , \Data_Mem/n5724 , \Data_Mem/n5723 ,
         \Data_Mem/n5722 , \Data_Mem/n5721 , \Data_Mem/n5720 ,
         \Data_Mem/n5719 , \Data_Mem/n5718 , \Data_Mem/n5717 ,
         \Data_Mem/n5716 , \Data_Mem/n5715 , \Data_Mem/n5714 ,
         \Data_Mem/n5713 , \Data_Mem/n5712 , \Data_Mem/n5711 ,
         \Data_Mem/n5710 , \Data_Mem/n5709 , \Data_Mem/n5708 ,
         \Data_Mem/n5707 , \Data_Mem/n5706 , \Data_Mem/n5705 ,
         \Data_Mem/n5704 , \Data_Mem/n5703 , \Data_Mem/n5702 ,
         \Data_Mem/n5701 , \Data_Mem/n5700 , \Data_Mem/n5699 ,
         \Data_Mem/n5698 , \Data_Mem/n5697 , \Data_Mem/n5696 ,
         \Data_Mem/n5695 , \Data_Mem/n5694 , \Data_Mem/n5693 ,
         \Data_Mem/n5692 , \Data_Mem/n5691 , \Data_Mem/n5690 ,
         \Data_Mem/n5689 , \Data_Mem/n5688 , \Data_Mem/n5687 ,
         \Data_Mem/n5686 , \Data_Mem/n5685 , \Data_Mem/n5684 ,
         \Data_Mem/n5683 , \Data_Mem/n5682 , \Data_Mem/n5681 ,
         \Data_Mem/n5680 , \Data_Mem/n5679 , \Data_Mem/n5678 ,
         \Data_Mem/n5677 , \Data_Mem/n5676 , \Data_Mem/n5675 ,
         \Data_Mem/n5674 , \Data_Mem/n5673 , \Data_Mem/n5672 ,
         \Data_Mem/n5671 , \Data_Mem/n5670 , \Data_Mem/n5669 ,
         \Data_Mem/n5668 , \Data_Mem/n5667 , \Data_Mem/n5666 ,
         \Data_Mem/n5665 , \Data_Mem/n5664 , \Data_Mem/n5663 ,
         \Data_Mem/n5662 , \Data_Mem/n5661 , \Data_Mem/n5660 ,
         \Data_Mem/n5659 , \Data_Mem/n5658 , \Data_Mem/n5657 ,
         \Data_Mem/n5656 , \Data_Mem/n5655 , \Data_Mem/n5654 ,
         \Data_Mem/n5653 , \Data_Mem/n5652 , \Data_Mem/n5651 ,
         \Data_Mem/n5650 , \Data_Mem/n5649 , \Data_Mem/n5648 ,
         \Data_Mem/n5647 , \Data_Mem/n5646 , \Data_Mem/n5645 ,
         \Data_Mem/n5644 , \Data_Mem/n5643 , \Data_Mem/n5642 ,
         \Data_Mem/n5641 , \Data_Mem/n5640 , \Data_Mem/n5639 ,
         \Data_Mem/n5638 , \Data_Mem/n5637 , \Data_Mem/n5636 ,
         \Data_Mem/n5635 , \Data_Mem/n5634 , \Data_Mem/n5633 ,
         \Data_Mem/n5632 , \Data_Mem/n5631 , \Data_Mem/n5630 ,
         \Data_Mem/n5629 , \Data_Mem/n5628 , \Data_Mem/n5627 ,
         \Data_Mem/n5626 , \Data_Mem/n5625 , \Data_Mem/n5624 ,
         \Data_Mem/n5623 , \Data_Mem/n5622 , \Data_Mem/n5621 ,
         \Data_Mem/n5620 , \Data_Mem/n5619 , \Data_Mem/n5618 ,
         \Data_Mem/n5617 , \Data_Mem/n5616 , \Data_Mem/n5615 ,
         \Data_Mem/n5614 , \Data_Mem/n5613 , \Data_Mem/n5612 ,
         \Data_Mem/n5611 , \Data_Mem/n5610 , \Data_Mem/n5609 ,
         \Data_Mem/n5608 , \Data_Mem/n5607 , \Data_Mem/n5606 ,
         \Data_Mem/n5605 , \Data_Mem/n5604 , \Data_Mem/n5603 ,
         \Data_Mem/n5602 , \Data_Mem/n5601 , \Data_Mem/n5600 ,
         \Data_Mem/n5599 , \Data_Mem/n5598 , \Data_Mem/n5597 ,
         \Data_Mem/n5596 , \Data_Mem/n5595 , \Data_Mem/n5594 ,
         \Data_Mem/n5593 , \Data_Mem/n5592 , \Data_Mem/n5591 ,
         \Data_Mem/n5590 , \Data_Mem/n5589 , \Data_Mem/n5588 ,
         \Data_Mem/n5587 , \Data_Mem/n5586 , \Data_Mem/n5585 ,
         \Data_Mem/n5584 , \Data_Mem/n5583 , \Data_Mem/n5582 ,
         \Data_Mem/n5581 , \Data_Mem/n5580 , \Data_Mem/n5579 ,
         \Data_Mem/n5578 , \Data_Mem/n5577 , \Data_Mem/n5576 ,
         \Data_Mem/n5575 , \Data_Mem/n5574 , \Data_Mem/n5573 ,
         \Data_Mem/n5572 , \Data_Mem/n5571 , \Data_Mem/n5570 ,
         \Data_Mem/n5569 , \Data_Mem/n5568 , \Data_Mem/n5567 ,
         \Data_Mem/n5566 , \Data_Mem/n5565 , \Data_Mem/n5564 ,
         \Data_Mem/n5563 , \Data_Mem/n5562 , \Data_Mem/n5561 ,
         \Data_Mem/n5560 , \Data_Mem/n5559 , \Data_Mem/n5558 ,
         \Data_Mem/n5557 , \Data_Mem/n5556 , \Data_Mem/n5555 ,
         \Data_Mem/n5554 , \Data_Mem/n5553 , \Data_Mem/n5552 ,
         \Data_Mem/n5551 , \Data_Mem/n5550 , \Data_Mem/n5549 ,
         \Data_Mem/n5548 , \Data_Mem/n5547 , \Data_Mem/n5546 ,
         \Data_Mem/n5545 , \Data_Mem/n5544 , \Data_Mem/n5543 ,
         \Data_Mem/n5542 , \Data_Mem/n5541 , \Data_Mem/n5540 ,
         \Data_Mem/n5539 , \Data_Mem/n5538 , \Data_Mem/n5537 ,
         \Data_Mem/n5536 , \Data_Mem/n5535 , \Data_Mem/n5534 ,
         \Data_Mem/n5533 , \Data_Mem/n5532 , \Data_Mem/n5531 ,
         \Data_Mem/n5530 , \Data_Mem/n5529 , \Data_Mem/n5528 ,
         \Data_Mem/n5527 , \Data_Mem/n5526 , \Data_Mem/n5525 ,
         \Data_Mem/n5524 , \Data_Mem/n5523 , \Data_Mem/n5522 ,
         \Data_Mem/n5521 , \Data_Mem/n5520 , \Data_Mem/n5519 ,
         \Data_Mem/n5518 , \Data_Mem/n5517 , \Data_Mem/n5516 ,
         \Data_Mem/n5515 , \Data_Mem/n5514 , \Data_Mem/n5513 ,
         \Data_Mem/n5512 , \Data_Mem/n5511 , \Data_Mem/n5510 ,
         \Data_Mem/n5509 , \Data_Mem/n5508 , \Data_Mem/n5507 ,
         \Data_Mem/n5506 , \Data_Mem/n5505 , \Data_Mem/n5504 ,
         \Data_Mem/n5503 , \Data_Mem/n5502 , \Data_Mem/n5501 ,
         \Data_Mem/n5500 , \Data_Mem/n5499 , \Data_Mem/n5498 ,
         \Data_Mem/n5497 , \Data_Mem/n5496 , \Data_Mem/n5495 ,
         \Data_Mem/n5494 , \Data_Mem/n5493 , \Data_Mem/n5492 ,
         \Data_Mem/n5491 , \Data_Mem/n5490 , \Data_Mem/n5489 ,
         \Data_Mem/n5488 , \Data_Mem/n5487 , \Data_Mem/n5486 ,
         \Data_Mem/n5485 , \Data_Mem/n5484 , \Data_Mem/n5483 ,
         \Data_Mem/n5482 , \Data_Mem/n5481 , \Data_Mem/n5480 ,
         \Data_Mem/n5479 , \Data_Mem/n5478 , \Data_Mem/n5477 ,
         \Data_Mem/n5476 , \Data_Mem/n5475 , \Data_Mem/n5474 ,
         \Data_Mem/n5473 , \Data_Mem/n5472 , \Data_Mem/n5471 ,
         \Data_Mem/n5470 , \Data_Mem/n5469 , \Data_Mem/n5468 ,
         \Data_Mem/n5467 , \Data_Mem/n5466 , \Data_Mem/n5465 ,
         \Data_Mem/n5464 , \Data_Mem/n5463 , \Data_Mem/n5462 ,
         \Data_Mem/n5461 , \Data_Mem/n5460 , \Data_Mem/n5459 ,
         \Data_Mem/n5458 , \Data_Mem/n5457 , \Data_Mem/n5456 ,
         \Data_Mem/n5455 , \Data_Mem/n5454 , \Data_Mem/n5453 ,
         \Data_Mem/n5452 , \Data_Mem/n5451 , \Data_Mem/n5450 ,
         \Data_Mem/n5449 , \Data_Mem/n5448 , \Data_Mem/n5447 ,
         \Data_Mem/n5446 , \Data_Mem/n5445 , \Data_Mem/n5444 ,
         \Data_Mem/n5443 , \Data_Mem/n5442 , \Data_Mem/n5441 ,
         \Data_Mem/n5440 , \Data_Mem/n5439 , \Data_Mem/n5438 ,
         \Data_Mem/n5437 , \Data_Mem/n5436 , \Data_Mem/n5435 ,
         \Data_Mem/n5434 , \Data_Mem/n5433 , \Data_Mem/n5432 ,
         \Data_Mem/n5431 , \Data_Mem/n5430 , \Data_Mem/n5429 ,
         \Data_Mem/n5428 , \Data_Mem/n5427 , \Data_Mem/n5426 ,
         \Data_Mem/n5425 , \Data_Mem/n5424 , \Data_Mem/n5423 ,
         \Data_Mem/n5422 , \Data_Mem/n5421 , \Data_Mem/n5420 ,
         \Data_Mem/n5419 , \Data_Mem/n5418 , \Data_Mem/n5417 ,
         \Data_Mem/n5416 , \Data_Mem/n5415 , \Data_Mem/n5414 ,
         \Data_Mem/n5413 , \Data_Mem/n5412 , \Data_Mem/n5411 ,
         \Data_Mem/n5410 , \Data_Mem/n5409 , \Data_Mem/n5408 ,
         \Data_Mem/n5407 , \Data_Mem/n5406 , \Data_Mem/n5405 ,
         \Data_Mem/n5404 , \Data_Mem/n5403 , \Data_Mem/n5402 ,
         \Data_Mem/n5401 , \Data_Mem/n5400 , \Data_Mem/n5399 ,
         \Data_Mem/n5398 , \Data_Mem/n5397 , \Data_Mem/n5396 ,
         \Data_Mem/n5395 , \Data_Mem/n5394 , \Data_Mem/n5393 ,
         \Data_Mem/n5392 , \Data_Mem/n5391 , \Data_Mem/n5390 ,
         \Data_Mem/n5389 , \Data_Mem/n5388 , \Data_Mem/n5387 ,
         \Data_Mem/n5386 , \Data_Mem/n5385 , \Data_Mem/n5384 ,
         \Data_Mem/n5383 , \Data_Mem/n5382 , \Data_Mem/n5381 ,
         \Data_Mem/n5380 , \Data_Mem/n5379 , \Data_Mem/n5378 ,
         \Data_Mem/n5377 , \Data_Mem/n5376 , \Data_Mem/n5375 ,
         \Data_Mem/n5374 , \Data_Mem/n5373 , \Data_Mem/n5372 ,
         \Data_Mem/n5371 , \Data_Mem/n5370 , \Data_Mem/n5369 ,
         \Data_Mem/n5368 , \Data_Mem/n5367 , \Data_Mem/n5366 ,
         \Data_Mem/n5365 , \Data_Mem/n5364 , \Data_Mem/n5363 ,
         \Data_Mem/n5362 , \Data_Mem/n5361 , \Data_Mem/n5360 ,
         \Data_Mem/n5359 , \Data_Mem/n5358 , \Data_Mem/n5357 ,
         \Data_Mem/n5356 , \Data_Mem/n5355 , \Data_Mem/n5354 ,
         \Data_Mem/n5353 , \Data_Mem/n5352 , \Data_Mem/n5351 ,
         \Data_Mem/n5350 , \Data_Mem/n5349 , \Data_Mem/n5348 ,
         \Data_Mem/n5347 , \Data_Mem/n5346 , \Data_Mem/n5345 ,
         \Data_Mem/n5344 , \Data_Mem/n5343 , \Data_Mem/n5342 ,
         \Data_Mem/n5341 , \Data_Mem/n5340 , \Data_Mem/n5339 ,
         \Data_Mem/n5338 , \Data_Mem/n5337 , \Data_Mem/n5336 ,
         \Data_Mem/n5335 , \Data_Mem/n5334 , \Data_Mem/n5333 ,
         \Data_Mem/n5332 , \Data_Mem/n5331 , \Data_Mem/n5330 ,
         \Data_Mem/n5329 , \Data_Mem/n5328 , \Data_Mem/n5327 ,
         \Data_Mem/n5326 , \Data_Mem/n5325 , \Data_Mem/n5324 ,
         \Data_Mem/n5323 , \Data_Mem/n5322 , \Data_Mem/n5321 ,
         \Data_Mem/n5320 , \Data_Mem/n5319 , \Data_Mem/n5318 ,
         \Data_Mem/n5317 , \Data_Mem/n5316 , \Data_Mem/n5315 ,
         \Data_Mem/n5314 , \Data_Mem/n5313 , \Data_Mem/n5312 ,
         \Data_Mem/n5311 , \Data_Mem/n5310 , \Data_Mem/n5309 ,
         \Data_Mem/n5308 , \Data_Mem/n5307 , \Data_Mem/n5306 ,
         \Data_Mem/n5305 , \Data_Mem/n5304 , \Data_Mem/n5303 ,
         \Data_Mem/n5302 , \Data_Mem/n5301 , \Data_Mem/n5300 ,
         \Data_Mem/n5299 , \Data_Mem/n5298 , \Data_Mem/n5297 ,
         \Data_Mem/n5296 , \Data_Mem/n5295 , \Data_Mem/n5294 ,
         \Data_Mem/n5293 , \Data_Mem/n5292 , \Data_Mem/n5291 ,
         \Data_Mem/n5290 , \Data_Mem/n5289 , \Data_Mem/n5288 ,
         \Data_Mem/n5287 , \Data_Mem/n5286 , \Data_Mem/n5285 ,
         \Data_Mem/n5284 , \Data_Mem/n5283 , \Data_Mem/n5282 ,
         \Data_Mem/n5281 , \Data_Mem/n5280 , \Data_Mem/n5279 ,
         \Data_Mem/n5278 , \Data_Mem/n5277 , \Data_Mem/n5276 ,
         \Data_Mem/n5275 , \Data_Mem/n5274 , \Data_Mem/n5273 ,
         \Data_Mem/n5272 , \Data_Mem/n5271 , \Data_Mem/n5270 ,
         \Data_Mem/n5269 , \Data_Mem/n5268 , \Data_Mem/n5267 ,
         \Data_Mem/n5266 , \Data_Mem/n5265 , \Data_Mem/n5264 ,
         \Data_Mem/n5263 , \Data_Mem/n5262 , \Data_Mem/n5261 ,
         \Data_Mem/n5260 , \Data_Mem/n5259 , \Data_Mem/n5258 ,
         \Data_Mem/n5257 , \Data_Mem/n5256 , \Data_Mem/n5255 ,
         \Data_Mem/n5254 , \Data_Mem/n5253 , \Data_Mem/n5252 ,
         \Data_Mem/n5251 , \Data_Mem/n5250 , \Data_Mem/n5249 ,
         \Data_Mem/n5248 , \Data_Mem/n5247 , \Data_Mem/n5246 ,
         \Data_Mem/n5245 , \Data_Mem/n5244 , \Data_Mem/n5243 ,
         \Data_Mem/n5242 , \Data_Mem/n5241 , \Data_Mem/n5240 ,
         \Data_Mem/n5239 , \Data_Mem/n5238 , \Data_Mem/n5237 ,
         \Data_Mem/n5236 , \Data_Mem/n5235 , \Data_Mem/n5234 ,
         \Data_Mem/n5233 , \Data_Mem/n5232 , \Data_Mem/n5231 ,
         \Data_Mem/n5230 , \Data_Mem/n5229 , \Data_Mem/n5228 ,
         \Data_Mem/n5227 , \Data_Mem/n5226 , \Data_Mem/n5225 ,
         \Data_Mem/n5224 , \Data_Mem/n5223 , \Data_Mem/n5222 ,
         \Data_Mem/n5221 , \Data_Mem/n5220 , \Data_Mem/n5219 ,
         \Data_Mem/n5218 , \Data_Mem/n5217 , \Data_Mem/n5216 ,
         \Data_Mem/n5215 , \Data_Mem/n5214 , \Data_Mem/n5213 ,
         \Data_Mem/n5212 , \Data_Mem/n5211 , \Data_Mem/n5210 ,
         \Data_Mem/n5209 , \Data_Mem/n5208 , \Data_Mem/n5207 ,
         \Data_Mem/n5206 , \Data_Mem/n5205 , \Data_Mem/n5204 ,
         \Data_Mem/n5203 , \Data_Mem/n5202 , \Data_Mem/n5201 ,
         \Data_Mem/n5200 , \Data_Mem/n5199 , \Data_Mem/n5198 ,
         \Data_Mem/n5197 , \Data_Mem/n5196 , \Data_Mem/n5195 ,
         \Data_Mem/n5194 , \Data_Mem/n5193 , \Data_Mem/n5192 ,
         \Data_Mem/n5191 , \Data_Mem/n5190 , \Data_Mem/n5189 ,
         \Data_Mem/n5188 , \Data_Mem/n5187 , \Data_Mem/n5186 ,
         \Data_Mem/n5185 , \Data_Mem/n5184 , \Data_Mem/n5183 ,
         \Data_Mem/n5182 , \Data_Mem/n5181 , \Data_Mem/n5180 ,
         \Data_Mem/n5179 , \Data_Mem/n5178 , \Data_Mem/n5177 ,
         \Data_Mem/n5176 , \Data_Mem/n5175 , \Data_Mem/n5174 ,
         \Data_Mem/n5173 , \Data_Mem/n5172 , \Data_Mem/n5171 ,
         \Data_Mem/n5170 , \Data_Mem/n5169 , \Data_Mem/n5168 ,
         \Data_Mem/n5167 , \Data_Mem/n5166 , \Data_Mem/n5165 ,
         \Data_Mem/n5164 , \Data_Mem/n5163 , \Data_Mem/n5162 ,
         \Data_Mem/n5161 , \Data_Mem/n5160 , \Data_Mem/n5159 ,
         \Data_Mem/n5158 , \Data_Mem/n5157 , \Data_Mem/n5156 ,
         \Data_Mem/n5155 , \Data_Mem/n5154 , \Data_Mem/n5153 ,
         \Data_Mem/n5152 , \Data_Mem/n5151 , \Data_Mem/n5150 ,
         \Data_Mem/n5149 , \Data_Mem/n5148 , \Data_Mem/n5147 ,
         \Data_Mem/n5146 , \Data_Mem/n5145 , \Data_Mem/n5144 ,
         \Data_Mem/n5143 , \Data_Mem/n5142 , \Data_Mem/n5141 ,
         \Data_Mem/n5140 , \Data_Mem/n5139 , \Data_Mem/n5138 ,
         \Data_Mem/n5137 , \Data_Mem/n5136 , \Data_Mem/n5135 ,
         \Data_Mem/n5134 , \Data_Mem/n5133 , \Data_Mem/n5132 ,
         \Data_Mem/n5131 , \Data_Mem/n5130 , \Data_Mem/n5129 ,
         \Data_Mem/n5128 , \Data_Mem/n5127 , \Data_Mem/n5126 ,
         \Data_Mem/n5125 , \Data_Mem/n5124 , \Data_Mem/n5123 ,
         \Data_Mem/n5122 , \Data_Mem/n5121 , \Data_Mem/n5120 ,
         \Data_Mem/n5119 , \Data_Mem/n5118 , \Data_Mem/n5117 ,
         \Data_Mem/n5116 , \Data_Mem/n5115 , \Data_Mem/n5114 ,
         \Data_Mem/n5113 , \Data_Mem/n5112 , \Data_Mem/n5111 ,
         \Data_Mem/n5110 , \Data_Mem/n5109 , \Data_Mem/n5108 ,
         \Data_Mem/n5107 , \Data_Mem/n5106 , \Data_Mem/n5105 ,
         \Data_Mem/n5104 , \Data_Mem/n5103 , \Data_Mem/n5102 ,
         \Data_Mem/n5101 , \Data_Mem/n5100 , \Data_Mem/n5099 ,
         \Data_Mem/n5098 , \Data_Mem/n5097 , \Data_Mem/n5096 ,
         \Data_Mem/n5095 , \Data_Mem/n5094 , \Data_Mem/n5093 ,
         \Data_Mem/n5092 , \Data_Mem/n5091 , \Data_Mem/n5090 ,
         \Data_Mem/n5089 , \Data_Mem/n5088 , \Data_Mem/n5087 ,
         \Data_Mem/n5086 , \Data_Mem/n5085 , \Data_Mem/n5084 ,
         \Data_Mem/n5083 , \Data_Mem/n5082 , \Data_Mem/n5081 ,
         \Data_Mem/n5080 , \Data_Mem/n5079 , \Data_Mem/n5078 ,
         \Data_Mem/n5077 , \Data_Mem/n5076 , \Data_Mem/n5075 ,
         \Data_Mem/n5074 , \Data_Mem/n5073 , \Data_Mem/n5072 ,
         \Data_Mem/n5071 , \Data_Mem/n5070 , \Data_Mem/n5069 ,
         \Data_Mem/n5068 , \Data_Mem/n5067 , \Data_Mem/n5066 ,
         \Data_Mem/n5065 , \Data_Mem/n5064 , \Data_Mem/n5063 ,
         \Data_Mem/n5062 , \Data_Mem/n5061 , \Data_Mem/n5060 ,
         \Data_Mem/n5059 , \Data_Mem/n5058 , \Data_Mem/n5057 ,
         \Data_Mem/n5056 , \Data_Mem/n5055 , \Data_Mem/n5054 ,
         \Data_Mem/n5053 , \Data_Mem/n5052 , \Data_Mem/n5051 ,
         \Data_Mem/n5050 , \Data_Mem/n5049 , \Data_Mem/n5048 ,
         \Data_Mem/n5047 , \Data_Mem/n5046 , \Data_Mem/n5045 ,
         \Data_Mem/n5044 , \Data_Mem/n5043 , \Data_Mem/n5042 ,
         \Data_Mem/n5041 , \Data_Mem/n5040 , \Data_Mem/n5039 ,
         \Data_Mem/n5038 , \Data_Mem/n5037 , \Data_Mem/n5036 ,
         \Data_Mem/n5035 , \Data_Mem/n5034 , \Data_Mem/n5033 ,
         \Data_Mem/n5032 , \Data_Mem/n5031 , \Data_Mem/n5030 ,
         \Data_Mem/n5029 , \Data_Mem/n5028 , \Data_Mem/n5027 ,
         \Data_Mem/n5026 , \Data_Mem/n5025 , \Data_Mem/n5024 ,
         \Data_Mem/n5023 , \Data_Mem/n5022 , \Data_Mem/n5021 ,
         \Data_Mem/n5020 , \Data_Mem/n5019 , \Data_Mem/n5018 ,
         \Data_Mem/n5017 , \Data_Mem/n5016 , \Data_Mem/n5015 ,
         \Data_Mem/n5014 , \Data_Mem/n5013 , \Data_Mem/n5012 ,
         \Data_Mem/n5011 , \Data_Mem/n5010 , \Data_Mem/n5009 ,
         \Data_Mem/n5008 , \Data_Mem/n5007 , \Data_Mem/n5006 ,
         \Data_Mem/n5005 , \Data_Mem/n5004 , \Data_Mem/n5003 ,
         \Data_Mem/n5002 , \Data_Mem/n5001 , \Data_Mem/n5000 ,
         \Data_Mem/n4999 , \Data_Mem/n4998 , \Data_Mem/n4997 ,
         \Data_Mem/n4996 , \Data_Mem/n4995 , \Data_Mem/n4994 ,
         \Data_Mem/n4993 , \Data_Mem/n4992 , \Data_Mem/n4991 ,
         \Data_Mem/n4990 , \Data_Mem/n4989 , \Data_Mem/n4988 ,
         \Data_Mem/n4987 , \Data_Mem/n4986 , \Data_Mem/n4985 ,
         \Data_Mem/n4984 , \Data_Mem/n4983 , \Data_Mem/n4982 ,
         \Data_Mem/n4981 , \Data_Mem/n4980 , \Data_Mem/n4979 ,
         \Data_Mem/n4978 , \Data_Mem/n4977 , \Data_Mem/n4976 ,
         \Data_Mem/n4975 , \Data_Mem/n4974 , \Data_Mem/n4973 ,
         \Data_Mem/n4972 , \Data_Mem/n4971 , \Data_Mem/n4970 ,
         \Data_Mem/n4969 , \Data_Mem/n4968 , \Data_Mem/n4967 ,
         \Data_Mem/n4966 , \Data_Mem/n4965 , \Data_Mem/n4964 ,
         \Data_Mem/n4963 , \Data_Mem/n4962 , \Data_Mem/n4961 ,
         \Data_Mem/n4960 , \Data_Mem/n4959 , \Data_Mem/n4958 ,
         \Data_Mem/n4957 , \Data_Mem/n4956 , \Data_Mem/n4955 ,
         \Data_Mem/n4954 , \Data_Mem/n4953 , \Data_Mem/n4952 ,
         \Data_Mem/n4951 , \Data_Mem/n4950 , \Data_Mem/n4949 ,
         \Data_Mem/n4948 , \Data_Mem/n4947 , \Data_Mem/n4946 ,
         \Data_Mem/n4945 , \Data_Mem/n4944 , \Data_Mem/n4943 ,
         \Data_Mem/n4942 , \Data_Mem/n4941 , \Data_Mem/n4940 ,
         \Data_Mem/n4939 , \Data_Mem/n4938 , \Data_Mem/n4937 ,
         \Data_Mem/n4936 , \Data_Mem/n4935 , \Data_Mem/n4934 ,
         \Data_Mem/n4933 , \Data_Mem/n4932 , \Data_Mem/n4931 ,
         \Data_Mem/n4930 , \Data_Mem/n4929 , \Data_Mem/n4928 ,
         \Data_Mem/n4927 , \Data_Mem/n4926 , \Data_Mem/n4925 ,
         \Data_Mem/n4924 , \Data_Mem/n4923 , \Data_Mem/n4922 ,
         \Data_Mem/n4921 , \Data_Mem/n4920 , \Data_Mem/n4919 ,
         \Data_Mem/n4918 , \Data_Mem/n4917 , \Data_Mem/n4916 ,
         \Data_Mem/n4915 , \Data_Mem/n4914 , \Data_Mem/n4913 ,
         \Data_Mem/n4912 , \Data_Mem/n4911 , \Data_Mem/n4910 ,
         \Data_Mem/n4909 , \Data_Mem/n4908 , \Data_Mem/n4907 ,
         \Data_Mem/n4906 , \Data_Mem/n4905 , \Data_Mem/n4904 ,
         \Data_Mem/n4903 , \Data_Mem/n4902 , \Data_Mem/n4901 ,
         \Data_Mem/n4900 , \Data_Mem/n4899 , \Data_Mem/n4898 ,
         \Data_Mem/n4897 , \Data_Mem/n4896 , \Data_Mem/n4895 ,
         \Data_Mem/n4894 , \Data_Mem/n4893 , \Data_Mem/n4892 ,
         \Data_Mem/n4891 , \Data_Mem/n4890 , \Data_Mem/n4889 ,
         \Data_Mem/n4888 , \Data_Mem/n4887 , \Data_Mem/n4886 ,
         \Data_Mem/n4885 , \Data_Mem/n4884 , \Data_Mem/n4883 ,
         \Data_Mem/n4882 , \Data_Mem/n4881 , \Data_Mem/n4880 ,
         \Data_Mem/n4879 , \Data_Mem/n4878 , \Data_Mem/n4877 ,
         \Data_Mem/n4876 , \Data_Mem/n4875 , \Data_Mem/n4874 ,
         \Data_Mem/n4873 , \Data_Mem/n4872 , \Data_Mem/n4871 ,
         \Data_Mem/n4870 , \Data_Mem/n4869 , \Data_Mem/n4868 ,
         \Data_Mem/n4867 , \Data_Mem/n4866 , \Data_Mem/n4865 ,
         \Data_Mem/n4864 , \Data_Mem/n4863 , \Data_Mem/n4862 ,
         \Data_Mem/n4861 , \Data_Mem/n4860 , \Data_Mem/n4859 ,
         \Data_Mem/n4858 , \Data_Mem/n4857 , \Data_Mem/n4856 ,
         \Data_Mem/n4855 , \Data_Mem/n4854 , \Data_Mem/n4853 ,
         \Data_Mem/n4852 , \Data_Mem/n4851 , \Data_Mem/n4850 ,
         \Data_Mem/n4849 , \Data_Mem/n4848 , \Data_Mem/n4847 ,
         \Data_Mem/n4846 , \Data_Mem/n4845 , \Data_Mem/n4844 ,
         \Data_Mem/n4843 , \Data_Mem/n4842 , \Data_Mem/n4841 ,
         \Data_Mem/n4840 , \Data_Mem/n4839 , \Data_Mem/n4838 ,
         \Data_Mem/n4837 , \Data_Mem/n4836 , \Data_Mem/n4835 ,
         \Data_Mem/n4834 , \Data_Mem/n4833 , \Data_Mem/n4832 ,
         \Data_Mem/n4831 , \Data_Mem/n4830 , \Data_Mem/n4829 ,
         \Data_Mem/n4828 , \Data_Mem/n4827 , \Data_Mem/n4826 ,
         \Data_Mem/n4825 , \Data_Mem/n4824 , \Data_Mem/n4823 ,
         \Data_Mem/n4822 , \Data_Mem/n4821 , \Data_Mem/n4820 ,
         \Data_Mem/n4819 , \Data_Mem/n4818 , \Data_Mem/n4817 ,
         \Data_Mem/n4816 , \Data_Mem/n4815 , \Data_Mem/n4814 ,
         \Data_Mem/n4813 , \Data_Mem/n4812 , \Data_Mem/n4811 ,
         \Data_Mem/n4810 , \Data_Mem/n4809 , \Data_Mem/n4808 ,
         \Data_Mem/n4807 , \Data_Mem/n4806 , \Data_Mem/n4805 ,
         \Data_Mem/n4804 , \Data_Mem/n4803 , \Data_Mem/n4802 ,
         \Data_Mem/n4801 , \Data_Mem/n4800 , \Data_Mem/n4799 ,
         \Data_Mem/n4798 , \Data_Mem/n4797 , \Data_Mem/n4796 ,
         \Data_Mem/n4795 , \Data_Mem/n4794 , \Data_Mem/n4793 ,
         \Data_Mem/n4792 , \Data_Mem/n4791 , \Data_Mem/n4790 ,
         \Data_Mem/n4789 , \Data_Mem/n4788 , \Data_Mem/n4787 ,
         \Data_Mem/n4786 , \Data_Mem/n4785 , \Data_Mem/n4784 ,
         \Data_Mem/n4783 , \Data_Mem/n4782 , \Data_Mem/n4781 ,
         \Data_Mem/n4780 , \Data_Mem/n4779 , \Data_Mem/n4778 ,
         \Data_Mem/n4777 , \Data_Mem/n4776 , \Data_Mem/n4775 ,
         \Data_Mem/n4774 , \Data_Mem/n4773 , \Data_Mem/n4772 ,
         \Data_Mem/n4771 , \Data_Mem/n4770 , \Data_Mem/n4769 ,
         \Data_Mem/n4768 , \Data_Mem/n4767 , \Data_Mem/n4766 ,
         \Data_Mem/n4765 , \Data_Mem/n4764 , \Data_Mem/n4763 ,
         \Data_Mem/n4762 , \Data_Mem/n4761 , \Data_Mem/n4760 ,
         \Data_Mem/n4759 , \Data_Mem/n4758 , \Data_Mem/n4757 ,
         \Data_Mem/n4756 , \Data_Mem/n4755 , \Data_Mem/n4754 ,
         \Data_Mem/n4753 , \Data_Mem/n4752 , \Data_Mem/n4751 ,
         \Data_Mem/n4750 , \Data_Mem/n4749 , \Data_Mem/n4748 ,
         \Data_Mem/n4747 , \Data_Mem/n4746 , \Data_Mem/n4745 ,
         \Data_Mem/n4744 , \Data_Mem/n4743 , \Data_Mem/n4742 ,
         \Data_Mem/n4741 , \Data_Mem/n4740 , \Data_Mem/n4739 ,
         \Data_Mem/n4738 , \Data_Mem/n4737 , \Data_Mem/n4736 ,
         \Data_Mem/n4735 , \Data_Mem/n4734 , \Data_Mem/n4733 ,
         \Data_Mem/n4732 , \Data_Mem/n4731 , \Data_Mem/n4730 ,
         \Data_Mem/n4729 , \Data_Mem/n4728 , \Data_Mem/n4727 ,
         \Data_Mem/n4726 , \Data_Mem/n4725 , \Data_Mem/n4724 ,
         \Data_Mem/n4723 , \Data_Mem/n4722 , \Data_Mem/n4721 ,
         \Data_Mem/n4720 , \Data_Mem/n4719 , \Data_Mem/n4718 ,
         \Data_Mem/n4717 , \Data_Mem/n4716 , \Data_Mem/n4715 ,
         \Data_Mem/n4714 , \Data_Mem/n4713 , \Data_Mem/n4712 ,
         \Data_Mem/n4711 , \Data_Mem/n4710 , \Data_Mem/n4709 ,
         \Data_Mem/n4708 , \Data_Mem/n4707 , \Data_Mem/n4706 ,
         \Data_Mem/n4705 , \Data_Mem/n4704 , \Data_Mem/n4703 ,
         \Data_Mem/n4702 , \Data_Mem/n4701 , \Data_Mem/n4700 ,
         \Data_Mem/n4699 , \Data_Mem/n4698 , \Data_Mem/n4697 ,
         \Data_Mem/n4696 , \Data_Mem/n4695 , \Data_Mem/n4694 ,
         \Data_Mem/n4693 , \Data_Mem/n4692 , \Data_Mem/n4691 ,
         \Data_Mem/n4690 , \Data_Mem/n4689 , \Data_Mem/n4688 ,
         \Data_Mem/n4687 , \Data_Mem/n4686 , \Data_Mem/n4685 ,
         \Data_Mem/n4684 , \Data_Mem/n4683 , \Data_Mem/n4682 ,
         \Data_Mem/n4681 , \Data_Mem/n4680 , \Data_Mem/n4679 ,
         \Data_Mem/n4678 , \Data_Mem/n4677 , \Data_Mem/n4676 ,
         \Data_Mem/n4675 , \Data_Mem/n4674 , \Data_Mem/n4673 ,
         \Data_Mem/n4672 , \Data_Mem/n4671 , \Data_Mem/n4670 ,
         \Data_Mem/n4669 , \Data_Mem/n4668 , \Data_Mem/n4667 ,
         \Data_Mem/n4666 , \Data_Mem/n4665 , \Data_Mem/n4664 ,
         \Data_Mem/n4663 , \Data_Mem/n4662 , \Data_Mem/n4661 ,
         \Data_Mem/n4660 , \Data_Mem/n4659 , \Data_Mem/n4658 ,
         \Data_Mem/n4657 , \Data_Mem/n4656 , \Data_Mem/n4655 ,
         \Data_Mem/n4654 , \Data_Mem/n4653 , \Data_Mem/n4652 ,
         \Data_Mem/n4651 , \Data_Mem/n4650 , \Data_Mem/n4649 ,
         \Data_Mem/n4648 , \Data_Mem/n4647 , \Data_Mem/n4646 ,
         \Data_Mem/n4645 , \Data_Mem/n4644 , \Data_Mem/n4643 ,
         \Data_Mem/n4642 , \Data_Mem/n4641 , \Data_Mem/n4640 ,
         \Data_Mem/n4639 , \Data_Mem/n4638 , \Data_Mem/n4637 ,
         \Data_Mem/n4636 , \Data_Mem/n4635 , \Data_Mem/n4634 ,
         \Data_Mem/n4633 , \Data_Mem/n4632 , \Data_Mem/n4631 ,
         \Data_Mem/n4630 , \Data_Mem/n4629 , \Data_Mem/n4628 ,
         \Data_Mem/n4627 , \Data_Mem/n4626 , \Data_Mem/n4625 ,
         \Data_Mem/n4624 , \Data_Mem/n4623 , \Data_Mem/n4622 ,
         \Data_Mem/n4621 , \Data_Mem/n4620 , \Data_Mem/n4619 ,
         \Data_Mem/n4618 , \Data_Mem/n4617 , \Data_Mem/n4616 ,
         \Data_Mem/n4615 , \Data_Mem/n4614 , \Data_Mem/n4613 ,
         \Data_Mem/n4612 , \Data_Mem/n4611 , \Data_Mem/n4610 ,
         \Data_Mem/n4609 , \Data_Mem/n4608 , \Data_Mem/n4607 ,
         \Data_Mem/n4606 , \Data_Mem/n4605 , \Data_Mem/n4604 ,
         \Data_Mem/n4603 , \Data_Mem/n4602 , \Data_Mem/n4601 ,
         \Data_Mem/n4600 , \Data_Mem/n4599 , \Data_Mem/n4598 ,
         \Data_Mem/n4597 , \Data_Mem/n4596 , \Data_Mem/n4595 ,
         \Data_Mem/n4594 , \Data_Mem/n4593 , \Data_Mem/n4592 ,
         \Data_Mem/n4591 , \Data_Mem/n4590 , \Data_Mem/n4589 ,
         \Data_Mem/n4588 , \Data_Mem/n4587 , \Data_Mem/n4586 ,
         \Data_Mem/n4585 , \Data_Mem/n4584 , \Data_Mem/n4583 ,
         \Data_Mem/n4582 , \Data_Mem/n4581 , \Data_Mem/n4580 ,
         \Data_Mem/n4579 , \Data_Mem/n4578 , \Data_Mem/n4577 ,
         \Data_Mem/n4576 , \Data_Mem/n4575 , \Data_Mem/n4574 ,
         \Data_Mem/n4573 , \Data_Mem/n4572 , \Data_Mem/n4571 ,
         \Data_Mem/n4570 , \Data_Mem/n4569 , \Data_Mem/n4568 ,
         \Data_Mem/n4567 , \Data_Mem/n4566 , \Data_Mem/n4565 ,
         \Data_Mem/n4564 , \Data_Mem/n4563 , \Data_Mem/n4562 ,
         \Data_Mem/n4561 , \Data_Mem/n4560 , \Data_Mem/n4559 ,
         \Data_Mem/n4558 , \Data_Mem/n4557 , \Data_Mem/n4556 ,
         \Data_Mem/n4555 , \Data_Mem/n4554 , \Data_Mem/n4553 ,
         \Data_Mem/n4552 , \Data_Mem/n4551 , \Data_Mem/n4550 ,
         \Data_Mem/n4549 , \Data_Mem/n4548 , \Data_Mem/n4547 ,
         \Data_Mem/n4546 , \Data_Mem/n4545 , \Data_Mem/n4544 ,
         \Data_Mem/n4543 , \Data_Mem/n4542 , \Data_Mem/n4541 ,
         \Data_Mem/n4540 , \Data_Mem/n4539 , \Data_Mem/n4538 ,
         \Data_Mem/n4537 , \Data_Mem/n4536 , \Data_Mem/n4535 ,
         \Data_Mem/n4534 , \Data_Mem/n4533 , \Data_Mem/n4532 ,
         \Data_Mem/n4531 , \Data_Mem/n4530 , \Data_Mem/n4529 ,
         \Data_Mem/n4528 , \Data_Mem/n4527 , \Data_Mem/n4526 ,
         \Data_Mem/n4525 , \Data_Mem/n4524 , \Data_Mem/n4523 ,
         \Data_Mem/n4522 , \Data_Mem/n4521 , \Data_Mem/n4520 ,
         \Data_Mem/n4519 , \Data_Mem/n4518 , \Data_Mem/n4517 ,
         \Data_Mem/n4516 , \Data_Mem/n4515 , \Data_Mem/n4514 ,
         \Data_Mem/n4513 , \Data_Mem/n4512 , \Data_Mem/n4511 ,
         \Data_Mem/n4510 , \Data_Mem/n4509 , \Data_Mem/n4508 ,
         \Data_Mem/n4507 , \Data_Mem/n4506 , \Data_Mem/n4505 ,
         \Data_Mem/n4504 , \Data_Mem/n4503 , \Data_Mem/n4502 ,
         \Data_Mem/n4501 , \Data_Mem/n4500 , \Data_Mem/n4499 ,
         \Data_Mem/n4498 , \Data_Mem/n4497 , \Data_Mem/n4496 ,
         \Data_Mem/n4495 , \Data_Mem/n4494 , \Data_Mem/n4493 ,
         \Data_Mem/n4492 , \Data_Mem/n4491 , \Data_Mem/n4490 ,
         \Data_Mem/n4489 , \Data_Mem/n4488 , \Data_Mem/n4487 ,
         \Data_Mem/n4486 , \Data_Mem/n4485 , \Data_Mem/n4484 ,
         \Data_Mem/n4483 , \Data_Mem/n4482 , \Data_Mem/n4481 ,
         \Data_Mem/n4480 , \Data_Mem/n4479 , \Data_Mem/n4478 ,
         \Data_Mem/n4477 , \Data_Mem/n4476 , \Data_Mem/n4475 ,
         \Data_Mem/n4474 , \Data_Mem/n4473 , \Data_Mem/n4472 ,
         \Data_Mem/n4471 , \Data_Mem/n4470 , \Data_Mem/n4469 ,
         \Data_Mem/n4468 , \Data_Mem/n4467 , \Data_Mem/n4466 ,
         \Data_Mem/n4465 , \Data_Mem/n4464 , \Data_Mem/n4463 ,
         \Data_Mem/n4462 , \Data_Mem/n4461 , \Data_Mem/n4460 ,
         \Data_Mem/n4459 , \Data_Mem/n4458 , \Data_Mem/n4457 ,
         \Data_Mem/n4456 , \Data_Mem/n4455 , \Data_Mem/n4454 ,
         \Data_Mem/n4453 , \Data_Mem/n4452 , \Data_Mem/n4451 ,
         \Data_Mem/n4450 , \Data_Mem/n4449 , \Data_Mem/n4448 ,
         \Data_Mem/n4447 , \Data_Mem/n4446 , \Data_Mem/n4445 ,
         \Data_Mem/n4444 , \Data_Mem/n4443 , \Data_Mem/n4442 ,
         \Data_Mem/n4441 , \Data_Mem/n4440 , \Data_Mem/n4439 ,
         \Data_Mem/n4438 , \Data_Mem/n4437 , \Data_Mem/n4436 ,
         \Data_Mem/n4435 , \Data_Mem/n4434 , \Data_Mem/n4433 ,
         \Data_Mem/n4432 , \Data_Mem/n4431 , \Data_Mem/n4430 ,
         \Data_Mem/n4429 , \Data_Mem/n4428 , \Data_Mem/n4427 ,
         \Data_Mem/n4426 , \Data_Mem/n4425 , \Data_Mem/n4424 ,
         \Data_Mem/n4423 , \Data_Mem/n4422 , \Data_Mem/n4421 ,
         \Data_Mem/n4420 , \Data_Mem/n4419 , \Data_Mem/n4418 ,
         \Data_Mem/n4417 , \Data_Mem/n4416 , \Data_Mem/n4415 ,
         \Data_Mem/n4414 , \Data_Mem/n4413 , \Data_Mem/n4412 ,
         \Data_Mem/n4411 , \Data_Mem/n4410 , \Data_Mem/n4409 ,
         \Data_Mem/n4408 , \Data_Mem/n4407 , \Data_Mem/n4406 ,
         \Data_Mem/n4405 , \Data_Mem/n4404 , \Data_Mem/n4403 ,
         \Data_Mem/n4402 , \Data_Mem/n4401 , \Data_Mem/n4400 ,
         \Data_Mem/n4399 , \Data_Mem/n4398 , \Data_Mem/n4397 ,
         \Data_Mem/n4396 , \Data_Mem/n4395 , \Data_Mem/n4394 ,
         \Data_Mem/n4393 , \Data_Mem/n4392 , \Data_Mem/n4391 ,
         \Data_Mem/n4390 , \Data_Mem/n4389 , \Data_Mem/n4388 ,
         \Data_Mem/n4387 , \Data_Mem/n4386 , \Data_Mem/n4385 ,
         \Data_Mem/n4384 , \Data_Mem/n4383 , \Data_Mem/n4382 ,
         \Data_Mem/n4381 , \Data_Mem/n4380 , \Data_Mem/n4379 ,
         \Data_Mem/n4378 , \Data_Mem/n4377 , \Data_Mem/n4376 ,
         \Data_Mem/n4375 , \Data_Mem/n4374 , \Data_Mem/n4373 ,
         \Data_Mem/n4372 , \Data_Mem/n4371 , \Data_Mem/n4370 ,
         \Data_Mem/n4369 , \Data_Mem/n4368 , \Data_Mem/n4367 ,
         \Data_Mem/n4366 , \Data_Mem/n4365 , \Data_Mem/n4364 ,
         \Data_Mem/n4363 , \Data_Mem/n4362 , \Data_Mem/n4361 ,
         \Data_Mem/n4360 , \Data_Mem/n4359 , \Data_Mem/n4358 ,
         \Data_Mem/n4357 , \Data_Mem/n4356 , \Data_Mem/n4355 ,
         \Data_Mem/n4354 , \Data_Mem/n4353 , \Data_Mem/n4352 ,
         \Data_Mem/n4351 , \Data_Mem/n4350 , \Data_Mem/n4349 ,
         \Data_Mem/n4348 , \Data_Mem/n4347 , \Data_Mem/n4346 ,
         \Data_Mem/n4345 , \Data_Mem/n4344 , \Data_Mem/n4343 ,
         \Data_Mem/n4342 , \Data_Mem/n4341 , \Data_Mem/n4340 ,
         \Data_Mem/n4339 , \Data_Mem/n4338 , \Data_Mem/n4337 ,
         \Data_Mem/n4336 , \Data_Mem/n4335 , \Data_Mem/n4334 ,
         \Data_Mem/n4333 , \Data_Mem/n4332 , \Data_Mem/n4331 ,
         \Data_Mem/n4330 , \Data_Mem/n4329 , \Data_Mem/n4328 ,
         \Data_Mem/n4327 , \Data_Mem/n4326 , \Data_Mem/n4325 ,
         \Data_Mem/n4324 , \Data_Mem/n4323 , \Data_Mem/n4322 ,
         \Data_Mem/n4321 , \Data_Mem/n4320 , \Data_Mem/n4319 ,
         \Data_Mem/n4318 , \Data_Mem/n4317 , \Data_Mem/n4316 ,
         \Data_Mem/n4315 , \Data_Mem/n4314 , \Data_Mem/n4313 ,
         \Data_Mem/n4312 , \Data_Mem/n4311 , \Data_Mem/n4310 ,
         \Data_Mem/n4309 , \Data_Mem/n4308 , \Data_Mem/n4307 ,
         \Data_Mem/n4306 , \Data_Mem/n4305 , \Data_Mem/n4304 ,
         \Data_Mem/n4303 , \Data_Mem/n4302 , \Data_Mem/n4301 ,
         \Data_Mem/n4300 , \Data_Mem/n4299 , \Data_Mem/n4298 ,
         \Data_Mem/n4297 , \Data_Mem/n4296 , \Data_Mem/n4295 ,
         \Data_Mem/n4294 , \Data_Mem/n4293 , \Data_Mem/n4292 ,
         \Data_Mem/n4291 , \Data_Mem/n4290 , \Data_Mem/n4289 ,
         \Data_Mem/n4288 , \Data_Mem/n4287 , \Data_Mem/n4286 ,
         \Data_Mem/n4285 , \Data_Mem/n4284 , \Data_Mem/n4283 ,
         \Data_Mem/n4282 , \Data_Mem/n4281 , \Data_Mem/n4280 ,
         \Data_Mem/n4279 , \Data_Mem/n4278 , \Data_Mem/n4277 ,
         \Data_Mem/n4276 , \Data_Mem/n4275 , \Data_Mem/n4274 ,
         \Data_Mem/n4273 , \Data_Mem/n4272 , \Data_Mem/n4271 ,
         \Data_Mem/n4270 , \Data_Mem/n4269 , \Data_Mem/n4268 ,
         \Data_Mem/n4267 , \Data_Mem/n4266 , \Data_Mem/n4265 ,
         \Data_Mem/n4264 , \Data_Mem/n4263 , \Data_Mem/n4262 ,
         \Data_Mem/n4261 , \Data_Mem/n4260 , \Data_Mem/n4259 ,
         \Data_Mem/n4258 , \Data_Mem/n4257 , \Data_Mem/n4256 ,
         \Data_Mem/n4255 , \Data_Mem/n4254 , \Data_Mem/n4253 ,
         \Data_Mem/n4252 , \Data_Mem/n4251 , \Data_Mem/n4250 ,
         \Data_Mem/n4249 , \Data_Mem/n4248 , \Data_Mem/n4247 ,
         \Data_Mem/n4246 , \Data_Mem/n4245 , \Data_Mem/n4244 ,
         \Data_Mem/n4243 , \Data_Mem/n4242 , \Data_Mem/n4241 ,
         \Data_Mem/n4240 , \Data_Mem/n4239 , \Data_Mem/n4238 ,
         \Data_Mem/n4237 , \Data_Mem/n4236 , \Data_Mem/n4235 ,
         \Data_Mem/n4234 , \Data_Mem/n4233 , \Data_Mem/n4232 ,
         \Data_Mem/n4231 , \Data_Mem/n4230 , \Data_Mem/n4229 ,
         \Data_Mem/n4228 , \Data_Mem/n4227 , \Data_Mem/n4226 ,
         \Data_Mem/n4225 , \Data_Mem/n4224 , \Data_Mem/n4223 ,
         \Data_Mem/n4222 , \Data_Mem/n4221 , \Data_Mem/n4220 ,
         \Data_Mem/n4219 , \Data_Mem/n4218 , \Data_Mem/n4217 ,
         \Data_Mem/n4216 , \Reg_Bank/n5941 , \Reg_Bank/n5940 ,
         \Reg_Bank/n5939 , \Reg_Bank/n5938 , \Reg_Bank/n5937 ,
         \Reg_Bank/n5936 , \Reg_Bank/n5935 , \Reg_Bank/n5934 ,
         \Reg_Bank/n5933 , \Reg_Bank/n5932 , \Reg_Bank/n5931 ,
         \Reg_Bank/n5930 , \Reg_Bank/n5929 , \Reg_Bank/n5928 ,
         \Reg_Bank/n5927 , \Reg_Bank/n5926 , \Reg_Bank/n5925 ,
         \Reg_Bank/n5924 , \Reg_Bank/n5923 , \Reg_Bank/n5922 ,
         \Reg_Bank/n5921 , \Reg_Bank/n5920 , \Reg_Bank/n5919 ,
         \Reg_Bank/n5918 , \Reg_Bank/n5917 , \Reg_Bank/n5916 ,
         \Reg_Bank/n5915 , \Reg_Bank/n5914 , \Reg_Bank/n5913 ,
         \Reg_Bank/n5912 , \Reg_Bank/n5911 , \Reg_Bank/n5910 ,
         \Reg_Bank/n5909 , \Reg_Bank/n5908 , \Reg_Bank/n5907 ,
         \Reg_Bank/n5906 , \Reg_Bank/n5905 , \Reg_Bank/n5904 ,
         \Reg_Bank/n5903 , \Reg_Bank/n5902 , \Reg_Bank/n5901 ,
         \Reg_Bank/n5900 , \Reg_Bank/n5899 , \Reg_Bank/n5898 ,
         \Reg_Bank/n5897 , \Reg_Bank/n5896 , \Reg_Bank/n5895 ,
         \Reg_Bank/n5894 , \Reg_Bank/n5893 , \Reg_Bank/n5892 ,
         \Reg_Bank/n5891 , \Reg_Bank/n5890 , \Reg_Bank/n5889 ,
         \Reg_Bank/n5888 , \Reg_Bank/n5887 , \Reg_Bank/n5886 ,
         \Reg_Bank/n5885 , \Reg_Bank/n5884 , \Reg_Bank/n5883 ,
         \Reg_Bank/n5882 , \Reg_Bank/n5881 , \Reg_Bank/n5880 ,
         \Reg_Bank/n5879 , \Reg_Bank/n5878 , \Reg_Bank/n5877 ,
         \Reg_Bank/n5876 , \Reg_Bank/n5875 , \Reg_Bank/n5874 ,
         \Reg_Bank/n5873 , \Reg_Bank/n5872 , \Reg_Bank/n5871 ,
         \Reg_Bank/n5870 , \Reg_Bank/n5869 , \Reg_Bank/n5868 ,
         \Reg_Bank/n5867 , \Reg_Bank/n5866 , \Reg_Bank/n5865 ,
         \Reg_Bank/n5864 , \Reg_Bank/n5863 , \Reg_Bank/n5862 ,
         \Reg_Bank/n5861 , \Reg_Bank/n5860 , \Reg_Bank/n5859 ,
         \Reg_Bank/n5858 , \Reg_Bank/n5857 , \Reg_Bank/n5856 ,
         \Reg_Bank/n5855 , \Reg_Bank/n5854 , \Reg_Bank/n5853 ,
         \Reg_Bank/n5852 , \Reg_Bank/n5851 , \Reg_Bank/n5850 ,
         \Reg_Bank/n5849 , \Reg_Bank/n5848 , \Reg_Bank/n5847 ,
         \Reg_Bank/n5846 , \Reg_Bank/n5845 , \Reg_Bank/n5844 ,
         \Reg_Bank/n5843 , \Reg_Bank/n5842 , \Reg_Bank/n5841 ,
         \Reg_Bank/n5840 , \Reg_Bank/n5839 , \Reg_Bank/n5838 ,
         \Reg_Bank/n5837 , \Reg_Bank/n5836 , \Reg_Bank/n5835 ,
         \Reg_Bank/n5834 , \Reg_Bank/n5833 , \Reg_Bank/n5832 ,
         \Reg_Bank/n5831 , \Reg_Bank/n5830 , \Reg_Bank/n5829 ,
         \Reg_Bank/n5828 , \Reg_Bank/n5827 , \Reg_Bank/n5826 ,
         \Reg_Bank/n5825 , \Reg_Bank/n5824 , \Reg_Bank/n5823 ,
         \Reg_Bank/n5822 , \Reg_Bank/n5821 , \Reg_Bank/n5820 ,
         \Reg_Bank/n5819 , \Reg_Bank/n5818 , \Reg_Bank/n5817 ,
         \Reg_Bank/n5816 , \Reg_Bank/n5815 , \Reg_Bank/n5814 ,
         \Reg_Bank/n5813 , \Reg_Bank/n5812 , \Reg_Bank/n5811 ,
         \Reg_Bank/n5810 , \Reg_Bank/n5809 , \Reg_Bank/n5808 ,
         \Reg_Bank/n5807 , \Reg_Bank/n5806 , \Reg_Bank/n5805 ,
         \Reg_Bank/n5804 , \Reg_Bank/n5803 , \Reg_Bank/n5802 ,
         \Reg_Bank/n5801 , \Reg_Bank/n5800 , \Reg_Bank/n5799 ,
         \Reg_Bank/n5798 , \Reg_Bank/n5797 , \Reg_Bank/n5796 ,
         \Reg_Bank/n5795 , \Reg_Bank/n5794 , \Reg_Bank/n5793 ,
         \Reg_Bank/n5792 , \Reg_Bank/n5791 , \Reg_Bank/n5790 ,
         \Reg_Bank/n5789 , \Reg_Bank/n5788 , \Reg_Bank/n5787 ,
         \Reg_Bank/n5786 , \Reg_Bank/n5785 , \Reg_Bank/n5784 ,
         \Reg_Bank/n5783 , \Reg_Bank/n5782 , \Reg_Bank/n5781 ,
         \Reg_Bank/n5780 , \Reg_Bank/n5779 , \Reg_Bank/n5778 ,
         \Reg_Bank/n5777 , \Reg_Bank/n5776 , \Reg_Bank/n5775 ,
         \Reg_Bank/n5774 , \Reg_Bank/n5773 , \Reg_Bank/n5772 ,
         \Reg_Bank/n5771 , \Reg_Bank/n5770 , \Reg_Bank/n5769 ,
         \Reg_Bank/n5768 , \Reg_Bank/n5767 , \Reg_Bank/n5766 ,
         \Reg_Bank/n5765 , \Reg_Bank/n5764 , \Reg_Bank/n5763 ,
         \Reg_Bank/n5762 , \Reg_Bank/n5761 , \Reg_Bank/n5760 ,
         \Reg_Bank/n5759 , \Reg_Bank/n5758 , \Reg_Bank/n5757 ,
         \Reg_Bank/n5756 , \Reg_Bank/n5755 , \Reg_Bank/n5754 ,
         \Reg_Bank/n5753 , \Reg_Bank/n5752 , \Reg_Bank/n5751 ,
         \Reg_Bank/n5750 , \Reg_Bank/n5749 , \Reg_Bank/n5748 ,
         \Reg_Bank/n5747 , \Reg_Bank/n5746 , \Reg_Bank/n5745 ,
         \Reg_Bank/n5744 , \Reg_Bank/n5743 , \Reg_Bank/n5742 ,
         \Reg_Bank/n5741 , \Reg_Bank/n5740 , \Reg_Bank/n5739 ,
         \Reg_Bank/n5738 , \Reg_Bank/n5737 , \Reg_Bank/n5736 ,
         \Reg_Bank/n5735 , \Reg_Bank/n5734 , \Reg_Bank/n5733 ,
         \Reg_Bank/n5732 , \Reg_Bank/n5731 , \Reg_Bank/n5730 ,
         \Reg_Bank/n5729 , \Reg_Bank/n5728 , \Reg_Bank/n5727 ,
         \Reg_Bank/n5726 , \Reg_Bank/n5725 , \Reg_Bank/n5724 ,
         \Reg_Bank/n5723 , \Reg_Bank/n5722 , \Reg_Bank/n5721 ,
         \Reg_Bank/n5720 , \Reg_Bank/n5719 , \Reg_Bank/n5718 ,
         \Reg_Bank/n5717 , \Reg_Bank/n5716 , \Reg_Bank/n5715 ,
         \Reg_Bank/n5714 , \Reg_Bank/n5713 , \Reg_Bank/n5712 ,
         \Reg_Bank/n5711 , \Reg_Bank/n5710 , \Reg_Bank/n5709 ,
         \Reg_Bank/n5708 , \Reg_Bank/n5707 , \Reg_Bank/n5706 ,
         \Reg_Bank/n5705 , \Reg_Bank/n5704 , \Reg_Bank/n5703 ,
         \Reg_Bank/n5702 , \Reg_Bank/n5701 , \Reg_Bank/n5700 ,
         \Reg_Bank/n5699 , \Reg_Bank/n5698 , \Reg_Bank/n5697 ,
         \Reg_Bank/n5696 , \Reg_Bank/n5695 , \Reg_Bank/n5694 ,
         \Reg_Bank/n5693 , \Reg_Bank/n5692 , \Reg_Bank/n5691 ,
         \Reg_Bank/n5690 , \Reg_Bank/n5689 , \Reg_Bank/n5688 ,
         \Reg_Bank/n5687 , \Reg_Bank/n5686 , \Reg_Bank/n5685 ,
         \Reg_Bank/n5684 , \Reg_Bank/n5683 , \Reg_Bank/n5682 ,
         \Reg_Bank/n5681 , \Reg_Bank/n5680 , \Reg_Bank/n5679 ,
         \Reg_Bank/n5678 , \Reg_Bank/n5677 , \Reg_Bank/n5676 ,
         \Reg_Bank/n5675 , \Reg_Bank/n5674 , \Reg_Bank/n5673 ,
         \Reg_Bank/n5672 , \Reg_Bank/n5671 , \Reg_Bank/n5670 ,
         \Reg_Bank/n5669 , \Reg_Bank/n5668 , \Reg_Bank/n5667 ,
         \Reg_Bank/n5666 , \Reg_Bank/n5665 , \Reg_Bank/n5664 ,
         \Reg_Bank/n5663 , \Reg_Bank/n5662 , \Reg_Bank/n5661 ,
         \Reg_Bank/n5660 , \Reg_Bank/n5659 , \Reg_Bank/n5658 ,
         \Reg_Bank/n5657 , \Reg_Bank/n5656 , \Reg_Bank/n5655 ,
         \Reg_Bank/n5654 , \Reg_Bank/n5653 , \Reg_Bank/n5652 ,
         \Reg_Bank/n5651 , \Reg_Bank/n5650 , \Reg_Bank/n5649 ,
         \Reg_Bank/n5648 , \Reg_Bank/n5647 , \Reg_Bank/n5646 ,
         \Reg_Bank/n5645 , \Reg_Bank/n5644 , \Reg_Bank/n5643 ,
         \Reg_Bank/n5642 , \Reg_Bank/n5641 , \Reg_Bank/n5640 ,
         \Reg_Bank/n5639 , \Reg_Bank/n5638 , \Reg_Bank/n5637 ,
         \Reg_Bank/n5636 , \Reg_Bank/n5635 , \Reg_Bank/n5634 ,
         \Reg_Bank/n5633 , \Reg_Bank/n5632 , \Reg_Bank/n5631 ,
         \Reg_Bank/n5630 , \Reg_Bank/n5629 , \Reg_Bank/n5628 ,
         \Reg_Bank/n5627 , \Reg_Bank/n5626 , \Reg_Bank/n5625 ,
         \Reg_Bank/n5624 , \Reg_Bank/n5623 , \Reg_Bank/n5622 ,
         \Reg_Bank/n5621 , \Reg_Bank/n5620 , \Reg_Bank/n5619 ,
         \Reg_Bank/n5618 , \Reg_Bank/n5617 , \Reg_Bank/n5616 ,
         \Reg_Bank/n5615 , \Reg_Bank/n5614 , \Reg_Bank/n5613 ,
         \Reg_Bank/n5612 , \Reg_Bank/n5611 , \Reg_Bank/n5610 ,
         \Reg_Bank/n5609 , \Reg_Bank/n5608 , \Reg_Bank/n5607 ,
         \Reg_Bank/n5606 , \Reg_Bank/n5605 , \Reg_Bank/n5604 ,
         \Reg_Bank/n5603 , \Reg_Bank/n5602 , \Reg_Bank/n5601 ,
         \Reg_Bank/n5600 , \Reg_Bank/n5599 , \Reg_Bank/n5598 ,
         \Reg_Bank/n5597 , \Reg_Bank/n5596 , \Reg_Bank/n5595 ,
         \Reg_Bank/n5594 , \Reg_Bank/n5593 , \Reg_Bank/n5592 ,
         \Reg_Bank/n5591 , \Reg_Bank/n5590 , \Reg_Bank/n5589 ,
         \Reg_Bank/n5588 , \Reg_Bank/n5587 , \Reg_Bank/n5586 ,
         \Reg_Bank/n5585 , \Reg_Bank/n5584 , \Reg_Bank/n5583 ,
         \Reg_Bank/n5582 , \Reg_Bank/n5581 , \Reg_Bank/n5580 ,
         \Reg_Bank/n5579 , \Reg_Bank/n5578 , \Reg_Bank/n5577 ,
         \Reg_Bank/n5576 , \Reg_Bank/n5575 , \Reg_Bank/n5574 ,
         \Reg_Bank/n5573 , \Reg_Bank/n5572 , \Reg_Bank/n5571 ,
         \Reg_Bank/n5570 , \Reg_Bank/n5569 , \Reg_Bank/n5568 ,
         \Reg_Bank/n5567 , \Reg_Bank/n5566 , \Reg_Bank/n5565 ,
         \Reg_Bank/n5564 , \Reg_Bank/n5563 , \Reg_Bank/n5562 ,
         \Reg_Bank/n5561 , \Reg_Bank/n5560 , \Reg_Bank/n5559 ,
         \Reg_Bank/n5558 , \Reg_Bank/n5557 , \Reg_Bank/n5556 ,
         \Reg_Bank/n5555 , \Reg_Bank/n5554 , \Reg_Bank/n5553 ,
         \Reg_Bank/n5552 , \Reg_Bank/n5551 , \Reg_Bank/n5550 ,
         \Reg_Bank/n5549 , \Reg_Bank/n5548 , \Reg_Bank/n5547 ,
         \Reg_Bank/n5546 , \Reg_Bank/n5545 , \Reg_Bank/n5544 ,
         \Reg_Bank/n5543 , \Reg_Bank/n5542 , \Reg_Bank/n5541 ,
         \Reg_Bank/n5540 , \Reg_Bank/n5539 , \Reg_Bank/n5538 ,
         \Reg_Bank/n5537 , \Reg_Bank/n5536 , \Reg_Bank/n5535 ,
         \Reg_Bank/n5534 , \Reg_Bank/n5533 , \Reg_Bank/n5532 ,
         \Reg_Bank/n5531 , \Reg_Bank/n5530 , \Reg_Bank/n5529 ,
         \Reg_Bank/n5528 , \Reg_Bank/n5527 , \Reg_Bank/n5526 ,
         \Reg_Bank/n5525 , \Reg_Bank/n5524 , \Reg_Bank/n5523 ,
         \Reg_Bank/n5522 , \Reg_Bank/n5521 , \Reg_Bank/n5520 ,
         \Reg_Bank/n5519 , \Reg_Bank/n5518 , \Reg_Bank/n5517 ,
         \Reg_Bank/n5516 , \Reg_Bank/n5515 , \Reg_Bank/n5514 ,
         \Reg_Bank/n5513 , \Reg_Bank/n5512 , \Reg_Bank/n5511 ,
         \Reg_Bank/n5510 , \Reg_Bank/n5509 , \Reg_Bank/n5508 ,
         \Reg_Bank/n5507 , \Reg_Bank/n5506 , \Reg_Bank/n5505 ,
         \Reg_Bank/n5504 , \Reg_Bank/n5503 , \Reg_Bank/n5502 ,
         \Reg_Bank/n5501 , \Reg_Bank/n5500 , \Reg_Bank/n5499 ,
         \Reg_Bank/n5498 , \Reg_Bank/n5497 , \Reg_Bank/n5496 ,
         \Reg_Bank/n5495 , \Reg_Bank/n5494 , \Reg_Bank/n5493 ,
         \Reg_Bank/n5492 , \Reg_Bank/n5491 , \Reg_Bank/n5490 ,
         \Reg_Bank/n5489 , \Reg_Bank/n5488 , \Reg_Bank/n5487 ,
         \Reg_Bank/n5486 , \Reg_Bank/n5485 , \Reg_Bank/n5484 ,
         \Reg_Bank/n5483 , \Reg_Bank/n5482 , \Reg_Bank/n5481 ,
         \Reg_Bank/n5480 , \Reg_Bank/n5479 , \Reg_Bank/n5478 ,
         \Reg_Bank/n5477 , \Reg_Bank/n5476 , \Reg_Bank/n5475 ,
         \Reg_Bank/n5474 , \Reg_Bank/n5473 , \Reg_Bank/n5472 ,
         \Reg_Bank/n5471 , \Reg_Bank/n5470 , \Reg_Bank/n5469 ,
         \Reg_Bank/n5468 , \Reg_Bank/n5467 , \Reg_Bank/n5466 ,
         \Reg_Bank/n5465 , \Reg_Bank/n5464 , \Reg_Bank/n5463 ,
         \Reg_Bank/n5462 , \Reg_Bank/n5461 , \Reg_Bank/n5460 ,
         \Reg_Bank/n5459 , \Reg_Bank/n5458 , \Reg_Bank/n5457 ,
         \Reg_Bank/n5456 , \Reg_Bank/n5455 , \Reg_Bank/n5454 ,
         \Reg_Bank/n5453 , \Reg_Bank/n5452 , \Reg_Bank/n5451 ,
         \Reg_Bank/n5450 , \Reg_Bank/n5449 , \Reg_Bank/n5448 ,
         \Reg_Bank/n5447 , \Reg_Bank/n5446 , \Reg_Bank/n5445 ,
         \Reg_Bank/n5444 , \Reg_Bank/n5443 , \Reg_Bank/n5442 ,
         \Reg_Bank/n5441 , \Reg_Bank/n5440 , \Reg_Bank/n5439 ,
         \Reg_Bank/n5438 , \Reg_Bank/n5437 , \Reg_Bank/n5436 ,
         \Reg_Bank/n5435 , \Reg_Bank/n5434 , \Reg_Bank/n5433 ,
         \Reg_Bank/n5432 , \Reg_Bank/n5431 , \Reg_Bank/n5430 ,
         \Reg_Bank/n5429 , \Reg_Bank/n5428 , \Reg_Bank/n5427 ,
         \Reg_Bank/n5426 , \Reg_Bank/n5425 , \Reg_Bank/n5424 ,
         \Reg_Bank/n5423 , \Reg_Bank/n5422 , \Reg_Bank/n5421 ,
         \Reg_Bank/n5420 , \Reg_Bank/n5419 , \Reg_Bank/n5418 ,
         \Reg_Bank/n5417 , \Reg_Bank/n5416 , \Reg_Bank/n5415 ,
         \Reg_Bank/n5414 , \Reg_Bank/n5413 , \Reg_Bank/n5412 ,
         \Reg_Bank/n5411 , \Reg_Bank/n5410 , \Reg_Bank/n5409 ,
         \Reg_Bank/n5408 , \Reg_Bank/n5407 , \Reg_Bank/n5406 ,
         \Reg_Bank/n5405 , \Reg_Bank/n5404 , \Reg_Bank/n5403 ,
         \Reg_Bank/n5402 , \Reg_Bank/n5401 , \Reg_Bank/n5400 ,
         \Reg_Bank/n5399 , \Reg_Bank/n5398 , \Reg_Bank/n5397 ,
         \Reg_Bank/n5396 , \Reg_Bank/n5395 , \Reg_Bank/n5394 ,
         \Reg_Bank/n5393 , \Reg_Bank/n5392 , \Reg_Bank/n5391 ,
         \Reg_Bank/n5390 , \Reg_Bank/n5389 , \Reg_Bank/n5388 ,
         \Reg_Bank/n5387 , \Reg_Bank/n5386 , \Reg_Bank/n5385 ,
         \Reg_Bank/n5384 , \Reg_Bank/n5383 , \Reg_Bank/n5382 ,
         \Reg_Bank/n5381 , \Reg_Bank/n5380 , \Reg_Bank/n5379 ,
         \Reg_Bank/n5378 , \Reg_Bank/n5377 , \Reg_Bank/n5376 ,
         \Reg_Bank/n5375 , \Reg_Bank/n5374 , \Reg_Bank/n5373 ,
         \Reg_Bank/n5372 , \Reg_Bank/n5371 , \Reg_Bank/n5370 ,
         \Reg_Bank/n5369 , \Reg_Bank/n5368 , \Reg_Bank/n5367 ,
         \Reg_Bank/n5366 , \Reg_Bank/n5365 , \Reg_Bank/n5364 ,
         \Reg_Bank/n5363 , \Reg_Bank/n5362 , \Reg_Bank/n5361 ,
         \Reg_Bank/n5360 , \Reg_Bank/n5359 , \Reg_Bank/n5358 ,
         \Reg_Bank/n5357 , \Reg_Bank/n5356 , \Reg_Bank/n5355 ,
         \Reg_Bank/n5354 , \Reg_Bank/n5353 , \Reg_Bank/n5352 ,
         \Reg_Bank/n5351 , \Reg_Bank/n5350 , \Reg_Bank/n5349 ,
         \Reg_Bank/n5348 , \Reg_Bank/n5347 , \Reg_Bank/n5346 ,
         \Reg_Bank/n5345 , \Reg_Bank/n5344 , \Reg_Bank/n5343 ,
         \Reg_Bank/n5342 , \Reg_Bank/n5341 , \Reg_Bank/n5340 ,
         \Reg_Bank/n5339 , \Reg_Bank/n5338 , \Reg_Bank/n5337 ,
         \Reg_Bank/n5336 , \Reg_Bank/n5335 , \Reg_Bank/n5334 ,
         \Reg_Bank/n5333 , \Reg_Bank/n5332 , \Reg_Bank/n5331 ,
         \Reg_Bank/n5330 , \Reg_Bank/n5329 , \Reg_Bank/n5328 ,
         \Reg_Bank/n5327 , \Reg_Bank/n5326 , \Reg_Bank/n5325 ,
         \Reg_Bank/n5324 , \Reg_Bank/n5323 , \Reg_Bank/n5322 ,
         \Reg_Bank/n5321 , \Reg_Bank/n5320 , \Reg_Bank/n5319 ,
         \Reg_Bank/n5318 , \Reg_Bank/n5317 , \Reg_Bank/n5316 ,
         \Reg_Bank/n5315 , \Reg_Bank/n5314 , \Reg_Bank/n5313 ,
         \Reg_Bank/n5312 , \Reg_Bank/n5311 , \Reg_Bank/n5310 ,
         \Reg_Bank/n5309 , \Reg_Bank/n5308 , \Reg_Bank/n5307 ,
         \Reg_Bank/n5306 , \Reg_Bank/n5305 , \Reg_Bank/n5304 ,
         \Reg_Bank/n5303 , \Reg_Bank/n5302 , \Reg_Bank/n5301 ,
         \Reg_Bank/n5300 , \Reg_Bank/n5299 , \Reg_Bank/n5298 ,
         \Reg_Bank/n5297 , \Reg_Bank/n5296 , \Reg_Bank/n5295 ,
         \Reg_Bank/n5294 , \Reg_Bank/n5293 , \Reg_Bank/n5292 ,
         \Reg_Bank/n5291 , \Reg_Bank/n5290 , \Reg_Bank/n5289 ,
         \Reg_Bank/n5288 , \Reg_Bank/n5287 , \Reg_Bank/n5286 ,
         \Reg_Bank/n5285 , \Reg_Bank/n5284 , \Reg_Bank/n5283 ,
         \Reg_Bank/n5282 , \Reg_Bank/n5281 , \Reg_Bank/n5280 ,
         \Reg_Bank/n5279 , \Reg_Bank/n5278 , \Reg_Bank/n5277 ,
         \Reg_Bank/n5276 , \Reg_Bank/n5275 , \Reg_Bank/n5274 ,
         \Reg_Bank/n5273 , \Reg_Bank/n5272 , \Reg_Bank/n5271 ,
         \Reg_Bank/n5270 , \Reg_Bank/n5269 , \Reg_Bank/n5268 ,
         \Reg_Bank/n5267 , \Reg_Bank/n5266 , \Reg_Bank/n5265 ,
         \Reg_Bank/n5264 , \Reg_Bank/n5263 , \Reg_Bank/n5262 ,
         \Reg_Bank/n5261 , \Reg_Bank/n5260 , \Reg_Bank/n5259 ,
         \Reg_Bank/n5258 , \Reg_Bank/n5257 , \Reg_Bank/n5256 ,
         \Reg_Bank/n5255 , \Reg_Bank/n5254 , \Reg_Bank/n5253 ,
         \Reg_Bank/n5252 , \Reg_Bank/n5251 , \Reg_Bank/n5250 ,
         \Reg_Bank/n5249 , \Reg_Bank/n5248 , \Reg_Bank/n5247 ,
         \Reg_Bank/n5246 , \Reg_Bank/n5245 , \Reg_Bank/n5244 ,
         \Reg_Bank/n5243 , \Reg_Bank/n5242 , \Reg_Bank/n5241 ,
         \Reg_Bank/n5240 , \Reg_Bank/n5239 , \Reg_Bank/n5238 ,
         \Reg_Bank/n5237 , \Reg_Bank/n5236 , \Reg_Bank/n5235 ,
         \Reg_Bank/n5234 , \Reg_Bank/n5233 , \Reg_Bank/n5232 ,
         \Reg_Bank/n5231 , \Reg_Bank/n5230 , \Reg_Bank/n5229 ,
         \Reg_Bank/n5228 , \Reg_Bank/n5227 , \Reg_Bank/n5226 ,
         \Reg_Bank/n5225 , \Reg_Bank/n5224 , \Reg_Bank/n5223 ,
         \Reg_Bank/n5222 , \Reg_Bank/n5221 , \Reg_Bank/n5220 ,
         \Reg_Bank/n5219 , \Reg_Bank/n5218 , \Reg_Bank/n5217 ,
         \Reg_Bank/n5216 , \Reg_Bank/n5215 , \Reg_Bank/n5214 ,
         \Reg_Bank/n5213 , \Reg_Bank/n5212 , \Reg_Bank/n5211 ,
         \Reg_Bank/n5210 , \Reg_Bank/n5209 , \Reg_Bank/n5208 ,
         \Reg_Bank/n5207 , \Reg_Bank/n5206 , \Reg_Bank/n5205 ,
         \Reg_Bank/n5204 , \Reg_Bank/n5203 , \Reg_Bank/n5202 ,
         \Reg_Bank/n5201 , \Reg_Bank/n5200 , \Reg_Bank/n5199 ,
         \Reg_Bank/n5198 , \Reg_Bank/n5197 , \Reg_Bank/n5196 ,
         \Reg_Bank/n5195 , \Reg_Bank/n5194 , \Reg_Bank/n5193 ,
         \Reg_Bank/n5192 , \Reg_Bank/n5191 , \Reg_Bank/n5190 ,
         \Reg_Bank/n5189 , \Reg_Bank/n5188 , \Reg_Bank/n5187 ,
         \Reg_Bank/n5186 , \Reg_Bank/n5185 , \Reg_Bank/n5184 ,
         \Reg_Bank/n5183 , \Reg_Bank/n5182 , \Reg_Bank/n5181 ,
         \Reg_Bank/n5180 , \Reg_Bank/n5179 , \Reg_Bank/n5178 ,
         \Reg_Bank/n5177 , \Reg_Bank/n5176 , \Reg_Bank/n5175 ,
         \Reg_Bank/n5174 , \Reg_Bank/n5173 , \Reg_Bank/n5172 ,
         \Reg_Bank/n5171 , \Reg_Bank/n5170 , \Reg_Bank/n5169 ,
         \Reg_Bank/n5168 , \Reg_Bank/n5167 , \Reg_Bank/n5166 ,
         \Reg_Bank/n5165 , \Reg_Bank/n5164 , \Reg_Bank/n5163 ,
         \Reg_Bank/n5162 , \Reg_Bank/n5161 , \Reg_Bank/n5160 ,
         \Reg_Bank/n5159 , \Reg_Bank/n5158 , \Reg_Bank/n5157 ,
         \Reg_Bank/n5156 , \Reg_Bank/n5155 , \Reg_Bank/n5154 ,
         \Reg_Bank/n5153 , \Reg_Bank/n5152 , \Reg_Bank/n5151 ,
         \Reg_Bank/n5150 , \Reg_Bank/n5149 , \Reg_Bank/n5148 ,
         \Reg_Bank/n5147 , \Reg_Bank/n5146 , \Reg_Bank/n5145 ,
         \Reg_Bank/n5144 , \Reg_Bank/n5143 , \Reg_Bank/n5142 ,
         \Reg_Bank/n5141 , \Reg_Bank/n5140 , \Reg_Bank/n5139 ,
         \Reg_Bank/n5138 , \Reg_Bank/n5137 , \Reg_Bank/n5136 ,
         \Reg_Bank/n5135 , \Reg_Bank/n5134 , \Reg_Bank/n5133 ,
         \Reg_Bank/n5132 , \Reg_Bank/n5131 , \Reg_Bank/n5130 ,
         \Reg_Bank/n5129 , \Reg_Bank/n5128 , \Reg_Bank/n5127 ,
         \Reg_Bank/n5126 , \Reg_Bank/n5125 , \Reg_Bank/n5124 ,
         \Reg_Bank/n5123 , \Reg_Bank/n5122 , \Reg_Bank/n5121 ,
         \Reg_Bank/n5120 , \Reg_Bank/n5119 , \Reg_Bank/n5118 ,
         \Reg_Bank/n5117 , \Reg_Bank/n5116 , \Reg_Bank/n5115 ,
         \Reg_Bank/n5114 , \Reg_Bank/n5113 , \Reg_Bank/n5112 ,
         \Reg_Bank/n5111 , \Reg_Bank/n5110 , \Reg_Bank/n5109 ,
         \Reg_Bank/n5108 , \Reg_Bank/n5107 , \Reg_Bank/n5106 ,
         \Reg_Bank/n5105 , \Reg_Bank/n5104 , \Reg_Bank/n5103 ,
         \Reg_Bank/n5102 , \Reg_Bank/n5101 , \Reg_Bank/n5100 ,
         \Reg_Bank/n5099 , \Reg_Bank/n5098 , \Reg_Bank/n5097 ,
         \Reg_Bank/n5096 , \Reg_Bank/n5095 , \Reg_Bank/n5094 ,
         \Reg_Bank/n5093 , \Reg_Bank/n5092 , \Reg_Bank/n5091 ,
         \Reg_Bank/n5090 , \Reg_Bank/n5089 , \Reg_Bank/n5088 ,
         \Reg_Bank/n5087 , \Reg_Bank/n5086 , \Reg_Bank/n5085 ,
         \Reg_Bank/n5084 , \Reg_Bank/n5083 , \Reg_Bank/n5082 ,
         \Reg_Bank/n5081 , \Reg_Bank/n5080 , \Reg_Bank/n5079 ,
         \Reg_Bank/n5078 , \Reg_Bank/n5077 , \Reg_Bank/n5076 ,
         \Reg_Bank/n5075 , \Reg_Bank/n5074 , \Reg_Bank/n5073 ,
         \Reg_Bank/n5072 , \Reg_Bank/n5071 , \Reg_Bank/n5070 ,
         \Reg_Bank/n5069 , \Reg_Bank/n5068 , \Reg_Bank/n5067 ,
         \Reg_Bank/n5066 , \Reg_Bank/n5065 , \Reg_Bank/n5064 ,
         \Reg_Bank/n5063 , \Reg_Bank/n5062 , \Reg_Bank/n5061 ,
         \Reg_Bank/n5060 , \Reg_Bank/n5059 , \Reg_Bank/n5058 ,
         \Reg_Bank/n5057 , \Reg_Bank/n5056 , \Reg_Bank/n5055 ,
         \Reg_Bank/n5054 , \Reg_Bank/n5053 , \Reg_Bank/n5052 ,
         \Reg_Bank/n5051 , \Reg_Bank/n5050 , \Reg_Bank/n5049 ,
         \Reg_Bank/n5048 , \Reg_Bank/n5047 , \Reg_Bank/n5046 ,
         \Reg_Bank/n5045 , \Reg_Bank/n5044 , \Reg_Bank/n5043 ,
         \Reg_Bank/n5042 , \Reg_Bank/n5041 , \Reg_Bank/n5040 ,
         \Reg_Bank/n5039 , \Reg_Bank/n5038 , \Reg_Bank/n5037 ,
         \Reg_Bank/n5036 , \Reg_Bank/n5035 , \Reg_Bank/n5034 ,
         \Reg_Bank/n5033 , \Reg_Bank/n5032 , \Reg_Bank/n5031 ,
         \Reg_Bank/n5030 , \Reg_Bank/n5029 , \Reg_Bank/n5028 ,
         \Reg_Bank/n5027 , \Reg_Bank/n5026 , \Reg_Bank/n5025 ,
         \Reg_Bank/n5024 , \Reg_Bank/n5023 , \Reg_Bank/n5022 ,
         \Reg_Bank/n5021 , \Reg_Bank/n5020 , \Reg_Bank/n5019 ,
         \Reg_Bank/n5018 , \Reg_Bank/n5017 , \Reg_Bank/n5016 ,
         \Reg_Bank/n5015 , \Reg_Bank/n5014 , \Reg_Bank/n5013 ,
         \Reg_Bank/n5012 , \Reg_Bank/n5011 , \Reg_Bank/n5010 ,
         \Reg_Bank/n5009 , \Reg_Bank/n5008 , \Reg_Bank/n5007 ,
         \Reg_Bank/n5006 , \Reg_Bank/n5005 , \Reg_Bank/n5004 ,
         \Reg_Bank/n5003 , \Reg_Bank/n5002 , \Reg_Bank/n5001 ,
         \Reg_Bank/n5000 , \Reg_Bank/n4999 , \Reg_Bank/n4998 ,
         \Reg_Bank/n4997 , \Reg_Bank/n4996 , \Reg_Bank/n4995 ,
         \Reg_Bank/n4994 , \Reg_Bank/n4993 , \Reg_Bank/n4992 ,
         \Reg_Bank/n4991 , \Reg_Bank/n4990 , \Reg_Bank/n4989 ,
         \Reg_Bank/n4988 , \Reg_Bank/n4987 , \Reg_Bank/n4986 ,
         \Reg_Bank/n4985 , \Reg_Bank/n4984 , \Reg_Bank/n4983 ,
         \Reg_Bank/n4982 , \Reg_Bank/n4981 , \Reg_Bank/n4980 ,
         \Reg_Bank/n4979 , \Reg_Bank/n4978 , \Reg_Bank/n4977 ,
         \Reg_Bank/n4976 , \Reg_Bank/n4975 , \Reg_Bank/n4974 ,
         \Reg_Bank/n4973 , \Reg_Bank/n4972 , \Reg_Bank/n4971 ,
         \Reg_Bank/n4970 , \Reg_Bank/n4969 , \Reg_Bank/n4968 ,
         \Reg_Bank/n4967 , \Reg_Bank/n4966 , \Reg_Bank/n4965 ,
         \Reg_Bank/n4964 , \Reg_Bank/n4963 , \Reg_Bank/n4962 ,
         \Reg_Bank/n4961 , \Reg_Bank/n4960 , \Reg_Bank/n4959 ,
         \Reg_Bank/n4958 , \Reg_Bank/n4957 , \Reg_Bank/n4956 ,
         \Reg_Bank/n4955 , \Reg_Bank/n4954 , \Reg_Bank/n4953 ,
         \Reg_Bank/n4952 , \Reg_Bank/n4951 , \Reg_Bank/n4950 ,
         \Reg_Bank/n4949 , \Reg_Bank/n4948 , \Reg_Bank/n4947 ,
         \Reg_Bank/n4946 , \Reg_Bank/n4945 , \Reg_Bank/n4944 ,
         \Reg_Bank/n4943 , \Reg_Bank/n4942 , \Reg_Bank/n4941 ,
         \Reg_Bank/n4940 , \Reg_Bank/n4939 , \Reg_Bank/n4938 ,
         \Reg_Bank/n4937 , \Reg_Bank/n4936 , \Reg_Bank/n4935 ,
         \Reg_Bank/n4934 , \Reg_Bank/n4933 , \Reg_Bank/n4932 ,
         \Reg_Bank/n4931 , \Reg_Bank/n4930 , \Reg_Bank/n4929 ,
         \Reg_Bank/n4928 , \Reg_Bank/n4927 , \Reg_Bank/n4926 ,
         \Reg_Bank/n4925 , \Reg_Bank/n4924 , \Reg_Bank/n4923 ,
         \Reg_Bank/n4922 , \Reg_Bank/n4921 , \Reg_Bank/n4920 ,
         \Reg_Bank/n4919 , \Reg_Bank/n4918 , \Reg_Bank/n4917 ,
         \Reg_Bank/n4916 , \Reg_Bank/n4915 , \Reg_Bank/n4914 ,
         \Reg_Bank/n4913 , \Reg_Bank/n4912 , \Reg_Bank/n4911 ,
         \Reg_Bank/n4910 , \Reg_Bank/n4909 , \Reg_Bank/n4908 ,
         \Reg_Bank/n4907 , \Reg_Bank/n4906 , \Reg_Bank/n4905 ,
         \Reg_Bank/n4904 , \Reg_Bank/n4903 , \Reg_Bank/n4902 ,
         \Reg_Bank/n4901 , \Reg_Bank/n4900 , \Reg_Bank/n4899 ,
         \Reg_Bank/n4898 , \Reg_Bank/n4897 , \Reg_Bank/n4896 ,
         \Reg_Bank/n4895 , \Reg_Bank/n4894 , \Reg_Bank/n4893 ,
         \Reg_Bank/n4892 , \Reg_Bank/n4891 , \Reg_Bank/n4890 ,
         \Reg_Bank/n4889 , \Reg_Bank/n4888 , \Reg_Bank/n4887 ,
         \Reg_Bank/n4886 , \Reg_Bank/n4885 , \Reg_Bank/n4884 ,
         \Reg_Bank/n4883 , \Reg_Bank/n4882 , \Reg_Bank/n4881 ,
         \Reg_Bank/n4880 , \Reg_Bank/n4879 , \Reg_Bank/n4878 ,
         \Reg_Bank/n4877 , \Reg_Bank/n4876 , \Reg_Bank/n4875 ,
         \Reg_Bank/n4874 , \Reg_Bank/n4873 , \Reg_Bank/n4872 ,
         \Reg_Bank/n4871 , \Reg_Bank/n4870 , \Reg_Bank/n4869 ,
         \Reg_Bank/n4868 , \Reg_Bank/n4867 , \Reg_Bank/n4866 ,
         \Reg_Bank/n4865 , \Reg_Bank/n4864 , \Reg_Bank/n4863 ,
         \Reg_Bank/n4862 , \Reg_Bank/n4861 , \Reg_Bank/n4860 ,
         \Reg_Bank/n4859 , \Reg_Bank/n4858 , \Reg_Bank/n4857 ,
         \Reg_Bank/n4856 , \Reg_Bank/n4855 , \Reg_Bank/n4854 ,
         \Reg_Bank/n4853 , \Reg_Bank/n4852 , \Reg_Bank/n4851 ,
         \Reg_Bank/n4850 , \Reg_Bank/n4849 , \Reg_Bank/n4848 ,
         \Reg_Bank/n4847 , \Reg_Bank/n4846 , \Reg_Bank/n4845 ,
         \Reg_Bank/n4844 , \Reg_Bank/n4843 , \Reg_Bank/n4842 ,
         \Reg_Bank/n4841 , \Reg_Bank/n4840 , \Reg_Bank/n4839 ,
         \Reg_Bank/n4838 , \Reg_Bank/n4837 , \Reg_Bank/n4836 ,
         \Reg_Bank/n4835 , \Reg_Bank/n4834 , \Reg_Bank/n4833 ,
         \Reg_Bank/n4832 , \Reg_Bank/n4831 , \Reg_Bank/n4830 ,
         \Reg_Bank/n4829 , \Reg_Bank/n4828 , \Reg_Bank/n4827 ,
         \Reg_Bank/n4826 , \Reg_Bank/n4825 , \Reg_Bank/n4824 ,
         \Reg_Bank/n4823 , \Reg_Bank/n4822 , \Reg_Bank/n4821 ,
         \Reg_Bank/n4820 , \Reg_Bank/n4819 , \Reg_Bank/n4818 ,
         \Reg_Bank/n4817 , \Reg_Bank/n4816 , \Reg_Bank/n4815 ,
         \Reg_Bank/n4814 , \Reg_Bank/n4813 , \Reg_Bank/n4812 ,
         \Reg_Bank/n4811 , \Reg_Bank/n4810 , \Reg_Bank/n4809 ,
         \Reg_Bank/n4808 , \Reg_Bank/n4807 , \Reg_Bank/n4806 ,
         \Reg_Bank/n4805 , \Reg_Bank/n4804 , \Reg_Bank/n4803 ,
         \Reg_Bank/n4802 , \Reg_Bank/n4801 , \Reg_Bank/n4800 ,
         \Reg_Bank/n4799 , \Reg_Bank/n4798 , \Reg_Bank/n4797 ,
         \Reg_Bank/n4796 , \Reg_Bank/n4795 , \Reg_Bank/n4794 ,
         \Reg_Bank/n4793 , \Reg_Bank/n4792 , \Reg_Bank/n4791 ,
         \Reg_Bank/n4790 , \Reg_Bank/n4789 , \Reg_Bank/n4788 ,
         \Reg_Bank/n4787 , \Reg_Bank/n4786 , \Reg_Bank/n4785 ,
         \Reg_Bank/n4784 , \Reg_Bank/n4783 , \Reg_Bank/n4782 ,
         \Reg_Bank/n4781 , \Reg_Bank/n4780 , \Reg_Bank/n4779 ,
         \Reg_Bank/n4778 , \Reg_Bank/n4777 , \Reg_Bank/n4776 ,
         \Reg_Bank/n4775 , \Reg_Bank/n4774 , \Reg_Bank/n4773 ,
         \Reg_Bank/n4772 , \Reg_Bank/n4771 , \Reg_Bank/n4770 ,
         \Reg_Bank/n4769 , \Reg_Bank/n4768 , \Reg_Bank/n4767 ,
         \Reg_Bank/n4766 , \Reg_Bank/n4765 , \Reg_Bank/n4764 ,
         \Reg_Bank/n4763 , \Reg_Bank/n4762 , \Reg_Bank/n4761 ,
         \Reg_Bank/n4760 , \Reg_Bank/n4759 , \Reg_Bank/n4758 ,
         \Reg_Bank/n4757 , \Reg_Bank/n4756 , \Reg_Bank/n4755 ,
         \Reg_Bank/n4754 , \Reg_Bank/n4753 , \Reg_Bank/n4752 ,
         \Reg_Bank/n4751 , \Reg_Bank/n4750 , \Reg_Bank/n4749 ,
         \Reg_Bank/n4748 , \Reg_Bank/n4747 , \Reg_Bank/n4746 ,
         \Reg_Bank/n4745 , \Reg_Bank/n4744 , \Reg_Bank/n4743 ,
         \Reg_Bank/n4742 , \Reg_Bank/n4741 , \Reg_Bank/n4740 ,
         \Reg_Bank/n4739 , \Reg_Bank/n4738 , \Reg_Bank/n4737 ,
         \Reg_Bank/n4736 , \Reg_Bank/n4735 , \Reg_Bank/n4734 ,
         \Reg_Bank/n4733 , \Reg_Bank/n4732 , \Reg_Bank/n4731 ,
         \Reg_Bank/n4730 , \Reg_Bank/n4729 , \Reg_Bank/n4728 ,
         \Reg_Bank/n4727 , \Reg_Bank/n4726 , \Reg_Bank/n4725 ,
         \Reg_Bank/n4724 , \Reg_Bank/n4723 , \Reg_Bank/n4722 ,
         \Reg_Bank/n4721 , \Reg_Bank/n4720 , \Reg_Bank/n4719 ,
         \Reg_Bank/n4718 , \Reg_Bank/n4717 , \Reg_Bank/n4716 ,
         \Reg_Bank/n4715 , \Reg_Bank/n4714 , \Reg_Bank/n4713 ,
         \Reg_Bank/n4712 , \Reg_Bank/n4711 , \Reg_Bank/n4710 ,
         \Reg_Bank/n4709 , \Reg_Bank/n4708 , \Reg_Bank/n4707 ,
         \Reg_Bank/n4706 , \Reg_Bank/n4705 , \Reg_Bank/n4704 ,
         \Reg_Bank/n4703 , \Reg_Bank/n4702 , \Reg_Bank/n4701 ,
         \Reg_Bank/n4700 , \Reg_Bank/n4699 , \Reg_Bank/n4698 ,
         \Reg_Bank/n4697 , \Reg_Bank/n4696 , \Reg_Bank/n4695 ,
         \Reg_Bank/n4694 , \Reg_Bank/n4693 , \Reg_Bank/n4692 ,
         \Reg_Bank/n4691 , \Reg_Bank/n4690 , \Reg_Bank/n4689 ,
         \Reg_Bank/n4688 , \Reg_Bank/n4687 , \Reg_Bank/n4686 ,
         \Reg_Bank/n4685 , \Reg_Bank/n4684 , \Reg_Bank/n4683 ,
         \Reg_Bank/n4682 , \Reg_Bank/n4681 , \Reg_Bank/n4680 ,
         \Reg_Bank/n4679 , \Reg_Bank/n4678 , \Reg_Bank/n4677 ,
         \Reg_Bank/n4676 , \Reg_Bank/n4675 , \Reg_Bank/n4674 ,
         \Reg_Bank/n4673 , \Reg_Bank/n4672 , \Reg_Bank/n4671 ,
         \Reg_Bank/n4670 , \Reg_Bank/n4669 , \Reg_Bank/n4668 ,
         \Reg_Bank/n4667 , \Reg_Bank/n4666 , \Reg_Bank/n4665 ,
         \Reg_Bank/n4664 , \Reg_Bank/n4663 , \Reg_Bank/n4662 ,
         \Reg_Bank/n4661 , \Reg_Bank/n4660 , \Reg_Bank/n4659 ,
         \Reg_Bank/n4658 , \Reg_Bank/n4657 , \Reg_Bank/n4656 ,
         \Reg_Bank/n4655 , \Reg_Bank/n4654 , \Reg_Bank/n4653 ,
         \Reg_Bank/n4652 , \Reg_Bank/n4651 , \Reg_Bank/n4650 ,
         \Reg_Bank/n4649 , \Reg_Bank/n4648 , \Reg_Bank/n4647 ,
         \Reg_Bank/n4646 , \Reg_Bank/n4645 , \Reg_Bank/n4644 ,
         \Reg_Bank/n4643 , \Reg_Bank/n4642 , \Reg_Bank/n4641 ,
         \Reg_Bank/n4640 , \Reg_Bank/n4639 , \Reg_Bank/n4638 ,
         \Reg_Bank/n4637 , \Reg_Bank/n4636 , \Reg_Bank/n4635 ,
         \Reg_Bank/n4634 , \Reg_Bank/n4633 , \Reg_Bank/n4632 ,
         \Reg_Bank/n4631 , \Reg_Bank/n4630 , \Reg_Bank/n4629 ,
         \Reg_Bank/n4628 , \Reg_Bank/n4627 , \Reg_Bank/n4626 ,
         \Reg_Bank/n4625 , \Reg_Bank/n4624 , \Reg_Bank/n4623 ,
         \Reg_Bank/n4622 , \Reg_Bank/n4621 , \Reg_Bank/n4620 ,
         \Reg_Bank/n4619 , \Reg_Bank/n4618 , \Reg_Bank/n4617 ,
         \Reg_Bank/n4616 , \Reg_Bank/n4615 , \Reg_Bank/n4614 ,
         \Reg_Bank/n4613 , \Reg_Bank/n4612 , \Reg_Bank/n4611 ,
         \Reg_Bank/n4610 , \Reg_Bank/n4609 , \Reg_Bank/n4608 ,
         \Reg_Bank/n4607 , \Reg_Bank/n4606 , \Reg_Bank/n4605 ,
         \Reg_Bank/n4604 , \Reg_Bank/n4603 , \Reg_Bank/n4602 ,
         \Reg_Bank/n4601 , \Reg_Bank/n4600 , \Reg_Bank/n4599 ,
         \Reg_Bank/n4598 , \Reg_Bank/n4597 , \Reg_Bank/n4596 ,
         \Reg_Bank/n4595 , \Reg_Bank/n4594 , \Reg_Bank/n4593 ,
         \Reg_Bank/n4592 , \Reg_Bank/n4591 , \Reg_Bank/n4590 ,
         \Reg_Bank/n4589 , \Reg_Bank/n4588 , \Reg_Bank/n4587 ,
         \Reg_Bank/n4586 , \Reg_Bank/n4585 , \Reg_Bank/n4584 ,
         \Reg_Bank/n4583 , \Reg_Bank/n4582 , \Reg_Bank/n4581 ,
         \Reg_Bank/n4580 , \Reg_Bank/n4579 , \Reg_Bank/n4578 ,
         \Reg_Bank/n4577 , \Reg_Bank/n4576 , \Reg_Bank/n4575 ,
         \Reg_Bank/n4574 , \Reg_Bank/n4573 , \Reg_Bank/n4572 ,
         \Reg_Bank/n4571 , \Reg_Bank/n4570 , \Reg_Bank/n4569 ,
         \Reg_Bank/n4568 , \Reg_Bank/n4567 , \Reg_Bank/n4566 ,
         \Reg_Bank/n4565 , \Reg_Bank/n4564 , \Reg_Bank/n4563 ,
         \Reg_Bank/n4562 , \Reg_Bank/n4561 , \Reg_Bank/n4560 ,
         \Reg_Bank/n4559 , \Reg_Bank/n4558 , \Reg_Bank/n4557 ,
         \Reg_Bank/n4556 , \Reg_Bank/n4555 , \Reg_Bank/n4554 ,
         \Reg_Bank/n4553 , \Reg_Bank/n4552 , \Reg_Bank/n4551 ,
         \Reg_Bank/n4550 , \Reg_Bank/n4549 , \Reg_Bank/n4548 ,
         \Reg_Bank/n4547 , \Reg_Bank/n4546 , \Reg_Bank/n4545 ,
         \Reg_Bank/n4544 , \Reg_Bank/n4543 , \Reg_Bank/n4542 ,
         \Reg_Bank/n4541 , \Reg_Bank/n4540 , \Reg_Bank/n4539 ,
         \Reg_Bank/n4538 , \Reg_Bank/n4537 , \Reg_Bank/n4536 ,
         \Reg_Bank/n4535 , \Reg_Bank/n4534 , \Reg_Bank/n4533 ,
         \Reg_Bank/n4532 , \Reg_Bank/n4531 , \Reg_Bank/n4530 ,
         \Reg_Bank/n4529 , \Reg_Bank/n4528 , \Reg_Bank/n4527 ,
         \Reg_Bank/n4526 , \Reg_Bank/n4525 , \Reg_Bank/n4524 ,
         \Reg_Bank/n4523 , \Reg_Bank/n4522 , \Reg_Bank/n4521 ,
         \Reg_Bank/n4520 , \Reg_Bank/n4519 , \Reg_Bank/n4518 ,
         \Reg_Bank/n4517 , \Reg_Bank/n4516 , \Reg_Bank/n4515 ,
         \Reg_Bank/n4514 , \Reg_Bank/n4513 , \Reg_Bank/n4512 ,
         \Reg_Bank/n4511 , \Reg_Bank/n4510 , \Reg_Bank/n4509 ,
         \Reg_Bank/n4508 , \Reg_Bank/n4507 , \Reg_Bank/n4506 ,
         \Reg_Bank/n4505 , \Reg_Bank/n4504 , \Reg_Bank/n4503 ,
         \Reg_Bank/n4502 , \Reg_Bank/n4501 , \Reg_Bank/n4500 ,
         \Reg_Bank/n4499 , \Reg_Bank/n4498 , \Reg_Bank/n4497 ,
         \Reg_Bank/n4496 , \Reg_Bank/n4495 , \Reg_Bank/n4494 ,
         \Reg_Bank/n4493 , \Reg_Bank/n4492 , \Reg_Bank/n4491 ,
         \Reg_Bank/n4490 , \Reg_Bank/n4489 , \Reg_Bank/n4488 ,
         \Reg_Bank/n4487 , \Reg_Bank/n4486 , \Reg_Bank/n4485 ,
         \Reg_Bank/n4484 , \Reg_Bank/n4483 , \Reg_Bank/n4482 ,
         \Reg_Bank/n4481 , \Reg_Bank/n4480 , \Reg_Bank/n4479 ,
         \Reg_Bank/n4478 , \Reg_Bank/n4477 , \Reg_Bank/n4476 ,
         \Reg_Bank/n4475 , \Reg_Bank/n4474 , \Reg_Bank/n4473 ,
         \Reg_Bank/n4472 , \Reg_Bank/n4471 , \Reg_Bank/n4470 ,
         \Reg_Bank/n4469 , \Reg_Bank/n4468 , \Reg_Bank/n4467 ,
         \Reg_Bank/n4466 , \Reg_Bank/n4465 , \Reg_Bank/n4464 ,
         \Reg_Bank/n4463 , \Reg_Bank/n4462 , \Reg_Bank/n4461 ,
         \Reg_Bank/n4460 , \Reg_Bank/n4459 , \Reg_Bank/n4458 ,
         \Reg_Bank/n4457 , \Reg_Bank/n4456 , \Reg_Bank/n4455 ,
         \Reg_Bank/n4454 , \Reg_Bank/n4453 , \Reg_Bank/n4452 ,
         \Reg_Bank/n4451 , \Reg_Bank/n4450 , \Reg_Bank/n4449 ,
         \Reg_Bank/n4448 , \Reg_Bank/n4447 , \Reg_Bank/n4446 ,
         \Reg_Bank/n4445 , \Reg_Bank/n4444 , \Reg_Bank/n4443 ,
         \Reg_Bank/n4442 , \Reg_Bank/n4441 , \Reg_Bank/n4440 ,
         \Reg_Bank/n4439 , \Reg_Bank/n4438 , \Reg_Bank/n4437 ,
         \Reg_Bank/n4436 , \Reg_Bank/n4435 , \Reg_Bank/n4434 ,
         \Reg_Bank/n4433 , \Reg_Bank/n4432 , \Reg_Bank/n4431 ,
         \Reg_Bank/n4430 , \Reg_Bank/n4429 , \Reg_Bank/n4428 ,
         \Reg_Bank/n4427 , \Reg_Bank/n4426 , \Reg_Bank/n4425 ,
         \Reg_Bank/n4424 , \Reg_Bank/n4423 , \Reg_Bank/n4422 ,
         \Reg_Bank/n4421 , \Reg_Bank/n4420 , \Reg_Bank/n4419 ,
         \Reg_Bank/n4418 , \Reg_Bank/n4417 , \Reg_Bank/n4416 ,
         \Reg_Bank/n4415 , \Reg_Bank/n4414 , \Reg_Bank/n4413 ,
         \Reg_Bank/n4412 , \Reg_Bank/n4411 , \Reg_Bank/n4410 ,
         \Reg_Bank/n4409 , \Reg_Bank/n4408 , \Reg_Bank/n4407 ,
         \Reg_Bank/n4406 , \Reg_Bank/n4405 , \Reg_Bank/n4404 ,
         \Reg_Bank/n4403 , \Reg_Bank/n4402 , \Reg_Bank/n4401 ,
         \Reg_Bank/n4400 , \Reg_Bank/n4399 , \Reg_Bank/n4398 ,
         \Reg_Bank/n4397 , \Reg_Bank/n4396 , \Reg_Bank/n4395 ,
         \Reg_Bank/n4394 , \Reg_Bank/n4393 , \Reg_Bank/n4392 ,
         \Reg_Bank/n4391 , \Reg_Bank/n4390 , \Reg_Bank/n4389 ,
         \Reg_Bank/n4388 , \Reg_Bank/n4387 , \Reg_Bank/n4386 ,
         \Reg_Bank/n4385 , \Reg_Bank/n4384 , \Reg_Bank/n4383 ,
         \Reg_Bank/n4382 , \Reg_Bank/n4381 , \Reg_Bank/n4380 ,
         \Reg_Bank/n4379 , \Reg_Bank/n4378 , \Reg_Bank/n4377 ,
         \Reg_Bank/n4376 , \Reg_Bank/n4375 , \Reg_Bank/n4374 ,
         \Reg_Bank/n4373 , \Reg_Bank/n4372 , \Reg_Bank/n4371 ,
         \Reg_Bank/n4370 , \Reg_Bank/n4369 , \Reg_Bank/n4368 ,
         \Reg_Bank/n4367 , \Reg_Bank/n4366 , \Reg_Bank/n4365 ,
         \Reg_Bank/n4364 , \Reg_Bank/n4363 , \Reg_Bank/n4362 ,
         \Reg_Bank/n4361 , \Reg_Bank/n4360 , \Reg_Bank/n4359 ,
         \Reg_Bank/n4358 , \Reg_Bank/n4357 , \Reg_Bank/n4356 ,
         \Reg_Bank/n4355 , \Reg_Bank/n4354 , \Reg_Bank/n4353 ,
         \Reg_Bank/n4352 , \Reg_Bank/n4351 , \Reg_Bank/n4350 ,
         \Reg_Bank/n4349 , \Reg_Bank/n4348 , \Reg_Bank/n4347 ,
         \Reg_Bank/n4346 , \Reg_Bank/n4345 , \Reg_Bank/n4344 ,
         \Reg_Bank/n4343 , \Reg_Bank/n4342 , \Reg_Bank/n4341 ,
         \Reg_Bank/n4340 , \Reg_Bank/n4339 , \Reg_Bank/n4338 ,
         \Reg_Bank/n4337 , \Reg_Bank/n4336 , \Reg_Bank/n4335 ,
         \Reg_Bank/n4334 , \Reg_Bank/n4333 , \Reg_Bank/n4332 ,
         \Reg_Bank/n4331 , \Reg_Bank/n4330 , \Reg_Bank/n4329 ,
         \Reg_Bank/n4328 , \Reg_Bank/n4327 , \Reg_Bank/n4326 ,
         \Reg_Bank/n4325 , \Reg_Bank/n4324 , \Reg_Bank/n4323 ,
         \Reg_Bank/n4322 , \Reg_Bank/n4321 , \Reg_Bank/n4320 ,
         \Reg_Bank/n4319 , \Reg_Bank/n4318 , \Reg_Bank/n4317 ,
         \Reg_Bank/n4316 , \Reg_Bank/n4315 , \Reg_Bank/n4314 ,
         \Reg_Bank/n4313 , \Reg_Bank/n4312 , \Reg_Bank/n4311 ,
         \Reg_Bank/n4310 , \Reg_Bank/n4309 , \Reg_Bank/n4308 ,
         \Reg_Bank/n4307 , \Reg_Bank/n4306 , \Reg_Bank/n4305 ,
         \Reg_Bank/n4304 , \Reg_Bank/n4303 , \Reg_Bank/n4302 ,
         \Reg_Bank/n4301 , \Reg_Bank/n4300 , \Reg_Bank/n4299 ,
         \Reg_Bank/n4298 , \Reg_Bank/n4297 , \Reg_Bank/n4296 ,
         \Reg_Bank/n4295 , \Reg_Bank/n4294 , \Reg_Bank/n4293 ,
         \Reg_Bank/n4292 , \Reg_Bank/n4291 , \Reg_Bank/n4290 ,
         \Reg_Bank/n4289 , \Reg_Bank/n4288 , \Reg_Bank/n4287 ,
         \Reg_Bank/n4286 , \Reg_Bank/n4285 , \Reg_Bank/n4284 ,
         \Reg_Bank/n4283 , \Reg_Bank/n4282 , \Reg_Bank/n4281 ,
         \Reg_Bank/n4280 , \Reg_Bank/n4279 , \Reg_Bank/n4278 ,
         \Reg_Bank/n4277 , \Reg_Bank/n4276 , \Reg_Bank/n4275 ,
         \Reg_Bank/n4274 , \Reg_Bank/n4273 , \Reg_Bank/n4272 ,
         \Reg_Bank/n4271 , \Reg_Bank/n4270 , \Reg_Bank/n4269 ,
         \Reg_Bank/n4268 , \Reg_Bank/n4267 , \Reg_Bank/n4266 ,
         \Reg_Bank/n4265 , \Reg_Bank/n4264 , \Reg_Bank/n4263 ,
         \Reg_Bank/n4262 , \Reg_Bank/n4261 , \Reg_Bank/n4260 ,
         \Reg_Bank/n4259 , \Reg_Bank/n4258 , \Reg_Bank/n4257 ,
         \Reg_Bank/n4256 , \Reg_Bank/n4255 , \Reg_Bank/n4254 ,
         \Reg_Bank/n4253 , \Reg_Bank/n4252 , \Reg_Bank/n4251 ,
         \Reg_Bank/n4250 , \Reg_Bank/n4249 , \Reg_Bank/n4248 ,
         \Reg_Bank/n4247 , \Reg_Bank/n4246 , \Reg_Bank/n4245 ,
         \Reg_Bank/n4244 , \Reg_Bank/n4243 , \Reg_Bank/n4242 ,
         \Reg_Bank/n4241 , \Reg_Bank/n4240 , \Reg_Bank/n4239 ,
         \Reg_Bank/n4238 , \Reg_Bank/n4237 , \Reg_Bank/n4236 ,
         \Reg_Bank/n4235 , \Reg_Bank/n4234 , \Reg_Bank/n4233 ,
         \Reg_Bank/n4232 , \Reg_Bank/n4231 , \Reg_Bank/n4230 ,
         \Reg_Bank/n4229 , \Reg_Bank/n4228 , \Reg_Bank/n4227 ,
         \Reg_Bank/n4226 , \Reg_Bank/n4225 , \Reg_Bank/n4224 ,
         \Reg_Bank/n4223 , \Reg_Bank/n4222 , \Reg_Bank/n4221 ,
         \Reg_Bank/n4220 , \Reg_Bank/n4219 , \Reg_Bank/n4218 ,
         \Reg_Bank/n4217 , \Reg_Bank/n4216 , \Reg_Bank/n4215 ,
         \Reg_Bank/n4214 , \Reg_Bank/n4213 , \Reg_Bank/n4212 ,
         \Reg_Bank/n4211 , \Reg_Bank/n4210 , \Reg_Bank/n4209 ,
         \Reg_Bank/n4208 , \Reg_Bank/n4207 , \Reg_Bank/n4206 ,
         \Reg_Bank/n4205 , \Reg_Bank/n4204 , \Reg_Bank/n4203 ,
         \Reg_Bank/n4202 , \Reg_Bank/n4201 , \Reg_Bank/n4200 ,
         \Reg_Bank/n4199 , \Reg_Bank/n4198 , \Reg_Bank/n4197 ,
         \Reg_Bank/n4196 , \Reg_Bank/n4195 , \Reg_Bank/n4194 ,
         \Reg_Bank/n4193 , \Reg_Bank/n4192 , \Reg_Bank/n4191 ,
         \Reg_Bank/n4190 , \Reg_Bank/n4189 , \Reg_Bank/n4188 ,
         \Reg_Bank/n4187 , \Reg_Bank/n4186 , \Reg_Bank/n4185 ,
         \Reg_Bank/n4184 , \Reg_Bank/n4183 , \Reg_Bank/n4182 ,
         \Reg_Bank/n4181 , \Reg_Bank/n4180 , \Reg_Bank/n4179 ,
         \Reg_Bank/n4178 , \Reg_Bank/n4177 , \Reg_Bank/n4176 ,
         \Reg_Bank/n4175 , \Reg_Bank/n4174 , \Reg_Bank/n4173 ,
         \Reg_Bank/n4172 , \Reg_Bank/n4171 , \Reg_Bank/n4170 ,
         \Reg_Bank/n4169 , \Reg_Bank/n4168 , \Reg_Bank/n4167 ,
         \Reg_Bank/n4166 , \Reg_Bank/n4165 , \Reg_Bank/n4164 ,
         \Reg_Bank/n4163 , \Reg_Bank/n4162 , \Reg_Bank/n4161 ,
         \Reg_Bank/n4160 , \Reg_Bank/n4159 , \Reg_Bank/n4158 ,
         \Reg_Bank/n4157 , \Reg_Bank/n4156 , \Reg_Bank/n4155 ,
         \Reg_Bank/n4154 , \Reg_Bank/n4153 , \Reg_Bank/n4152 ,
         \Reg_Bank/n4151 , \Reg_Bank/n4150 , \Reg_Bank/n4149 ,
         \Reg_Bank/n4148 , \Reg_Bank/n4147 , \Reg_Bank/n4146 ,
         \Reg_Bank/n4145 , \Reg_Bank/n4144 , \Reg_Bank/n4143 ,
         \Reg_Bank/n4142 , \Reg_Bank/n4141 , \Reg_Bank/n4140 ,
         \Reg_Bank/n4139 , \Reg_Bank/n4138 , \Reg_Bank/n4137 ,
         \Reg_Bank/n4136 , \Reg_Bank/n4135 , \Reg_Bank/n4134 ,
         \Reg_Bank/n4133 , \Reg_Bank/n4132 , \Reg_Bank/n4131 ,
         \Reg_Bank/n4130 , \Reg_Bank/n4129 , \Reg_Bank/n4128 ,
         \Reg_Bank/n4127 , \Reg_Bank/n4126 , \Reg_Bank/n4125 ,
         \Reg_Bank/n4124 , \Reg_Bank/n4123 , \Reg_Bank/n4122 ,
         \Reg_Bank/n4121 , \Reg_Bank/n4120 , \Reg_Bank/n4119 ,
         \Reg_Bank/n4118 , \Reg_Bank/n4117 , \Reg_Bank/n4116 ,
         \Reg_Bank/n4115 , \Reg_Bank/n4114 , \Reg_Bank/n4113 ,
         \Reg_Bank/n4112 , \Reg_Bank/n4111 , \Reg_Bank/n4110 ,
         \Reg_Bank/n4109 , \Reg_Bank/n4108 , \Reg_Bank/n4107 ,
         \Reg_Bank/n4106 , \Reg_Bank/n4105 , \Reg_Bank/n4104 ,
         \Reg_Bank/n4103 , \Reg_Bank/n4102 , \Reg_Bank/n4101 ,
         \Reg_Bank/n4100 , \Reg_Bank/n4099 , \Reg_Bank/n4098 ,
         \Reg_Bank/n4097 , \Reg_Bank/n4096 , \Reg_Bank/n4095 ,
         \Reg_Bank/n4094 , \Reg_Bank/n4093 , \Reg_Bank/n4092 ,
         \Reg_Bank/n4091 , \Reg_Bank/n4090 , \Reg_Bank/n4089 ,
         \Reg_Bank/n4088 , \Reg_Bank/n4087 , \Reg_Bank/n4086 ,
         \Reg_Bank/n4085 , \Reg_Bank/n4084 , \Reg_Bank/n4083 ,
         \Reg_Bank/n4082 , \Reg_Bank/n4081 , \Reg_Bank/n4080 ,
         \Reg_Bank/n4079 , \Reg_Bank/n4078 , \Reg_Bank/n4077 ,
         \Reg_Bank/n4076 , \Reg_Bank/n4075 , \Reg_Bank/n4074 ,
         \Reg_Bank/n4073 , \Reg_Bank/n4072 , \Reg_Bank/n4071 ,
         \Reg_Bank/n4070 , \Reg_Bank/n4069 , \Reg_Bank/n4068 ,
         \Reg_Bank/n4067 , \Reg_Bank/n4066 , \Reg_Bank/n4065 ,
         \Reg_Bank/n4064 , \Reg_Bank/n4063 , \Reg_Bank/n4062 ,
         \Reg_Bank/n4061 , \Reg_Bank/n4060 , \Reg_Bank/n4059 ,
         \Reg_Bank/n4058 , \Reg_Bank/n4057 , \Reg_Bank/n4056 ,
         \Reg_Bank/n4055 , \Reg_Bank/n4054 , \Reg_Bank/n4053 ,
         \Reg_Bank/n4052 , \Reg_Bank/n4051 , \Reg_Bank/n4050 ,
         \Reg_Bank/n4049 , \Reg_Bank/n4048 , \Reg_Bank/n4047 ,
         \Reg_Bank/n4046 , \Reg_Bank/n4045 , \Reg_Bank/n4044 ,
         \Reg_Bank/n4043 , \Reg_Bank/n4042 , \Reg_Bank/n4041 ,
         \Reg_Bank/n4040 , \Reg_Bank/n4039 , \Reg_Bank/n4038 ,
         \Reg_Bank/n4037 , \Reg_Bank/n4036 , \Reg_Bank/n4035 ,
         \Reg_Bank/n4034 , \Reg_Bank/n4033 , \Reg_Bank/n4032 ,
         \Reg_Bank/n4031 , \Reg_Bank/n4030 , \Reg_Bank/n4029 ,
         \Reg_Bank/n4028 , \Reg_Bank/n4027 , \Reg_Bank/n4026 ,
         \Reg_Bank/n4025 , \Reg_Bank/n4024 , \Reg_Bank/n4023 ,
         \Reg_Bank/n4022 , \Reg_Bank/n4021 , \Reg_Bank/n4020 ,
         \Reg_Bank/n4019 , \Reg_Bank/n4018 , \Reg_Bank/n4017 ,
         \Reg_Bank/n4016 , \Reg_Bank/n4015 , \Reg_Bank/n4014 ,
         \Reg_Bank/n4013 , \Reg_Bank/n4012 , \Reg_Bank/n4011 ,
         \Reg_Bank/n4010 , \Reg_Bank/n4009 , \Reg_Bank/n4008 ,
         \Reg_Bank/n4007 , \Reg_Bank/n4006 , \Reg_Bank/n4005 ,
         \Reg_Bank/n4004 , \Reg_Bank/n4003 , \Reg_Bank/n4002 ,
         \Reg_Bank/n4001 , \Reg_Bank/n4000 , \Reg_Bank/n3999 ,
         \Reg_Bank/n3998 , \Reg_Bank/n3997 , \Reg_Bank/n3996 ,
         \Reg_Bank/n3995 , \Reg_Bank/n3994 , \Reg_Bank/n3993 ,
         \Reg_Bank/n3992 , \Reg_Bank/n3991 , \Reg_Bank/n3990 ,
         \Reg_Bank/n3989 , \Reg_Bank/n3988 , \Reg_Bank/n3987 ,
         \Reg_Bank/n3986 , \Reg_Bank/n3985 , \Reg_Bank/n3984 ,
         \Reg_Bank/n3983 , \Reg_Bank/n3982 , \Reg_Bank/n3981 ,
         \Reg_Bank/n3980 , \Reg_Bank/n3979 , \Reg_Bank/n3978 ,
         \Reg_Bank/n3977 , \Reg_Bank/n3976 , \Reg_Bank/n3975 ,
         \Reg_Bank/n3974 , \Reg_Bank/n3973 , \Reg_Bank/n3972 ,
         \Reg_Bank/n3971 , \Reg_Bank/n3970 , \Reg_Bank/n3969 ,
         \Reg_Bank/n3968 , \Reg_Bank/n3967 , \Reg_Bank/n3966 ,
         \Reg_Bank/n3965 , \Reg_Bank/n3964 , \Reg_Bank/n3963 ,
         \Reg_Bank/n3962 , \Reg_Bank/n3961 , \Reg_Bank/n3960 ,
         \Reg_Bank/n3959 , \Reg_Bank/n3958 , \Reg_Bank/n3957 ,
         \Reg_Bank/n3956 , \Reg_Bank/n3955 , \Reg_Bank/n3954 ,
         \Reg_Bank/n3953 , \Reg_Bank/n3952 , \Reg_Bank/n3951 ,
         \Reg_Bank/n3950 , \Reg_Bank/n3949 , \Reg_Bank/n3948 ,
         \Reg_Bank/n3947 , \Reg_Bank/n3946 , \Reg_Bank/n3945 ,
         \Reg_Bank/n3944 , \Reg_Bank/n3943 , \Reg_Bank/n3942 ,
         \Reg_Bank/n3941 , \Reg_Bank/n3940 , \Reg_Bank/n3939 ,
         \Reg_Bank/n3938 , \Reg_Bank/n3937 , \Reg_Bank/n3936 ,
         \Reg_Bank/n3935 , \Reg_Bank/n3934 , \Reg_Bank/n3933 ,
         \Reg_Bank/n3932 , \Reg_Bank/n3931 , \Reg_Bank/n3930 ,
         \Reg_Bank/n3929 , \Reg_Bank/n3928 , \Reg_Bank/n3927 ,
         \Reg_Bank/n3926 , \Reg_Bank/n3925 , \Reg_Bank/n3924 ,
         \Reg_Bank/n3923 , \Reg_Bank/n3922 , \Reg_Bank/n3921 ,
         \Reg_Bank/n3920 , \Reg_Bank/n3919 , \Reg_Bank/n3918 ,
         \Reg_Bank/n3917 , \Reg_Bank/n3916 , \Reg_Bank/n3915 ,
         \Reg_Bank/n3914 , \Reg_Bank/n3913 , \Reg_Bank/n3912 ,
         \Reg_Bank/n3911 , \Reg_Bank/n3910 , \Reg_Bank/n3909 ,
         \Reg_Bank/n3908 , \Reg_Bank/n3907 , \Reg_Bank/n3906 ,
         \Reg_Bank/n3905 , \Reg_Bank/n3904 , \Reg_Bank/n3903 ,
         \Reg_Bank/n3902 , \Reg_Bank/n3901 , \Reg_Bank/n3900 ,
         \Reg_Bank/n3899 , \Reg_Bank/n3898 , \Reg_Bank/n3897 ,
         \Reg_Bank/n3896 , \Reg_Bank/n3895 , \Reg_Bank/n3894 ,
         \Reg_Bank/n3893 , \Reg_Bank/n3892 , \Reg_Bank/n3891 ,
         \Reg_Bank/n3890 , \Reg_Bank/n3889 , \Reg_Bank/n3888 ,
         \Reg_Bank/n3887 , \Reg_Bank/n3886 , \Reg_Bank/n3885 ,
         \Reg_Bank/n3884 , \Reg_Bank/n3883 , \Reg_Bank/n3882 ,
         \Reg_Bank/n3881 , \Reg_Bank/n3880 , \Reg_Bank/n3879 ,
         \Reg_Bank/n3878 , \Reg_Bank/n3877 , \Reg_Bank/n3876 ,
         \Reg_Bank/n3875 , \Reg_Bank/n3874 , \Reg_Bank/n3873 ,
         \Reg_Bank/n3872 , \Reg_Bank/n3871 , \Reg_Bank/n3870 ,
         \Reg_Bank/n3869 , \Reg_Bank/n3868 , \Reg_Bank/n3867 ,
         \Reg_Bank/n3866 , \Reg_Bank/n3865 , \Reg_Bank/n3864 ,
         \Reg_Bank/n3863 , \Reg_Bank/n3862 , \Reg_Bank/n3861 ,
         \Reg_Bank/n3860 , \Reg_Bank/n3859 , \Reg_Bank/n3858 ,
         \Reg_Bank/n3857 , \Reg_Bank/n3856 , \Reg_Bank/n3855 ,
         \Reg_Bank/n3854 , \Reg_Bank/n3853 , \Reg_Bank/n3852 ,
         \Reg_Bank/n3851 , \Reg_Bank/n3850 , \Reg_Bank/n3849 ,
         \Reg_Bank/n3848 , \Reg_Bank/n3847 , \Reg_Bank/n3846 ,
         \Reg_Bank/n3845 , \Reg_Bank/n3844 , \Reg_Bank/n3843 ,
         \Reg_Bank/n3842 , \Reg_Bank/n3841 , \Reg_Bank/n3840 ,
         \Reg_Bank/n3839 , \Reg_Bank/n3838 , \Reg_Bank/n3837 ,
         \Reg_Bank/n3836 , \Reg_Bank/n3835 , \Reg_Bank/n3834 ,
         \Reg_Bank/n3833 , \Reg_Bank/n3832 , \Reg_Bank/n3831 ,
         \Reg_Bank/n3830 , \Reg_Bank/n3829 , \Reg_Bank/n3828 ,
         \Reg_Bank/n3827 , \Reg_Bank/n3826 , \Reg_Bank/n3825 ,
         \Reg_Bank/n3824 , \Reg_Bank/n3823 , \Reg_Bank/n3822 ,
         \Reg_Bank/n3821 , \Reg_Bank/n3820 , \Reg_Bank/n3819 ,
         \Reg_Bank/n3818 , \Reg_Bank/n3817 , \Reg_Bank/n3816 ,
         \Reg_Bank/n3815 , \Reg_Bank/n3814 , \Reg_Bank/n3813 ,
         \Reg_Bank/n3812 , \Reg_Bank/n3811 , \Reg_Bank/n3810 ,
         \Reg_Bank/n3809 , \Reg_Bank/n3808 , \Reg_Bank/n3807 ,
         \Reg_Bank/n3806 , \Reg_Bank/n3805 , \Reg_Bank/n3804 ,
         \Reg_Bank/n3803 , \Reg_Bank/n3802 , \Reg_Bank/n3801 ,
         \Reg_Bank/n3800 , \Reg_Bank/n3799 , \Reg_Bank/n3798 ,
         \Reg_Bank/n3797 , \Reg_Bank/n3796 , \Reg_Bank/n3795 ,
         \Reg_Bank/n3794 , \Reg_Bank/n3793 , \Reg_Bank/n3792 ,
         \Reg_Bank/n3791 , \Reg_Bank/n3790 , \Reg_Bank/n3789 ,
         \Reg_Bank/n3788 , \Reg_Bank/n3787 , \Reg_Bank/n3786 ,
         \Reg_Bank/n3785 , \Reg_Bank/n3784 , \Reg_Bank/n3783 ,
         \Reg_Bank/n3782 , \Reg_Bank/n3781 , \Reg_Bank/n3780 ,
         \Reg_Bank/n3779 , \Reg_Bank/n3778 , \Reg_Bank/n3777 ,
         \Reg_Bank/n3776 , \Reg_Bank/n3775 , \Reg_Bank/n3774 ,
         \Reg_Bank/n3773 , \Reg_Bank/n3772 , \Reg_Bank/n3771 ,
         \Reg_Bank/n3770 , \Reg_Bank/n3769 , \Reg_Bank/n3768 ,
         \Reg_Bank/n3767 , \Reg_Bank/n3766 , \Reg_Bank/n3765 ,
         \Reg_Bank/n3764 , \Reg_Bank/n3763 , \Reg_Bank/n3762 ,
         \Reg_Bank/n3761 , \Reg_Bank/n3760 , \Reg_Bank/n3759 ,
         \Reg_Bank/n3758 , \Reg_Bank/n3757 , \Reg_Bank/n3756 ,
         \Reg_Bank/n3755 , \Reg_Bank/n3754 , \Reg_Bank/n3753 ,
         \Reg_Bank/n3752 , \Reg_Bank/n3751 , \Reg_Bank/n3750 ,
         \Reg_Bank/n3749 , \Reg_Bank/n3748 , \Reg_Bank/n3747 ,
         \Reg_Bank/n3746 , \Reg_Bank/n3745 , \Reg_Bank/n3744 ,
         \Reg_Bank/n3743 , \Reg_Bank/n3742 , \Reg_Bank/n3741 ,
         \Reg_Bank/n3740 , \Reg_Bank/n3739 , \Reg_Bank/n3738 ,
         \Reg_Bank/n3737 , \Reg_Bank/n3736 , \Reg_Bank/n3735 ,
         \Reg_Bank/n3734 , \Reg_Bank/n3733 , \Reg_Bank/n3732 ,
         \Reg_Bank/n3731 , \Reg_Bank/n3730 , \Reg_Bank/n3729 ,
         \Reg_Bank/n3728 , \Reg_Bank/n3727 , \Reg_Bank/n3726 ,
         \Reg_Bank/n3725 , \Reg_Bank/n3724 , \Reg_Bank/n3723 ,
         \Reg_Bank/n3722 , \Reg_Bank/n3721 , \Reg_Bank/n3720 ,
         \Reg_Bank/n3719 , \Reg_Bank/n3718 , \Reg_Bank/n3717 ,
         \Reg_Bank/n3716 , \Reg_Bank/n3715 , \Reg_Bank/n3714 ,
         \Reg_Bank/n3713 , \Reg_Bank/n3712 , \Reg_Bank/n3711 ,
         \Reg_Bank/n3710 , \Reg_Bank/n3709 , \Reg_Bank/n3708 ,
         \Reg_Bank/n3707 , \Reg_Bank/n3706 , \Reg_Bank/n3705 ,
         \Reg_Bank/n3704 , \Reg_Bank/n3703 , \Reg_Bank/n3702 ,
         \Reg_Bank/n3701 , \Reg_Bank/n3700 , \Reg_Bank/n3699 ,
         \Reg_Bank/n3698 , \Reg_Bank/n3697 , \Reg_Bank/n3696 ,
         \Reg_Bank/n3695 , \Reg_Bank/n3694 , \Reg_Bank/n3693 ,
         \Reg_Bank/n3692 , \Reg_Bank/n3691 , \Reg_Bank/n3690 ,
         \Reg_Bank/n3689 , \Reg_Bank/n3688 , \Reg_Bank/n3687 ,
         \Reg_Bank/n3686 , \Reg_Bank/n3685 , \Reg_Bank/n3684 ,
         \Reg_Bank/n3683 , \Reg_Bank/n3682 , \Reg_Bank/n3681 ,
         \Reg_Bank/n3680 , \Reg_Bank/n3679 , \Reg_Bank/n3678 ,
         \Reg_Bank/n3677 , \Reg_Bank/n3676 , \Reg_Bank/n3675 ,
         \Reg_Bank/n3674 , \Reg_Bank/n3673 , \Reg_Bank/n3672 ,
         \Reg_Bank/n3671 , \Reg_Bank/n3670 , \Reg_Bank/n3669 ,
         \Reg_Bank/n3668 , \Reg_Bank/n3667 , \Reg_Bank/n3666 ,
         \Reg_Bank/n3665 , \Reg_Bank/n3664 , \Reg_Bank/n3663 ,
         \Reg_Bank/n3662 , \Reg_Bank/n3661 , \Reg_Bank/n3660 ,
         \Reg_Bank/n3659 , \Reg_Bank/n3658 , \Reg_Bank/n3657 ,
         \Reg_Bank/n3656 , \Reg_Bank/n3655 , \Reg_Bank/n3654 ,
         \Reg_Bank/n3653 , \Reg_Bank/n3652 , \Reg_Bank/n3651 ,
         \Reg_Bank/n3650 , \Reg_Bank/n3649 , \Reg_Bank/n3648 ,
         \Reg_Bank/n3647 , \Reg_Bank/n3646 , \Reg_Bank/n3645 ,
         \Reg_Bank/n3644 , \Reg_Bank/n3643 , \Reg_Bank/n3642 ,
         \Reg_Bank/n3641 , \Reg_Bank/n3640 , \Reg_Bank/n3639 ,
         \Reg_Bank/n3638 , \Reg_Bank/n3637 , \Reg_Bank/n3636 ,
         \Reg_Bank/n3635 , \Reg_Bank/n3634 , \Reg_Bank/n3633 ,
         \Reg_Bank/n3632 , \Reg_Bank/n3631 , \Reg_Bank/n3630 ,
         \Reg_Bank/n3629 , \Reg_Bank/n3628 , \Reg_Bank/n3627 ,
         \Reg_Bank/n3626 , \Reg_Bank/n3625 , \Reg_Bank/n3624 ,
         \Reg_Bank/n3623 , \Reg_Bank/n3622 , \Reg_Bank/n3621 ,
         \Reg_Bank/n3620 , \Reg_Bank/n3619 , \Reg_Bank/n3618 ,
         \Reg_Bank/n3617 , \Reg_Bank/n3616 , \Reg_Bank/n3615 ,
         \Reg_Bank/n3614 , \Reg_Bank/n3613 , \Reg_Bank/n3612 ,
         \Reg_Bank/n3611 , \Reg_Bank/n3610 , \Reg_Bank/n3609 ,
         \Reg_Bank/n3608 , \Reg_Bank/n3607 , \Reg_Bank/n3606 ,
         \Reg_Bank/n3605 , \Reg_Bank/n3604 , \Reg_Bank/n3603 ,
         \Reg_Bank/n3602 , \Reg_Bank/n3601 , \Reg_Bank/n3600 ,
         \Reg_Bank/n3599 , \Reg_Bank/n3598 , \Reg_Bank/n3597 ,
         \Reg_Bank/n3596 , \Reg_Bank/n3595 , \Reg_Bank/n3594 ,
         \Reg_Bank/n3593 , \Reg_Bank/n3592 , \Reg_Bank/n3591 ,
         \Reg_Bank/n3590 , \Reg_Bank/n3589 , \Reg_Bank/n3588 ,
         \Reg_Bank/n3587 , \Reg_Bank/n3586 , \Reg_Bank/n3585 ,
         \Reg_Bank/n3584 , \Reg_Bank/n3583 , \Reg_Bank/n3582 ,
         \Reg_Bank/n3581 , \Reg_Bank/n3580 , \Reg_Bank/n3579 ,
         \Reg_Bank/n3578 , \Reg_Bank/n3577 , \Reg_Bank/n3576 ,
         \Reg_Bank/n3575 , \Reg_Bank/n3574 , \Reg_Bank/n3573 ,
         \Reg_Bank/n3572 , \Reg_Bank/n3571 , \Reg_Bank/n3570 ,
         \Reg_Bank/n3569 , \Reg_Bank/n3568 , \Reg_Bank/n3567 ,
         \Reg_Bank/n3566 , \Reg_Bank/n3565 , \Reg_Bank/n3564 ,
         \Reg_Bank/n3563 , \Reg_Bank/n3562 , \Reg_Bank/n3561 ,
         \Reg_Bank/n3560 , \Reg_Bank/n3559 , \Reg_Bank/n3558 ,
         \Reg_Bank/n3557 , \Reg_Bank/n3556 , \Reg_Bank/n3555 ,
         \Reg_Bank/n3554 , \Reg_Bank/n3553 , \Reg_Bank/n3552 ,
         \Reg_Bank/n3551 , \Reg_Bank/n3550 , \Reg_Bank/n3549 ,
         \Reg_Bank/n3548 , \Reg_Bank/n3547 , \Reg_Bank/n3546 ,
         \Reg_Bank/n3545 , \Reg_Bank/n3544 , \Reg_Bank/n3543 ,
         \Reg_Bank/n3542 , \Reg_Bank/n3541 , \Reg_Bank/n3540 ,
         \Reg_Bank/n3539 , \Reg_Bank/n3538 , \Reg_Bank/n3537 ,
         \Reg_Bank/n3536 , \Reg_Bank/n3535 , \Reg_Bank/n3534 ,
         \Reg_Bank/n3533 , \Reg_Bank/n3532 , \Reg_Bank/n3531 ,
         \Reg_Bank/n3530 , \Reg_Bank/n3529 , \Reg_Bank/n3528 ,
         \Reg_Bank/n3527 , \Reg_Bank/n3526 , \Reg_Bank/n3525 ,
         \Reg_Bank/n3524 , \Reg_Bank/n3523 , \Reg_Bank/n3522 ,
         \Reg_Bank/n3521 , \Reg_Bank/n3520 , \Reg_Bank/n3519 ,
         \Reg_Bank/n3518 , \Reg_Bank/n3517 , \Reg_Bank/n3516 ,
         \Reg_Bank/n3515 , \Reg_Bank/n3514 , \Reg_Bank/n3513 ,
         \Reg_Bank/n3512 , \Reg_Bank/n3511 , \Reg_Bank/n3510 ,
         \Reg_Bank/n3509 , \Reg_Bank/n3508 , \Reg_Bank/n3507 ,
         \Reg_Bank/n3506 , \Reg_Bank/n3505 , \Reg_Bank/n3504 ,
         \Reg_Bank/n3503 , \Reg_Bank/n3502 , \Reg_Bank/n3501 ,
         \Reg_Bank/n3500 , \Reg_Bank/n3499 , \Reg_Bank/n3498 ,
         \Reg_Bank/n3497 , \Reg_Bank/n3496 , \Reg_Bank/n3495 ,
         \Reg_Bank/n3494 , \Reg_Bank/n3493 , \Reg_Bank/n3492 ,
         \Reg_Bank/n3491 , \Reg_Bank/n3490 , \Reg_Bank/n3489 ,
         \Reg_Bank/n3488 , \Reg_Bank/n3487 , \Reg_Bank/n3486 ,
         \Reg_Bank/n3485 , \Reg_Bank/n3484 , \Reg_Bank/n3483 ,
         \Reg_Bank/n3482 , \Reg_Bank/n3481 , \Reg_Bank/n3480 ,
         \Reg_Bank/n3479 , \Reg_Bank/n3478 , \Reg_Bank/n3477 ,
         \Reg_Bank/n3476 , \Reg_Bank/n3475 , \Reg_Bank/n3474 ,
         \Reg_Bank/n3473 , \Reg_Bank/n3472 , \Reg_Bank/n3471 ,
         \Reg_Bank/n3470 , \Reg_Bank/n3469 , \Reg_Bank/n3468 ,
         \Reg_Bank/n3467 , \Reg_Bank/n3466 , \Reg_Bank/n3465 ,
         \Reg_Bank/n3464 , \Reg_Bank/n3463 , \Reg_Bank/n3462 ,
         \Reg_Bank/n3461 , \Reg_Bank/n3460 , \Reg_Bank/n3459 ,
         \Reg_Bank/n3458 , \Reg_Bank/n3457 , \Reg_Bank/n3456 ,
         \Reg_Bank/n3455 , \Reg_Bank/n3454 , \Reg_Bank/n3453 ,
         \Reg_Bank/n3452 , \Reg_Bank/n3451 , \Reg_Bank/n3450 ,
         \Reg_Bank/n3449 , \Reg_Bank/n3448 , \Reg_Bank/n3447 ,
         \Reg_Bank/n3446 , \Reg_Bank/n3445 , \Reg_Bank/n3444 ,
         \Reg_Bank/n3443 , \Reg_Bank/n3442 , \Reg_Bank/n3441 ,
         \Reg_Bank/n3440 , \Reg_Bank/n3439 , \Reg_Bank/n3438 ,
         \Reg_Bank/n3437 , \Reg_Bank/n3436 , \Reg_Bank/n3435 ,
         \Reg_Bank/n3434 , \Reg_Bank/n3433 , \Reg_Bank/n3432 ,
         \Reg_Bank/n3431 , \Reg_Bank/n3430 , \Reg_Bank/n3429 ,
         \Reg_Bank/n3428 , \Reg_Bank/n3427 , \Reg_Bank/n3426 ,
         \Reg_Bank/n3425 , \Reg_Bank/n3424 , \Reg_Bank/n3423 ,
         \Reg_Bank/n3422 , \Reg_Bank/n3421 , \Reg_Bank/n3420 ,
         \Reg_Bank/n3419 , \Reg_Bank/n3418 , \Reg_Bank/n3417 ,
         \Reg_Bank/n3416 , \Reg_Bank/n3415 , \Reg_Bank/n3414 ,
         \Reg_Bank/n3413 , \Reg_Bank/n3412 , \Reg_Bank/n3411 ,
         \Reg_Bank/n3410 , \Reg_Bank/n3409 , \Reg_Bank/n3408 ,
         \Reg_Bank/n3407 , \Reg_Bank/n3406 , \Reg_Bank/n3405 ,
         \Reg_Bank/n3404 , \Reg_Bank/n3403 , \Reg_Bank/n3402 ,
         \Reg_Bank/n3401 , \Reg_Bank/n3400 , \Reg_Bank/n3399 ,
         \Reg_Bank/n3398 , \Reg_Bank/n3397 , \Reg_Bank/n3396 ,
         \Reg_Bank/n3395 , \Reg_Bank/n3394 , \Reg_Bank/n3393 ,
         \Reg_Bank/n3392 , \Reg_Bank/n3391 , \Reg_Bank/n3390 ,
         \Reg_Bank/n3389 , \Reg_Bank/n3388 , \Reg_Bank/n3387 ,
         \Reg_Bank/n3386 , \Reg_Bank/n3385 , \Reg_Bank/n3384 ,
         \Reg_Bank/n3383 , \Reg_Bank/n3382 , \Reg_Bank/n3381 ,
         \Reg_Bank/n3380 , \Reg_Bank/n3379 , \Reg_Bank/n3378 ,
         \Reg_Bank/n3377 , \Reg_Bank/n3376 , \Reg_Bank/n3375 ,
         \Reg_Bank/n3374 , \Reg_Bank/n3373 , \Reg_Bank/n3372 ,
         \Reg_Bank/n3371 , \Reg_Bank/n3370 , \Reg_Bank/n3369 ,
         \Reg_Bank/n3368 , \Reg_Bank/n3367 , \Reg_Bank/n3366 ,
         \Reg_Bank/n3365 , \Reg_Bank/n3364 , \Reg_Bank/n3363 ,
         \Reg_Bank/n3362 , \Reg_Bank/n3361 , \Reg_Bank/n3360 ,
         \Reg_Bank/n3359 , \Reg_Bank/n3358 , \Reg_Bank/n3357 ,
         \Reg_Bank/n3356 , \Reg_Bank/n3355 , \Reg_Bank/n3354 ,
         \Reg_Bank/n3353 , \Reg_Bank/n3352 , \Reg_Bank/n3351 ,
         \Reg_Bank/n3350 , \Reg_Bank/n3349 , \Reg_Bank/n3348 ,
         \Reg_Bank/n3347 , \Reg_Bank/n3346 , \Reg_Bank/n3345 ,
         \Reg_Bank/n3344 , \Reg_Bank/n3343 , \Reg_Bank/n3342 ,
         \Reg_Bank/n3341 , \Reg_Bank/n3340 , \Reg_Bank/n3339 ,
         \Reg_Bank/n3338 , \Reg_Bank/n3337 , \Reg_Bank/n3336 ,
         \Reg_Bank/n3335 , \Reg_Bank/n3334 , \Reg_Bank/n3333 ,
         \Reg_Bank/n3332 , \Reg_Bank/n3331 , \Reg_Bank/n3330 ,
         \Reg_Bank/n3329 , \Reg_Bank/n3328 , \Reg_Bank/n3327 ,
         \Reg_Bank/n3326 , \Reg_Bank/n3325 , \Reg_Bank/n3324 ,
         \Reg_Bank/n3323 , \Reg_Bank/n3322 , \Reg_Bank/n3321 ,
         \Reg_Bank/n3320 , \Reg_Bank/n3319 , \Reg_Bank/n3318 ,
         \Reg_Bank/n3317 , \Reg_Bank/n3316 , \Reg_Bank/n3315 ,
         \Reg_Bank/n3314 , \Reg_Bank/n3313 , \Reg_Bank/n3312 ,
         \Reg_Bank/n3311 , \Reg_Bank/n3310 , \Reg_Bank/n3309 ,
         \Reg_Bank/n3308 , \Reg_Bank/n3307 , \Reg_Bank/n3306 ,
         \Reg_Bank/n3305 , \Reg_Bank/n3304 , \Reg_Bank/n3303 ,
         \Reg_Bank/n3302 , \Reg_Bank/n3301 , \Reg_Bank/n3300 ,
         \Reg_Bank/n3299 , \Reg_Bank/n3298 , \Reg_Bank/n3297 ,
         \Reg_Bank/n3296 , \Reg_Bank/n3295 , \Reg_Bank/n3294 ,
         \Reg_Bank/n3293 , \Reg_Bank/n3292 , \Reg_Bank/n3291 ,
         \Reg_Bank/n3290 , \Reg_Bank/n3289 , \Reg_Bank/n3288 ,
         \Reg_Bank/n3287 , \Reg_Bank/n3286 , \Reg_Bank/n3285 ,
         \Reg_Bank/n3284 , \Reg_Bank/n3283 , \Reg_Bank/n3282 ,
         \Reg_Bank/n3281 , \Reg_Bank/n3280 , \Reg_Bank/n3279 ,
         \Reg_Bank/n3278 , \Reg_Bank/n3277 , \Reg_Bank/n3276 ,
         \Reg_Bank/n3275 , \Reg_Bank/n3274 , \Reg_Bank/n3273 ,
         \Reg_Bank/n3272 , \Reg_Bank/n3271 , \Reg_Bank/n3270 ,
         \Reg_Bank/n3269 , \Reg_Bank/n3268 , \Reg_Bank/n3267 ,
         \Reg_Bank/n3266 , \Reg_Bank/n3265 , \Reg_Bank/n3264 ,
         \Reg_Bank/n3263 , \Reg_Bank/n3262 , \Reg_Bank/n3261 ,
         \Reg_Bank/n3260 , \Reg_Bank/n3259 , \Reg_Bank/n3258 ,
         \Reg_Bank/n3257 , \Reg_Bank/n3256 , \Reg_Bank/n3255 ,
         \Reg_Bank/n3254 , \Reg_Bank/n3253 , \Reg_Bank/n3252 ,
         \Reg_Bank/n3251 , \Reg_Bank/n3250 , \Reg_Bank/n3249 ,
         \Reg_Bank/n3248 , \Reg_Bank/n3247 , \Reg_Bank/n3246 ,
         \Reg_Bank/n3245 , \Reg_Bank/n3244 , \Reg_Bank/n3243 ,
         \Reg_Bank/n3242 , \Reg_Bank/n3241 , \Reg_Bank/n3240 ,
         \Reg_Bank/n3239 , \Reg_Bank/n3238 , \Reg_Bank/n3237 ,
         \Reg_Bank/n3236 , \Reg_Bank/n3235 , \Reg_Bank/n3234 ,
         \Reg_Bank/n3233 , \Reg_Bank/n3232 , \Reg_Bank/n3231 ,
         \Reg_Bank/n3230 , \Reg_Bank/n3229 , \Reg_Bank/n3228 ,
         \Reg_Bank/n3227 , \Reg_Bank/n3226 , \Reg_Bank/n3225 ,
         \Reg_Bank/n3224 , \Reg_Bank/n3223 , \Reg_Bank/n3222 ,
         \Reg_Bank/n3221 , \Reg_Bank/n3220 , \Reg_Bank/n3219 ,
         \Reg_Bank/n3218 , \Reg_Bank/n3217 , \Reg_Bank/n3216 ,
         \Reg_Bank/n3215 , \Reg_Bank/n3214 , \Reg_Bank/n3213 ,
         \Reg_Bank/n3212 , \Reg_Bank/n3211 , \Reg_Bank/n3210 ,
         \Reg_Bank/n3209 , \Reg_Bank/n3208 , \Reg_Bank/n3207 ,
         \Reg_Bank/n3206 , \Reg_Bank/n3205 , \Reg_Bank/n3204 ,
         \Reg_Bank/n3203 , \Reg_Bank/n3202 , \Reg_Bank/n3201 ,
         \Reg_Bank/n3200 , \Reg_Bank/n3199 , \Reg_Bank/n3198 ,
         \Reg_Bank/n3197 , \Reg_Bank/n3196 , \Reg_Bank/n3195 ,
         \Reg_Bank/n3194 , \Reg_Bank/n3193 , \Reg_Bank/n3192 ,
         \Reg_Bank/n3191 , \Reg_Bank/n3190 , \Reg_Bank/n3189 ,
         \Reg_Bank/n3188 , \Reg_Bank/n3187 , \Reg_Bank/n3186 ,
         \Reg_Bank/n3185 , \Reg_Bank/n3184 , \Reg_Bank/n3183 ,
         \Reg_Bank/n3182 , \Reg_Bank/n3181 , \Reg_Bank/n3180 ,
         \Reg_Bank/n3179 , \Reg_Bank/n3178 , \Reg_Bank/n3177 ,
         \Reg_Bank/n3176 , \Reg_Bank/n3175 , \Reg_Bank/n3174 ,
         \Reg_Bank/n3173 , \Reg_Bank/n3172 , \Reg_Bank/n3171 ,
         \Reg_Bank/n3170 , \Reg_Bank/n3169 , \Reg_Bank/n3168 ,
         \Reg_Bank/n3167 , \Reg_Bank/n3166 , \Reg_Bank/n3165 ,
         \Reg_Bank/n3164 , \Reg_Bank/n3163 , \Reg_Bank/n3162 ,
         \Reg_Bank/n3161 , \Reg_Bank/n3160 , \Reg_Bank/n3159 ,
         \Reg_Bank/n3158 , \Reg_Bank/n3157 , \Reg_Bank/n3156 ,
         \Reg_Bank/n3155 , \Reg_Bank/n3154 , \Reg_Bank/n3153 ,
         \Reg_Bank/n3152 , \Reg_Bank/n3151 , \Reg_Bank/n3150 ,
         \Reg_Bank/n3149 , \Reg_Bank/n3148 , \Reg_Bank/n3147 ,
         \Reg_Bank/n3146 , \Reg_Bank/n3145 , \Reg_Bank/n3144 ,
         \Reg_Bank/n3143 , \Reg_Bank/n3142 , \Reg_Bank/n3141 ,
         \Reg_Bank/n3140 , \Reg_Bank/n3139 , \Reg_Bank/n3138 ,
         \Reg_Bank/n3137 , \Reg_Bank/n3136 , \Reg_Bank/n3135 ,
         \Reg_Bank/n3134 , \Reg_Bank/n3133 , \Reg_Bank/n3132 ,
         \Reg_Bank/n3131 , \Reg_Bank/n3130 , \Reg_Bank/n3129 ,
         \Reg_Bank/n3128 , \Reg_Bank/n3127 , \Reg_Bank/n3126 ,
         \Reg_Bank/n3125 , \Reg_Bank/n3124 , \Reg_Bank/n3123 ,
         \Reg_Bank/n3122 , \Reg_Bank/n3121 , \Reg_Bank/n3120 ,
         \Reg_Bank/n3119 , \Reg_Bank/n3118 , \Reg_Bank/n3117 ,
         \Reg_Bank/n3116 , \Reg_Bank/n3115 , \Reg_Bank/n3114 ,
         \Reg_Bank/n3113 , \Reg_Bank/n3112 , \Reg_Bank/n3111 ,
         \Reg_Bank/n3110 , \Reg_Bank/n3109 , \Reg_Bank/n3108 ,
         \Reg_Bank/n3107 , \Reg_Bank/n3106 , \Reg_Bank/n3105 ,
         \Reg_Bank/n3104 , \Reg_Bank/n3103 , \Reg_Bank/n3102 ,
         \Reg_Bank/n3101 , \Reg_Bank/n3100 , \Reg_Bank/n3099 ,
         \Reg_Bank/n3098 , \Reg_Bank/n3097 , \Reg_Bank/n3096 ,
         \Reg_Bank/n3095 , \Reg_Bank/n3094 , \Reg_Bank/n3093 ,
         \Reg_Bank/n3092 , \Reg_Bank/n3091 , \Reg_Bank/n3090 ,
         \Reg_Bank/n3089 , \Reg_Bank/n3088 , \Reg_Bank/n3087 ,
         \Reg_Bank/n3086 , \Reg_Bank/n3085 , \Reg_Bank/n3084 ,
         \Reg_Bank/n3083 , \Reg_Bank/n3082 , \Reg_Bank/n3081 ,
         \Reg_Bank/n3080 , \Reg_Bank/n3079 , \Reg_Bank/n3078 ,
         \Reg_Bank/n3077 , \Reg_Bank/n3076 , \Reg_Bank/n3075 ,
         \Reg_Bank/n3074 , \Reg_Bank/n3073 , \Reg_Bank/n3072 ,
         \Reg_Bank/n3071 , \Reg_Bank/n3070 , \Reg_Bank/n3069 ,
         \Reg_Bank/n3068 , \Reg_Bank/n3067 , \Reg_Bank/n3066 ,
         \Reg_Bank/n3065 , \Reg_Bank/n3064 , \Reg_Bank/n3063 ,
         \Reg_Bank/n3062 , \Reg_Bank/n3061 , \Reg_Bank/n3060 ,
         \Reg_Bank/n3059 , \Reg_Bank/n3058 , \Reg_Bank/n3057 ,
         \Reg_Bank/n3056 , \Reg_Bank/n3055 , \Reg_Bank/n3054 ,
         \Reg_Bank/n3053 , \Reg_Bank/n3052 , \Reg_Bank/n3051 ,
         \Reg_Bank/n3050 , \Reg_Bank/n3049 , \Reg_Bank/n3048 ,
         \Reg_Bank/n3047 , \Reg_Bank/n3046 , \Reg_Bank/n3045 ,
         \Reg_Bank/n3044 , \Reg_Bank/n3043 , \Reg_Bank/n3042 ,
         \Reg_Bank/n3041 , \Reg_Bank/n3040 , \Reg_Bank/n3039 ,
         \Reg_Bank/n3038 , \Reg_Bank/n3037 , \Reg_Bank/n3036 ,
         \Reg_Bank/n3035 , \Reg_Bank/n3034 , \Reg_Bank/n3033 ,
         \Reg_Bank/n3032 , \Reg_Bank/n3031 , \Reg_Bank/n3030 ,
         \Reg_Bank/registers[1][0] , \Reg_Bank/registers[1][1] ,
         \Reg_Bank/registers[1][2] , \Reg_Bank/registers[1][3] ,
         \Reg_Bank/registers[1][4] , \Reg_Bank/registers[1][5] ,
         \Reg_Bank/registers[1][6] , \Reg_Bank/registers[1][7] ,
         \Reg_Bank/registers[1][8] , \Reg_Bank/registers[1][9] ,
         \Reg_Bank/registers[1][10] , \Reg_Bank/registers[1][11] ,
         \Reg_Bank/registers[1][12] , \Reg_Bank/registers[1][13] ,
         \Reg_Bank/registers[1][14] , \Reg_Bank/registers[1][15] ,
         \Reg_Bank/registers[1][16] , \Reg_Bank/registers[1][17] ,
         \Reg_Bank/registers[1][18] , \Reg_Bank/registers[1][19] ,
         \Reg_Bank/registers[1][20] , \Reg_Bank/registers[1][21] ,
         \Reg_Bank/registers[1][22] , \Reg_Bank/registers[1][23] ,
         \Reg_Bank/registers[1][24] , \Reg_Bank/registers[1][25] ,
         \Reg_Bank/registers[1][26] , \Reg_Bank/registers[1][27] ,
         \Reg_Bank/registers[1][28] , \Reg_Bank/registers[1][29] ,
         \Reg_Bank/registers[1][30] , \Reg_Bank/registers[1][31] ,
         \Reg_Bank/registers[2][0] , \Reg_Bank/registers[2][1] ,
         \Reg_Bank/registers[2][2] , \Reg_Bank/registers[2][3] ,
         \Reg_Bank/registers[2][4] , \Reg_Bank/registers[2][5] ,
         \Reg_Bank/registers[2][6] , \Reg_Bank/registers[2][7] ,
         \Reg_Bank/registers[2][8] , \Reg_Bank/registers[2][9] ,
         \Reg_Bank/registers[2][10] , \Reg_Bank/registers[2][11] ,
         \Reg_Bank/registers[2][12] , \Reg_Bank/registers[2][13] ,
         \Reg_Bank/registers[2][14] , \Reg_Bank/registers[2][15] ,
         \Reg_Bank/registers[2][16] , \Reg_Bank/registers[2][17] ,
         \Reg_Bank/registers[2][18] , \Reg_Bank/registers[2][19] ,
         \Reg_Bank/registers[2][20] , \Reg_Bank/registers[2][21] ,
         \Reg_Bank/registers[2][22] , \Reg_Bank/registers[2][23] ,
         \Reg_Bank/registers[2][24] , \Reg_Bank/registers[2][25] ,
         \Reg_Bank/registers[2][26] , \Reg_Bank/registers[2][27] ,
         \Reg_Bank/registers[2][28] , \Reg_Bank/registers[2][29] ,
         \Reg_Bank/registers[2][30] , \Reg_Bank/registers[2][31] ,
         \Reg_Bank/registers[3][0] , \Reg_Bank/registers[3][1] ,
         \Reg_Bank/registers[3][2] , \Reg_Bank/registers[3][3] ,
         \Reg_Bank/registers[3][4] , \Reg_Bank/registers[3][5] ,
         \Reg_Bank/registers[3][6] , \Reg_Bank/registers[3][7] ,
         \Reg_Bank/registers[3][8] , \Reg_Bank/registers[3][9] ,
         \Reg_Bank/registers[3][10] , \Reg_Bank/registers[3][11] ,
         \Reg_Bank/registers[3][12] , \Reg_Bank/registers[3][13] ,
         \Reg_Bank/registers[3][14] , \Reg_Bank/registers[3][15] ,
         \Reg_Bank/registers[3][16] , \Reg_Bank/registers[3][17] ,
         \Reg_Bank/registers[3][18] , \Reg_Bank/registers[3][19] ,
         \Reg_Bank/registers[3][20] , \Reg_Bank/registers[3][21] ,
         \Reg_Bank/registers[3][22] , \Reg_Bank/registers[3][23] ,
         \Reg_Bank/registers[3][24] , \Reg_Bank/registers[3][25] ,
         \Reg_Bank/registers[3][26] , \Reg_Bank/registers[3][27] ,
         \Reg_Bank/registers[3][28] , \Reg_Bank/registers[3][29] ,
         \Reg_Bank/registers[3][30] , \Reg_Bank/registers[3][31] ,
         \Reg_Bank/registers[4][0] , \Reg_Bank/registers[4][1] ,
         \Reg_Bank/registers[4][2] , \Reg_Bank/registers[4][3] ,
         \Reg_Bank/registers[4][4] , \Reg_Bank/registers[4][5] ,
         \Reg_Bank/registers[4][6] , \Reg_Bank/registers[4][7] ,
         \Reg_Bank/registers[4][8] , \Reg_Bank/registers[4][9] ,
         \Reg_Bank/registers[4][10] , \Reg_Bank/registers[4][11] ,
         \Reg_Bank/registers[4][12] , \Reg_Bank/registers[4][13] ,
         \Reg_Bank/registers[4][14] , \Reg_Bank/registers[4][15] ,
         \Reg_Bank/registers[4][16] , \Reg_Bank/registers[4][17] ,
         \Reg_Bank/registers[4][18] , \Reg_Bank/registers[4][19] ,
         \Reg_Bank/registers[4][20] , \Reg_Bank/registers[4][21] ,
         \Reg_Bank/registers[4][22] , \Reg_Bank/registers[4][23] ,
         \Reg_Bank/registers[4][24] , \Reg_Bank/registers[4][25] ,
         \Reg_Bank/registers[4][26] , \Reg_Bank/registers[4][27] ,
         \Reg_Bank/registers[4][28] , \Reg_Bank/registers[4][29] ,
         \Reg_Bank/registers[4][30] , \Reg_Bank/registers[4][31] ,
         \Reg_Bank/registers[5][0] , \Reg_Bank/registers[5][1] ,
         \Reg_Bank/registers[5][2] , \Reg_Bank/registers[5][3] ,
         \Reg_Bank/registers[5][4] , \Reg_Bank/registers[5][5] ,
         \Reg_Bank/registers[5][6] , \Reg_Bank/registers[5][7] ,
         \Reg_Bank/registers[5][8] , \Reg_Bank/registers[5][9] ,
         \Reg_Bank/registers[5][10] , \Reg_Bank/registers[5][11] ,
         \Reg_Bank/registers[5][12] , \Reg_Bank/registers[5][13] ,
         \Reg_Bank/registers[5][14] , \Reg_Bank/registers[5][15] ,
         \Reg_Bank/registers[5][16] , \Reg_Bank/registers[5][17] ,
         \Reg_Bank/registers[5][18] , \Reg_Bank/registers[5][19] ,
         \Reg_Bank/registers[5][20] , \Reg_Bank/registers[5][21] ,
         \Reg_Bank/registers[5][22] , \Reg_Bank/registers[5][23] ,
         \Reg_Bank/registers[5][24] , \Reg_Bank/registers[5][25] ,
         \Reg_Bank/registers[5][26] , \Reg_Bank/registers[5][27] ,
         \Reg_Bank/registers[5][28] , \Reg_Bank/registers[5][29] ,
         \Reg_Bank/registers[5][30] , \Reg_Bank/registers[5][31] ,
         \Reg_Bank/registers[6][0] , \Reg_Bank/registers[6][1] ,
         \Reg_Bank/registers[6][2] , \Reg_Bank/registers[6][3] ,
         \Reg_Bank/registers[6][4] , \Reg_Bank/registers[6][5] ,
         \Reg_Bank/registers[6][6] , \Reg_Bank/registers[6][7] ,
         \Reg_Bank/registers[6][8] , \Reg_Bank/registers[6][9] ,
         \Reg_Bank/registers[6][10] , \Reg_Bank/registers[6][11] ,
         \Reg_Bank/registers[6][12] , \Reg_Bank/registers[6][13] ,
         \Reg_Bank/registers[6][14] , \Reg_Bank/registers[6][15] ,
         \Reg_Bank/registers[6][16] , \Reg_Bank/registers[6][17] ,
         \Reg_Bank/registers[6][18] , \Reg_Bank/registers[6][19] ,
         \Reg_Bank/registers[6][20] , \Reg_Bank/registers[6][21] ,
         \Reg_Bank/registers[6][22] , \Reg_Bank/registers[6][23] ,
         \Reg_Bank/registers[6][24] , \Reg_Bank/registers[6][25] ,
         \Reg_Bank/registers[6][26] , \Reg_Bank/registers[6][27] ,
         \Reg_Bank/registers[6][28] , \Reg_Bank/registers[6][29] ,
         \Reg_Bank/registers[6][30] , \Reg_Bank/registers[6][31] ,
         \Reg_Bank/registers[7][0] , \Reg_Bank/registers[7][1] ,
         \Reg_Bank/registers[7][2] , \Reg_Bank/registers[7][3] ,
         \Reg_Bank/registers[7][4] , \Reg_Bank/registers[7][5] ,
         \Reg_Bank/registers[7][6] , \Reg_Bank/registers[7][7] ,
         \Reg_Bank/registers[7][8] , \Reg_Bank/registers[7][9] ,
         \Reg_Bank/registers[7][10] , \Reg_Bank/registers[7][11] ,
         \Reg_Bank/registers[7][12] , \Reg_Bank/registers[7][13] ,
         \Reg_Bank/registers[7][14] , \Reg_Bank/registers[7][15] ,
         \Reg_Bank/registers[7][16] , \Reg_Bank/registers[7][17] ,
         \Reg_Bank/registers[7][18] , \Reg_Bank/registers[7][19] ,
         \Reg_Bank/registers[7][20] , \Reg_Bank/registers[7][21] ,
         \Reg_Bank/registers[7][22] , \Reg_Bank/registers[7][23] ,
         \Reg_Bank/registers[7][24] , \Reg_Bank/registers[7][25] ,
         \Reg_Bank/registers[7][26] , \Reg_Bank/registers[7][27] ,
         \Reg_Bank/registers[7][28] , \Reg_Bank/registers[7][29] ,
         \Reg_Bank/registers[7][30] , \Reg_Bank/registers[7][31] ,
         \Reg_Bank/registers[8][0] , \Reg_Bank/registers[8][1] ,
         \Reg_Bank/registers[8][2] , \Reg_Bank/registers[8][3] ,
         \Reg_Bank/registers[8][4] , \Reg_Bank/registers[8][5] ,
         \Reg_Bank/registers[8][6] , \Reg_Bank/registers[8][7] ,
         \Reg_Bank/registers[8][8] , \Reg_Bank/registers[8][9] ,
         \Reg_Bank/registers[8][10] , \Reg_Bank/registers[8][11] ,
         \Reg_Bank/registers[8][12] , \Reg_Bank/registers[8][13] ,
         \Reg_Bank/registers[8][14] , \Reg_Bank/registers[8][15] ,
         \Reg_Bank/registers[8][16] , \Reg_Bank/registers[8][17] ,
         \Reg_Bank/registers[8][18] , \Reg_Bank/registers[8][19] ,
         \Reg_Bank/registers[8][20] , \Reg_Bank/registers[8][21] ,
         \Reg_Bank/registers[8][22] , \Reg_Bank/registers[8][23] ,
         \Reg_Bank/registers[8][24] , \Reg_Bank/registers[8][25] ,
         \Reg_Bank/registers[8][26] , \Reg_Bank/registers[8][27] ,
         \Reg_Bank/registers[8][28] , \Reg_Bank/registers[8][29] ,
         \Reg_Bank/registers[8][30] , \Reg_Bank/registers[8][31] ,
         \Reg_Bank/registers[9][0] , \Reg_Bank/registers[9][1] ,
         \Reg_Bank/registers[9][2] , \Reg_Bank/registers[9][3] ,
         \Reg_Bank/registers[9][4] , \Reg_Bank/registers[9][5] ,
         \Reg_Bank/registers[9][6] , \Reg_Bank/registers[9][7] ,
         \Reg_Bank/registers[9][8] , \Reg_Bank/registers[9][9] ,
         \Reg_Bank/registers[9][10] , \Reg_Bank/registers[9][11] ,
         \Reg_Bank/registers[9][12] , \Reg_Bank/registers[9][13] ,
         \Reg_Bank/registers[9][14] , \Reg_Bank/registers[9][15] ,
         \Reg_Bank/registers[9][16] , \Reg_Bank/registers[9][17] ,
         \Reg_Bank/registers[9][18] , \Reg_Bank/registers[9][19] ,
         \Reg_Bank/registers[9][20] , \Reg_Bank/registers[9][21] ,
         \Reg_Bank/registers[9][22] , \Reg_Bank/registers[9][23] ,
         \Reg_Bank/registers[9][24] , \Reg_Bank/registers[9][25] ,
         \Reg_Bank/registers[9][26] , \Reg_Bank/registers[9][27] ,
         \Reg_Bank/registers[9][28] , \Reg_Bank/registers[9][29] ,
         \Reg_Bank/registers[9][30] , \Reg_Bank/registers[9][31] ,
         \Reg_Bank/registers[10][0] , \Reg_Bank/registers[10][1] ,
         \Reg_Bank/registers[10][2] , \Reg_Bank/registers[10][3] ,
         \Reg_Bank/registers[10][4] , \Reg_Bank/registers[10][5] ,
         \Reg_Bank/registers[10][6] , \Reg_Bank/registers[10][7] ,
         \Reg_Bank/registers[10][8] , \Reg_Bank/registers[10][9] ,
         \Reg_Bank/registers[10][10] , \Reg_Bank/registers[10][11] ,
         \Reg_Bank/registers[10][12] , \Reg_Bank/registers[10][13] ,
         \Reg_Bank/registers[10][14] , \Reg_Bank/registers[10][15] ,
         \Reg_Bank/registers[10][16] , \Reg_Bank/registers[10][17] ,
         \Reg_Bank/registers[10][18] , \Reg_Bank/registers[10][19] ,
         \Reg_Bank/registers[10][20] , \Reg_Bank/registers[10][21] ,
         \Reg_Bank/registers[10][22] , \Reg_Bank/registers[10][23] ,
         \Reg_Bank/registers[10][24] , \Reg_Bank/registers[10][25] ,
         \Reg_Bank/registers[10][26] , \Reg_Bank/registers[10][27] ,
         \Reg_Bank/registers[10][28] , \Reg_Bank/registers[10][29] ,
         \Reg_Bank/registers[10][30] , \Reg_Bank/registers[10][31] ,
         \Reg_Bank/registers[11][0] , \Reg_Bank/registers[11][1] ,
         \Reg_Bank/registers[11][2] , \Reg_Bank/registers[11][3] ,
         \Reg_Bank/registers[11][4] , \Reg_Bank/registers[11][5] ,
         \Reg_Bank/registers[11][6] , \Reg_Bank/registers[11][7] ,
         \Reg_Bank/registers[11][8] , \Reg_Bank/registers[11][9] ,
         \Reg_Bank/registers[11][10] , \Reg_Bank/registers[11][11] ,
         \Reg_Bank/registers[11][12] , \Reg_Bank/registers[11][13] ,
         \Reg_Bank/registers[11][14] , \Reg_Bank/registers[11][15] ,
         \Reg_Bank/registers[11][16] , \Reg_Bank/registers[11][17] ,
         \Reg_Bank/registers[11][18] , \Reg_Bank/registers[11][19] ,
         \Reg_Bank/registers[11][20] , \Reg_Bank/registers[11][21] ,
         \Reg_Bank/registers[11][22] , \Reg_Bank/registers[11][23] ,
         \Reg_Bank/registers[11][24] , \Reg_Bank/registers[11][25] ,
         \Reg_Bank/registers[11][26] , \Reg_Bank/registers[11][27] ,
         \Reg_Bank/registers[11][28] , \Reg_Bank/registers[11][29] ,
         \Reg_Bank/registers[11][30] , \Reg_Bank/registers[11][31] ,
         \Reg_Bank/registers[12][0] , \Reg_Bank/registers[12][1] ,
         \Reg_Bank/registers[12][2] , \Reg_Bank/registers[12][3] ,
         \Reg_Bank/registers[12][4] , \Reg_Bank/registers[12][5] ,
         \Reg_Bank/registers[12][6] , \Reg_Bank/registers[12][7] ,
         \Reg_Bank/registers[12][8] , \Reg_Bank/registers[12][9] ,
         \Reg_Bank/registers[12][10] , \Reg_Bank/registers[12][11] ,
         \Reg_Bank/registers[12][12] , \Reg_Bank/registers[12][13] ,
         \Reg_Bank/registers[12][14] , \Reg_Bank/registers[12][15] ,
         \Reg_Bank/registers[12][16] , \Reg_Bank/registers[12][17] ,
         \Reg_Bank/registers[12][18] , \Reg_Bank/registers[12][19] ,
         \Reg_Bank/registers[12][20] , \Reg_Bank/registers[12][21] ,
         \Reg_Bank/registers[12][22] , \Reg_Bank/registers[12][23] ,
         \Reg_Bank/registers[12][24] , \Reg_Bank/registers[12][25] ,
         \Reg_Bank/registers[12][26] , \Reg_Bank/registers[12][27] ,
         \Reg_Bank/registers[12][28] , \Reg_Bank/registers[12][29] ,
         \Reg_Bank/registers[12][30] , \Reg_Bank/registers[12][31] ,
         \Reg_Bank/registers[13][0] , \Reg_Bank/registers[13][1] ,
         \Reg_Bank/registers[13][2] , \Reg_Bank/registers[13][3] ,
         \Reg_Bank/registers[13][4] , \Reg_Bank/registers[13][5] ,
         \Reg_Bank/registers[13][6] , \Reg_Bank/registers[13][7] ,
         \Reg_Bank/registers[13][8] , \Reg_Bank/registers[13][9] ,
         \Reg_Bank/registers[13][10] , \Reg_Bank/registers[13][11] ,
         \Reg_Bank/registers[13][12] , \Reg_Bank/registers[13][13] ,
         \Reg_Bank/registers[13][14] , \Reg_Bank/registers[13][15] ,
         \Reg_Bank/registers[13][16] , \Reg_Bank/registers[13][17] ,
         \Reg_Bank/registers[13][18] , \Reg_Bank/registers[13][19] ,
         \Reg_Bank/registers[13][20] , \Reg_Bank/registers[13][21] ,
         \Reg_Bank/registers[13][22] , \Reg_Bank/registers[13][23] ,
         \Reg_Bank/registers[13][24] , \Reg_Bank/registers[13][25] ,
         \Reg_Bank/registers[13][26] , \Reg_Bank/registers[13][27] ,
         \Reg_Bank/registers[13][28] , \Reg_Bank/registers[13][29] ,
         \Reg_Bank/registers[13][30] , \Reg_Bank/registers[13][31] ,
         \Reg_Bank/registers[14][0] , \Reg_Bank/registers[14][1] ,
         \Reg_Bank/registers[14][2] , \Reg_Bank/registers[14][3] ,
         \Reg_Bank/registers[14][4] , \Reg_Bank/registers[14][5] ,
         \Reg_Bank/registers[14][6] , \Reg_Bank/registers[14][7] ,
         \Reg_Bank/registers[14][8] , \Reg_Bank/registers[14][9] ,
         \Reg_Bank/registers[14][10] , \Reg_Bank/registers[14][11] ,
         \Reg_Bank/registers[14][12] , \Reg_Bank/registers[14][13] ,
         \Reg_Bank/registers[14][14] , \Reg_Bank/registers[14][15] ,
         \Reg_Bank/registers[14][16] , \Reg_Bank/registers[14][17] ,
         \Reg_Bank/registers[14][18] , \Reg_Bank/registers[14][19] ,
         \Reg_Bank/registers[14][20] , \Reg_Bank/registers[14][21] ,
         \Reg_Bank/registers[14][22] , \Reg_Bank/registers[14][23] ,
         \Reg_Bank/registers[14][24] , \Reg_Bank/registers[14][25] ,
         \Reg_Bank/registers[14][26] , \Reg_Bank/registers[14][27] ,
         \Reg_Bank/registers[14][28] , \Reg_Bank/registers[14][29] ,
         \Reg_Bank/registers[14][30] , \Reg_Bank/registers[14][31] ,
         \Reg_Bank/registers[15][0] , \Reg_Bank/registers[15][1] ,
         \Reg_Bank/registers[15][2] , \Reg_Bank/registers[15][3] ,
         \Reg_Bank/registers[15][4] , \Reg_Bank/registers[15][5] ,
         \Reg_Bank/registers[15][6] , \Reg_Bank/registers[15][7] ,
         \Reg_Bank/registers[15][8] , \Reg_Bank/registers[15][9] ,
         \Reg_Bank/registers[15][10] , \Reg_Bank/registers[15][11] ,
         \Reg_Bank/registers[15][12] , \Reg_Bank/registers[15][13] ,
         \Reg_Bank/registers[15][14] , \Reg_Bank/registers[15][15] ,
         \Reg_Bank/registers[15][16] , \Reg_Bank/registers[15][17] ,
         \Reg_Bank/registers[15][18] , \Reg_Bank/registers[15][19] ,
         \Reg_Bank/registers[15][20] , \Reg_Bank/registers[15][21] ,
         \Reg_Bank/registers[15][22] , \Reg_Bank/registers[15][23] ,
         \Reg_Bank/registers[15][24] , \Reg_Bank/registers[15][25] ,
         \Reg_Bank/registers[15][26] , \Reg_Bank/registers[15][27] ,
         \Reg_Bank/registers[15][28] , \Reg_Bank/registers[15][29] ,
         \Reg_Bank/registers[15][30] , \Reg_Bank/registers[15][31] ,
         \Reg_Bank/registers[16][0] , \Reg_Bank/registers[16][1] ,
         \Reg_Bank/registers[16][2] , \Reg_Bank/registers[16][3] ,
         \Reg_Bank/registers[16][4] , \Reg_Bank/registers[16][5] ,
         \Reg_Bank/registers[16][6] , \Reg_Bank/registers[16][7] ,
         \Reg_Bank/registers[16][8] , \Reg_Bank/registers[16][9] ,
         \Reg_Bank/registers[16][10] , \Reg_Bank/registers[16][11] ,
         \Reg_Bank/registers[16][12] , \Reg_Bank/registers[16][13] ,
         \Reg_Bank/registers[16][14] , \Reg_Bank/registers[16][15] ,
         \Reg_Bank/registers[16][16] , \Reg_Bank/registers[16][17] ,
         \Reg_Bank/registers[16][18] , \Reg_Bank/registers[16][19] ,
         \Reg_Bank/registers[16][20] , \Reg_Bank/registers[16][21] ,
         \Reg_Bank/registers[16][22] , \Reg_Bank/registers[16][23] ,
         \Reg_Bank/registers[16][24] , \Reg_Bank/registers[16][25] ,
         \Reg_Bank/registers[16][26] , \Reg_Bank/registers[16][27] ,
         \Reg_Bank/registers[16][28] , \Reg_Bank/registers[16][29] ,
         \Reg_Bank/registers[16][30] , \Reg_Bank/registers[16][31] ,
         \Reg_Bank/registers[17][0] , \Reg_Bank/registers[17][1] ,
         \Reg_Bank/registers[17][2] , \Reg_Bank/registers[17][3] ,
         \Reg_Bank/registers[17][4] , \Reg_Bank/registers[17][5] ,
         \Reg_Bank/registers[17][6] , \Reg_Bank/registers[17][7] ,
         \Reg_Bank/registers[17][8] , \Reg_Bank/registers[17][9] ,
         \Reg_Bank/registers[17][10] , \Reg_Bank/registers[17][11] ,
         \Reg_Bank/registers[17][12] , \Reg_Bank/registers[17][13] ,
         \Reg_Bank/registers[17][14] , \Reg_Bank/registers[17][15] ,
         \Reg_Bank/registers[17][16] , \Reg_Bank/registers[17][17] ,
         \Reg_Bank/registers[17][18] , \Reg_Bank/registers[17][19] ,
         \Reg_Bank/registers[17][20] , \Reg_Bank/registers[17][21] ,
         \Reg_Bank/registers[17][22] , \Reg_Bank/registers[17][23] ,
         \Reg_Bank/registers[17][24] , \Reg_Bank/registers[17][25] ,
         \Reg_Bank/registers[17][26] , \Reg_Bank/registers[17][27] ,
         \Reg_Bank/registers[17][28] , \Reg_Bank/registers[17][29] ,
         \Reg_Bank/registers[17][30] , \Reg_Bank/registers[17][31] ,
         \Reg_Bank/registers[18][0] , \Reg_Bank/registers[18][1] ,
         \Reg_Bank/registers[18][2] , \Reg_Bank/registers[18][3] ,
         \Reg_Bank/registers[18][4] , \Reg_Bank/registers[18][5] ,
         \Reg_Bank/registers[18][6] , \Reg_Bank/registers[18][7] ,
         \Reg_Bank/registers[18][8] , \Reg_Bank/registers[18][9] ,
         \Reg_Bank/registers[18][10] , \Reg_Bank/registers[18][11] ,
         \Reg_Bank/registers[18][12] , \Reg_Bank/registers[18][13] ,
         \Reg_Bank/registers[18][14] , \Reg_Bank/registers[18][15] ,
         \Reg_Bank/registers[18][16] , \Reg_Bank/registers[18][17] ,
         \Reg_Bank/registers[18][18] , \Reg_Bank/registers[18][19] ,
         \Reg_Bank/registers[18][20] , \Reg_Bank/registers[18][21] ,
         \Reg_Bank/registers[18][22] , \Reg_Bank/registers[18][23] ,
         \Reg_Bank/registers[18][24] , \Reg_Bank/registers[18][25] ,
         \Reg_Bank/registers[18][26] , \Reg_Bank/registers[18][27] ,
         \Reg_Bank/registers[18][28] , \Reg_Bank/registers[18][29] ,
         \Reg_Bank/registers[18][30] , \Reg_Bank/registers[18][31] ,
         \Reg_Bank/registers[19][0] , \Reg_Bank/registers[19][1] ,
         \Reg_Bank/registers[19][2] , \Reg_Bank/registers[19][3] ,
         \Reg_Bank/registers[19][4] , \Reg_Bank/registers[19][5] ,
         \Reg_Bank/registers[19][6] , \Reg_Bank/registers[19][7] ,
         \Reg_Bank/registers[19][8] , \Reg_Bank/registers[19][9] ,
         \Reg_Bank/registers[19][10] , \Reg_Bank/registers[19][11] ,
         \Reg_Bank/registers[19][12] , \Reg_Bank/registers[19][13] ,
         \Reg_Bank/registers[19][14] , \Reg_Bank/registers[19][15] ,
         \Reg_Bank/registers[19][16] , \Reg_Bank/registers[19][17] ,
         \Reg_Bank/registers[19][18] , \Reg_Bank/registers[19][19] ,
         \Reg_Bank/registers[19][20] , \Reg_Bank/registers[19][21] ,
         \Reg_Bank/registers[19][22] , \Reg_Bank/registers[19][23] ,
         \Reg_Bank/registers[19][24] , \Reg_Bank/registers[19][25] ,
         \Reg_Bank/registers[19][26] , \Reg_Bank/registers[19][27] ,
         \Reg_Bank/registers[19][28] , \Reg_Bank/registers[19][29] ,
         \Reg_Bank/registers[19][30] , \Reg_Bank/registers[19][31] ,
         \Reg_Bank/registers[20][0] , \Reg_Bank/registers[20][1] ,
         \Reg_Bank/registers[20][2] , \Reg_Bank/registers[20][3] ,
         \Reg_Bank/registers[20][4] , \Reg_Bank/registers[20][5] ,
         \Reg_Bank/registers[20][6] , \Reg_Bank/registers[20][7] ,
         \Reg_Bank/registers[20][8] , \Reg_Bank/registers[20][9] ,
         \Reg_Bank/registers[20][10] , \Reg_Bank/registers[20][11] ,
         \Reg_Bank/registers[20][12] , \Reg_Bank/registers[20][13] ,
         \Reg_Bank/registers[20][14] , \Reg_Bank/registers[20][15] ,
         \Reg_Bank/registers[20][16] , \Reg_Bank/registers[20][17] ,
         \Reg_Bank/registers[20][18] , \Reg_Bank/registers[20][19] ,
         \Reg_Bank/registers[20][20] , \Reg_Bank/registers[20][21] ,
         \Reg_Bank/registers[20][22] , \Reg_Bank/registers[20][23] ,
         \Reg_Bank/registers[20][24] , \Reg_Bank/registers[20][25] ,
         \Reg_Bank/registers[20][26] , \Reg_Bank/registers[20][27] ,
         \Reg_Bank/registers[20][28] , \Reg_Bank/registers[20][29] ,
         \Reg_Bank/registers[20][30] , \Reg_Bank/registers[20][31] ,
         \Reg_Bank/registers[21][0] , \Reg_Bank/registers[21][1] ,
         \Reg_Bank/registers[21][2] , \Reg_Bank/registers[21][3] ,
         \Reg_Bank/registers[21][4] , \Reg_Bank/registers[21][5] ,
         \Reg_Bank/registers[21][6] , \Reg_Bank/registers[21][7] ,
         \Reg_Bank/registers[21][8] , \Reg_Bank/registers[21][9] ,
         \Reg_Bank/registers[21][10] , \Reg_Bank/registers[21][11] ,
         \Reg_Bank/registers[21][12] , \Reg_Bank/registers[21][13] ,
         \Reg_Bank/registers[21][14] , \Reg_Bank/registers[21][15] ,
         \Reg_Bank/registers[21][16] , \Reg_Bank/registers[21][17] ,
         \Reg_Bank/registers[21][18] , \Reg_Bank/registers[21][19] ,
         \Reg_Bank/registers[21][20] , \Reg_Bank/registers[21][21] ,
         \Reg_Bank/registers[21][22] , \Reg_Bank/registers[21][23] ,
         \Reg_Bank/registers[21][24] , \Reg_Bank/registers[21][25] ,
         \Reg_Bank/registers[21][26] , \Reg_Bank/registers[21][27] ,
         \Reg_Bank/registers[21][28] , \Reg_Bank/registers[21][29] ,
         \Reg_Bank/registers[21][30] , \Reg_Bank/registers[21][31] ,
         \Reg_Bank/registers[22][0] , \Reg_Bank/registers[22][1] ,
         \Reg_Bank/registers[22][2] , \Reg_Bank/registers[22][3] ,
         \Reg_Bank/registers[22][4] , \Reg_Bank/registers[22][5] ,
         \Reg_Bank/registers[22][6] , \Reg_Bank/registers[22][7] ,
         \Reg_Bank/registers[22][8] , \Reg_Bank/registers[22][9] ,
         \Reg_Bank/registers[22][10] , \Reg_Bank/registers[22][11] ,
         \Reg_Bank/registers[22][12] , \Reg_Bank/registers[22][13] ,
         \Reg_Bank/registers[22][14] , \Reg_Bank/registers[22][15] ,
         \Reg_Bank/registers[22][16] , \Reg_Bank/registers[22][17] ,
         \Reg_Bank/registers[22][18] , \Reg_Bank/registers[22][19] ,
         \Reg_Bank/registers[22][20] , \Reg_Bank/registers[22][21] ,
         \Reg_Bank/registers[22][22] , \Reg_Bank/registers[22][23] ,
         \Reg_Bank/registers[22][24] , \Reg_Bank/registers[22][25] ,
         \Reg_Bank/registers[22][26] , \Reg_Bank/registers[22][27] ,
         \Reg_Bank/registers[22][28] , \Reg_Bank/registers[22][29] ,
         \Reg_Bank/registers[22][30] , \Reg_Bank/registers[22][31] ,
         \Reg_Bank/registers[23][0] , \Reg_Bank/registers[23][1] ,
         \Reg_Bank/registers[23][2] , \Reg_Bank/registers[23][3] ,
         \Reg_Bank/registers[23][4] , \Reg_Bank/registers[23][5] ,
         \Reg_Bank/registers[23][6] , \Reg_Bank/registers[23][7] ,
         \Reg_Bank/registers[23][8] , \Reg_Bank/registers[23][9] ,
         \Reg_Bank/registers[23][10] , \Reg_Bank/registers[23][11] ,
         \Reg_Bank/registers[23][12] , \Reg_Bank/registers[23][13] ,
         \Reg_Bank/registers[23][14] , \Reg_Bank/registers[23][15] ,
         \Reg_Bank/registers[23][16] , \Reg_Bank/registers[23][17] ,
         \Reg_Bank/registers[23][18] , \Reg_Bank/registers[23][19] ,
         \Reg_Bank/registers[23][20] , \Reg_Bank/registers[23][21] ,
         \Reg_Bank/registers[23][22] , \Reg_Bank/registers[23][23] ,
         \Reg_Bank/registers[23][24] , \Reg_Bank/registers[23][25] ,
         \Reg_Bank/registers[23][26] , \Reg_Bank/registers[23][27] ,
         \Reg_Bank/registers[23][28] , \Reg_Bank/registers[23][29] ,
         \Reg_Bank/registers[23][30] , \Reg_Bank/registers[23][31] ,
         \Reg_Bank/registers[24][0] , \Reg_Bank/registers[24][1] ,
         \Reg_Bank/registers[24][2] , \Reg_Bank/registers[24][3] ,
         \Reg_Bank/registers[24][4] , \Reg_Bank/registers[24][5] ,
         \Reg_Bank/registers[24][6] , \Reg_Bank/registers[24][7] ,
         \Reg_Bank/registers[24][8] , \Reg_Bank/registers[24][9] ,
         \Reg_Bank/registers[24][10] , \Reg_Bank/registers[24][11] ,
         \Reg_Bank/registers[24][12] , \Reg_Bank/registers[24][13] ,
         \Reg_Bank/registers[24][14] , \Reg_Bank/registers[24][15] ,
         \Reg_Bank/registers[24][16] , \Reg_Bank/registers[24][17] ,
         \Reg_Bank/registers[24][18] , \Reg_Bank/registers[24][19] ,
         \Reg_Bank/registers[24][20] , \Reg_Bank/registers[24][21] ,
         \Reg_Bank/registers[24][22] , \Reg_Bank/registers[24][23] ,
         \Reg_Bank/registers[24][24] , \Reg_Bank/registers[24][25] ,
         \Reg_Bank/registers[24][26] , \Reg_Bank/registers[24][27] ,
         \Reg_Bank/registers[24][28] , \Reg_Bank/registers[24][29] ,
         \Reg_Bank/registers[24][30] , \Reg_Bank/registers[24][31] ,
         \Reg_Bank/registers[25][0] , \Reg_Bank/registers[25][1] ,
         \Reg_Bank/registers[25][2] , \Reg_Bank/registers[25][3] ,
         \Reg_Bank/registers[25][4] , \Reg_Bank/registers[25][5] ,
         \Reg_Bank/registers[25][6] , \Reg_Bank/registers[25][7] ,
         \Reg_Bank/registers[25][8] , \Reg_Bank/registers[25][9] ,
         \Reg_Bank/registers[25][10] , \Reg_Bank/registers[25][11] ,
         \Reg_Bank/registers[25][12] , \Reg_Bank/registers[25][13] ,
         \Reg_Bank/registers[25][14] , \Reg_Bank/registers[25][15] ,
         \Reg_Bank/registers[25][16] , \Reg_Bank/registers[25][17] ,
         \Reg_Bank/registers[25][18] , \Reg_Bank/registers[25][19] ,
         \Reg_Bank/registers[25][20] , \Reg_Bank/registers[25][21] ,
         \Reg_Bank/registers[25][22] , \Reg_Bank/registers[25][23] ,
         \Reg_Bank/registers[25][24] , \Reg_Bank/registers[25][25] ,
         \Reg_Bank/registers[25][26] , \Reg_Bank/registers[25][27] ,
         \Reg_Bank/registers[25][28] , \Reg_Bank/registers[25][29] ,
         \Reg_Bank/registers[25][30] , \Reg_Bank/registers[25][31] ,
         \Reg_Bank/registers[26][0] , \Reg_Bank/registers[26][1] ,
         \Reg_Bank/registers[26][2] , \Reg_Bank/registers[26][3] ,
         \Reg_Bank/registers[26][4] , \Reg_Bank/registers[26][5] ,
         \Reg_Bank/registers[26][6] , \Reg_Bank/registers[26][7] ,
         \Reg_Bank/registers[26][8] , \Reg_Bank/registers[26][9] ,
         \Reg_Bank/registers[26][10] , \Reg_Bank/registers[26][11] ,
         \Reg_Bank/registers[26][12] , \Reg_Bank/registers[26][13] ,
         \Reg_Bank/registers[26][14] , \Reg_Bank/registers[26][15] ,
         \Reg_Bank/registers[26][16] , \Reg_Bank/registers[26][17] ,
         \Reg_Bank/registers[26][18] , \Reg_Bank/registers[26][19] ,
         \Reg_Bank/registers[26][20] , \Reg_Bank/registers[26][21] ,
         \Reg_Bank/registers[26][22] , \Reg_Bank/registers[26][23] ,
         \Reg_Bank/registers[26][24] , \Reg_Bank/registers[26][25] ,
         \Reg_Bank/registers[26][26] , \Reg_Bank/registers[26][27] ,
         \Reg_Bank/registers[26][28] , \Reg_Bank/registers[26][29] ,
         \Reg_Bank/registers[26][30] , \Reg_Bank/registers[26][31] ,
         \Reg_Bank/registers[27][0] , \Reg_Bank/registers[27][1] ,
         \Reg_Bank/registers[27][2] , \Reg_Bank/registers[27][3] ,
         \Reg_Bank/registers[27][4] , \Reg_Bank/registers[27][5] ,
         \Reg_Bank/registers[27][6] , \Reg_Bank/registers[27][7] ,
         \Reg_Bank/registers[27][8] , \Reg_Bank/registers[27][9] ,
         \Reg_Bank/registers[27][10] , \Reg_Bank/registers[27][11] ,
         \Reg_Bank/registers[27][12] , \Reg_Bank/registers[27][13] ,
         \Reg_Bank/registers[27][14] , \Reg_Bank/registers[27][15] ,
         \Reg_Bank/registers[27][16] , \Reg_Bank/registers[27][17] ,
         \Reg_Bank/registers[27][18] , \Reg_Bank/registers[27][19] ,
         \Reg_Bank/registers[27][20] , \Reg_Bank/registers[27][21] ,
         \Reg_Bank/registers[27][22] , \Reg_Bank/registers[27][23] ,
         \Reg_Bank/registers[27][24] , \Reg_Bank/registers[27][25] ,
         \Reg_Bank/registers[27][26] , \Reg_Bank/registers[27][27] ,
         \Reg_Bank/registers[27][28] , \Reg_Bank/registers[27][29] ,
         \Reg_Bank/registers[27][30] , \Reg_Bank/registers[27][31] ,
         \Reg_Bank/registers[28][0] , \Reg_Bank/registers[28][1] ,
         \Reg_Bank/registers[28][2] , \Reg_Bank/registers[28][3] ,
         \Reg_Bank/registers[28][4] , \Reg_Bank/registers[28][5] ,
         \Reg_Bank/registers[28][6] , \Reg_Bank/registers[28][7] ,
         \Reg_Bank/registers[28][8] , \Reg_Bank/registers[28][9] ,
         \Reg_Bank/registers[28][10] , \Reg_Bank/registers[28][11] ,
         \Reg_Bank/registers[28][12] , \Reg_Bank/registers[28][13] ,
         \Reg_Bank/registers[28][14] , \Reg_Bank/registers[28][15] ,
         \Reg_Bank/registers[28][16] , \Reg_Bank/registers[28][17] ,
         \Reg_Bank/registers[28][18] , \Reg_Bank/registers[28][19] ,
         \Reg_Bank/registers[28][20] , \Reg_Bank/registers[28][21] ,
         \Reg_Bank/registers[28][22] , \Reg_Bank/registers[28][23] ,
         \Reg_Bank/registers[28][24] , \Reg_Bank/registers[28][25] ,
         \Reg_Bank/registers[28][26] , \Reg_Bank/registers[28][27] ,
         \Reg_Bank/registers[28][28] , \Reg_Bank/registers[28][29] ,
         \Reg_Bank/registers[28][30] , \Reg_Bank/registers[28][31] ,
         \Reg_Bank/registers[29][0] , \Reg_Bank/registers[29][1] ,
         \Reg_Bank/registers[29][2] , \Reg_Bank/registers[29][3] ,
         \Reg_Bank/registers[29][4] , \Reg_Bank/registers[29][5] ,
         \Reg_Bank/registers[29][6] , \Reg_Bank/registers[29][7] ,
         \Reg_Bank/registers[29][8] , \Reg_Bank/registers[29][9] ,
         \Reg_Bank/registers[29][10] , \Reg_Bank/registers[29][11] ,
         \Reg_Bank/registers[29][12] , \Reg_Bank/registers[29][13] ,
         \Reg_Bank/registers[29][14] , \Reg_Bank/registers[29][15] ,
         \Reg_Bank/registers[29][16] , \Reg_Bank/registers[29][17] ,
         \Reg_Bank/registers[29][18] , \Reg_Bank/registers[29][19] ,
         \Reg_Bank/registers[29][20] , \Reg_Bank/registers[29][21] ,
         \Reg_Bank/registers[29][22] , \Reg_Bank/registers[29][23] ,
         \Reg_Bank/registers[29][24] , \Reg_Bank/registers[29][25] ,
         \Reg_Bank/registers[29][26] , \Reg_Bank/registers[29][27] ,
         \Reg_Bank/registers[29][28] , \Reg_Bank/registers[29][29] ,
         \Reg_Bank/registers[29][30] , \Reg_Bank/registers[29][31] ,
         \Reg_Bank/registers[30][0] , \Reg_Bank/registers[30][1] ,
         \Reg_Bank/registers[30][2] , \Reg_Bank/registers[30][3] ,
         \Reg_Bank/registers[30][4] , \Reg_Bank/registers[30][5] ,
         \Reg_Bank/registers[30][6] , \Reg_Bank/registers[30][7] ,
         \Reg_Bank/registers[30][8] , \Reg_Bank/registers[30][9] ,
         \Reg_Bank/registers[30][10] , \Reg_Bank/registers[30][11] ,
         \Reg_Bank/registers[30][12] , \Reg_Bank/registers[30][13] ,
         \Reg_Bank/registers[30][14] , \Reg_Bank/registers[30][15] ,
         \Reg_Bank/registers[30][16] , \Reg_Bank/registers[30][17] ,
         \Reg_Bank/registers[30][18] , \Reg_Bank/registers[30][19] ,
         \Reg_Bank/registers[30][20] , \Reg_Bank/registers[30][21] ,
         \Reg_Bank/registers[30][22] , \Reg_Bank/registers[30][23] ,
         \Reg_Bank/registers[30][24] , \Reg_Bank/registers[30][25] ,
         \Reg_Bank/registers[30][26] , \Reg_Bank/registers[30][27] ,
         \Reg_Bank/registers[30][28] , \Reg_Bank/registers[30][29] ,
         \Reg_Bank/registers[30][30] , \Reg_Bank/registers[30][31] ,
         \Reg_Bank/registers[31][0] , \Reg_Bank/registers[31][1] ,
         \Reg_Bank/registers[31][2] , \Reg_Bank/registers[31][3] ,
         \Reg_Bank/registers[31][4] , \Reg_Bank/registers[31][5] ,
         \Reg_Bank/registers[31][6] , \Reg_Bank/registers[31][7] ,
         \Reg_Bank/registers[31][8] , \Reg_Bank/registers[31][9] ,
         \Reg_Bank/registers[31][10] , \Reg_Bank/registers[31][11] ,
         \Reg_Bank/registers[31][12] , \Reg_Bank/registers[31][13] ,
         \Reg_Bank/registers[31][14] , \Reg_Bank/registers[31][15] ,
         \Reg_Bank/registers[31][16] , \Reg_Bank/registers[31][17] ,
         \Reg_Bank/registers[31][18] , \Reg_Bank/registers[31][19] ,
         \Reg_Bank/registers[31][20] , \Reg_Bank/registers[31][21] ,
         \Reg_Bank/registers[31][22] , \Reg_Bank/registers[31][23] ,
         \Reg_Bank/registers[31][24] , \Reg_Bank/registers[31][25] ,
         \Reg_Bank/registers[31][26] , \Reg_Bank/registers[31][27] ,
         \Reg_Bank/registers[31][28] , \Reg_Bank/registers[31][29] ,
         \Reg_Bank/registers[31][30] , \Reg_Bank/registers[31][31] ,
         \ALU/U2/U1/Z_0 , \ALU/N139 , \ALU/N138 , \ALU/N137 , \ALU/N136 ,
         \ALU/N135 , \ALU/N134 , \ALU/N133 , \ALU/N132 , \ALU/N131 ,
         \ALU/N130 , \ALU/N129 , \ALU/N128 , \ALU/N127 , \ALU/N126 ,
         \ALU/N125 , \ALU/N124 , \ALU/N123 , \ALU/N122 , \ALU/N121 ,
         \ALU/N120 , \ALU/N119 , \ALU/N118 , \ALU/N117 , \ALU/N116 ,
         \ALU/N115 , \ALU/N114 , \ALU/N113 , \ALU/N112 , \ALU/N111 ,
         \ALU/N110 , \ALU/N109 , \ALU/N108 , \Shifter/N75 ,
         \Shifter/sll_27/ML_int[5][16] , \Shifter/sll_27/ML_int[5][17] ,
         \Shifter/sll_27/ML_int[5][18] , \Shifter/sll_27/ML_int[5][19] ,
         \Shifter/sll_27/ML_int[5][20] , \Shifter/sll_27/ML_int[5][21] ,
         \Shifter/sll_27/ML_int[5][22] , \Shifter/sll_27/ML_int[5][23] ,
         \Shifter/sll_27/ML_int[5][24] , \Shifter/sll_27/ML_int[5][25] ,
         \Shifter/sll_27/ML_int[5][26] , \Shifter/sll_27/ML_int[5][27] ,
         \Shifter/sll_27/ML_int[5][28] , \Shifter/sll_27/ML_int[5][29] ,
         \Shifter/sll_27/ML_int[5][30] , \Shifter/sll_27/ML_int[5][31] ,
         \Shifter/sll_27/ML_int[4][0] , \Shifter/sll_27/ML_int[4][1] ,
         \Shifter/sll_27/ML_int[4][2] , \Shifter/sll_27/ML_int[4][3] ,
         \Shifter/sll_27/ML_int[4][4] , \Shifter/sll_27/ML_int[4][5] ,
         \Shifter/sll_27/ML_int[4][6] , \Shifter/sll_27/ML_int[4][7] ,
         \Shifter/sll_27/ML_int[4][8] , \Shifter/sll_27/ML_int[4][9] ,
         \Shifter/sll_27/ML_int[4][10] , \Shifter/sll_27/ML_int[4][11] ,
         \Shifter/sll_27/ML_int[4][12] , \Shifter/sll_27/ML_int[4][13] ,
         \Shifter/sll_27/ML_int[4][14] , \Shifter/sll_27/ML_int[4][15] ,
         \Shifter/sll_27/ML_int[4][16] , \Shifter/sll_27/ML_int[4][17] ,
         \Shifter/sll_27/ML_int[4][18] , \Shifter/sll_27/ML_int[4][19] ,
         \Shifter/sll_27/ML_int[4][20] , \Shifter/sll_27/ML_int[4][21] ,
         \Shifter/sll_27/ML_int[4][22] , \Shifter/sll_27/ML_int[4][23] ,
         \Shifter/sll_27/ML_int[4][24] , \Shifter/sll_27/ML_int[4][25] ,
         \Shifter/sll_27/ML_int[4][26] , \Shifter/sll_27/ML_int[4][27] ,
         \Shifter/sll_27/ML_int[4][28] , \Shifter/sll_27/ML_int[4][29] ,
         \Shifter/sll_27/ML_int[4][30] , \Shifter/sll_27/ML_int[4][31] ,
         \Shifter/sll_27/ML_int[3][0] , \Shifter/sll_27/ML_int[3][1] ,
         \Shifter/sll_27/ML_int[3][2] , \Shifter/sll_27/ML_int[3][3] ,
         \Shifter/sll_27/ML_int[3][4] , \Shifter/sll_27/ML_int[3][5] ,
         \Shifter/sll_27/ML_int[3][6] , \Shifter/sll_27/ML_int[3][7] ,
         \Shifter/sll_27/ML_int[3][8] , \Shifter/sll_27/ML_int[3][9] ,
         \Shifter/sll_27/ML_int[3][10] , \Shifter/sll_27/ML_int[3][11] ,
         \Shifter/sll_27/ML_int[3][12] , \Shifter/sll_27/ML_int[3][13] ,
         \Shifter/sll_27/ML_int[3][14] , \Shifter/sll_27/ML_int[3][15] ,
         \Shifter/sll_27/ML_int[3][16] , \Shifter/sll_27/ML_int[3][17] ,
         \Shifter/sll_27/ML_int[3][18] , \Shifter/sll_27/ML_int[3][19] ,
         \Shifter/sll_27/ML_int[3][20] , \Shifter/sll_27/ML_int[3][21] ,
         \Shifter/sll_27/ML_int[3][22] , \Shifter/sll_27/ML_int[3][23] ,
         \Shifter/sll_27/ML_int[3][24] , \Shifter/sll_27/ML_int[3][25] ,
         \Shifter/sll_27/ML_int[3][26] , \Shifter/sll_27/ML_int[3][27] ,
         \Shifter/sll_27/ML_int[3][28] , \Shifter/sll_27/ML_int[3][29] ,
         \Shifter/sll_27/ML_int[3][30] , \Shifter/sll_27/ML_int[3][31] ,
         \Shifter/sll_27/ML_int[2][0] , \Shifter/sll_27/ML_int[2][1] ,
         \Shifter/sll_27/ML_int[2][2] , \Shifter/sll_27/ML_int[2][3] ,
         \Shifter/sll_27/ML_int[2][4] , \Shifter/sll_27/ML_int[2][5] ,
         \Shifter/sll_27/ML_int[2][6] , \Shifter/sll_27/ML_int[2][7] ,
         \Shifter/sll_27/ML_int[2][8] , \Shifter/sll_27/ML_int[2][9] ,
         \Shifter/sll_27/ML_int[2][10] , \Shifter/sll_27/ML_int[2][11] ,
         \Shifter/sll_27/ML_int[2][12] , \Shifter/sll_27/ML_int[2][13] ,
         \Shifter/sll_27/ML_int[2][14] , \Shifter/sll_27/ML_int[2][15] ,
         \Shifter/sll_27/ML_int[2][16] , \Shifter/sll_27/ML_int[2][17] ,
         \Shifter/sll_27/ML_int[2][18] , \Shifter/sll_27/ML_int[2][19] ,
         \Shifter/sll_27/ML_int[2][20] , \Shifter/sll_27/ML_int[2][21] ,
         \Shifter/sll_27/ML_int[2][22] , \Shifter/sll_27/ML_int[2][23] ,
         \Shifter/sll_27/ML_int[2][24] , \Shifter/sll_27/ML_int[2][25] ,
         \Shifter/sll_27/ML_int[2][26] , \Shifter/sll_27/ML_int[2][27] ,
         \Shifter/sll_27/ML_int[2][28] , \Shifter/sll_27/ML_int[2][29] ,
         \Shifter/sll_27/ML_int[2][30] , \Shifter/sll_27/ML_int[2][31] ,
         \Shifter/sll_27/ML_int[1][0] , \Shifter/sll_27/ML_int[1][1] ,
         \Shifter/sll_27/ML_int[1][2] , \Shifter/sll_27/ML_int[1][3] ,
         \Shifter/sll_27/ML_int[1][4] , \Shifter/sll_27/ML_int[1][5] ,
         \Shifter/sll_27/ML_int[1][6] , \Shifter/sll_27/ML_int[1][7] ,
         \Shifter/sll_27/ML_int[1][8] , \Shifter/sll_27/ML_int[1][9] ,
         \Shifter/sll_27/ML_int[1][10] , \Shifter/sll_27/ML_int[1][11] ,
         \Shifter/sll_27/ML_int[1][12] , \Shifter/sll_27/ML_int[1][13] ,
         \Shifter/sll_27/ML_int[1][14] , \Shifter/sll_27/ML_int[1][15] ,
         \Shifter/sll_27/ML_int[1][16] , \Shifter/sll_27/ML_int[1][17] ,
         \Shifter/sll_27/ML_int[1][18] , \Shifter/sll_27/ML_int[1][19] ,
         \Shifter/sll_27/ML_int[1][20] , \Shifter/sll_27/ML_int[1][21] ,
         \Shifter/sll_27/ML_int[1][22] , \Shifter/sll_27/ML_int[1][23] ,
         \Shifter/sll_27/ML_int[1][24] , \Shifter/sll_27/ML_int[1][25] ,
         \Shifter/sll_27/ML_int[1][26] , \Shifter/sll_27/ML_int[1][27] ,
         \Shifter/sll_27/ML_int[1][28] , \Shifter/sll_27/ML_int[1][29] ,
         \Shifter/sll_27/ML_int[1][30] , \Shifter/sll_27/ML_int[1][31] ,
         \ALU/r67/B_AS[31] , \ALU/r67/B_AS[30] , \ALU/r67/B_AS[29] ,
         \ALU/r67/B_AS[28] , \ALU/r67/B_AS[27] , \ALU/r67/B_AS[26] ,
         \ALU/r67/B_AS[25] , \ALU/r67/B_AS[24] , \ALU/r67/B_AS[23] ,
         \ALU/r67/B_AS[22] , \ALU/r67/B_AS[21] , \ALU/r67/B_AS[20] ,
         \ALU/r67/B_AS[19] , \ALU/r67/B_AS[18] , \ALU/r67/B_AS[17] ,
         \ALU/r67/B_AS[16] , \ALU/r67/B_AS[15] , \ALU/r67/B_AS[14] ,
         \ALU/r67/B_AS[13] , \ALU/r67/B_AS[12] , \ALU/r67/B_AS[11] ,
         \ALU/r67/B_AS[10] , \ALU/r67/B_AS[9] , \ALU/r67/B_AS[8] ,
         \ALU/r67/B_AS[7] , \ALU/r67/B_AS[6] , \ALU/r67/B_AS[5] ,
         \ALU/r67/B_AS[4] , \ALU/r67/B_AS[3] , \ALU/r67/B_AS[2] ,
         \ALU/r67/B_AS[1] , \ALU/r67/B_AS[0] , \ALU/r67/carry[1] ,
         \ALU/r67/carry[2] , \ALU/r67/carry[3] , \ALU/r67/carry[4] ,
         \ALU/r67/carry[5] , \ALU/r67/carry[6] , \ALU/r67/carry[7] ,
         \ALU/r67/carry[8] , \ALU/r67/carry[9] , \ALU/r67/carry[10] ,
         \ALU/r67/carry[11] , \ALU/r67/carry[12] , \ALU/r67/carry[13] ,
         \ALU/r67/carry[14] , \ALU/r67/carry[15] , \ALU/r67/carry[16] ,
         \ALU/r67/carry[17] , \ALU/r67/carry[18] , \ALU/r67/carry[19] ,
         \ALU/r67/carry[20] , \ALU/r67/carry[21] , \ALU/r67/carry[22] ,
         \ALU/r67/carry[23] , \ALU/r67/carry[24] , \ALU/r67/carry[25] ,
         \ALU/r67/carry[26] , \ALU/r67/carry[27] , \ALU/r67/carry[28] ,
         \ALU/r67/carry[29] , \ALU/r67/carry[30] , \ALU/r67/carry[31] ,
         \PC_Next/add_30/carry[29] , \PC_Next/add_30/carry[28] ,
         \PC_Next/add_30/carry[27] , \PC_Next/add_30/carry[26] ,
         \PC_Next/add_30/carry[25] , \PC_Next/add_30/carry[24] ,
         \PC_Next/add_30/carry[23] , \PC_Next/add_30/carry[22] ,
         \PC_Next/add_30/carry[21] , \PC_Next/add_30/carry[20] ,
         \PC_Next/add_30/carry[19] , \PC_Next/add_30/carry[18] ,
         \PC_Next/add_30/carry[17] , \PC_Next/add_30/carry[16] ,
         \PC_Next/add_30/carry[15] , \PC_Next/add_30/carry[14] ,
         \PC_Next/add_30/carry[13] , \PC_Next/add_30/carry[12] ,
         \PC_Next/add_30/carry[11] , \PC_Next/add_30/carry[10] ,
         \PC_Next/add_30/carry[9] , \PC_Next/add_30/carry[8] ,
         \PC_Next/add_30/carry[7] , \PC_Next/add_30/carry[6] ,
         \PC_Next/add_30/carry[5] , \PC_Next/add_30/carry[4] ,
         \PC_Next/add_30/carry[3] , \PC_Next/add_30/carry[2] ,
         \PC_Next/add_41/carry[29] , \PC_Next/add_41/carry[28] ,
         \PC_Next/add_41/carry[27] , \PC_Next/add_41/carry[26] ,
         \PC_Next/add_41/carry[25] , \PC_Next/add_41/carry[24] ,
         \PC_Next/add_41/carry[23] , \PC_Next/add_41/carry[22] ,
         \PC_Next/add_41/carry[21] , \PC_Next/add_41/carry[20] ,
         \PC_Next/add_41/carry[19] , \PC_Next/add_41/carry[18] ,
         \PC_Next/add_41/carry[17] , \PC_Next/add_41/carry[16] ,
         \PC_Next/add_41/carry[15] , \PC_Next/add_41/carry[14] ,
         \PC_Next/add_41/carry[13] , \PC_Next/add_41/carry[12] ,
         \PC_Next/add_41/carry[11] , \PC_Next/add_41/carry[10] ,
         \PC_Next/add_41/carry[9] , \PC_Next/add_41/carry[8] ,
         \PC_Next/add_41/carry[7] , \PC_Next/add_41/carry[6] ,
         \PC_Next/add_41/carry[5] , \PC_Next/add_41/carry[4] ,
         \PC_Next/add_41/carry[3] , \PC_Next/add_41/carry[2] ,
         \PC_Next/add_41/carry[1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507;
  wire   [31:0] opcode;
  wire   [31:2] pc_current;
  wire   [31:2] pc_plus4;
  wire   [31:0] reg_target;
  wire   [31:0] c_memory;
  wire   [4:0] rs_index;
  wire   [4:0] rt_index;
  wire   [15:0] imm;
  wire   [31:0] reg_source;
  wire   [31:0] a_bus;
  wire   [31:0] b_bus;

  DFF \PC_Next/pc_reg[30]  ( .D(\PC_Next/n309 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[30]) );
  DFF \PC_Next/pc_reg[29]  ( .D(\PC_Next/n310 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[29]) );
  DFF \PC_Next/pc_reg[28]  ( .D(\PC_Next/n311 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[28]) );
  DFF \PC_Next/pc_reg[27]  ( .D(\PC_Next/pc_future[27] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[27]) );
  DFF \PC_Next/pc_reg[26]  ( .D(\PC_Next/pc_future[26] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[26]) );
  DFF \PC_Next/pc_reg[25]  ( .D(\PC_Next/pc_future[25] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[25]) );
  DFF \PC_Next/pc_reg[24]  ( .D(\PC_Next/pc_future[24] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[24]) );
  DFF \PC_Next/pc_reg[23]  ( .D(\PC_Next/pc_future[23] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[23]) );
  DFF \PC_Next/pc_reg[22]  ( .D(\PC_Next/pc_future[22] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[22]) );
  DFF \PC_Next/pc_reg[21]  ( .D(\PC_Next/pc_future[21] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[21]) );
  DFF \PC_Next/pc_reg[20]  ( .D(\PC_Next/pc_future[20] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[20]) );
  DFF \PC_Next/pc_reg[19]  ( .D(\PC_Next/pc_future[19] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[19]) );
  DFF \PC_Next/pc_reg[18]  ( .D(\PC_Next/pc_future[18] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[18]) );
  DFF \PC_Next/pc_reg[17]  ( .D(\PC_Next/pc_future[17] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[17]) );
  DFF \PC_Next/pc_reg[16]  ( .D(\PC_Next/pc_future[16] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[16]) );
  DFF \PC_Next/pc_reg[15]  ( .D(\PC_Next/pc_future[15] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[15]) );
  DFF \PC_Next/pc_reg[14]  ( .D(\PC_Next/pc_future[14] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[14]) );
  DFF \PC_Next/pc_reg[13]  ( .D(\PC_Next/pc_future[13] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[13]) );
  DFF \PC_Next/pc_reg[12]  ( .D(\PC_Next/pc_future[12] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[12]) );
  DFF \PC_Next/pc_reg[11]  ( .D(\PC_Next/pc_future[11] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[11]) );
  DFF \PC_Next/pc_reg[10]  ( .D(\PC_Next/pc_future[10] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[10]) );
  DFF \PC_Next/pc_reg[9]  ( .D(\PC_Next/pc_future[9] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[9]) );
  DFF \PC_Next/pc_reg[8]  ( .D(\PC_Next/pc_future[8] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[8]) );
  DFF \PC_Next/pc_reg[7]  ( .D(\PC_Next/pc_future[7] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[7]) );
  DFF \PC_Next/pc_reg[6]  ( .D(\PC_Next/pc_future[6] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[6]) );
  DFF \PC_Next/pc_reg[5]  ( .D(\PC_Next/pc_future[5] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[5]) );
  DFF \PC_Next/pc_reg[4]  ( .D(\PC_Next/pc_future[4] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[4]) );
  DFF \PC_Next/pc_reg[3]  ( .D(\PC_Next/pc_future[3] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[3]) );
  DFF \PC_Next/pc_reg[31]  ( .D(\PC_Next/n308 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[31]) );
  DFF \PC_Next/pc_reg[2]  ( .D(\PC_Next/pc_future[2] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[2]) );
  MUX \Inst_Mem/U2016  ( .A(\Inst_Mem/n1984 ), .B(\Inst_Mem/n1953 ), .S(
        pc_current[7]), .Z(opcode[31]) );
  MUX \Inst_Mem/U2015  ( .A(\Inst_Mem/n1983 ), .B(\Inst_Mem/n1968 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1984 ) );
  MUX \Inst_Mem/U2014  ( .A(\Inst_Mem/n1982 ), .B(\Inst_Mem/n1975 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1983 ) );
  MUX \Inst_Mem/U2013  ( .A(\Inst_Mem/n1981 ), .B(\Inst_Mem/n1978 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1982 ) );
  MUX \Inst_Mem/U2012  ( .A(\Inst_Mem/n1980 ), .B(\Inst_Mem/n1979 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1981 ) );
  MUX \Inst_Mem/U2011  ( .A(inst_mem_in_wire[31]), .B(inst_mem_in_wire[63]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1980 ) );
  MUX \Inst_Mem/U2010  ( .A(inst_mem_in_wire[95]), .B(inst_mem_in_wire[127]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1979 ) );
  MUX \Inst_Mem/U2009  ( .A(\Inst_Mem/n1977 ), .B(\Inst_Mem/n1976 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1978 ) );
  MUX \Inst_Mem/U2008  ( .A(inst_mem_in_wire[159]), .B(inst_mem_in_wire[191]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1977 ) );
  MUX \Inst_Mem/U2007  ( .A(inst_mem_in_wire[223]), .B(inst_mem_in_wire[255]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1976 ) );
  MUX \Inst_Mem/U2006  ( .A(\Inst_Mem/n1974 ), .B(\Inst_Mem/n1971 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1975 ) );
  MUX \Inst_Mem/U2005  ( .A(\Inst_Mem/n1973 ), .B(\Inst_Mem/n1972 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1974 ) );
  MUX \Inst_Mem/U2004  ( .A(inst_mem_in_wire[287]), .B(inst_mem_in_wire[319]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1973 ) );
  MUX \Inst_Mem/U2003  ( .A(inst_mem_in_wire[351]), .B(inst_mem_in_wire[383]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1972 ) );
  MUX \Inst_Mem/U2002  ( .A(\Inst_Mem/n1970 ), .B(\Inst_Mem/n1969 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1971 ) );
  MUX \Inst_Mem/U2001  ( .A(inst_mem_in_wire[415]), .B(inst_mem_in_wire[447]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1970 ) );
  MUX \Inst_Mem/U2000  ( .A(inst_mem_in_wire[479]), .B(inst_mem_in_wire[511]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1969 ) );
  MUX \Inst_Mem/U1999  ( .A(\Inst_Mem/n1967 ), .B(\Inst_Mem/n1960 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1968 ) );
  MUX \Inst_Mem/U1998  ( .A(\Inst_Mem/n1966 ), .B(\Inst_Mem/n1963 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1967 ) );
  MUX \Inst_Mem/U1997  ( .A(\Inst_Mem/n1965 ), .B(\Inst_Mem/n1964 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1966 ) );
  MUX \Inst_Mem/U1996  ( .A(inst_mem_in_wire[543]), .B(inst_mem_in_wire[575]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1965 ) );
  MUX \Inst_Mem/U1995  ( .A(inst_mem_in_wire[607]), .B(inst_mem_in_wire[639]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1964 ) );
  MUX \Inst_Mem/U1994  ( .A(\Inst_Mem/n1962 ), .B(\Inst_Mem/n1961 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1963 ) );
  MUX \Inst_Mem/U1993  ( .A(inst_mem_in_wire[671]), .B(inst_mem_in_wire[703]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1962 ) );
  MUX \Inst_Mem/U1992  ( .A(inst_mem_in_wire[735]), .B(inst_mem_in_wire[767]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1961 ) );
  MUX \Inst_Mem/U1991  ( .A(\Inst_Mem/n1959 ), .B(\Inst_Mem/n1956 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1960 ) );
  MUX \Inst_Mem/U1990  ( .A(\Inst_Mem/n1958 ), .B(\Inst_Mem/n1957 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1959 ) );
  MUX \Inst_Mem/U1989  ( .A(inst_mem_in_wire[799]), .B(inst_mem_in_wire[831]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1958 ) );
  MUX \Inst_Mem/U1988  ( .A(inst_mem_in_wire[863]), .B(inst_mem_in_wire[895]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1957 ) );
  MUX \Inst_Mem/U1987  ( .A(\Inst_Mem/n1955 ), .B(\Inst_Mem/n1954 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1956 ) );
  MUX \Inst_Mem/U1986  ( .A(inst_mem_in_wire[927]), .B(inst_mem_in_wire[959]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1955 ) );
  MUX \Inst_Mem/U1985  ( .A(inst_mem_in_wire[991]), .B(inst_mem_in_wire[1023]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1954 ) );
  MUX \Inst_Mem/U1984  ( .A(\Inst_Mem/n1952 ), .B(\Inst_Mem/n1937 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1953 ) );
  MUX \Inst_Mem/U1983  ( .A(\Inst_Mem/n1951 ), .B(\Inst_Mem/n1944 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1952 ) );
  MUX \Inst_Mem/U1982  ( .A(\Inst_Mem/n1950 ), .B(\Inst_Mem/n1947 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1951 ) );
  MUX \Inst_Mem/U1981  ( .A(\Inst_Mem/n1949 ), .B(\Inst_Mem/n1948 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1950 ) );
  MUX \Inst_Mem/U1980  ( .A(inst_mem_in_wire[1055]), .B(inst_mem_in_wire[1087]), .S(pc_current[2]), .Z(\Inst_Mem/n1949 ) );
  MUX \Inst_Mem/U1979  ( .A(inst_mem_in_wire[1119]), .B(inst_mem_in_wire[1151]), .S(pc_current[2]), .Z(\Inst_Mem/n1948 ) );
  MUX \Inst_Mem/U1978  ( .A(\Inst_Mem/n1946 ), .B(\Inst_Mem/n1945 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1947 ) );
  MUX \Inst_Mem/U1977  ( .A(inst_mem_in_wire[1183]), .B(inst_mem_in_wire[1215]), .S(pc_current[2]), .Z(\Inst_Mem/n1946 ) );
  MUX \Inst_Mem/U1976  ( .A(inst_mem_in_wire[1247]), .B(inst_mem_in_wire[1279]), .S(pc_current[2]), .Z(\Inst_Mem/n1945 ) );
  MUX \Inst_Mem/U1975  ( .A(\Inst_Mem/n1943 ), .B(\Inst_Mem/n1940 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1944 ) );
  MUX \Inst_Mem/U1974  ( .A(\Inst_Mem/n1942 ), .B(\Inst_Mem/n1941 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1943 ) );
  MUX \Inst_Mem/U1973  ( .A(inst_mem_in_wire[1311]), .B(inst_mem_in_wire[1343]), .S(pc_current[2]), .Z(\Inst_Mem/n1942 ) );
  MUX \Inst_Mem/U1972  ( .A(inst_mem_in_wire[1375]), .B(inst_mem_in_wire[1407]), .S(pc_current[2]), .Z(\Inst_Mem/n1941 ) );
  MUX \Inst_Mem/U1971  ( .A(\Inst_Mem/n1939 ), .B(\Inst_Mem/n1938 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1940 ) );
  MUX \Inst_Mem/U1970  ( .A(inst_mem_in_wire[1439]), .B(inst_mem_in_wire[1471]), .S(pc_current[2]), .Z(\Inst_Mem/n1939 ) );
  MUX \Inst_Mem/U1969  ( .A(inst_mem_in_wire[1503]), .B(inst_mem_in_wire[1535]), .S(pc_current[2]), .Z(\Inst_Mem/n1938 ) );
  MUX \Inst_Mem/U1968  ( .A(\Inst_Mem/n1936 ), .B(\Inst_Mem/n1929 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1937 ) );
  MUX \Inst_Mem/U1967  ( .A(\Inst_Mem/n1935 ), .B(\Inst_Mem/n1932 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1936 ) );
  MUX \Inst_Mem/U1966  ( .A(\Inst_Mem/n1934 ), .B(\Inst_Mem/n1933 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1935 ) );
  MUX \Inst_Mem/U1965  ( .A(inst_mem_in_wire[1567]), .B(inst_mem_in_wire[1599]), .S(pc_current[2]), .Z(\Inst_Mem/n1934 ) );
  MUX \Inst_Mem/U1964  ( .A(inst_mem_in_wire[1631]), .B(inst_mem_in_wire[1663]), .S(pc_current[2]), .Z(\Inst_Mem/n1933 ) );
  MUX \Inst_Mem/U1963  ( .A(\Inst_Mem/n1931 ), .B(\Inst_Mem/n1930 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1932 ) );
  MUX \Inst_Mem/U1962  ( .A(inst_mem_in_wire[1695]), .B(inst_mem_in_wire[1727]), .S(pc_current[2]), .Z(\Inst_Mem/n1931 ) );
  MUX \Inst_Mem/U1961  ( .A(inst_mem_in_wire[1759]), .B(inst_mem_in_wire[1791]), .S(pc_current[2]), .Z(\Inst_Mem/n1930 ) );
  MUX \Inst_Mem/U1960  ( .A(\Inst_Mem/n1928 ), .B(\Inst_Mem/n1925 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1929 ) );
  MUX \Inst_Mem/U1959  ( .A(\Inst_Mem/n1927 ), .B(\Inst_Mem/n1926 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1928 ) );
  MUX \Inst_Mem/U1958  ( .A(inst_mem_in_wire[1823]), .B(inst_mem_in_wire[1855]), .S(pc_current[2]), .Z(\Inst_Mem/n1927 ) );
  MUX \Inst_Mem/U1957  ( .A(inst_mem_in_wire[1887]), .B(inst_mem_in_wire[1919]), .S(pc_current[2]), .Z(\Inst_Mem/n1926 ) );
  MUX \Inst_Mem/U1956  ( .A(\Inst_Mem/n1924 ), .B(\Inst_Mem/n1923 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1925 ) );
  MUX \Inst_Mem/U1955  ( .A(inst_mem_in_wire[1951]), .B(inst_mem_in_wire[1983]), .S(pc_current[2]), .Z(\Inst_Mem/n1924 ) );
  MUX \Inst_Mem/U1954  ( .A(inst_mem_in_wire[2015]), .B(inst_mem_in_wire[2047]), .S(pc_current[2]), .Z(\Inst_Mem/n1923 ) );
  MUX \Inst_Mem/U1953  ( .A(\Inst_Mem/n1922 ), .B(\Inst_Mem/n1891 ), .S(
        pc_current[7]), .Z(opcode[30]) );
  MUX \Inst_Mem/U1952  ( .A(\Inst_Mem/n1921 ), .B(\Inst_Mem/n1906 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1922 ) );
  MUX \Inst_Mem/U1951  ( .A(\Inst_Mem/n1920 ), .B(\Inst_Mem/n1913 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1921 ) );
  MUX \Inst_Mem/U1950  ( .A(\Inst_Mem/n1919 ), .B(\Inst_Mem/n1916 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1920 ) );
  MUX \Inst_Mem/U1949  ( .A(\Inst_Mem/n1918 ), .B(\Inst_Mem/n1917 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1919 ) );
  MUX \Inst_Mem/U1948  ( .A(inst_mem_in_wire[30]), .B(inst_mem_in_wire[62]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1918 ) );
  MUX \Inst_Mem/U1947  ( .A(inst_mem_in_wire[94]), .B(inst_mem_in_wire[126]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1917 ) );
  MUX \Inst_Mem/U1946  ( .A(\Inst_Mem/n1915 ), .B(\Inst_Mem/n1914 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1916 ) );
  MUX \Inst_Mem/U1945  ( .A(inst_mem_in_wire[158]), .B(inst_mem_in_wire[190]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1915 ) );
  MUX \Inst_Mem/U1944  ( .A(inst_mem_in_wire[222]), .B(inst_mem_in_wire[254]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1914 ) );
  MUX \Inst_Mem/U1943  ( .A(\Inst_Mem/n1912 ), .B(\Inst_Mem/n1909 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1913 ) );
  MUX \Inst_Mem/U1942  ( .A(\Inst_Mem/n1911 ), .B(\Inst_Mem/n1910 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1912 ) );
  MUX \Inst_Mem/U1941  ( .A(inst_mem_in_wire[286]), .B(inst_mem_in_wire[318]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1911 ) );
  MUX \Inst_Mem/U1940  ( .A(inst_mem_in_wire[350]), .B(inst_mem_in_wire[382]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1910 ) );
  MUX \Inst_Mem/U1939  ( .A(\Inst_Mem/n1908 ), .B(\Inst_Mem/n1907 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1909 ) );
  MUX \Inst_Mem/U1938  ( .A(inst_mem_in_wire[414]), .B(inst_mem_in_wire[446]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1908 ) );
  MUX \Inst_Mem/U1937  ( .A(inst_mem_in_wire[478]), .B(inst_mem_in_wire[510]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1907 ) );
  MUX \Inst_Mem/U1936  ( .A(\Inst_Mem/n1905 ), .B(\Inst_Mem/n1898 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1906 ) );
  MUX \Inst_Mem/U1935  ( .A(\Inst_Mem/n1904 ), .B(\Inst_Mem/n1901 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1905 ) );
  MUX \Inst_Mem/U1934  ( .A(\Inst_Mem/n1903 ), .B(\Inst_Mem/n1902 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1904 ) );
  MUX \Inst_Mem/U1933  ( .A(inst_mem_in_wire[542]), .B(inst_mem_in_wire[574]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1903 ) );
  MUX \Inst_Mem/U1932  ( .A(inst_mem_in_wire[606]), .B(inst_mem_in_wire[638]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1902 ) );
  MUX \Inst_Mem/U1931  ( .A(\Inst_Mem/n1900 ), .B(\Inst_Mem/n1899 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1901 ) );
  MUX \Inst_Mem/U1930  ( .A(inst_mem_in_wire[670]), .B(inst_mem_in_wire[702]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1900 ) );
  MUX \Inst_Mem/U1929  ( .A(inst_mem_in_wire[734]), .B(inst_mem_in_wire[766]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1899 ) );
  MUX \Inst_Mem/U1928  ( .A(\Inst_Mem/n1897 ), .B(\Inst_Mem/n1894 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1898 ) );
  MUX \Inst_Mem/U1927  ( .A(\Inst_Mem/n1896 ), .B(\Inst_Mem/n1895 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1897 ) );
  MUX \Inst_Mem/U1926  ( .A(inst_mem_in_wire[798]), .B(inst_mem_in_wire[830]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1896 ) );
  MUX \Inst_Mem/U1925  ( .A(inst_mem_in_wire[862]), .B(inst_mem_in_wire[894]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1895 ) );
  MUX \Inst_Mem/U1924  ( .A(\Inst_Mem/n1893 ), .B(\Inst_Mem/n1892 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1894 ) );
  MUX \Inst_Mem/U1923  ( .A(inst_mem_in_wire[926]), .B(inst_mem_in_wire[958]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1893 ) );
  MUX \Inst_Mem/U1922  ( .A(inst_mem_in_wire[990]), .B(inst_mem_in_wire[1022]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1892 ) );
  MUX \Inst_Mem/U1921  ( .A(\Inst_Mem/n1890 ), .B(\Inst_Mem/n1875 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1891 ) );
  MUX \Inst_Mem/U1920  ( .A(\Inst_Mem/n1889 ), .B(\Inst_Mem/n1882 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1890 ) );
  MUX \Inst_Mem/U1919  ( .A(\Inst_Mem/n1888 ), .B(\Inst_Mem/n1885 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1889 ) );
  MUX \Inst_Mem/U1918  ( .A(\Inst_Mem/n1887 ), .B(\Inst_Mem/n1886 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1888 ) );
  MUX \Inst_Mem/U1917  ( .A(inst_mem_in_wire[1054]), .B(inst_mem_in_wire[1086]), .S(pc_current[2]), .Z(\Inst_Mem/n1887 ) );
  MUX \Inst_Mem/U1916  ( .A(inst_mem_in_wire[1118]), .B(inst_mem_in_wire[1150]), .S(pc_current[2]), .Z(\Inst_Mem/n1886 ) );
  MUX \Inst_Mem/U1915  ( .A(\Inst_Mem/n1884 ), .B(\Inst_Mem/n1883 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1885 ) );
  MUX \Inst_Mem/U1914  ( .A(inst_mem_in_wire[1182]), .B(inst_mem_in_wire[1214]), .S(pc_current[2]), .Z(\Inst_Mem/n1884 ) );
  MUX \Inst_Mem/U1913  ( .A(inst_mem_in_wire[1246]), .B(inst_mem_in_wire[1278]), .S(pc_current[2]), .Z(\Inst_Mem/n1883 ) );
  MUX \Inst_Mem/U1912  ( .A(\Inst_Mem/n1881 ), .B(\Inst_Mem/n1878 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1882 ) );
  MUX \Inst_Mem/U1911  ( .A(\Inst_Mem/n1880 ), .B(\Inst_Mem/n1879 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1881 ) );
  MUX \Inst_Mem/U1910  ( .A(inst_mem_in_wire[1310]), .B(inst_mem_in_wire[1342]), .S(pc_current[2]), .Z(\Inst_Mem/n1880 ) );
  MUX \Inst_Mem/U1909  ( .A(inst_mem_in_wire[1374]), .B(inst_mem_in_wire[1406]), .S(pc_current[2]), .Z(\Inst_Mem/n1879 ) );
  MUX \Inst_Mem/U1908  ( .A(\Inst_Mem/n1877 ), .B(\Inst_Mem/n1876 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1878 ) );
  MUX \Inst_Mem/U1907  ( .A(inst_mem_in_wire[1438]), .B(inst_mem_in_wire[1470]), .S(pc_current[2]), .Z(\Inst_Mem/n1877 ) );
  MUX \Inst_Mem/U1906  ( .A(inst_mem_in_wire[1502]), .B(inst_mem_in_wire[1534]), .S(pc_current[2]), .Z(\Inst_Mem/n1876 ) );
  MUX \Inst_Mem/U1905  ( .A(\Inst_Mem/n1874 ), .B(\Inst_Mem/n1867 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1875 ) );
  MUX \Inst_Mem/U1904  ( .A(\Inst_Mem/n1873 ), .B(\Inst_Mem/n1870 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1874 ) );
  MUX \Inst_Mem/U1903  ( .A(\Inst_Mem/n1872 ), .B(\Inst_Mem/n1871 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1873 ) );
  MUX \Inst_Mem/U1902  ( .A(inst_mem_in_wire[1566]), .B(inst_mem_in_wire[1598]), .S(pc_current[2]), .Z(\Inst_Mem/n1872 ) );
  MUX \Inst_Mem/U1901  ( .A(inst_mem_in_wire[1630]), .B(inst_mem_in_wire[1662]), .S(pc_current[2]), .Z(\Inst_Mem/n1871 ) );
  MUX \Inst_Mem/U1900  ( .A(\Inst_Mem/n1869 ), .B(\Inst_Mem/n1868 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1870 ) );
  MUX \Inst_Mem/U1899  ( .A(inst_mem_in_wire[1694]), .B(inst_mem_in_wire[1726]), .S(pc_current[2]), .Z(\Inst_Mem/n1869 ) );
  MUX \Inst_Mem/U1898  ( .A(inst_mem_in_wire[1758]), .B(inst_mem_in_wire[1790]), .S(pc_current[2]), .Z(\Inst_Mem/n1868 ) );
  MUX \Inst_Mem/U1897  ( .A(\Inst_Mem/n1866 ), .B(\Inst_Mem/n1863 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1867 ) );
  MUX \Inst_Mem/U1896  ( .A(\Inst_Mem/n1865 ), .B(\Inst_Mem/n1864 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1866 ) );
  MUX \Inst_Mem/U1895  ( .A(inst_mem_in_wire[1822]), .B(inst_mem_in_wire[1854]), .S(pc_current[2]), .Z(\Inst_Mem/n1865 ) );
  MUX \Inst_Mem/U1894  ( .A(inst_mem_in_wire[1886]), .B(inst_mem_in_wire[1918]), .S(pc_current[2]), .Z(\Inst_Mem/n1864 ) );
  MUX \Inst_Mem/U1893  ( .A(\Inst_Mem/n1862 ), .B(\Inst_Mem/n1861 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1863 ) );
  MUX \Inst_Mem/U1892  ( .A(inst_mem_in_wire[1950]), .B(inst_mem_in_wire[1982]), .S(pc_current[2]), .Z(\Inst_Mem/n1862 ) );
  MUX \Inst_Mem/U1891  ( .A(inst_mem_in_wire[2014]), .B(inst_mem_in_wire[2046]), .S(pc_current[2]), .Z(\Inst_Mem/n1861 ) );
  MUX \Inst_Mem/U1890  ( .A(\Inst_Mem/n1860 ), .B(\Inst_Mem/n1829 ), .S(
        pc_current[7]), .Z(opcode[29]) );
  MUX \Inst_Mem/U1889  ( .A(\Inst_Mem/n1859 ), .B(\Inst_Mem/n1844 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1860 ) );
  MUX \Inst_Mem/U1888  ( .A(\Inst_Mem/n1858 ), .B(\Inst_Mem/n1851 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1859 ) );
  MUX \Inst_Mem/U1887  ( .A(\Inst_Mem/n1857 ), .B(\Inst_Mem/n1854 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1858 ) );
  MUX \Inst_Mem/U1886  ( .A(\Inst_Mem/n1856 ), .B(\Inst_Mem/n1855 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1857 ) );
  MUX \Inst_Mem/U1885  ( .A(inst_mem_in_wire[29]), .B(inst_mem_in_wire[61]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1856 ) );
  MUX \Inst_Mem/U1884  ( .A(inst_mem_in_wire[93]), .B(inst_mem_in_wire[125]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1855 ) );
  MUX \Inst_Mem/U1883  ( .A(\Inst_Mem/n1853 ), .B(\Inst_Mem/n1852 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1854 ) );
  MUX \Inst_Mem/U1882  ( .A(inst_mem_in_wire[157]), .B(inst_mem_in_wire[189]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1853 ) );
  MUX \Inst_Mem/U1881  ( .A(inst_mem_in_wire[221]), .B(inst_mem_in_wire[253]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1852 ) );
  MUX \Inst_Mem/U1880  ( .A(\Inst_Mem/n1850 ), .B(\Inst_Mem/n1847 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1851 ) );
  MUX \Inst_Mem/U1879  ( .A(\Inst_Mem/n1849 ), .B(\Inst_Mem/n1848 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1850 ) );
  MUX \Inst_Mem/U1878  ( .A(inst_mem_in_wire[285]), .B(inst_mem_in_wire[317]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1849 ) );
  MUX \Inst_Mem/U1877  ( .A(inst_mem_in_wire[349]), .B(inst_mem_in_wire[381]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1848 ) );
  MUX \Inst_Mem/U1876  ( .A(\Inst_Mem/n1846 ), .B(\Inst_Mem/n1845 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1847 ) );
  MUX \Inst_Mem/U1875  ( .A(inst_mem_in_wire[413]), .B(inst_mem_in_wire[445]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1846 ) );
  MUX \Inst_Mem/U1874  ( .A(inst_mem_in_wire[477]), .B(inst_mem_in_wire[509]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1845 ) );
  MUX \Inst_Mem/U1873  ( .A(\Inst_Mem/n1843 ), .B(\Inst_Mem/n1836 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1844 ) );
  MUX \Inst_Mem/U1872  ( .A(\Inst_Mem/n1842 ), .B(\Inst_Mem/n1839 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1843 ) );
  MUX \Inst_Mem/U1871  ( .A(\Inst_Mem/n1841 ), .B(\Inst_Mem/n1840 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1842 ) );
  MUX \Inst_Mem/U1870  ( .A(inst_mem_in_wire[541]), .B(inst_mem_in_wire[573]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1841 ) );
  MUX \Inst_Mem/U1869  ( .A(inst_mem_in_wire[605]), .B(inst_mem_in_wire[637]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1840 ) );
  MUX \Inst_Mem/U1868  ( .A(\Inst_Mem/n1838 ), .B(\Inst_Mem/n1837 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1839 ) );
  MUX \Inst_Mem/U1867  ( .A(inst_mem_in_wire[669]), .B(inst_mem_in_wire[701]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1838 ) );
  MUX \Inst_Mem/U1866  ( .A(inst_mem_in_wire[733]), .B(inst_mem_in_wire[765]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1837 ) );
  MUX \Inst_Mem/U1865  ( .A(\Inst_Mem/n1835 ), .B(\Inst_Mem/n1832 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1836 ) );
  MUX \Inst_Mem/U1864  ( .A(\Inst_Mem/n1834 ), .B(\Inst_Mem/n1833 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1835 ) );
  MUX \Inst_Mem/U1863  ( .A(inst_mem_in_wire[797]), .B(inst_mem_in_wire[829]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1834 ) );
  MUX \Inst_Mem/U1862  ( .A(inst_mem_in_wire[861]), .B(inst_mem_in_wire[893]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1833 ) );
  MUX \Inst_Mem/U1861  ( .A(\Inst_Mem/n1831 ), .B(\Inst_Mem/n1830 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1832 ) );
  MUX \Inst_Mem/U1860  ( .A(inst_mem_in_wire[925]), .B(inst_mem_in_wire[957]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1831 ) );
  MUX \Inst_Mem/U1859  ( .A(inst_mem_in_wire[989]), .B(inst_mem_in_wire[1021]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1830 ) );
  MUX \Inst_Mem/U1858  ( .A(\Inst_Mem/n1828 ), .B(\Inst_Mem/n1813 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1829 ) );
  MUX \Inst_Mem/U1857  ( .A(\Inst_Mem/n1827 ), .B(\Inst_Mem/n1820 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1828 ) );
  MUX \Inst_Mem/U1856  ( .A(\Inst_Mem/n1826 ), .B(\Inst_Mem/n1823 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1827 ) );
  MUX \Inst_Mem/U1855  ( .A(\Inst_Mem/n1825 ), .B(\Inst_Mem/n1824 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1826 ) );
  MUX \Inst_Mem/U1854  ( .A(inst_mem_in_wire[1053]), .B(inst_mem_in_wire[1085]), .S(pc_current[2]), .Z(\Inst_Mem/n1825 ) );
  MUX \Inst_Mem/U1853  ( .A(inst_mem_in_wire[1117]), .B(inst_mem_in_wire[1149]), .S(pc_current[2]), .Z(\Inst_Mem/n1824 ) );
  MUX \Inst_Mem/U1852  ( .A(\Inst_Mem/n1822 ), .B(\Inst_Mem/n1821 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1823 ) );
  MUX \Inst_Mem/U1851  ( .A(inst_mem_in_wire[1181]), .B(inst_mem_in_wire[1213]), .S(pc_current[2]), .Z(\Inst_Mem/n1822 ) );
  MUX \Inst_Mem/U1850  ( .A(inst_mem_in_wire[1245]), .B(inst_mem_in_wire[1277]), .S(pc_current[2]), .Z(\Inst_Mem/n1821 ) );
  MUX \Inst_Mem/U1849  ( .A(\Inst_Mem/n1819 ), .B(\Inst_Mem/n1816 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1820 ) );
  MUX \Inst_Mem/U1848  ( .A(\Inst_Mem/n1818 ), .B(\Inst_Mem/n1817 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1819 ) );
  MUX \Inst_Mem/U1847  ( .A(inst_mem_in_wire[1309]), .B(inst_mem_in_wire[1341]), .S(pc_current[2]), .Z(\Inst_Mem/n1818 ) );
  MUX \Inst_Mem/U1846  ( .A(inst_mem_in_wire[1373]), .B(inst_mem_in_wire[1405]), .S(pc_current[2]), .Z(\Inst_Mem/n1817 ) );
  MUX \Inst_Mem/U1845  ( .A(\Inst_Mem/n1815 ), .B(\Inst_Mem/n1814 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1816 ) );
  MUX \Inst_Mem/U1844  ( .A(inst_mem_in_wire[1437]), .B(inst_mem_in_wire[1469]), .S(pc_current[2]), .Z(\Inst_Mem/n1815 ) );
  MUX \Inst_Mem/U1843  ( .A(inst_mem_in_wire[1501]), .B(inst_mem_in_wire[1533]), .S(pc_current[2]), .Z(\Inst_Mem/n1814 ) );
  MUX \Inst_Mem/U1842  ( .A(\Inst_Mem/n1812 ), .B(\Inst_Mem/n1805 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1813 ) );
  MUX \Inst_Mem/U1841  ( .A(\Inst_Mem/n1811 ), .B(\Inst_Mem/n1808 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1812 ) );
  MUX \Inst_Mem/U1840  ( .A(\Inst_Mem/n1810 ), .B(\Inst_Mem/n1809 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1811 ) );
  MUX \Inst_Mem/U1839  ( .A(inst_mem_in_wire[1565]), .B(inst_mem_in_wire[1597]), .S(pc_current[2]), .Z(\Inst_Mem/n1810 ) );
  MUX \Inst_Mem/U1838  ( .A(inst_mem_in_wire[1629]), .B(inst_mem_in_wire[1661]), .S(pc_current[2]), .Z(\Inst_Mem/n1809 ) );
  MUX \Inst_Mem/U1837  ( .A(\Inst_Mem/n1807 ), .B(\Inst_Mem/n1806 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1808 ) );
  MUX \Inst_Mem/U1836  ( .A(inst_mem_in_wire[1693]), .B(inst_mem_in_wire[1725]), .S(pc_current[2]), .Z(\Inst_Mem/n1807 ) );
  MUX \Inst_Mem/U1835  ( .A(inst_mem_in_wire[1757]), .B(inst_mem_in_wire[1789]), .S(pc_current[2]), .Z(\Inst_Mem/n1806 ) );
  MUX \Inst_Mem/U1834  ( .A(\Inst_Mem/n1804 ), .B(\Inst_Mem/n1801 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1805 ) );
  MUX \Inst_Mem/U1833  ( .A(\Inst_Mem/n1803 ), .B(\Inst_Mem/n1802 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1804 ) );
  MUX \Inst_Mem/U1832  ( .A(inst_mem_in_wire[1821]), .B(inst_mem_in_wire[1853]), .S(pc_current[2]), .Z(\Inst_Mem/n1803 ) );
  MUX \Inst_Mem/U1831  ( .A(inst_mem_in_wire[1885]), .B(inst_mem_in_wire[1917]), .S(pc_current[2]), .Z(\Inst_Mem/n1802 ) );
  MUX \Inst_Mem/U1830  ( .A(\Inst_Mem/n1800 ), .B(\Inst_Mem/n1799 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1801 ) );
  MUX \Inst_Mem/U1829  ( .A(inst_mem_in_wire[1949]), .B(inst_mem_in_wire[1981]), .S(pc_current[2]), .Z(\Inst_Mem/n1800 ) );
  MUX \Inst_Mem/U1828  ( .A(inst_mem_in_wire[2013]), .B(inst_mem_in_wire[2045]), .S(pc_current[2]), .Z(\Inst_Mem/n1799 ) );
  MUX \Inst_Mem/U1827  ( .A(\Inst_Mem/n1798 ), .B(\Inst_Mem/n1767 ), .S(
        pc_current[7]), .Z(opcode[28]) );
  MUX \Inst_Mem/U1826  ( .A(\Inst_Mem/n1797 ), .B(\Inst_Mem/n1782 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1798 ) );
  MUX \Inst_Mem/U1825  ( .A(\Inst_Mem/n1796 ), .B(\Inst_Mem/n1789 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1797 ) );
  MUX \Inst_Mem/U1824  ( .A(\Inst_Mem/n1795 ), .B(\Inst_Mem/n1792 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1796 ) );
  MUX \Inst_Mem/U1823  ( .A(\Inst_Mem/n1794 ), .B(\Inst_Mem/n1793 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1795 ) );
  MUX \Inst_Mem/U1822  ( .A(inst_mem_in_wire[28]), .B(inst_mem_in_wire[60]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1794 ) );
  MUX \Inst_Mem/U1821  ( .A(inst_mem_in_wire[92]), .B(inst_mem_in_wire[124]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1793 ) );
  MUX \Inst_Mem/U1820  ( .A(\Inst_Mem/n1791 ), .B(\Inst_Mem/n1790 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1792 ) );
  MUX \Inst_Mem/U1819  ( .A(inst_mem_in_wire[156]), .B(inst_mem_in_wire[188]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1791 ) );
  MUX \Inst_Mem/U1818  ( .A(inst_mem_in_wire[220]), .B(inst_mem_in_wire[252]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1790 ) );
  MUX \Inst_Mem/U1817  ( .A(\Inst_Mem/n1788 ), .B(\Inst_Mem/n1785 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1789 ) );
  MUX \Inst_Mem/U1816  ( .A(\Inst_Mem/n1787 ), .B(\Inst_Mem/n1786 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1788 ) );
  MUX \Inst_Mem/U1815  ( .A(inst_mem_in_wire[284]), .B(inst_mem_in_wire[316]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1787 ) );
  MUX \Inst_Mem/U1814  ( .A(inst_mem_in_wire[348]), .B(inst_mem_in_wire[380]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1786 ) );
  MUX \Inst_Mem/U1813  ( .A(\Inst_Mem/n1784 ), .B(\Inst_Mem/n1783 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1785 ) );
  MUX \Inst_Mem/U1812  ( .A(inst_mem_in_wire[412]), .B(inst_mem_in_wire[444]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1784 ) );
  MUX \Inst_Mem/U1811  ( .A(inst_mem_in_wire[476]), .B(inst_mem_in_wire[508]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1783 ) );
  MUX \Inst_Mem/U1810  ( .A(\Inst_Mem/n1781 ), .B(\Inst_Mem/n1774 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1782 ) );
  MUX \Inst_Mem/U1809  ( .A(\Inst_Mem/n1780 ), .B(\Inst_Mem/n1777 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1781 ) );
  MUX \Inst_Mem/U1808  ( .A(\Inst_Mem/n1779 ), .B(\Inst_Mem/n1778 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1780 ) );
  MUX \Inst_Mem/U1807  ( .A(inst_mem_in_wire[540]), .B(inst_mem_in_wire[572]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1779 ) );
  MUX \Inst_Mem/U1806  ( .A(inst_mem_in_wire[604]), .B(inst_mem_in_wire[636]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1778 ) );
  MUX \Inst_Mem/U1805  ( .A(\Inst_Mem/n1776 ), .B(\Inst_Mem/n1775 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1777 ) );
  MUX \Inst_Mem/U1804  ( .A(inst_mem_in_wire[668]), .B(inst_mem_in_wire[700]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1776 ) );
  MUX \Inst_Mem/U1803  ( .A(inst_mem_in_wire[732]), .B(inst_mem_in_wire[764]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1775 ) );
  MUX \Inst_Mem/U1802  ( .A(\Inst_Mem/n1773 ), .B(\Inst_Mem/n1770 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1774 ) );
  MUX \Inst_Mem/U1801  ( .A(\Inst_Mem/n1772 ), .B(\Inst_Mem/n1771 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1773 ) );
  MUX \Inst_Mem/U1800  ( .A(inst_mem_in_wire[796]), .B(inst_mem_in_wire[828]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1772 ) );
  MUX \Inst_Mem/U1799  ( .A(inst_mem_in_wire[860]), .B(inst_mem_in_wire[892]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1771 ) );
  MUX \Inst_Mem/U1798  ( .A(\Inst_Mem/n1769 ), .B(\Inst_Mem/n1768 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1770 ) );
  MUX \Inst_Mem/U1797  ( .A(inst_mem_in_wire[924]), .B(inst_mem_in_wire[956]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1769 ) );
  MUX \Inst_Mem/U1796  ( .A(inst_mem_in_wire[988]), .B(inst_mem_in_wire[1020]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1768 ) );
  MUX \Inst_Mem/U1795  ( .A(\Inst_Mem/n1766 ), .B(\Inst_Mem/n1751 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1767 ) );
  MUX \Inst_Mem/U1794  ( .A(\Inst_Mem/n1765 ), .B(\Inst_Mem/n1758 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1766 ) );
  MUX \Inst_Mem/U1793  ( .A(\Inst_Mem/n1764 ), .B(\Inst_Mem/n1761 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1765 ) );
  MUX \Inst_Mem/U1792  ( .A(\Inst_Mem/n1763 ), .B(\Inst_Mem/n1762 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1764 ) );
  MUX \Inst_Mem/U1791  ( .A(inst_mem_in_wire[1052]), .B(inst_mem_in_wire[1084]), .S(pc_current[2]), .Z(\Inst_Mem/n1763 ) );
  MUX \Inst_Mem/U1790  ( .A(inst_mem_in_wire[1116]), .B(inst_mem_in_wire[1148]), .S(pc_current[2]), .Z(\Inst_Mem/n1762 ) );
  MUX \Inst_Mem/U1789  ( .A(\Inst_Mem/n1760 ), .B(\Inst_Mem/n1759 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1761 ) );
  MUX \Inst_Mem/U1788  ( .A(inst_mem_in_wire[1180]), .B(inst_mem_in_wire[1212]), .S(pc_current[2]), .Z(\Inst_Mem/n1760 ) );
  MUX \Inst_Mem/U1787  ( .A(inst_mem_in_wire[1244]), .B(inst_mem_in_wire[1276]), .S(pc_current[2]), .Z(\Inst_Mem/n1759 ) );
  MUX \Inst_Mem/U1786  ( .A(\Inst_Mem/n1757 ), .B(\Inst_Mem/n1754 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1758 ) );
  MUX \Inst_Mem/U1785  ( .A(\Inst_Mem/n1756 ), .B(\Inst_Mem/n1755 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1757 ) );
  MUX \Inst_Mem/U1784  ( .A(inst_mem_in_wire[1308]), .B(inst_mem_in_wire[1340]), .S(pc_current[2]), .Z(\Inst_Mem/n1756 ) );
  MUX \Inst_Mem/U1783  ( .A(inst_mem_in_wire[1372]), .B(inst_mem_in_wire[1404]), .S(pc_current[2]), .Z(\Inst_Mem/n1755 ) );
  MUX \Inst_Mem/U1782  ( .A(\Inst_Mem/n1753 ), .B(\Inst_Mem/n1752 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1754 ) );
  MUX \Inst_Mem/U1781  ( .A(inst_mem_in_wire[1436]), .B(inst_mem_in_wire[1468]), .S(pc_current[2]), .Z(\Inst_Mem/n1753 ) );
  MUX \Inst_Mem/U1780  ( .A(inst_mem_in_wire[1500]), .B(inst_mem_in_wire[1532]), .S(pc_current[2]), .Z(\Inst_Mem/n1752 ) );
  MUX \Inst_Mem/U1779  ( .A(\Inst_Mem/n1750 ), .B(\Inst_Mem/n1743 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1751 ) );
  MUX \Inst_Mem/U1778  ( .A(\Inst_Mem/n1749 ), .B(\Inst_Mem/n1746 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1750 ) );
  MUX \Inst_Mem/U1777  ( .A(\Inst_Mem/n1748 ), .B(\Inst_Mem/n1747 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1749 ) );
  MUX \Inst_Mem/U1776  ( .A(inst_mem_in_wire[1564]), .B(inst_mem_in_wire[1596]), .S(pc_current[2]), .Z(\Inst_Mem/n1748 ) );
  MUX \Inst_Mem/U1775  ( .A(inst_mem_in_wire[1628]), .B(inst_mem_in_wire[1660]), .S(pc_current[2]), .Z(\Inst_Mem/n1747 ) );
  MUX \Inst_Mem/U1774  ( .A(\Inst_Mem/n1745 ), .B(\Inst_Mem/n1744 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1746 ) );
  MUX \Inst_Mem/U1773  ( .A(inst_mem_in_wire[1692]), .B(inst_mem_in_wire[1724]), .S(pc_current[2]), .Z(\Inst_Mem/n1745 ) );
  MUX \Inst_Mem/U1772  ( .A(inst_mem_in_wire[1756]), .B(inst_mem_in_wire[1788]), .S(pc_current[2]), .Z(\Inst_Mem/n1744 ) );
  MUX \Inst_Mem/U1771  ( .A(\Inst_Mem/n1742 ), .B(\Inst_Mem/n1739 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1743 ) );
  MUX \Inst_Mem/U1770  ( .A(\Inst_Mem/n1741 ), .B(\Inst_Mem/n1740 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1742 ) );
  MUX \Inst_Mem/U1769  ( .A(inst_mem_in_wire[1820]), .B(inst_mem_in_wire[1852]), .S(pc_current[2]), .Z(\Inst_Mem/n1741 ) );
  MUX \Inst_Mem/U1768  ( .A(inst_mem_in_wire[1884]), .B(inst_mem_in_wire[1916]), .S(pc_current[2]), .Z(\Inst_Mem/n1740 ) );
  MUX \Inst_Mem/U1767  ( .A(\Inst_Mem/n1738 ), .B(\Inst_Mem/n1737 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1739 ) );
  MUX \Inst_Mem/U1766  ( .A(inst_mem_in_wire[1948]), .B(inst_mem_in_wire[1980]), .S(pc_current[2]), .Z(\Inst_Mem/n1738 ) );
  MUX \Inst_Mem/U1765  ( .A(inst_mem_in_wire[2012]), .B(inst_mem_in_wire[2044]), .S(pc_current[2]), .Z(\Inst_Mem/n1737 ) );
  MUX \Inst_Mem/U1764  ( .A(\Inst_Mem/n1736 ), .B(\Inst_Mem/n1705 ), .S(
        pc_current[7]), .Z(opcode[27]) );
  MUX \Inst_Mem/U1763  ( .A(\Inst_Mem/n1735 ), .B(\Inst_Mem/n1720 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1736 ) );
  MUX \Inst_Mem/U1762  ( .A(\Inst_Mem/n1734 ), .B(\Inst_Mem/n1727 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1735 ) );
  MUX \Inst_Mem/U1761  ( .A(\Inst_Mem/n1733 ), .B(\Inst_Mem/n1730 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1734 ) );
  MUX \Inst_Mem/U1760  ( .A(\Inst_Mem/n1732 ), .B(\Inst_Mem/n1731 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1733 ) );
  MUX \Inst_Mem/U1759  ( .A(inst_mem_in_wire[27]), .B(inst_mem_in_wire[59]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1732 ) );
  MUX \Inst_Mem/U1758  ( .A(inst_mem_in_wire[91]), .B(inst_mem_in_wire[123]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1731 ) );
  MUX \Inst_Mem/U1757  ( .A(\Inst_Mem/n1729 ), .B(\Inst_Mem/n1728 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1730 ) );
  MUX \Inst_Mem/U1756  ( .A(inst_mem_in_wire[155]), .B(inst_mem_in_wire[187]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1729 ) );
  MUX \Inst_Mem/U1755  ( .A(inst_mem_in_wire[219]), .B(inst_mem_in_wire[251]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1728 ) );
  MUX \Inst_Mem/U1754  ( .A(\Inst_Mem/n1726 ), .B(\Inst_Mem/n1723 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1727 ) );
  MUX \Inst_Mem/U1753  ( .A(\Inst_Mem/n1725 ), .B(\Inst_Mem/n1724 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1726 ) );
  MUX \Inst_Mem/U1752  ( .A(inst_mem_in_wire[283]), .B(inst_mem_in_wire[315]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1725 ) );
  MUX \Inst_Mem/U1751  ( .A(inst_mem_in_wire[347]), .B(inst_mem_in_wire[379]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1724 ) );
  MUX \Inst_Mem/U1750  ( .A(\Inst_Mem/n1722 ), .B(\Inst_Mem/n1721 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1723 ) );
  MUX \Inst_Mem/U1749  ( .A(inst_mem_in_wire[411]), .B(inst_mem_in_wire[443]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1722 ) );
  MUX \Inst_Mem/U1748  ( .A(inst_mem_in_wire[475]), .B(inst_mem_in_wire[507]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1721 ) );
  MUX \Inst_Mem/U1747  ( .A(\Inst_Mem/n1719 ), .B(\Inst_Mem/n1712 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1720 ) );
  MUX \Inst_Mem/U1746  ( .A(\Inst_Mem/n1718 ), .B(\Inst_Mem/n1715 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1719 ) );
  MUX \Inst_Mem/U1745  ( .A(\Inst_Mem/n1717 ), .B(\Inst_Mem/n1716 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1718 ) );
  MUX \Inst_Mem/U1744  ( .A(inst_mem_in_wire[539]), .B(inst_mem_in_wire[571]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1717 ) );
  MUX \Inst_Mem/U1743  ( .A(inst_mem_in_wire[603]), .B(inst_mem_in_wire[635]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1716 ) );
  MUX \Inst_Mem/U1742  ( .A(\Inst_Mem/n1714 ), .B(\Inst_Mem/n1713 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1715 ) );
  MUX \Inst_Mem/U1741  ( .A(inst_mem_in_wire[667]), .B(inst_mem_in_wire[699]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1714 ) );
  MUX \Inst_Mem/U1740  ( .A(inst_mem_in_wire[731]), .B(inst_mem_in_wire[763]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1713 ) );
  MUX \Inst_Mem/U1739  ( .A(\Inst_Mem/n1711 ), .B(\Inst_Mem/n1708 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1712 ) );
  MUX \Inst_Mem/U1738  ( .A(\Inst_Mem/n1710 ), .B(\Inst_Mem/n1709 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1711 ) );
  MUX \Inst_Mem/U1737  ( .A(inst_mem_in_wire[795]), .B(inst_mem_in_wire[827]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1710 ) );
  MUX \Inst_Mem/U1736  ( .A(inst_mem_in_wire[859]), .B(inst_mem_in_wire[891]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1709 ) );
  MUX \Inst_Mem/U1735  ( .A(\Inst_Mem/n1707 ), .B(\Inst_Mem/n1706 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1708 ) );
  MUX \Inst_Mem/U1734  ( .A(inst_mem_in_wire[923]), .B(inst_mem_in_wire[955]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1707 ) );
  MUX \Inst_Mem/U1733  ( .A(inst_mem_in_wire[987]), .B(inst_mem_in_wire[1019]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1706 ) );
  MUX \Inst_Mem/U1732  ( .A(\Inst_Mem/n1704 ), .B(\Inst_Mem/n1689 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1705 ) );
  MUX \Inst_Mem/U1731  ( .A(\Inst_Mem/n1703 ), .B(\Inst_Mem/n1696 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1704 ) );
  MUX \Inst_Mem/U1730  ( .A(\Inst_Mem/n1702 ), .B(\Inst_Mem/n1699 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1703 ) );
  MUX \Inst_Mem/U1729  ( .A(\Inst_Mem/n1701 ), .B(\Inst_Mem/n1700 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1702 ) );
  MUX \Inst_Mem/U1728  ( .A(inst_mem_in_wire[1051]), .B(inst_mem_in_wire[1083]), .S(pc_current[2]), .Z(\Inst_Mem/n1701 ) );
  MUX \Inst_Mem/U1727  ( .A(inst_mem_in_wire[1115]), .B(inst_mem_in_wire[1147]), .S(pc_current[2]), .Z(\Inst_Mem/n1700 ) );
  MUX \Inst_Mem/U1726  ( .A(\Inst_Mem/n1698 ), .B(\Inst_Mem/n1697 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1699 ) );
  MUX \Inst_Mem/U1725  ( .A(inst_mem_in_wire[1179]), .B(inst_mem_in_wire[1211]), .S(pc_current[2]), .Z(\Inst_Mem/n1698 ) );
  MUX \Inst_Mem/U1724  ( .A(inst_mem_in_wire[1243]), .B(inst_mem_in_wire[1275]), .S(pc_current[2]), .Z(\Inst_Mem/n1697 ) );
  MUX \Inst_Mem/U1723  ( .A(\Inst_Mem/n1695 ), .B(\Inst_Mem/n1692 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1696 ) );
  MUX \Inst_Mem/U1722  ( .A(\Inst_Mem/n1694 ), .B(\Inst_Mem/n1693 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1695 ) );
  MUX \Inst_Mem/U1721  ( .A(inst_mem_in_wire[1307]), .B(inst_mem_in_wire[1339]), .S(pc_current[2]), .Z(\Inst_Mem/n1694 ) );
  MUX \Inst_Mem/U1720  ( .A(inst_mem_in_wire[1371]), .B(inst_mem_in_wire[1403]), .S(pc_current[2]), .Z(\Inst_Mem/n1693 ) );
  MUX \Inst_Mem/U1719  ( .A(\Inst_Mem/n1691 ), .B(\Inst_Mem/n1690 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1692 ) );
  MUX \Inst_Mem/U1718  ( .A(inst_mem_in_wire[1435]), .B(inst_mem_in_wire[1467]), .S(pc_current[2]), .Z(\Inst_Mem/n1691 ) );
  MUX \Inst_Mem/U1717  ( .A(inst_mem_in_wire[1499]), .B(inst_mem_in_wire[1531]), .S(pc_current[2]), .Z(\Inst_Mem/n1690 ) );
  MUX \Inst_Mem/U1716  ( .A(\Inst_Mem/n1688 ), .B(\Inst_Mem/n1681 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1689 ) );
  MUX \Inst_Mem/U1715  ( .A(\Inst_Mem/n1687 ), .B(\Inst_Mem/n1684 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1688 ) );
  MUX \Inst_Mem/U1714  ( .A(\Inst_Mem/n1686 ), .B(\Inst_Mem/n1685 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1687 ) );
  MUX \Inst_Mem/U1713  ( .A(inst_mem_in_wire[1563]), .B(inst_mem_in_wire[1595]), .S(pc_current[2]), .Z(\Inst_Mem/n1686 ) );
  MUX \Inst_Mem/U1712  ( .A(inst_mem_in_wire[1627]), .B(inst_mem_in_wire[1659]), .S(pc_current[2]), .Z(\Inst_Mem/n1685 ) );
  MUX \Inst_Mem/U1711  ( .A(\Inst_Mem/n1683 ), .B(\Inst_Mem/n1682 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1684 ) );
  MUX \Inst_Mem/U1710  ( .A(inst_mem_in_wire[1691]), .B(inst_mem_in_wire[1723]), .S(pc_current[2]), .Z(\Inst_Mem/n1683 ) );
  MUX \Inst_Mem/U1709  ( .A(inst_mem_in_wire[1755]), .B(inst_mem_in_wire[1787]), .S(pc_current[2]), .Z(\Inst_Mem/n1682 ) );
  MUX \Inst_Mem/U1708  ( .A(\Inst_Mem/n1680 ), .B(\Inst_Mem/n1677 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1681 ) );
  MUX \Inst_Mem/U1707  ( .A(\Inst_Mem/n1679 ), .B(\Inst_Mem/n1678 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1680 ) );
  MUX \Inst_Mem/U1706  ( .A(inst_mem_in_wire[1819]), .B(inst_mem_in_wire[1851]), .S(pc_current[2]), .Z(\Inst_Mem/n1679 ) );
  MUX \Inst_Mem/U1705  ( .A(inst_mem_in_wire[1883]), .B(inst_mem_in_wire[1915]), .S(pc_current[2]), .Z(\Inst_Mem/n1678 ) );
  MUX \Inst_Mem/U1704  ( .A(\Inst_Mem/n1676 ), .B(\Inst_Mem/n1675 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1677 ) );
  MUX \Inst_Mem/U1703  ( .A(inst_mem_in_wire[1947]), .B(inst_mem_in_wire[1979]), .S(pc_current[2]), .Z(\Inst_Mem/n1676 ) );
  MUX \Inst_Mem/U1702  ( .A(inst_mem_in_wire[2011]), .B(inst_mem_in_wire[2043]), .S(pc_current[2]), .Z(\Inst_Mem/n1675 ) );
  MUX \Inst_Mem/U1701  ( .A(\Inst_Mem/n1674 ), .B(\Inst_Mem/n1643 ), .S(
        pc_current[7]), .Z(opcode[26]) );
  MUX \Inst_Mem/U1700  ( .A(\Inst_Mem/n1673 ), .B(\Inst_Mem/n1658 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1674 ) );
  MUX \Inst_Mem/U1699  ( .A(\Inst_Mem/n1672 ), .B(\Inst_Mem/n1665 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1673 ) );
  MUX \Inst_Mem/U1698  ( .A(\Inst_Mem/n1671 ), .B(\Inst_Mem/n1668 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1672 ) );
  MUX \Inst_Mem/U1697  ( .A(\Inst_Mem/n1670 ), .B(\Inst_Mem/n1669 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1671 ) );
  MUX \Inst_Mem/U1696  ( .A(inst_mem_in_wire[26]), .B(inst_mem_in_wire[58]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1670 ) );
  MUX \Inst_Mem/U1695  ( .A(inst_mem_in_wire[90]), .B(inst_mem_in_wire[122]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1669 ) );
  MUX \Inst_Mem/U1694  ( .A(\Inst_Mem/n1667 ), .B(\Inst_Mem/n1666 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1668 ) );
  MUX \Inst_Mem/U1693  ( .A(inst_mem_in_wire[154]), .B(inst_mem_in_wire[186]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1667 ) );
  MUX \Inst_Mem/U1692  ( .A(inst_mem_in_wire[218]), .B(inst_mem_in_wire[250]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1666 ) );
  MUX \Inst_Mem/U1691  ( .A(\Inst_Mem/n1664 ), .B(\Inst_Mem/n1661 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1665 ) );
  MUX \Inst_Mem/U1690  ( .A(\Inst_Mem/n1663 ), .B(\Inst_Mem/n1662 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1664 ) );
  MUX \Inst_Mem/U1689  ( .A(inst_mem_in_wire[282]), .B(inst_mem_in_wire[314]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1663 ) );
  MUX \Inst_Mem/U1688  ( .A(inst_mem_in_wire[346]), .B(inst_mem_in_wire[378]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1662 ) );
  MUX \Inst_Mem/U1687  ( .A(\Inst_Mem/n1660 ), .B(\Inst_Mem/n1659 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1661 ) );
  MUX \Inst_Mem/U1686  ( .A(inst_mem_in_wire[410]), .B(inst_mem_in_wire[442]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1660 ) );
  MUX \Inst_Mem/U1685  ( .A(inst_mem_in_wire[474]), .B(inst_mem_in_wire[506]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1659 ) );
  MUX \Inst_Mem/U1684  ( .A(\Inst_Mem/n1657 ), .B(\Inst_Mem/n1650 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1658 ) );
  MUX \Inst_Mem/U1683  ( .A(\Inst_Mem/n1656 ), .B(\Inst_Mem/n1653 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1657 ) );
  MUX \Inst_Mem/U1682  ( .A(\Inst_Mem/n1655 ), .B(\Inst_Mem/n1654 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1656 ) );
  MUX \Inst_Mem/U1681  ( .A(inst_mem_in_wire[538]), .B(inst_mem_in_wire[570]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1655 ) );
  MUX \Inst_Mem/U1680  ( .A(inst_mem_in_wire[602]), .B(inst_mem_in_wire[634]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1654 ) );
  MUX \Inst_Mem/U1679  ( .A(\Inst_Mem/n1652 ), .B(\Inst_Mem/n1651 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1653 ) );
  MUX \Inst_Mem/U1678  ( .A(inst_mem_in_wire[666]), .B(inst_mem_in_wire[698]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1652 ) );
  MUX \Inst_Mem/U1677  ( .A(inst_mem_in_wire[730]), .B(inst_mem_in_wire[762]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1651 ) );
  MUX \Inst_Mem/U1676  ( .A(\Inst_Mem/n1649 ), .B(\Inst_Mem/n1646 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1650 ) );
  MUX \Inst_Mem/U1675  ( .A(\Inst_Mem/n1648 ), .B(\Inst_Mem/n1647 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1649 ) );
  MUX \Inst_Mem/U1674  ( .A(inst_mem_in_wire[794]), .B(inst_mem_in_wire[826]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1648 ) );
  MUX \Inst_Mem/U1673  ( .A(inst_mem_in_wire[858]), .B(inst_mem_in_wire[890]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1647 ) );
  MUX \Inst_Mem/U1672  ( .A(\Inst_Mem/n1645 ), .B(\Inst_Mem/n1644 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1646 ) );
  MUX \Inst_Mem/U1671  ( .A(inst_mem_in_wire[922]), .B(inst_mem_in_wire[954]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1645 ) );
  MUX \Inst_Mem/U1670  ( .A(inst_mem_in_wire[986]), .B(inst_mem_in_wire[1018]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1644 ) );
  MUX \Inst_Mem/U1669  ( .A(\Inst_Mem/n1642 ), .B(\Inst_Mem/n1627 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1643 ) );
  MUX \Inst_Mem/U1668  ( .A(\Inst_Mem/n1641 ), .B(\Inst_Mem/n1634 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1642 ) );
  MUX \Inst_Mem/U1667  ( .A(\Inst_Mem/n1640 ), .B(\Inst_Mem/n1637 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1641 ) );
  MUX \Inst_Mem/U1666  ( .A(\Inst_Mem/n1639 ), .B(\Inst_Mem/n1638 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1640 ) );
  MUX \Inst_Mem/U1665  ( .A(inst_mem_in_wire[1050]), .B(inst_mem_in_wire[1082]), .S(pc_current[2]), .Z(\Inst_Mem/n1639 ) );
  MUX \Inst_Mem/U1664  ( .A(inst_mem_in_wire[1114]), .B(inst_mem_in_wire[1146]), .S(pc_current[2]), .Z(\Inst_Mem/n1638 ) );
  MUX \Inst_Mem/U1663  ( .A(\Inst_Mem/n1636 ), .B(\Inst_Mem/n1635 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1637 ) );
  MUX \Inst_Mem/U1662  ( .A(inst_mem_in_wire[1178]), .B(inst_mem_in_wire[1210]), .S(pc_current[2]), .Z(\Inst_Mem/n1636 ) );
  MUX \Inst_Mem/U1661  ( .A(inst_mem_in_wire[1242]), .B(inst_mem_in_wire[1274]), .S(pc_current[2]), .Z(\Inst_Mem/n1635 ) );
  MUX \Inst_Mem/U1660  ( .A(\Inst_Mem/n1633 ), .B(\Inst_Mem/n1630 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1634 ) );
  MUX \Inst_Mem/U1659  ( .A(\Inst_Mem/n1632 ), .B(\Inst_Mem/n1631 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1633 ) );
  MUX \Inst_Mem/U1658  ( .A(inst_mem_in_wire[1306]), .B(inst_mem_in_wire[1338]), .S(pc_current[2]), .Z(\Inst_Mem/n1632 ) );
  MUX \Inst_Mem/U1657  ( .A(inst_mem_in_wire[1370]), .B(inst_mem_in_wire[1402]), .S(pc_current[2]), .Z(\Inst_Mem/n1631 ) );
  MUX \Inst_Mem/U1656  ( .A(\Inst_Mem/n1629 ), .B(\Inst_Mem/n1628 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1630 ) );
  MUX \Inst_Mem/U1655  ( .A(inst_mem_in_wire[1434]), .B(inst_mem_in_wire[1466]), .S(pc_current[2]), .Z(\Inst_Mem/n1629 ) );
  MUX \Inst_Mem/U1654  ( .A(inst_mem_in_wire[1498]), .B(inst_mem_in_wire[1530]), .S(pc_current[2]), .Z(\Inst_Mem/n1628 ) );
  MUX \Inst_Mem/U1653  ( .A(\Inst_Mem/n1626 ), .B(\Inst_Mem/n1619 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1627 ) );
  MUX \Inst_Mem/U1652  ( .A(\Inst_Mem/n1625 ), .B(\Inst_Mem/n1622 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1626 ) );
  MUX \Inst_Mem/U1651  ( .A(\Inst_Mem/n1624 ), .B(\Inst_Mem/n1623 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1625 ) );
  MUX \Inst_Mem/U1650  ( .A(inst_mem_in_wire[1562]), .B(inst_mem_in_wire[1594]), .S(pc_current[2]), .Z(\Inst_Mem/n1624 ) );
  MUX \Inst_Mem/U1649  ( .A(inst_mem_in_wire[1626]), .B(inst_mem_in_wire[1658]), .S(pc_current[2]), .Z(\Inst_Mem/n1623 ) );
  MUX \Inst_Mem/U1648  ( .A(\Inst_Mem/n1621 ), .B(\Inst_Mem/n1620 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1622 ) );
  MUX \Inst_Mem/U1647  ( .A(inst_mem_in_wire[1690]), .B(inst_mem_in_wire[1722]), .S(pc_current[2]), .Z(\Inst_Mem/n1621 ) );
  MUX \Inst_Mem/U1646  ( .A(inst_mem_in_wire[1754]), .B(inst_mem_in_wire[1786]), .S(pc_current[2]), .Z(\Inst_Mem/n1620 ) );
  MUX \Inst_Mem/U1645  ( .A(\Inst_Mem/n1618 ), .B(\Inst_Mem/n1615 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1619 ) );
  MUX \Inst_Mem/U1644  ( .A(\Inst_Mem/n1617 ), .B(\Inst_Mem/n1616 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1618 ) );
  MUX \Inst_Mem/U1643  ( .A(inst_mem_in_wire[1818]), .B(inst_mem_in_wire[1850]), .S(pc_current[2]), .Z(\Inst_Mem/n1617 ) );
  MUX \Inst_Mem/U1642  ( .A(inst_mem_in_wire[1882]), .B(inst_mem_in_wire[1914]), .S(pc_current[2]), .Z(\Inst_Mem/n1616 ) );
  MUX \Inst_Mem/U1641  ( .A(\Inst_Mem/n1614 ), .B(\Inst_Mem/n1613 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1615 ) );
  MUX \Inst_Mem/U1640  ( .A(inst_mem_in_wire[1946]), .B(inst_mem_in_wire[1978]), .S(pc_current[2]), .Z(\Inst_Mem/n1614 ) );
  MUX \Inst_Mem/U1639  ( .A(inst_mem_in_wire[2010]), .B(inst_mem_in_wire[2042]), .S(pc_current[2]), .Z(\Inst_Mem/n1613 ) );
  MUX \Inst_Mem/U1638  ( .A(\Inst_Mem/n1612 ), .B(\Inst_Mem/n1581 ), .S(
        pc_current[7]), .Z(opcode[25]) );
  MUX \Inst_Mem/U1637  ( .A(\Inst_Mem/n1611 ), .B(\Inst_Mem/n1596 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1612 ) );
  MUX \Inst_Mem/U1636  ( .A(\Inst_Mem/n1610 ), .B(\Inst_Mem/n1603 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1611 ) );
  MUX \Inst_Mem/U1635  ( .A(\Inst_Mem/n1609 ), .B(\Inst_Mem/n1606 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1610 ) );
  MUX \Inst_Mem/U1634  ( .A(\Inst_Mem/n1608 ), .B(\Inst_Mem/n1607 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1609 ) );
  MUX \Inst_Mem/U1633  ( .A(inst_mem_in_wire[25]), .B(inst_mem_in_wire[57]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1608 ) );
  MUX \Inst_Mem/U1632  ( .A(inst_mem_in_wire[89]), .B(inst_mem_in_wire[121]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1607 ) );
  MUX \Inst_Mem/U1631  ( .A(\Inst_Mem/n1605 ), .B(\Inst_Mem/n1604 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1606 ) );
  MUX \Inst_Mem/U1630  ( .A(inst_mem_in_wire[153]), .B(inst_mem_in_wire[185]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1605 ) );
  MUX \Inst_Mem/U1629  ( .A(inst_mem_in_wire[217]), .B(inst_mem_in_wire[249]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1604 ) );
  MUX \Inst_Mem/U1628  ( .A(\Inst_Mem/n1602 ), .B(\Inst_Mem/n1599 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1603 ) );
  MUX \Inst_Mem/U1627  ( .A(\Inst_Mem/n1601 ), .B(\Inst_Mem/n1600 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1602 ) );
  MUX \Inst_Mem/U1626  ( .A(inst_mem_in_wire[281]), .B(inst_mem_in_wire[313]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1601 ) );
  MUX \Inst_Mem/U1625  ( .A(inst_mem_in_wire[345]), .B(inst_mem_in_wire[377]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1600 ) );
  MUX \Inst_Mem/U1624  ( .A(\Inst_Mem/n1598 ), .B(\Inst_Mem/n1597 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1599 ) );
  MUX \Inst_Mem/U1623  ( .A(inst_mem_in_wire[409]), .B(inst_mem_in_wire[441]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1598 ) );
  MUX \Inst_Mem/U1622  ( .A(inst_mem_in_wire[473]), .B(inst_mem_in_wire[505]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1597 ) );
  MUX \Inst_Mem/U1621  ( .A(\Inst_Mem/n1595 ), .B(\Inst_Mem/n1588 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1596 ) );
  MUX \Inst_Mem/U1620  ( .A(\Inst_Mem/n1594 ), .B(\Inst_Mem/n1591 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1595 ) );
  MUX \Inst_Mem/U1619  ( .A(\Inst_Mem/n1593 ), .B(\Inst_Mem/n1592 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1594 ) );
  MUX \Inst_Mem/U1618  ( .A(inst_mem_in_wire[537]), .B(inst_mem_in_wire[569]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1593 ) );
  MUX \Inst_Mem/U1617  ( .A(inst_mem_in_wire[601]), .B(inst_mem_in_wire[633]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1592 ) );
  MUX \Inst_Mem/U1616  ( .A(\Inst_Mem/n1590 ), .B(\Inst_Mem/n1589 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1591 ) );
  MUX \Inst_Mem/U1615  ( .A(inst_mem_in_wire[665]), .B(inst_mem_in_wire[697]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1590 ) );
  MUX \Inst_Mem/U1614  ( .A(inst_mem_in_wire[729]), .B(inst_mem_in_wire[761]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1589 ) );
  MUX \Inst_Mem/U1613  ( .A(\Inst_Mem/n1587 ), .B(\Inst_Mem/n1584 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1588 ) );
  MUX \Inst_Mem/U1612  ( .A(\Inst_Mem/n1586 ), .B(\Inst_Mem/n1585 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1587 ) );
  MUX \Inst_Mem/U1611  ( .A(inst_mem_in_wire[793]), .B(inst_mem_in_wire[825]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1586 ) );
  MUX \Inst_Mem/U1610  ( .A(inst_mem_in_wire[857]), .B(inst_mem_in_wire[889]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1585 ) );
  MUX \Inst_Mem/U1609  ( .A(\Inst_Mem/n1583 ), .B(\Inst_Mem/n1582 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1584 ) );
  MUX \Inst_Mem/U1608  ( .A(inst_mem_in_wire[921]), .B(inst_mem_in_wire[953]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1583 ) );
  MUX \Inst_Mem/U1607  ( .A(inst_mem_in_wire[985]), .B(inst_mem_in_wire[1017]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1582 ) );
  MUX \Inst_Mem/U1606  ( .A(\Inst_Mem/n1580 ), .B(\Inst_Mem/n1565 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1581 ) );
  MUX \Inst_Mem/U1605  ( .A(\Inst_Mem/n1579 ), .B(\Inst_Mem/n1572 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1580 ) );
  MUX \Inst_Mem/U1604  ( .A(\Inst_Mem/n1578 ), .B(\Inst_Mem/n1575 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1579 ) );
  MUX \Inst_Mem/U1603  ( .A(\Inst_Mem/n1577 ), .B(\Inst_Mem/n1576 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1578 ) );
  MUX \Inst_Mem/U1602  ( .A(inst_mem_in_wire[1049]), .B(inst_mem_in_wire[1081]), .S(pc_current[2]), .Z(\Inst_Mem/n1577 ) );
  MUX \Inst_Mem/U1601  ( .A(inst_mem_in_wire[1113]), .B(inst_mem_in_wire[1145]), .S(pc_current[2]), .Z(\Inst_Mem/n1576 ) );
  MUX \Inst_Mem/U1600  ( .A(\Inst_Mem/n1574 ), .B(\Inst_Mem/n1573 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1575 ) );
  MUX \Inst_Mem/U1599  ( .A(inst_mem_in_wire[1177]), .B(inst_mem_in_wire[1209]), .S(pc_current[2]), .Z(\Inst_Mem/n1574 ) );
  MUX \Inst_Mem/U1598  ( .A(inst_mem_in_wire[1241]), .B(inst_mem_in_wire[1273]), .S(pc_current[2]), .Z(\Inst_Mem/n1573 ) );
  MUX \Inst_Mem/U1597  ( .A(\Inst_Mem/n1571 ), .B(\Inst_Mem/n1568 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1572 ) );
  MUX \Inst_Mem/U1596  ( .A(\Inst_Mem/n1570 ), .B(\Inst_Mem/n1569 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1571 ) );
  MUX \Inst_Mem/U1595  ( .A(inst_mem_in_wire[1305]), .B(inst_mem_in_wire[1337]), .S(pc_current[2]), .Z(\Inst_Mem/n1570 ) );
  MUX \Inst_Mem/U1594  ( .A(inst_mem_in_wire[1369]), .B(inst_mem_in_wire[1401]), .S(pc_current[2]), .Z(\Inst_Mem/n1569 ) );
  MUX \Inst_Mem/U1593  ( .A(\Inst_Mem/n1567 ), .B(\Inst_Mem/n1566 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1568 ) );
  MUX \Inst_Mem/U1592  ( .A(inst_mem_in_wire[1433]), .B(inst_mem_in_wire[1465]), .S(pc_current[2]), .Z(\Inst_Mem/n1567 ) );
  MUX \Inst_Mem/U1591  ( .A(inst_mem_in_wire[1497]), .B(inst_mem_in_wire[1529]), .S(pc_current[2]), .Z(\Inst_Mem/n1566 ) );
  MUX \Inst_Mem/U1590  ( .A(\Inst_Mem/n1564 ), .B(\Inst_Mem/n1557 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1565 ) );
  MUX \Inst_Mem/U1589  ( .A(\Inst_Mem/n1563 ), .B(\Inst_Mem/n1560 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1564 ) );
  MUX \Inst_Mem/U1588  ( .A(\Inst_Mem/n1562 ), .B(\Inst_Mem/n1561 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1563 ) );
  MUX \Inst_Mem/U1587  ( .A(inst_mem_in_wire[1561]), .B(inst_mem_in_wire[1593]), .S(pc_current[2]), .Z(\Inst_Mem/n1562 ) );
  MUX \Inst_Mem/U1586  ( .A(inst_mem_in_wire[1625]), .B(inst_mem_in_wire[1657]), .S(pc_current[2]), .Z(\Inst_Mem/n1561 ) );
  MUX \Inst_Mem/U1585  ( .A(\Inst_Mem/n1559 ), .B(\Inst_Mem/n1558 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1560 ) );
  MUX \Inst_Mem/U1584  ( .A(inst_mem_in_wire[1689]), .B(inst_mem_in_wire[1721]), .S(pc_current[2]), .Z(\Inst_Mem/n1559 ) );
  MUX \Inst_Mem/U1583  ( .A(inst_mem_in_wire[1753]), .B(inst_mem_in_wire[1785]), .S(pc_current[2]), .Z(\Inst_Mem/n1558 ) );
  MUX \Inst_Mem/U1582  ( .A(\Inst_Mem/n1556 ), .B(\Inst_Mem/n1553 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1557 ) );
  MUX \Inst_Mem/U1581  ( .A(\Inst_Mem/n1555 ), .B(\Inst_Mem/n1554 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1556 ) );
  MUX \Inst_Mem/U1580  ( .A(inst_mem_in_wire[1817]), .B(inst_mem_in_wire[1849]), .S(pc_current[2]), .Z(\Inst_Mem/n1555 ) );
  MUX \Inst_Mem/U1579  ( .A(inst_mem_in_wire[1881]), .B(inst_mem_in_wire[1913]), .S(pc_current[2]), .Z(\Inst_Mem/n1554 ) );
  MUX \Inst_Mem/U1578  ( .A(\Inst_Mem/n1552 ), .B(\Inst_Mem/n1551 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1553 ) );
  MUX \Inst_Mem/U1577  ( .A(inst_mem_in_wire[1945]), .B(inst_mem_in_wire[1977]), .S(pc_current[2]), .Z(\Inst_Mem/n1552 ) );
  MUX \Inst_Mem/U1576  ( .A(inst_mem_in_wire[2009]), .B(inst_mem_in_wire[2041]), .S(pc_current[2]), .Z(\Inst_Mem/n1551 ) );
  MUX \Inst_Mem/U1575  ( .A(\Inst_Mem/n1550 ), .B(\Inst_Mem/n1519 ), .S(
        pc_current[7]), .Z(opcode[24]) );
  MUX \Inst_Mem/U1574  ( .A(\Inst_Mem/n1549 ), .B(\Inst_Mem/n1534 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1550 ) );
  MUX \Inst_Mem/U1573  ( .A(\Inst_Mem/n1548 ), .B(\Inst_Mem/n1541 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1549 ) );
  MUX \Inst_Mem/U1572  ( .A(\Inst_Mem/n1547 ), .B(\Inst_Mem/n1544 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1548 ) );
  MUX \Inst_Mem/U1571  ( .A(\Inst_Mem/n1546 ), .B(\Inst_Mem/n1545 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1547 ) );
  MUX \Inst_Mem/U1570  ( .A(inst_mem_in_wire[24]), .B(inst_mem_in_wire[56]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1546 ) );
  MUX \Inst_Mem/U1569  ( .A(inst_mem_in_wire[88]), .B(inst_mem_in_wire[120]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1545 ) );
  MUX \Inst_Mem/U1568  ( .A(\Inst_Mem/n1543 ), .B(\Inst_Mem/n1542 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1544 ) );
  MUX \Inst_Mem/U1567  ( .A(inst_mem_in_wire[152]), .B(inst_mem_in_wire[184]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1543 ) );
  MUX \Inst_Mem/U1566  ( .A(inst_mem_in_wire[216]), .B(inst_mem_in_wire[248]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1542 ) );
  MUX \Inst_Mem/U1565  ( .A(\Inst_Mem/n1540 ), .B(\Inst_Mem/n1537 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1541 ) );
  MUX \Inst_Mem/U1564  ( .A(\Inst_Mem/n1539 ), .B(\Inst_Mem/n1538 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1540 ) );
  MUX \Inst_Mem/U1563  ( .A(inst_mem_in_wire[280]), .B(inst_mem_in_wire[312]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1539 ) );
  MUX \Inst_Mem/U1562  ( .A(inst_mem_in_wire[344]), .B(inst_mem_in_wire[376]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1538 ) );
  MUX \Inst_Mem/U1561  ( .A(\Inst_Mem/n1536 ), .B(\Inst_Mem/n1535 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1537 ) );
  MUX \Inst_Mem/U1560  ( .A(inst_mem_in_wire[408]), .B(inst_mem_in_wire[440]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1536 ) );
  MUX \Inst_Mem/U1559  ( .A(inst_mem_in_wire[472]), .B(inst_mem_in_wire[504]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1535 ) );
  MUX \Inst_Mem/U1558  ( .A(\Inst_Mem/n1533 ), .B(\Inst_Mem/n1526 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1534 ) );
  MUX \Inst_Mem/U1557  ( .A(\Inst_Mem/n1532 ), .B(\Inst_Mem/n1529 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1533 ) );
  MUX \Inst_Mem/U1556  ( .A(\Inst_Mem/n1531 ), .B(\Inst_Mem/n1530 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1532 ) );
  MUX \Inst_Mem/U1555  ( .A(inst_mem_in_wire[536]), .B(inst_mem_in_wire[568]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1531 ) );
  MUX \Inst_Mem/U1554  ( .A(inst_mem_in_wire[600]), .B(inst_mem_in_wire[632]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1530 ) );
  MUX \Inst_Mem/U1553  ( .A(\Inst_Mem/n1528 ), .B(\Inst_Mem/n1527 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1529 ) );
  MUX \Inst_Mem/U1552  ( .A(inst_mem_in_wire[664]), .B(inst_mem_in_wire[696]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1528 ) );
  MUX \Inst_Mem/U1551  ( .A(inst_mem_in_wire[728]), .B(inst_mem_in_wire[760]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1527 ) );
  MUX \Inst_Mem/U1550  ( .A(\Inst_Mem/n1525 ), .B(\Inst_Mem/n1522 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1526 ) );
  MUX \Inst_Mem/U1549  ( .A(\Inst_Mem/n1524 ), .B(\Inst_Mem/n1523 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1525 ) );
  MUX \Inst_Mem/U1548  ( .A(inst_mem_in_wire[792]), .B(inst_mem_in_wire[824]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1524 ) );
  MUX \Inst_Mem/U1547  ( .A(inst_mem_in_wire[856]), .B(inst_mem_in_wire[888]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1523 ) );
  MUX \Inst_Mem/U1546  ( .A(\Inst_Mem/n1521 ), .B(\Inst_Mem/n1520 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1522 ) );
  MUX \Inst_Mem/U1545  ( .A(inst_mem_in_wire[920]), .B(inst_mem_in_wire[952]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1521 ) );
  MUX \Inst_Mem/U1544  ( .A(inst_mem_in_wire[984]), .B(inst_mem_in_wire[1016]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1520 ) );
  MUX \Inst_Mem/U1543  ( .A(\Inst_Mem/n1518 ), .B(\Inst_Mem/n1503 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1519 ) );
  MUX \Inst_Mem/U1542  ( .A(\Inst_Mem/n1517 ), .B(\Inst_Mem/n1510 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1518 ) );
  MUX \Inst_Mem/U1541  ( .A(\Inst_Mem/n1516 ), .B(\Inst_Mem/n1513 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1517 ) );
  MUX \Inst_Mem/U1540  ( .A(\Inst_Mem/n1515 ), .B(\Inst_Mem/n1514 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1516 ) );
  MUX \Inst_Mem/U1539  ( .A(inst_mem_in_wire[1048]), .B(inst_mem_in_wire[1080]), .S(pc_current[2]), .Z(\Inst_Mem/n1515 ) );
  MUX \Inst_Mem/U1538  ( .A(inst_mem_in_wire[1112]), .B(inst_mem_in_wire[1144]), .S(pc_current[2]), .Z(\Inst_Mem/n1514 ) );
  MUX \Inst_Mem/U1537  ( .A(\Inst_Mem/n1512 ), .B(\Inst_Mem/n1511 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1513 ) );
  MUX \Inst_Mem/U1536  ( .A(inst_mem_in_wire[1176]), .B(inst_mem_in_wire[1208]), .S(pc_current[2]), .Z(\Inst_Mem/n1512 ) );
  MUX \Inst_Mem/U1535  ( .A(inst_mem_in_wire[1240]), .B(inst_mem_in_wire[1272]), .S(pc_current[2]), .Z(\Inst_Mem/n1511 ) );
  MUX \Inst_Mem/U1534  ( .A(\Inst_Mem/n1509 ), .B(\Inst_Mem/n1506 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1510 ) );
  MUX \Inst_Mem/U1533  ( .A(\Inst_Mem/n1508 ), .B(\Inst_Mem/n1507 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1509 ) );
  MUX \Inst_Mem/U1532  ( .A(inst_mem_in_wire[1304]), .B(inst_mem_in_wire[1336]), .S(pc_current[2]), .Z(\Inst_Mem/n1508 ) );
  MUX \Inst_Mem/U1531  ( .A(inst_mem_in_wire[1368]), .B(inst_mem_in_wire[1400]), .S(pc_current[2]), .Z(\Inst_Mem/n1507 ) );
  MUX \Inst_Mem/U1530  ( .A(\Inst_Mem/n1505 ), .B(\Inst_Mem/n1504 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1506 ) );
  MUX \Inst_Mem/U1529  ( .A(inst_mem_in_wire[1432]), .B(inst_mem_in_wire[1464]), .S(pc_current[2]), .Z(\Inst_Mem/n1505 ) );
  MUX \Inst_Mem/U1528  ( .A(inst_mem_in_wire[1496]), .B(inst_mem_in_wire[1528]), .S(pc_current[2]), .Z(\Inst_Mem/n1504 ) );
  MUX \Inst_Mem/U1527  ( .A(\Inst_Mem/n1502 ), .B(\Inst_Mem/n1495 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1503 ) );
  MUX \Inst_Mem/U1526  ( .A(\Inst_Mem/n1501 ), .B(\Inst_Mem/n1498 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1502 ) );
  MUX \Inst_Mem/U1525  ( .A(\Inst_Mem/n1500 ), .B(\Inst_Mem/n1499 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1501 ) );
  MUX \Inst_Mem/U1524  ( .A(inst_mem_in_wire[1560]), .B(inst_mem_in_wire[1592]), .S(pc_current[2]), .Z(\Inst_Mem/n1500 ) );
  MUX \Inst_Mem/U1523  ( .A(inst_mem_in_wire[1624]), .B(inst_mem_in_wire[1656]), .S(pc_current[2]), .Z(\Inst_Mem/n1499 ) );
  MUX \Inst_Mem/U1522  ( .A(\Inst_Mem/n1497 ), .B(\Inst_Mem/n1496 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1498 ) );
  MUX \Inst_Mem/U1521  ( .A(inst_mem_in_wire[1688]), .B(inst_mem_in_wire[1720]), .S(pc_current[2]), .Z(\Inst_Mem/n1497 ) );
  MUX \Inst_Mem/U1520  ( .A(inst_mem_in_wire[1752]), .B(inst_mem_in_wire[1784]), .S(pc_current[2]), .Z(\Inst_Mem/n1496 ) );
  MUX \Inst_Mem/U1519  ( .A(\Inst_Mem/n1494 ), .B(\Inst_Mem/n1491 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1495 ) );
  MUX \Inst_Mem/U1518  ( .A(\Inst_Mem/n1493 ), .B(\Inst_Mem/n1492 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1494 ) );
  MUX \Inst_Mem/U1517  ( .A(inst_mem_in_wire[1816]), .B(inst_mem_in_wire[1848]), .S(pc_current[2]), .Z(\Inst_Mem/n1493 ) );
  MUX \Inst_Mem/U1516  ( .A(inst_mem_in_wire[1880]), .B(inst_mem_in_wire[1912]), .S(pc_current[2]), .Z(\Inst_Mem/n1492 ) );
  MUX \Inst_Mem/U1515  ( .A(\Inst_Mem/n1490 ), .B(\Inst_Mem/n1489 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1491 ) );
  MUX \Inst_Mem/U1514  ( .A(inst_mem_in_wire[1944]), .B(inst_mem_in_wire[1976]), .S(pc_current[2]), .Z(\Inst_Mem/n1490 ) );
  MUX \Inst_Mem/U1513  ( .A(inst_mem_in_wire[2008]), .B(inst_mem_in_wire[2040]), .S(pc_current[2]), .Z(\Inst_Mem/n1489 ) );
  MUX \Inst_Mem/U1512  ( .A(\Inst_Mem/n1488 ), .B(\Inst_Mem/n1457 ), .S(
        pc_current[7]), .Z(opcode[23]) );
  MUX \Inst_Mem/U1511  ( .A(\Inst_Mem/n1487 ), .B(\Inst_Mem/n1472 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1488 ) );
  MUX \Inst_Mem/U1510  ( .A(\Inst_Mem/n1486 ), .B(\Inst_Mem/n1479 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1487 ) );
  MUX \Inst_Mem/U1509  ( .A(\Inst_Mem/n1485 ), .B(\Inst_Mem/n1482 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1486 ) );
  MUX \Inst_Mem/U1508  ( .A(\Inst_Mem/n1484 ), .B(\Inst_Mem/n1483 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1485 ) );
  MUX \Inst_Mem/U1507  ( .A(inst_mem_in_wire[23]), .B(inst_mem_in_wire[55]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1484 ) );
  MUX \Inst_Mem/U1506  ( .A(inst_mem_in_wire[87]), .B(inst_mem_in_wire[119]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1483 ) );
  MUX \Inst_Mem/U1505  ( .A(\Inst_Mem/n1481 ), .B(\Inst_Mem/n1480 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1482 ) );
  MUX \Inst_Mem/U1504  ( .A(inst_mem_in_wire[151]), .B(inst_mem_in_wire[183]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1481 ) );
  MUX \Inst_Mem/U1503  ( .A(inst_mem_in_wire[215]), .B(inst_mem_in_wire[247]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1480 ) );
  MUX \Inst_Mem/U1502  ( .A(\Inst_Mem/n1478 ), .B(\Inst_Mem/n1475 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1479 ) );
  MUX \Inst_Mem/U1501  ( .A(\Inst_Mem/n1477 ), .B(\Inst_Mem/n1476 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1478 ) );
  MUX \Inst_Mem/U1500  ( .A(inst_mem_in_wire[279]), .B(inst_mem_in_wire[311]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1477 ) );
  MUX \Inst_Mem/U1499  ( .A(inst_mem_in_wire[343]), .B(inst_mem_in_wire[375]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1476 ) );
  MUX \Inst_Mem/U1498  ( .A(\Inst_Mem/n1474 ), .B(\Inst_Mem/n1473 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1475 ) );
  MUX \Inst_Mem/U1497  ( .A(inst_mem_in_wire[407]), .B(inst_mem_in_wire[439]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1474 ) );
  MUX \Inst_Mem/U1496  ( .A(inst_mem_in_wire[471]), .B(inst_mem_in_wire[503]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1473 ) );
  MUX \Inst_Mem/U1495  ( .A(\Inst_Mem/n1471 ), .B(\Inst_Mem/n1464 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1472 ) );
  MUX \Inst_Mem/U1494  ( .A(\Inst_Mem/n1470 ), .B(\Inst_Mem/n1467 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1471 ) );
  MUX \Inst_Mem/U1493  ( .A(\Inst_Mem/n1469 ), .B(\Inst_Mem/n1468 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1470 ) );
  MUX \Inst_Mem/U1492  ( .A(inst_mem_in_wire[535]), .B(inst_mem_in_wire[567]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1469 ) );
  MUX \Inst_Mem/U1491  ( .A(inst_mem_in_wire[599]), .B(inst_mem_in_wire[631]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1468 ) );
  MUX \Inst_Mem/U1490  ( .A(\Inst_Mem/n1466 ), .B(\Inst_Mem/n1465 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1467 ) );
  MUX \Inst_Mem/U1489  ( .A(inst_mem_in_wire[663]), .B(inst_mem_in_wire[695]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1466 ) );
  MUX \Inst_Mem/U1488  ( .A(inst_mem_in_wire[727]), .B(inst_mem_in_wire[759]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1465 ) );
  MUX \Inst_Mem/U1487  ( .A(\Inst_Mem/n1463 ), .B(\Inst_Mem/n1460 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1464 ) );
  MUX \Inst_Mem/U1486  ( .A(\Inst_Mem/n1462 ), .B(\Inst_Mem/n1461 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1463 ) );
  MUX \Inst_Mem/U1485  ( .A(inst_mem_in_wire[791]), .B(inst_mem_in_wire[823]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1462 ) );
  MUX \Inst_Mem/U1484  ( .A(inst_mem_in_wire[855]), .B(inst_mem_in_wire[887]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1461 ) );
  MUX \Inst_Mem/U1483  ( .A(\Inst_Mem/n1459 ), .B(\Inst_Mem/n1458 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1460 ) );
  MUX \Inst_Mem/U1482  ( .A(inst_mem_in_wire[919]), .B(inst_mem_in_wire[951]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1459 ) );
  MUX \Inst_Mem/U1481  ( .A(inst_mem_in_wire[983]), .B(inst_mem_in_wire[1015]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1458 ) );
  MUX \Inst_Mem/U1480  ( .A(\Inst_Mem/n1456 ), .B(\Inst_Mem/n1441 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1457 ) );
  MUX \Inst_Mem/U1479  ( .A(\Inst_Mem/n1455 ), .B(\Inst_Mem/n1448 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1456 ) );
  MUX \Inst_Mem/U1478  ( .A(\Inst_Mem/n1454 ), .B(\Inst_Mem/n1451 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1455 ) );
  MUX \Inst_Mem/U1477  ( .A(\Inst_Mem/n1453 ), .B(\Inst_Mem/n1452 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1454 ) );
  MUX \Inst_Mem/U1476  ( .A(inst_mem_in_wire[1047]), .B(inst_mem_in_wire[1079]), .S(pc_current[2]), .Z(\Inst_Mem/n1453 ) );
  MUX \Inst_Mem/U1475  ( .A(inst_mem_in_wire[1111]), .B(inst_mem_in_wire[1143]), .S(pc_current[2]), .Z(\Inst_Mem/n1452 ) );
  MUX \Inst_Mem/U1474  ( .A(\Inst_Mem/n1450 ), .B(\Inst_Mem/n1449 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1451 ) );
  MUX \Inst_Mem/U1473  ( .A(inst_mem_in_wire[1175]), .B(inst_mem_in_wire[1207]), .S(pc_current[2]), .Z(\Inst_Mem/n1450 ) );
  MUX \Inst_Mem/U1472  ( .A(inst_mem_in_wire[1239]), .B(inst_mem_in_wire[1271]), .S(pc_current[2]), .Z(\Inst_Mem/n1449 ) );
  MUX \Inst_Mem/U1471  ( .A(\Inst_Mem/n1447 ), .B(\Inst_Mem/n1444 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1448 ) );
  MUX \Inst_Mem/U1470  ( .A(\Inst_Mem/n1446 ), .B(\Inst_Mem/n1445 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1447 ) );
  MUX \Inst_Mem/U1469  ( .A(inst_mem_in_wire[1303]), .B(inst_mem_in_wire[1335]), .S(pc_current[2]), .Z(\Inst_Mem/n1446 ) );
  MUX \Inst_Mem/U1468  ( .A(inst_mem_in_wire[1367]), .B(inst_mem_in_wire[1399]), .S(pc_current[2]), .Z(\Inst_Mem/n1445 ) );
  MUX \Inst_Mem/U1467  ( .A(\Inst_Mem/n1443 ), .B(\Inst_Mem/n1442 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1444 ) );
  MUX \Inst_Mem/U1466  ( .A(inst_mem_in_wire[1431]), .B(inst_mem_in_wire[1463]), .S(pc_current[2]), .Z(\Inst_Mem/n1443 ) );
  MUX \Inst_Mem/U1465  ( .A(inst_mem_in_wire[1495]), .B(inst_mem_in_wire[1527]), .S(pc_current[2]), .Z(\Inst_Mem/n1442 ) );
  MUX \Inst_Mem/U1464  ( .A(\Inst_Mem/n1440 ), .B(\Inst_Mem/n1433 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1441 ) );
  MUX \Inst_Mem/U1463  ( .A(\Inst_Mem/n1439 ), .B(\Inst_Mem/n1436 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1440 ) );
  MUX \Inst_Mem/U1462  ( .A(\Inst_Mem/n1438 ), .B(\Inst_Mem/n1437 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1439 ) );
  MUX \Inst_Mem/U1461  ( .A(inst_mem_in_wire[1559]), .B(inst_mem_in_wire[1591]), .S(pc_current[2]), .Z(\Inst_Mem/n1438 ) );
  MUX \Inst_Mem/U1460  ( .A(inst_mem_in_wire[1623]), .B(inst_mem_in_wire[1655]), .S(pc_current[2]), .Z(\Inst_Mem/n1437 ) );
  MUX \Inst_Mem/U1459  ( .A(\Inst_Mem/n1435 ), .B(\Inst_Mem/n1434 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1436 ) );
  MUX \Inst_Mem/U1458  ( .A(inst_mem_in_wire[1687]), .B(inst_mem_in_wire[1719]), .S(pc_current[2]), .Z(\Inst_Mem/n1435 ) );
  MUX \Inst_Mem/U1457  ( .A(inst_mem_in_wire[1751]), .B(inst_mem_in_wire[1783]), .S(pc_current[2]), .Z(\Inst_Mem/n1434 ) );
  MUX \Inst_Mem/U1456  ( .A(\Inst_Mem/n1432 ), .B(\Inst_Mem/n1429 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1433 ) );
  MUX \Inst_Mem/U1455  ( .A(\Inst_Mem/n1431 ), .B(\Inst_Mem/n1430 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1432 ) );
  MUX \Inst_Mem/U1454  ( .A(inst_mem_in_wire[1815]), .B(inst_mem_in_wire[1847]), .S(pc_current[2]), .Z(\Inst_Mem/n1431 ) );
  MUX \Inst_Mem/U1453  ( .A(inst_mem_in_wire[1879]), .B(inst_mem_in_wire[1911]), .S(pc_current[2]), .Z(\Inst_Mem/n1430 ) );
  MUX \Inst_Mem/U1452  ( .A(\Inst_Mem/n1428 ), .B(\Inst_Mem/n1427 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1429 ) );
  MUX \Inst_Mem/U1451  ( .A(inst_mem_in_wire[1943]), .B(inst_mem_in_wire[1975]), .S(pc_current[2]), .Z(\Inst_Mem/n1428 ) );
  MUX \Inst_Mem/U1450  ( .A(inst_mem_in_wire[2007]), .B(inst_mem_in_wire[2039]), .S(pc_current[2]), .Z(\Inst_Mem/n1427 ) );
  MUX \Inst_Mem/U1449  ( .A(\Inst_Mem/n1426 ), .B(\Inst_Mem/n1395 ), .S(
        pc_current[7]), .Z(opcode[22]) );
  MUX \Inst_Mem/U1448  ( .A(\Inst_Mem/n1425 ), .B(\Inst_Mem/n1410 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1426 ) );
  MUX \Inst_Mem/U1447  ( .A(\Inst_Mem/n1424 ), .B(\Inst_Mem/n1417 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1425 ) );
  MUX \Inst_Mem/U1446  ( .A(\Inst_Mem/n1423 ), .B(\Inst_Mem/n1420 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1424 ) );
  MUX \Inst_Mem/U1445  ( .A(\Inst_Mem/n1422 ), .B(\Inst_Mem/n1421 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1423 ) );
  MUX \Inst_Mem/U1444  ( .A(inst_mem_in_wire[22]), .B(inst_mem_in_wire[54]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1422 ) );
  MUX \Inst_Mem/U1443  ( .A(inst_mem_in_wire[86]), .B(inst_mem_in_wire[118]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1421 ) );
  MUX \Inst_Mem/U1442  ( .A(\Inst_Mem/n1419 ), .B(\Inst_Mem/n1418 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1420 ) );
  MUX \Inst_Mem/U1441  ( .A(inst_mem_in_wire[150]), .B(inst_mem_in_wire[182]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1419 ) );
  MUX \Inst_Mem/U1440  ( .A(inst_mem_in_wire[214]), .B(inst_mem_in_wire[246]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1418 ) );
  MUX \Inst_Mem/U1439  ( .A(\Inst_Mem/n1416 ), .B(\Inst_Mem/n1413 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1417 ) );
  MUX \Inst_Mem/U1438  ( .A(\Inst_Mem/n1415 ), .B(\Inst_Mem/n1414 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1416 ) );
  MUX \Inst_Mem/U1437  ( .A(inst_mem_in_wire[278]), .B(inst_mem_in_wire[310]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1415 ) );
  MUX \Inst_Mem/U1436  ( .A(inst_mem_in_wire[342]), .B(inst_mem_in_wire[374]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1414 ) );
  MUX \Inst_Mem/U1435  ( .A(\Inst_Mem/n1412 ), .B(\Inst_Mem/n1411 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1413 ) );
  MUX \Inst_Mem/U1434  ( .A(inst_mem_in_wire[406]), .B(inst_mem_in_wire[438]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1412 ) );
  MUX \Inst_Mem/U1433  ( .A(inst_mem_in_wire[470]), .B(inst_mem_in_wire[502]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1411 ) );
  MUX \Inst_Mem/U1432  ( .A(\Inst_Mem/n1409 ), .B(\Inst_Mem/n1402 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1410 ) );
  MUX \Inst_Mem/U1431  ( .A(\Inst_Mem/n1408 ), .B(\Inst_Mem/n1405 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1409 ) );
  MUX \Inst_Mem/U1430  ( .A(\Inst_Mem/n1407 ), .B(\Inst_Mem/n1406 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1408 ) );
  MUX \Inst_Mem/U1429  ( .A(inst_mem_in_wire[534]), .B(inst_mem_in_wire[566]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1407 ) );
  MUX \Inst_Mem/U1428  ( .A(inst_mem_in_wire[598]), .B(inst_mem_in_wire[630]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1406 ) );
  MUX \Inst_Mem/U1427  ( .A(\Inst_Mem/n1404 ), .B(\Inst_Mem/n1403 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1405 ) );
  MUX \Inst_Mem/U1426  ( .A(inst_mem_in_wire[662]), .B(inst_mem_in_wire[694]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1404 ) );
  MUX \Inst_Mem/U1425  ( .A(inst_mem_in_wire[726]), .B(inst_mem_in_wire[758]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1403 ) );
  MUX \Inst_Mem/U1424  ( .A(\Inst_Mem/n1401 ), .B(\Inst_Mem/n1398 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1402 ) );
  MUX \Inst_Mem/U1423  ( .A(\Inst_Mem/n1400 ), .B(\Inst_Mem/n1399 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1401 ) );
  MUX \Inst_Mem/U1422  ( .A(inst_mem_in_wire[790]), .B(inst_mem_in_wire[822]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1400 ) );
  MUX \Inst_Mem/U1421  ( .A(inst_mem_in_wire[854]), .B(inst_mem_in_wire[886]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1399 ) );
  MUX \Inst_Mem/U1420  ( .A(\Inst_Mem/n1397 ), .B(\Inst_Mem/n1396 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1398 ) );
  MUX \Inst_Mem/U1419  ( .A(inst_mem_in_wire[918]), .B(inst_mem_in_wire[950]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1397 ) );
  MUX \Inst_Mem/U1418  ( .A(inst_mem_in_wire[982]), .B(inst_mem_in_wire[1014]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1396 ) );
  MUX \Inst_Mem/U1417  ( .A(\Inst_Mem/n1394 ), .B(\Inst_Mem/n1379 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1395 ) );
  MUX \Inst_Mem/U1416  ( .A(\Inst_Mem/n1393 ), .B(\Inst_Mem/n1386 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1394 ) );
  MUX \Inst_Mem/U1415  ( .A(\Inst_Mem/n1392 ), .B(\Inst_Mem/n1389 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1393 ) );
  MUX \Inst_Mem/U1414  ( .A(\Inst_Mem/n1391 ), .B(\Inst_Mem/n1390 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1392 ) );
  MUX \Inst_Mem/U1413  ( .A(inst_mem_in_wire[1046]), .B(inst_mem_in_wire[1078]), .S(pc_current[2]), .Z(\Inst_Mem/n1391 ) );
  MUX \Inst_Mem/U1412  ( .A(inst_mem_in_wire[1110]), .B(inst_mem_in_wire[1142]), .S(pc_current[2]), .Z(\Inst_Mem/n1390 ) );
  MUX \Inst_Mem/U1411  ( .A(\Inst_Mem/n1388 ), .B(\Inst_Mem/n1387 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1389 ) );
  MUX \Inst_Mem/U1410  ( .A(inst_mem_in_wire[1174]), .B(inst_mem_in_wire[1206]), .S(pc_current[2]), .Z(\Inst_Mem/n1388 ) );
  MUX \Inst_Mem/U1409  ( .A(inst_mem_in_wire[1238]), .B(inst_mem_in_wire[1270]), .S(pc_current[2]), .Z(\Inst_Mem/n1387 ) );
  MUX \Inst_Mem/U1408  ( .A(\Inst_Mem/n1385 ), .B(\Inst_Mem/n1382 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1386 ) );
  MUX \Inst_Mem/U1407  ( .A(\Inst_Mem/n1384 ), .B(\Inst_Mem/n1383 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1385 ) );
  MUX \Inst_Mem/U1406  ( .A(inst_mem_in_wire[1302]), .B(inst_mem_in_wire[1334]), .S(pc_current[2]), .Z(\Inst_Mem/n1384 ) );
  MUX \Inst_Mem/U1405  ( .A(inst_mem_in_wire[1366]), .B(inst_mem_in_wire[1398]), .S(pc_current[2]), .Z(\Inst_Mem/n1383 ) );
  MUX \Inst_Mem/U1404  ( .A(\Inst_Mem/n1381 ), .B(\Inst_Mem/n1380 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1382 ) );
  MUX \Inst_Mem/U1403  ( .A(inst_mem_in_wire[1430]), .B(inst_mem_in_wire[1462]), .S(pc_current[2]), .Z(\Inst_Mem/n1381 ) );
  MUX \Inst_Mem/U1402  ( .A(inst_mem_in_wire[1494]), .B(inst_mem_in_wire[1526]), .S(pc_current[2]), .Z(\Inst_Mem/n1380 ) );
  MUX \Inst_Mem/U1401  ( .A(\Inst_Mem/n1378 ), .B(\Inst_Mem/n1371 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1379 ) );
  MUX \Inst_Mem/U1400  ( .A(\Inst_Mem/n1377 ), .B(\Inst_Mem/n1374 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1378 ) );
  MUX \Inst_Mem/U1399  ( .A(\Inst_Mem/n1376 ), .B(\Inst_Mem/n1375 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1377 ) );
  MUX \Inst_Mem/U1398  ( .A(inst_mem_in_wire[1558]), .B(inst_mem_in_wire[1590]), .S(pc_current[2]), .Z(\Inst_Mem/n1376 ) );
  MUX \Inst_Mem/U1397  ( .A(inst_mem_in_wire[1622]), .B(inst_mem_in_wire[1654]), .S(pc_current[2]), .Z(\Inst_Mem/n1375 ) );
  MUX \Inst_Mem/U1396  ( .A(\Inst_Mem/n1373 ), .B(\Inst_Mem/n1372 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1374 ) );
  MUX \Inst_Mem/U1395  ( .A(inst_mem_in_wire[1686]), .B(inst_mem_in_wire[1718]), .S(pc_current[2]), .Z(\Inst_Mem/n1373 ) );
  MUX \Inst_Mem/U1394  ( .A(inst_mem_in_wire[1750]), .B(inst_mem_in_wire[1782]), .S(pc_current[2]), .Z(\Inst_Mem/n1372 ) );
  MUX \Inst_Mem/U1393  ( .A(\Inst_Mem/n1370 ), .B(\Inst_Mem/n1367 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1371 ) );
  MUX \Inst_Mem/U1392  ( .A(\Inst_Mem/n1369 ), .B(\Inst_Mem/n1368 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1370 ) );
  MUX \Inst_Mem/U1391  ( .A(inst_mem_in_wire[1814]), .B(inst_mem_in_wire[1846]), .S(pc_current[2]), .Z(\Inst_Mem/n1369 ) );
  MUX \Inst_Mem/U1390  ( .A(inst_mem_in_wire[1878]), .B(inst_mem_in_wire[1910]), .S(pc_current[2]), .Z(\Inst_Mem/n1368 ) );
  MUX \Inst_Mem/U1389  ( .A(\Inst_Mem/n1366 ), .B(\Inst_Mem/n1365 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1367 ) );
  MUX \Inst_Mem/U1388  ( .A(inst_mem_in_wire[1942]), .B(inst_mem_in_wire[1974]), .S(pc_current[2]), .Z(\Inst_Mem/n1366 ) );
  MUX \Inst_Mem/U1387  ( .A(inst_mem_in_wire[2006]), .B(inst_mem_in_wire[2038]), .S(pc_current[2]), .Z(\Inst_Mem/n1365 ) );
  MUX \Inst_Mem/U1386  ( .A(\Inst_Mem/n1364 ), .B(\Inst_Mem/n1333 ), .S(
        pc_current[7]), .Z(opcode[21]) );
  MUX \Inst_Mem/U1385  ( .A(\Inst_Mem/n1363 ), .B(\Inst_Mem/n1348 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1364 ) );
  MUX \Inst_Mem/U1384  ( .A(\Inst_Mem/n1362 ), .B(\Inst_Mem/n1355 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1363 ) );
  MUX \Inst_Mem/U1383  ( .A(\Inst_Mem/n1361 ), .B(\Inst_Mem/n1358 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1362 ) );
  MUX \Inst_Mem/U1382  ( .A(\Inst_Mem/n1360 ), .B(\Inst_Mem/n1359 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1361 ) );
  MUX \Inst_Mem/U1381  ( .A(inst_mem_in_wire[21]), .B(inst_mem_in_wire[53]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1360 ) );
  MUX \Inst_Mem/U1380  ( .A(inst_mem_in_wire[85]), .B(inst_mem_in_wire[117]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1359 ) );
  MUX \Inst_Mem/U1379  ( .A(\Inst_Mem/n1357 ), .B(\Inst_Mem/n1356 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1358 ) );
  MUX \Inst_Mem/U1378  ( .A(inst_mem_in_wire[149]), .B(inst_mem_in_wire[181]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1357 ) );
  MUX \Inst_Mem/U1377  ( .A(inst_mem_in_wire[213]), .B(inst_mem_in_wire[245]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1356 ) );
  MUX \Inst_Mem/U1376  ( .A(\Inst_Mem/n1354 ), .B(\Inst_Mem/n1351 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1355 ) );
  MUX \Inst_Mem/U1375  ( .A(\Inst_Mem/n1353 ), .B(\Inst_Mem/n1352 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1354 ) );
  MUX \Inst_Mem/U1374  ( .A(inst_mem_in_wire[277]), .B(inst_mem_in_wire[309]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1353 ) );
  MUX \Inst_Mem/U1373  ( .A(inst_mem_in_wire[341]), .B(inst_mem_in_wire[373]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1352 ) );
  MUX \Inst_Mem/U1372  ( .A(\Inst_Mem/n1350 ), .B(\Inst_Mem/n1349 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1351 ) );
  MUX \Inst_Mem/U1371  ( .A(inst_mem_in_wire[405]), .B(inst_mem_in_wire[437]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1350 ) );
  MUX \Inst_Mem/U1370  ( .A(inst_mem_in_wire[469]), .B(inst_mem_in_wire[501]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1349 ) );
  MUX \Inst_Mem/U1369  ( .A(\Inst_Mem/n1347 ), .B(\Inst_Mem/n1340 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1348 ) );
  MUX \Inst_Mem/U1368  ( .A(\Inst_Mem/n1346 ), .B(\Inst_Mem/n1343 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1347 ) );
  MUX \Inst_Mem/U1367  ( .A(\Inst_Mem/n1345 ), .B(\Inst_Mem/n1344 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1346 ) );
  MUX \Inst_Mem/U1366  ( .A(inst_mem_in_wire[533]), .B(inst_mem_in_wire[565]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1345 ) );
  MUX \Inst_Mem/U1365  ( .A(inst_mem_in_wire[597]), .B(inst_mem_in_wire[629]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1344 ) );
  MUX \Inst_Mem/U1364  ( .A(\Inst_Mem/n1342 ), .B(\Inst_Mem/n1341 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1343 ) );
  MUX \Inst_Mem/U1363  ( .A(inst_mem_in_wire[661]), .B(inst_mem_in_wire[693]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1342 ) );
  MUX \Inst_Mem/U1362  ( .A(inst_mem_in_wire[725]), .B(inst_mem_in_wire[757]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1341 ) );
  MUX \Inst_Mem/U1361  ( .A(\Inst_Mem/n1339 ), .B(\Inst_Mem/n1336 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1340 ) );
  MUX \Inst_Mem/U1360  ( .A(\Inst_Mem/n1338 ), .B(\Inst_Mem/n1337 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1339 ) );
  MUX \Inst_Mem/U1359  ( .A(inst_mem_in_wire[789]), .B(inst_mem_in_wire[821]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1338 ) );
  MUX \Inst_Mem/U1358  ( .A(inst_mem_in_wire[853]), .B(inst_mem_in_wire[885]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1337 ) );
  MUX \Inst_Mem/U1357  ( .A(\Inst_Mem/n1335 ), .B(\Inst_Mem/n1334 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1336 ) );
  MUX \Inst_Mem/U1356  ( .A(inst_mem_in_wire[917]), .B(inst_mem_in_wire[949]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1335 ) );
  MUX \Inst_Mem/U1355  ( .A(inst_mem_in_wire[981]), .B(inst_mem_in_wire[1013]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1334 ) );
  MUX \Inst_Mem/U1354  ( .A(\Inst_Mem/n1332 ), .B(\Inst_Mem/n1317 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1333 ) );
  MUX \Inst_Mem/U1353  ( .A(\Inst_Mem/n1331 ), .B(\Inst_Mem/n1324 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1332 ) );
  MUX \Inst_Mem/U1352  ( .A(\Inst_Mem/n1330 ), .B(\Inst_Mem/n1327 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1331 ) );
  MUX \Inst_Mem/U1351  ( .A(\Inst_Mem/n1329 ), .B(\Inst_Mem/n1328 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1330 ) );
  MUX \Inst_Mem/U1350  ( .A(inst_mem_in_wire[1045]), .B(inst_mem_in_wire[1077]), .S(pc_current[2]), .Z(\Inst_Mem/n1329 ) );
  MUX \Inst_Mem/U1349  ( .A(inst_mem_in_wire[1109]), .B(inst_mem_in_wire[1141]), .S(pc_current[2]), .Z(\Inst_Mem/n1328 ) );
  MUX \Inst_Mem/U1348  ( .A(\Inst_Mem/n1326 ), .B(\Inst_Mem/n1325 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1327 ) );
  MUX \Inst_Mem/U1347  ( .A(inst_mem_in_wire[1173]), .B(inst_mem_in_wire[1205]), .S(pc_current[2]), .Z(\Inst_Mem/n1326 ) );
  MUX \Inst_Mem/U1346  ( .A(inst_mem_in_wire[1237]), .B(inst_mem_in_wire[1269]), .S(pc_current[2]), .Z(\Inst_Mem/n1325 ) );
  MUX \Inst_Mem/U1345  ( .A(\Inst_Mem/n1323 ), .B(\Inst_Mem/n1320 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1324 ) );
  MUX \Inst_Mem/U1344  ( .A(\Inst_Mem/n1322 ), .B(\Inst_Mem/n1321 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1323 ) );
  MUX \Inst_Mem/U1343  ( .A(inst_mem_in_wire[1301]), .B(inst_mem_in_wire[1333]), .S(pc_current[2]), .Z(\Inst_Mem/n1322 ) );
  MUX \Inst_Mem/U1342  ( .A(inst_mem_in_wire[1365]), .B(inst_mem_in_wire[1397]), .S(pc_current[2]), .Z(\Inst_Mem/n1321 ) );
  MUX \Inst_Mem/U1341  ( .A(\Inst_Mem/n1319 ), .B(\Inst_Mem/n1318 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1320 ) );
  MUX \Inst_Mem/U1340  ( .A(inst_mem_in_wire[1429]), .B(inst_mem_in_wire[1461]), .S(pc_current[2]), .Z(\Inst_Mem/n1319 ) );
  MUX \Inst_Mem/U1339  ( .A(inst_mem_in_wire[1493]), .B(inst_mem_in_wire[1525]), .S(pc_current[2]), .Z(\Inst_Mem/n1318 ) );
  MUX \Inst_Mem/U1338  ( .A(\Inst_Mem/n1316 ), .B(\Inst_Mem/n1309 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1317 ) );
  MUX \Inst_Mem/U1337  ( .A(\Inst_Mem/n1315 ), .B(\Inst_Mem/n1312 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1316 ) );
  MUX \Inst_Mem/U1336  ( .A(\Inst_Mem/n1314 ), .B(\Inst_Mem/n1313 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1315 ) );
  MUX \Inst_Mem/U1335  ( .A(inst_mem_in_wire[1557]), .B(inst_mem_in_wire[1589]), .S(pc_current[2]), .Z(\Inst_Mem/n1314 ) );
  MUX \Inst_Mem/U1334  ( .A(inst_mem_in_wire[1621]), .B(inst_mem_in_wire[1653]), .S(pc_current[2]), .Z(\Inst_Mem/n1313 ) );
  MUX \Inst_Mem/U1333  ( .A(\Inst_Mem/n1311 ), .B(\Inst_Mem/n1310 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1312 ) );
  MUX \Inst_Mem/U1332  ( .A(inst_mem_in_wire[1685]), .B(inst_mem_in_wire[1717]), .S(pc_current[2]), .Z(\Inst_Mem/n1311 ) );
  MUX \Inst_Mem/U1331  ( .A(inst_mem_in_wire[1749]), .B(inst_mem_in_wire[1781]), .S(pc_current[2]), .Z(\Inst_Mem/n1310 ) );
  MUX \Inst_Mem/U1330  ( .A(\Inst_Mem/n1308 ), .B(\Inst_Mem/n1305 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1309 ) );
  MUX \Inst_Mem/U1329  ( .A(\Inst_Mem/n1307 ), .B(\Inst_Mem/n1306 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1308 ) );
  MUX \Inst_Mem/U1328  ( .A(inst_mem_in_wire[1813]), .B(inst_mem_in_wire[1845]), .S(pc_current[2]), .Z(\Inst_Mem/n1307 ) );
  MUX \Inst_Mem/U1327  ( .A(inst_mem_in_wire[1877]), .B(inst_mem_in_wire[1909]), .S(pc_current[2]), .Z(\Inst_Mem/n1306 ) );
  MUX \Inst_Mem/U1326  ( .A(\Inst_Mem/n1304 ), .B(\Inst_Mem/n1303 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1305 ) );
  MUX \Inst_Mem/U1325  ( .A(inst_mem_in_wire[1941]), .B(inst_mem_in_wire[1973]), .S(pc_current[2]), .Z(\Inst_Mem/n1304 ) );
  MUX \Inst_Mem/U1324  ( .A(inst_mem_in_wire[2005]), .B(inst_mem_in_wire[2037]), .S(pc_current[2]), .Z(\Inst_Mem/n1303 ) );
  MUX \Inst_Mem/U1323  ( .A(\Inst_Mem/n1302 ), .B(\Inst_Mem/n1271 ), .S(
        pc_current[7]), .Z(opcode[20]) );
  MUX \Inst_Mem/U1322  ( .A(\Inst_Mem/n1301 ), .B(\Inst_Mem/n1286 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1302 ) );
  MUX \Inst_Mem/U1321  ( .A(\Inst_Mem/n1300 ), .B(\Inst_Mem/n1293 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1301 ) );
  MUX \Inst_Mem/U1320  ( .A(\Inst_Mem/n1299 ), .B(\Inst_Mem/n1296 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1300 ) );
  MUX \Inst_Mem/U1319  ( .A(\Inst_Mem/n1298 ), .B(\Inst_Mem/n1297 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1299 ) );
  MUX \Inst_Mem/U1318  ( .A(inst_mem_in_wire[20]), .B(inst_mem_in_wire[52]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1298 ) );
  MUX \Inst_Mem/U1317  ( .A(inst_mem_in_wire[84]), .B(inst_mem_in_wire[116]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1297 ) );
  MUX \Inst_Mem/U1316  ( .A(\Inst_Mem/n1295 ), .B(\Inst_Mem/n1294 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1296 ) );
  MUX \Inst_Mem/U1315  ( .A(inst_mem_in_wire[148]), .B(inst_mem_in_wire[180]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1295 ) );
  MUX \Inst_Mem/U1314  ( .A(inst_mem_in_wire[212]), .B(inst_mem_in_wire[244]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1294 ) );
  MUX \Inst_Mem/U1313  ( .A(\Inst_Mem/n1292 ), .B(\Inst_Mem/n1289 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1293 ) );
  MUX \Inst_Mem/U1312  ( .A(\Inst_Mem/n1291 ), .B(\Inst_Mem/n1290 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1292 ) );
  MUX \Inst_Mem/U1311  ( .A(inst_mem_in_wire[276]), .B(inst_mem_in_wire[308]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1291 ) );
  MUX \Inst_Mem/U1310  ( .A(inst_mem_in_wire[340]), .B(inst_mem_in_wire[372]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1290 ) );
  MUX \Inst_Mem/U1309  ( .A(\Inst_Mem/n1288 ), .B(\Inst_Mem/n1287 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1289 ) );
  MUX \Inst_Mem/U1308  ( .A(inst_mem_in_wire[404]), .B(inst_mem_in_wire[436]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1288 ) );
  MUX \Inst_Mem/U1307  ( .A(inst_mem_in_wire[468]), .B(inst_mem_in_wire[500]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1287 ) );
  MUX \Inst_Mem/U1306  ( .A(\Inst_Mem/n1285 ), .B(\Inst_Mem/n1278 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1286 ) );
  MUX \Inst_Mem/U1305  ( .A(\Inst_Mem/n1284 ), .B(\Inst_Mem/n1281 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1285 ) );
  MUX \Inst_Mem/U1304  ( .A(\Inst_Mem/n1283 ), .B(\Inst_Mem/n1282 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1284 ) );
  MUX \Inst_Mem/U1303  ( .A(inst_mem_in_wire[532]), .B(inst_mem_in_wire[564]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1283 ) );
  MUX \Inst_Mem/U1302  ( .A(inst_mem_in_wire[596]), .B(inst_mem_in_wire[628]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1282 ) );
  MUX \Inst_Mem/U1301  ( .A(\Inst_Mem/n1280 ), .B(\Inst_Mem/n1279 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1281 ) );
  MUX \Inst_Mem/U1300  ( .A(inst_mem_in_wire[660]), .B(inst_mem_in_wire[692]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1280 ) );
  MUX \Inst_Mem/U1299  ( .A(inst_mem_in_wire[724]), .B(inst_mem_in_wire[756]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1279 ) );
  MUX \Inst_Mem/U1298  ( .A(\Inst_Mem/n1277 ), .B(\Inst_Mem/n1274 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1278 ) );
  MUX \Inst_Mem/U1297  ( .A(\Inst_Mem/n1276 ), .B(\Inst_Mem/n1275 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1277 ) );
  MUX \Inst_Mem/U1296  ( .A(inst_mem_in_wire[788]), .B(inst_mem_in_wire[820]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1276 ) );
  MUX \Inst_Mem/U1295  ( .A(inst_mem_in_wire[852]), .B(inst_mem_in_wire[884]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1275 ) );
  MUX \Inst_Mem/U1294  ( .A(\Inst_Mem/n1273 ), .B(\Inst_Mem/n1272 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1274 ) );
  MUX \Inst_Mem/U1293  ( .A(inst_mem_in_wire[916]), .B(inst_mem_in_wire[948]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1273 ) );
  MUX \Inst_Mem/U1292  ( .A(inst_mem_in_wire[980]), .B(inst_mem_in_wire[1012]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1272 ) );
  MUX \Inst_Mem/U1291  ( .A(\Inst_Mem/n1270 ), .B(\Inst_Mem/n1255 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1271 ) );
  MUX \Inst_Mem/U1290  ( .A(\Inst_Mem/n1269 ), .B(\Inst_Mem/n1262 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1270 ) );
  MUX \Inst_Mem/U1289  ( .A(\Inst_Mem/n1268 ), .B(\Inst_Mem/n1265 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1269 ) );
  MUX \Inst_Mem/U1288  ( .A(\Inst_Mem/n1267 ), .B(\Inst_Mem/n1266 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1268 ) );
  MUX \Inst_Mem/U1287  ( .A(inst_mem_in_wire[1044]), .B(inst_mem_in_wire[1076]), .S(pc_current[2]), .Z(\Inst_Mem/n1267 ) );
  MUX \Inst_Mem/U1286  ( .A(inst_mem_in_wire[1108]), .B(inst_mem_in_wire[1140]), .S(pc_current[2]), .Z(\Inst_Mem/n1266 ) );
  MUX \Inst_Mem/U1285  ( .A(\Inst_Mem/n1264 ), .B(\Inst_Mem/n1263 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1265 ) );
  MUX \Inst_Mem/U1284  ( .A(inst_mem_in_wire[1172]), .B(inst_mem_in_wire[1204]), .S(pc_current[2]), .Z(\Inst_Mem/n1264 ) );
  MUX \Inst_Mem/U1283  ( .A(inst_mem_in_wire[1236]), .B(inst_mem_in_wire[1268]), .S(pc_current[2]), .Z(\Inst_Mem/n1263 ) );
  MUX \Inst_Mem/U1282  ( .A(\Inst_Mem/n1261 ), .B(\Inst_Mem/n1258 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1262 ) );
  MUX \Inst_Mem/U1281  ( .A(\Inst_Mem/n1260 ), .B(\Inst_Mem/n1259 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1261 ) );
  MUX \Inst_Mem/U1280  ( .A(inst_mem_in_wire[1300]), .B(inst_mem_in_wire[1332]), .S(pc_current[2]), .Z(\Inst_Mem/n1260 ) );
  MUX \Inst_Mem/U1279  ( .A(inst_mem_in_wire[1364]), .B(inst_mem_in_wire[1396]), .S(pc_current[2]), .Z(\Inst_Mem/n1259 ) );
  MUX \Inst_Mem/U1278  ( .A(\Inst_Mem/n1257 ), .B(\Inst_Mem/n1256 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1258 ) );
  MUX \Inst_Mem/U1277  ( .A(inst_mem_in_wire[1428]), .B(inst_mem_in_wire[1460]), .S(pc_current[2]), .Z(\Inst_Mem/n1257 ) );
  MUX \Inst_Mem/U1276  ( .A(inst_mem_in_wire[1492]), .B(inst_mem_in_wire[1524]), .S(pc_current[2]), .Z(\Inst_Mem/n1256 ) );
  MUX \Inst_Mem/U1275  ( .A(\Inst_Mem/n1254 ), .B(\Inst_Mem/n1247 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1255 ) );
  MUX \Inst_Mem/U1274  ( .A(\Inst_Mem/n1253 ), .B(\Inst_Mem/n1250 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1254 ) );
  MUX \Inst_Mem/U1273  ( .A(\Inst_Mem/n1252 ), .B(\Inst_Mem/n1251 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1253 ) );
  MUX \Inst_Mem/U1272  ( .A(inst_mem_in_wire[1556]), .B(inst_mem_in_wire[1588]), .S(pc_current[2]), .Z(\Inst_Mem/n1252 ) );
  MUX \Inst_Mem/U1271  ( .A(inst_mem_in_wire[1620]), .B(inst_mem_in_wire[1652]), .S(pc_current[2]), .Z(\Inst_Mem/n1251 ) );
  MUX \Inst_Mem/U1270  ( .A(\Inst_Mem/n1249 ), .B(\Inst_Mem/n1248 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1250 ) );
  MUX \Inst_Mem/U1269  ( .A(inst_mem_in_wire[1684]), .B(inst_mem_in_wire[1716]), .S(pc_current[2]), .Z(\Inst_Mem/n1249 ) );
  MUX \Inst_Mem/U1268  ( .A(inst_mem_in_wire[1748]), .B(inst_mem_in_wire[1780]), .S(pc_current[2]), .Z(\Inst_Mem/n1248 ) );
  MUX \Inst_Mem/U1267  ( .A(\Inst_Mem/n1246 ), .B(\Inst_Mem/n1243 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1247 ) );
  MUX \Inst_Mem/U1266  ( .A(\Inst_Mem/n1245 ), .B(\Inst_Mem/n1244 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1246 ) );
  MUX \Inst_Mem/U1265  ( .A(inst_mem_in_wire[1812]), .B(inst_mem_in_wire[1844]), .S(pc_current[2]), .Z(\Inst_Mem/n1245 ) );
  MUX \Inst_Mem/U1264  ( .A(inst_mem_in_wire[1876]), .B(inst_mem_in_wire[1908]), .S(pc_current[2]), .Z(\Inst_Mem/n1244 ) );
  MUX \Inst_Mem/U1263  ( .A(\Inst_Mem/n1242 ), .B(\Inst_Mem/n1241 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1243 ) );
  MUX \Inst_Mem/U1262  ( .A(inst_mem_in_wire[1940]), .B(inst_mem_in_wire[1972]), .S(pc_current[2]), .Z(\Inst_Mem/n1242 ) );
  MUX \Inst_Mem/U1261  ( .A(inst_mem_in_wire[2004]), .B(inst_mem_in_wire[2036]), .S(pc_current[2]), .Z(\Inst_Mem/n1241 ) );
  MUX \Inst_Mem/U1260  ( .A(\Inst_Mem/n1240 ), .B(\Inst_Mem/n1209 ), .S(
        pc_current[7]), .Z(opcode[19]) );
  MUX \Inst_Mem/U1259  ( .A(\Inst_Mem/n1239 ), .B(\Inst_Mem/n1224 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1240 ) );
  MUX \Inst_Mem/U1258  ( .A(\Inst_Mem/n1238 ), .B(\Inst_Mem/n1231 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1239 ) );
  MUX \Inst_Mem/U1257  ( .A(\Inst_Mem/n1237 ), .B(\Inst_Mem/n1234 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1238 ) );
  MUX \Inst_Mem/U1256  ( .A(\Inst_Mem/n1236 ), .B(\Inst_Mem/n1235 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1237 ) );
  MUX \Inst_Mem/U1255  ( .A(inst_mem_in_wire[19]), .B(inst_mem_in_wire[51]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1236 ) );
  MUX \Inst_Mem/U1254  ( .A(inst_mem_in_wire[83]), .B(inst_mem_in_wire[115]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1235 ) );
  MUX \Inst_Mem/U1253  ( .A(\Inst_Mem/n1233 ), .B(\Inst_Mem/n1232 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1234 ) );
  MUX \Inst_Mem/U1252  ( .A(inst_mem_in_wire[147]), .B(inst_mem_in_wire[179]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1233 ) );
  MUX \Inst_Mem/U1251  ( .A(inst_mem_in_wire[211]), .B(inst_mem_in_wire[243]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1232 ) );
  MUX \Inst_Mem/U1250  ( .A(\Inst_Mem/n1230 ), .B(\Inst_Mem/n1227 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1231 ) );
  MUX \Inst_Mem/U1249  ( .A(\Inst_Mem/n1229 ), .B(\Inst_Mem/n1228 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1230 ) );
  MUX \Inst_Mem/U1248  ( .A(inst_mem_in_wire[275]), .B(inst_mem_in_wire[307]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1229 ) );
  MUX \Inst_Mem/U1247  ( .A(inst_mem_in_wire[339]), .B(inst_mem_in_wire[371]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1228 ) );
  MUX \Inst_Mem/U1246  ( .A(\Inst_Mem/n1226 ), .B(\Inst_Mem/n1225 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1227 ) );
  MUX \Inst_Mem/U1245  ( .A(inst_mem_in_wire[403]), .B(inst_mem_in_wire[435]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1226 ) );
  MUX \Inst_Mem/U1244  ( .A(inst_mem_in_wire[467]), .B(inst_mem_in_wire[499]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1225 ) );
  MUX \Inst_Mem/U1243  ( .A(\Inst_Mem/n1223 ), .B(\Inst_Mem/n1216 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1224 ) );
  MUX \Inst_Mem/U1242  ( .A(\Inst_Mem/n1222 ), .B(\Inst_Mem/n1219 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1223 ) );
  MUX \Inst_Mem/U1241  ( .A(\Inst_Mem/n1221 ), .B(\Inst_Mem/n1220 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1222 ) );
  MUX \Inst_Mem/U1240  ( .A(inst_mem_in_wire[531]), .B(inst_mem_in_wire[563]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1221 ) );
  MUX \Inst_Mem/U1239  ( .A(inst_mem_in_wire[595]), .B(inst_mem_in_wire[627]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1220 ) );
  MUX \Inst_Mem/U1238  ( .A(\Inst_Mem/n1218 ), .B(\Inst_Mem/n1217 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1219 ) );
  MUX \Inst_Mem/U1237  ( .A(inst_mem_in_wire[659]), .B(inst_mem_in_wire[691]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1218 ) );
  MUX \Inst_Mem/U1236  ( .A(inst_mem_in_wire[723]), .B(inst_mem_in_wire[755]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1217 ) );
  MUX \Inst_Mem/U1235  ( .A(\Inst_Mem/n1215 ), .B(\Inst_Mem/n1212 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1216 ) );
  MUX \Inst_Mem/U1234  ( .A(\Inst_Mem/n1214 ), .B(\Inst_Mem/n1213 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1215 ) );
  MUX \Inst_Mem/U1233  ( .A(inst_mem_in_wire[787]), .B(inst_mem_in_wire[819]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1214 ) );
  MUX \Inst_Mem/U1232  ( .A(inst_mem_in_wire[851]), .B(inst_mem_in_wire[883]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1213 ) );
  MUX \Inst_Mem/U1231  ( .A(\Inst_Mem/n1211 ), .B(\Inst_Mem/n1210 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1212 ) );
  MUX \Inst_Mem/U1230  ( .A(inst_mem_in_wire[915]), .B(inst_mem_in_wire[947]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1211 ) );
  MUX \Inst_Mem/U1229  ( .A(inst_mem_in_wire[979]), .B(inst_mem_in_wire[1011]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1210 ) );
  MUX \Inst_Mem/U1228  ( .A(\Inst_Mem/n1208 ), .B(\Inst_Mem/n1193 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1209 ) );
  MUX \Inst_Mem/U1227  ( .A(\Inst_Mem/n1207 ), .B(\Inst_Mem/n1200 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1208 ) );
  MUX \Inst_Mem/U1226  ( .A(\Inst_Mem/n1206 ), .B(\Inst_Mem/n1203 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1207 ) );
  MUX \Inst_Mem/U1225  ( .A(\Inst_Mem/n1205 ), .B(\Inst_Mem/n1204 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1206 ) );
  MUX \Inst_Mem/U1224  ( .A(inst_mem_in_wire[1043]), .B(inst_mem_in_wire[1075]), .S(pc_current[2]), .Z(\Inst_Mem/n1205 ) );
  MUX \Inst_Mem/U1223  ( .A(inst_mem_in_wire[1107]), .B(inst_mem_in_wire[1139]), .S(pc_current[2]), .Z(\Inst_Mem/n1204 ) );
  MUX \Inst_Mem/U1222  ( .A(\Inst_Mem/n1202 ), .B(\Inst_Mem/n1201 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1203 ) );
  MUX \Inst_Mem/U1221  ( .A(inst_mem_in_wire[1171]), .B(inst_mem_in_wire[1203]), .S(pc_current[2]), .Z(\Inst_Mem/n1202 ) );
  MUX \Inst_Mem/U1220  ( .A(inst_mem_in_wire[1235]), .B(inst_mem_in_wire[1267]), .S(pc_current[2]), .Z(\Inst_Mem/n1201 ) );
  MUX \Inst_Mem/U1219  ( .A(\Inst_Mem/n1199 ), .B(\Inst_Mem/n1196 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1200 ) );
  MUX \Inst_Mem/U1218  ( .A(\Inst_Mem/n1198 ), .B(\Inst_Mem/n1197 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1199 ) );
  MUX \Inst_Mem/U1217  ( .A(inst_mem_in_wire[1299]), .B(inst_mem_in_wire[1331]), .S(pc_current[2]), .Z(\Inst_Mem/n1198 ) );
  MUX \Inst_Mem/U1216  ( .A(inst_mem_in_wire[1363]), .B(inst_mem_in_wire[1395]), .S(pc_current[2]), .Z(\Inst_Mem/n1197 ) );
  MUX \Inst_Mem/U1215  ( .A(\Inst_Mem/n1195 ), .B(\Inst_Mem/n1194 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1196 ) );
  MUX \Inst_Mem/U1214  ( .A(inst_mem_in_wire[1427]), .B(inst_mem_in_wire[1459]), .S(pc_current[2]), .Z(\Inst_Mem/n1195 ) );
  MUX \Inst_Mem/U1213  ( .A(inst_mem_in_wire[1491]), .B(inst_mem_in_wire[1523]), .S(pc_current[2]), .Z(\Inst_Mem/n1194 ) );
  MUX \Inst_Mem/U1212  ( .A(\Inst_Mem/n1192 ), .B(\Inst_Mem/n1185 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1193 ) );
  MUX \Inst_Mem/U1211  ( .A(\Inst_Mem/n1191 ), .B(\Inst_Mem/n1188 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1192 ) );
  MUX \Inst_Mem/U1210  ( .A(\Inst_Mem/n1190 ), .B(\Inst_Mem/n1189 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1191 ) );
  MUX \Inst_Mem/U1209  ( .A(inst_mem_in_wire[1555]), .B(inst_mem_in_wire[1587]), .S(pc_current[2]), .Z(\Inst_Mem/n1190 ) );
  MUX \Inst_Mem/U1208  ( .A(inst_mem_in_wire[1619]), .B(inst_mem_in_wire[1651]), .S(pc_current[2]), .Z(\Inst_Mem/n1189 ) );
  MUX \Inst_Mem/U1207  ( .A(\Inst_Mem/n1187 ), .B(\Inst_Mem/n1186 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1188 ) );
  MUX \Inst_Mem/U1206  ( .A(inst_mem_in_wire[1683]), .B(inst_mem_in_wire[1715]), .S(pc_current[2]), .Z(\Inst_Mem/n1187 ) );
  MUX \Inst_Mem/U1205  ( .A(inst_mem_in_wire[1747]), .B(inst_mem_in_wire[1779]), .S(pc_current[2]), .Z(\Inst_Mem/n1186 ) );
  MUX \Inst_Mem/U1204  ( .A(\Inst_Mem/n1184 ), .B(\Inst_Mem/n1181 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1185 ) );
  MUX \Inst_Mem/U1203  ( .A(\Inst_Mem/n1183 ), .B(\Inst_Mem/n1182 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1184 ) );
  MUX \Inst_Mem/U1202  ( .A(inst_mem_in_wire[1811]), .B(inst_mem_in_wire[1843]), .S(pc_current[2]), .Z(\Inst_Mem/n1183 ) );
  MUX \Inst_Mem/U1201  ( .A(inst_mem_in_wire[1875]), .B(inst_mem_in_wire[1907]), .S(pc_current[2]), .Z(\Inst_Mem/n1182 ) );
  MUX \Inst_Mem/U1200  ( .A(\Inst_Mem/n1180 ), .B(\Inst_Mem/n1179 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1181 ) );
  MUX \Inst_Mem/U1199  ( .A(inst_mem_in_wire[1939]), .B(inst_mem_in_wire[1971]), .S(pc_current[2]), .Z(\Inst_Mem/n1180 ) );
  MUX \Inst_Mem/U1198  ( .A(inst_mem_in_wire[2003]), .B(inst_mem_in_wire[2035]), .S(pc_current[2]), .Z(\Inst_Mem/n1179 ) );
  MUX \Inst_Mem/U1197  ( .A(\Inst_Mem/n1178 ), .B(\Inst_Mem/n1147 ), .S(
        pc_current[7]), .Z(opcode[18]) );
  MUX \Inst_Mem/U1196  ( .A(\Inst_Mem/n1177 ), .B(\Inst_Mem/n1162 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1178 ) );
  MUX \Inst_Mem/U1195  ( .A(\Inst_Mem/n1176 ), .B(\Inst_Mem/n1169 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1177 ) );
  MUX \Inst_Mem/U1194  ( .A(\Inst_Mem/n1175 ), .B(\Inst_Mem/n1172 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1176 ) );
  MUX \Inst_Mem/U1193  ( .A(\Inst_Mem/n1174 ), .B(\Inst_Mem/n1173 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1175 ) );
  MUX \Inst_Mem/U1192  ( .A(inst_mem_in_wire[18]), .B(inst_mem_in_wire[50]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1174 ) );
  MUX \Inst_Mem/U1191  ( .A(inst_mem_in_wire[82]), .B(inst_mem_in_wire[114]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1173 ) );
  MUX \Inst_Mem/U1190  ( .A(\Inst_Mem/n1171 ), .B(\Inst_Mem/n1170 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1172 ) );
  MUX \Inst_Mem/U1189  ( .A(inst_mem_in_wire[146]), .B(inst_mem_in_wire[178]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1171 ) );
  MUX \Inst_Mem/U1188  ( .A(inst_mem_in_wire[210]), .B(inst_mem_in_wire[242]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1170 ) );
  MUX \Inst_Mem/U1187  ( .A(\Inst_Mem/n1168 ), .B(\Inst_Mem/n1165 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1169 ) );
  MUX \Inst_Mem/U1186  ( .A(\Inst_Mem/n1167 ), .B(\Inst_Mem/n1166 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1168 ) );
  MUX \Inst_Mem/U1185  ( .A(inst_mem_in_wire[274]), .B(inst_mem_in_wire[306]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1167 ) );
  MUX \Inst_Mem/U1184  ( .A(inst_mem_in_wire[338]), .B(inst_mem_in_wire[370]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1166 ) );
  MUX \Inst_Mem/U1183  ( .A(\Inst_Mem/n1164 ), .B(\Inst_Mem/n1163 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1165 ) );
  MUX \Inst_Mem/U1182  ( .A(inst_mem_in_wire[402]), .B(inst_mem_in_wire[434]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1164 ) );
  MUX \Inst_Mem/U1181  ( .A(inst_mem_in_wire[466]), .B(inst_mem_in_wire[498]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1163 ) );
  MUX \Inst_Mem/U1180  ( .A(\Inst_Mem/n1161 ), .B(\Inst_Mem/n1154 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1162 ) );
  MUX \Inst_Mem/U1179  ( .A(\Inst_Mem/n1160 ), .B(\Inst_Mem/n1157 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1161 ) );
  MUX \Inst_Mem/U1178  ( .A(\Inst_Mem/n1159 ), .B(\Inst_Mem/n1158 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1160 ) );
  MUX \Inst_Mem/U1177  ( .A(inst_mem_in_wire[530]), .B(inst_mem_in_wire[562]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1159 ) );
  MUX \Inst_Mem/U1176  ( .A(inst_mem_in_wire[594]), .B(inst_mem_in_wire[626]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1158 ) );
  MUX \Inst_Mem/U1175  ( .A(\Inst_Mem/n1156 ), .B(\Inst_Mem/n1155 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1157 ) );
  MUX \Inst_Mem/U1174  ( .A(inst_mem_in_wire[658]), .B(inst_mem_in_wire[690]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1156 ) );
  MUX \Inst_Mem/U1173  ( .A(inst_mem_in_wire[722]), .B(inst_mem_in_wire[754]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1155 ) );
  MUX \Inst_Mem/U1172  ( .A(\Inst_Mem/n1153 ), .B(\Inst_Mem/n1150 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1154 ) );
  MUX \Inst_Mem/U1171  ( .A(\Inst_Mem/n1152 ), .B(\Inst_Mem/n1151 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1153 ) );
  MUX \Inst_Mem/U1170  ( .A(inst_mem_in_wire[786]), .B(inst_mem_in_wire[818]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1152 ) );
  MUX \Inst_Mem/U1169  ( .A(inst_mem_in_wire[850]), .B(inst_mem_in_wire[882]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1151 ) );
  MUX \Inst_Mem/U1168  ( .A(\Inst_Mem/n1149 ), .B(\Inst_Mem/n1148 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1150 ) );
  MUX \Inst_Mem/U1167  ( .A(inst_mem_in_wire[914]), .B(inst_mem_in_wire[946]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1149 ) );
  MUX \Inst_Mem/U1166  ( .A(inst_mem_in_wire[978]), .B(inst_mem_in_wire[1010]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1148 ) );
  MUX \Inst_Mem/U1165  ( .A(\Inst_Mem/n1146 ), .B(\Inst_Mem/n1131 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1147 ) );
  MUX \Inst_Mem/U1164  ( .A(\Inst_Mem/n1145 ), .B(\Inst_Mem/n1138 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1146 ) );
  MUX \Inst_Mem/U1163  ( .A(\Inst_Mem/n1144 ), .B(\Inst_Mem/n1141 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1145 ) );
  MUX \Inst_Mem/U1162  ( .A(\Inst_Mem/n1143 ), .B(\Inst_Mem/n1142 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1144 ) );
  MUX \Inst_Mem/U1161  ( .A(inst_mem_in_wire[1042]), .B(inst_mem_in_wire[1074]), .S(pc_current[2]), .Z(\Inst_Mem/n1143 ) );
  MUX \Inst_Mem/U1160  ( .A(inst_mem_in_wire[1106]), .B(inst_mem_in_wire[1138]), .S(pc_current[2]), .Z(\Inst_Mem/n1142 ) );
  MUX \Inst_Mem/U1159  ( .A(\Inst_Mem/n1140 ), .B(\Inst_Mem/n1139 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1141 ) );
  MUX \Inst_Mem/U1158  ( .A(inst_mem_in_wire[1170]), .B(inst_mem_in_wire[1202]), .S(pc_current[2]), .Z(\Inst_Mem/n1140 ) );
  MUX \Inst_Mem/U1157  ( .A(inst_mem_in_wire[1234]), .B(inst_mem_in_wire[1266]), .S(pc_current[2]), .Z(\Inst_Mem/n1139 ) );
  MUX \Inst_Mem/U1156  ( .A(\Inst_Mem/n1137 ), .B(\Inst_Mem/n1134 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1138 ) );
  MUX \Inst_Mem/U1155  ( .A(\Inst_Mem/n1136 ), .B(\Inst_Mem/n1135 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1137 ) );
  MUX \Inst_Mem/U1154  ( .A(inst_mem_in_wire[1298]), .B(inst_mem_in_wire[1330]), .S(pc_current[2]), .Z(\Inst_Mem/n1136 ) );
  MUX \Inst_Mem/U1153  ( .A(inst_mem_in_wire[1362]), .B(inst_mem_in_wire[1394]), .S(pc_current[2]), .Z(\Inst_Mem/n1135 ) );
  MUX \Inst_Mem/U1152  ( .A(\Inst_Mem/n1133 ), .B(\Inst_Mem/n1132 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1134 ) );
  MUX \Inst_Mem/U1151  ( .A(inst_mem_in_wire[1426]), .B(inst_mem_in_wire[1458]), .S(pc_current[2]), .Z(\Inst_Mem/n1133 ) );
  MUX \Inst_Mem/U1150  ( .A(inst_mem_in_wire[1490]), .B(inst_mem_in_wire[1522]), .S(pc_current[2]), .Z(\Inst_Mem/n1132 ) );
  MUX \Inst_Mem/U1149  ( .A(\Inst_Mem/n1130 ), .B(\Inst_Mem/n1123 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1131 ) );
  MUX \Inst_Mem/U1148  ( .A(\Inst_Mem/n1129 ), .B(\Inst_Mem/n1126 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1130 ) );
  MUX \Inst_Mem/U1147  ( .A(\Inst_Mem/n1128 ), .B(\Inst_Mem/n1127 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1129 ) );
  MUX \Inst_Mem/U1146  ( .A(inst_mem_in_wire[1554]), .B(inst_mem_in_wire[1586]), .S(pc_current[2]), .Z(\Inst_Mem/n1128 ) );
  MUX \Inst_Mem/U1145  ( .A(inst_mem_in_wire[1618]), .B(inst_mem_in_wire[1650]), .S(pc_current[2]), .Z(\Inst_Mem/n1127 ) );
  MUX \Inst_Mem/U1144  ( .A(\Inst_Mem/n1125 ), .B(\Inst_Mem/n1124 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1126 ) );
  MUX \Inst_Mem/U1143  ( .A(inst_mem_in_wire[1682]), .B(inst_mem_in_wire[1714]), .S(pc_current[2]), .Z(\Inst_Mem/n1125 ) );
  MUX \Inst_Mem/U1142  ( .A(inst_mem_in_wire[1746]), .B(inst_mem_in_wire[1778]), .S(pc_current[2]), .Z(\Inst_Mem/n1124 ) );
  MUX \Inst_Mem/U1141  ( .A(\Inst_Mem/n1122 ), .B(\Inst_Mem/n1119 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1123 ) );
  MUX \Inst_Mem/U1140  ( .A(\Inst_Mem/n1121 ), .B(\Inst_Mem/n1120 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1122 ) );
  MUX \Inst_Mem/U1139  ( .A(inst_mem_in_wire[1810]), .B(inst_mem_in_wire[1842]), .S(pc_current[2]), .Z(\Inst_Mem/n1121 ) );
  MUX \Inst_Mem/U1138  ( .A(inst_mem_in_wire[1874]), .B(inst_mem_in_wire[1906]), .S(pc_current[2]), .Z(\Inst_Mem/n1120 ) );
  MUX \Inst_Mem/U1137  ( .A(\Inst_Mem/n1118 ), .B(\Inst_Mem/n1117 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1119 ) );
  MUX \Inst_Mem/U1136  ( .A(inst_mem_in_wire[1938]), .B(inst_mem_in_wire[1970]), .S(pc_current[2]), .Z(\Inst_Mem/n1118 ) );
  MUX \Inst_Mem/U1135  ( .A(inst_mem_in_wire[2002]), .B(inst_mem_in_wire[2034]), .S(pc_current[2]), .Z(\Inst_Mem/n1117 ) );
  MUX \Inst_Mem/U1134  ( .A(\Inst_Mem/n1116 ), .B(\Inst_Mem/n1085 ), .S(
        pc_current[7]), .Z(opcode[17]) );
  MUX \Inst_Mem/U1133  ( .A(\Inst_Mem/n1115 ), .B(\Inst_Mem/n1100 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1116 ) );
  MUX \Inst_Mem/U1132  ( .A(\Inst_Mem/n1114 ), .B(\Inst_Mem/n1107 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1115 ) );
  MUX \Inst_Mem/U1131  ( .A(\Inst_Mem/n1113 ), .B(\Inst_Mem/n1110 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1114 ) );
  MUX \Inst_Mem/U1130  ( .A(\Inst_Mem/n1112 ), .B(\Inst_Mem/n1111 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1113 ) );
  MUX \Inst_Mem/U1129  ( .A(inst_mem_in_wire[17]), .B(inst_mem_in_wire[49]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1112 ) );
  MUX \Inst_Mem/U1128  ( .A(inst_mem_in_wire[81]), .B(inst_mem_in_wire[113]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1111 ) );
  MUX \Inst_Mem/U1127  ( .A(\Inst_Mem/n1109 ), .B(\Inst_Mem/n1108 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1110 ) );
  MUX \Inst_Mem/U1126  ( .A(inst_mem_in_wire[145]), .B(inst_mem_in_wire[177]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1109 ) );
  MUX \Inst_Mem/U1125  ( .A(inst_mem_in_wire[209]), .B(inst_mem_in_wire[241]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1108 ) );
  MUX \Inst_Mem/U1124  ( .A(\Inst_Mem/n1106 ), .B(\Inst_Mem/n1103 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1107 ) );
  MUX \Inst_Mem/U1123  ( .A(\Inst_Mem/n1105 ), .B(\Inst_Mem/n1104 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1106 ) );
  MUX \Inst_Mem/U1122  ( .A(inst_mem_in_wire[273]), .B(inst_mem_in_wire[305]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1105 ) );
  MUX \Inst_Mem/U1121  ( .A(inst_mem_in_wire[337]), .B(inst_mem_in_wire[369]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1104 ) );
  MUX \Inst_Mem/U1120  ( .A(\Inst_Mem/n1102 ), .B(\Inst_Mem/n1101 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1103 ) );
  MUX \Inst_Mem/U1119  ( .A(inst_mem_in_wire[401]), .B(inst_mem_in_wire[433]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1102 ) );
  MUX \Inst_Mem/U1118  ( .A(inst_mem_in_wire[465]), .B(inst_mem_in_wire[497]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1101 ) );
  MUX \Inst_Mem/U1117  ( .A(\Inst_Mem/n1099 ), .B(\Inst_Mem/n1092 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1100 ) );
  MUX \Inst_Mem/U1116  ( .A(\Inst_Mem/n1098 ), .B(\Inst_Mem/n1095 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1099 ) );
  MUX \Inst_Mem/U1115  ( .A(\Inst_Mem/n1097 ), .B(\Inst_Mem/n1096 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1098 ) );
  MUX \Inst_Mem/U1114  ( .A(inst_mem_in_wire[529]), .B(inst_mem_in_wire[561]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1097 ) );
  MUX \Inst_Mem/U1113  ( .A(inst_mem_in_wire[593]), .B(inst_mem_in_wire[625]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1096 ) );
  MUX \Inst_Mem/U1112  ( .A(\Inst_Mem/n1094 ), .B(\Inst_Mem/n1093 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1095 ) );
  MUX \Inst_Mem/U1111  ( .A(inst_mem_in_wire[657]), .B(inst_mem_in_wire[689]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1094 ) );
  MUX \Inst_Mem/U1110  ( .A(inst_mem_in_wire[721]), .B(inst_mem_in_wire[753]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1093 ) );
  MUX \Inst_Mem/U1109  ( .A(\Inst_Mem/n1091 ), .B(\Inst_Mem/n1088 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1092 ) );
  MUX \Inst_Mem/U1108  ( .A(\Inst_Mem/n1090 ), .B(\Inst_Mem/n1089 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1091 ) );
  MUX \Inst_Mem/U1107  ( .A(inst_mem_in_wire[785]), .B(inst_mem_in_wire[817]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1090 ) );
  MUX \Inst_Mem/U1106  ( .A(inst_mem_in_wire[849]), .B(inst_mem_in_wire[881]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1089 ) );
  MUX \Inst_Mem/U1105  ( .A(\Inst_Mem/n1087 ), .B(\Inst_Mem/n1086 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1088 ) );
  MUX \Inst_Mem/U1104  ( .A(inst_mem_in_wire[913]), .B(inst_mem_in_wire[945]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1087 ) );
  MUX \Inst_Mem/U1103  ( .A(inst_mem_in_wire[977]), .B(inst_mem_in_wire[1009]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1086 ) );
  MUX \Inst_Mem/U1102  ( .A(\Inst_Mem/n1084 ), .B(\Inst_Mem/n1069 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1085 ) );
  MUX \Inst_Mem/U1101  ( .A(\Inst_Mem/n1083 ), .B(\Inst_Mem/n1076 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1084 ) );
  MUX \Inst_Mem/U1100  ( .A(\Inst_Mem/n1082 ), .B(\Inst_Mem/n1079 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1083 ) );
  MUX \Inst_Mem/U1099  ( .A(\Inst_Mem/n1081 ), .B(\Inst_Mem/n1080 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1082 ) );
  MUX \Inst_Mem/U1098  ( .A(inst_mem_in_wire[1041]), .B(inst_mem_in_wire[1073]), .S(pc_current[2]), .Z(\Inst_Mem/n1081 ) );
  MUX \Inst_Mem/U1097  ( .A(inst_mem_in_wire[1105]), .B(inst_mem_in_wire[1137]), .S(pc_current[2]), .Z(\Inst_Mem/n1080 ) );
  MUX \Inst_Mem/U1096  ( .A(\Inst_Mem/n1078 ), .B(\Inst_Mem/n1077 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1079 ) );
  MUX \Inst_Mem/U1095  ( .A(inst_mem_in_wire[1169]), .B(inst_mem_in_wire[1201]), .S(pc_current[2]), .Z(\Inst_Mem/n1078 ) );
  MUX \Inst_Mem/U1094  ( .A(inst_mem_in_wire[1233]), .B(inst_mem_in_wire[1265]), .S(pc_current[2]), .Z(\Inst_Mem/n1077 ) );
  MUX \Inst_Mem/U1093  ( .A(\Inst_Mem/n1075 ), .B(\Inst_Mem/n1072 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1076 ) );
  MUX \Inst_Mem/U1092  ( .A(\Inst_Mem/n1074 ), .B(\Inst_Mem/n1073 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1075 ) );
  MUX \Inst_Mem/U1091  ( .A(inst_mem_in_wire[1297]), .B(inst_mem_in_wire[1329]), .S(pc_current[2]), .Z(\Inst_Mem/n1074 ) );
  MUX \Inst_Mem/U1090  ( .A(inst_mem_in_wire[1361]), .B(inst_mem_in_wire[1393]), .S(pc_current[2]), .Z(\Inst_Mem/n1073 ) );
  MUX \Inst_Mem/U1089  ( .A(\Inst_Mem/n1071 ), .B(\Inst_Mem/n1070 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1072 ) );
  MUX \Inst_Mem/U1088  ( .A(inst_mem_in_wire[1425]), .B(inst_mem_in_wire[1457]), .S(pc_current[2]), .Z(\Inst_Mem/n1071 ) );
  MUX \Inst_Mem/U1087  ( .A(inst_mem_in_wire[1489]), .B(inst_mem_in_wire[1521]), .S(pc_current[2]), .Z(\Inst_Mem/n1070 ) );
  MUX \Inst_Mem/U1086  ( .A(\Inst_Mem/n1068 ), .B(\Inst_Mem/n1061 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1069 ) );
  MUX \Inst_Mem/U1085  ( .A(\Inst_Mem/n1067 ), .B(\Inst_Mem/n1064 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1068 ) );
  MUX \Inst_Mem/U1084  ( .A(\Inst_Mem/n1066 ), .B(\Inst_Mem/n1065 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1067 ) );
  MUX \Inst_Mem/U1083  ( .A(inst_mem_in_wire[1553]), .B(inst_mem_in_wire[1585]), .S(pc_current[2]), .Z(\Inst_Mem/n1066 ) );
  MUX \Inst_Mem/U1082  ( .A(inst_mem_in_wire[1617]), .B(inst_mem_in_wire[1649]), .S(pc_current[2]), .Z(\Inst_Mem/n1065 ) );
  MUX \Inst_Mem/U1081  ( .A(\Inst_Mem/n1063 ), .B(\Inst_Mem/n1062 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1064 ) );
  MUX \Inst_Mem/U1080  ( .A(inst_mem_in_wire[1681]), .B(inst_mem_in_wire[1713]), .S(pc_current[2]), .Z(\Inst_Mem/n1063 ) );
  MUX \Inst_Mem/U1079  ( .A(inst_mem_in_wire[1745]), .B(inst_mem_in_wire[1777]), .S(pc_current[2]), .Z(\Inst_Mem/n1062 ) );
  MUX \Inst_Mem/U1078  ( .A(\Inst_Mem/n1060 ), .B(\Inst_Mem/n1057 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1061 ) );
  MUX \Inst_Mem/U1077  ( .A(\Inst_Mem/n1059 ), .B(\Inst_Mem/n1058 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1060 ) );
  MUX \Inst_Mem/U1076  ( .A(inst_mem_in_wire[1809]), .B(inst_mem_in_wire[1841]), .S(pc_current[2]), .Z(\Inst_Mem/n1059 ) );
  MUX \Inst_Mem/U1075  ( .A(inst_mem_in_wire[1873]), .B(inst_mem_in_wire[1905]), .S(pc_current[2]), .Z(\Inst_Mem/n1058 ) );
  MUX \Inst_Mem/U1074  ( .A(\Inst_Mem/n1056 ), .B(\Inst_Mem/n1055 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1057 ) );
  MUX \Inst_Mem/U1073  ( .A(inst_mem_in_wire[1937]), .B(inst_mem_in_wire[1969]), .S(pc_current[2]), .Z(\Inst_Mem/n1056 ) );
  MUX \Inst_Mem/U1072  ( .A(inst_mem_in_wire[2001]), .B(inst_mem_in_wire[2033]), .S(pc_current[2]), .Z(\Inst_Mem/n1055 ) );
  MUX \Inst_Mem/U1071  ( .A(\Inst_Mem/n1054 ), .B(\Inst_Mem/n1023 ), .S(
        pc_current[7]), .Z(opcode[16]) );
  MUX \Inst_Mem/U1070  ( .A(\Inst_Mem/n1053 ), .B(\Inst_Mem/n1038 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1054 ) );
  MUX \Inst_Mem/U1069  ( .A(\Inst_Mem/n1052 ), .B(\Inst_Mem/n1045 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1053 ) );
  MUX \Inst_Mem/U1068  ( .A(\Inst_Mem/n1051 ), .B(\Inst_Mem/n1048 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1052 ) );
  MUX \Inst_Mem/U1067  ( .A(\Inst_Mem/n1050 ), .B(\Inst_Mem/n1049 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1051 ) );
  MUX \Inst_Mem/U1066  ( .A(inst_mem_in_wire[16]), .B(inst_mem_in_wire[48]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1050 ) );
  MUX \Inst_Mem/U1065  ( .A(inst_mem_in_wire[80]), .B(inst_mem_in_wire[112]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1049 ) );
  MUX \Inst_Mem/U1064  ( .A(\Inst_Mem/n1047 ), .B(\Inst_Mem/n1046 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1048 ) );
  MUX \Inst_Mem/U1063  ( .A(inst_mem_in_wire[144]), .B(inst_mem_in_wire[176]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1047 ) );
  MUX \Inst_Mem/U1062  ( .A(inst_mem_in_wire[208]), .B(inst_mem_in_wire[240]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1046 ) );
  MUX \Inst_Mem/U1061  ( .A(\Inst_Mem/n1044 ), .B(\Inst_Mem/n1041 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1045 ) );
  MUX \Inst_Mem/U1060  ( .A(\Inst_Mem/n1043 ), .B(\Inst_Mem/n1042 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1044 ) );
  MUX \Inst_Mem/U1059  ( .A(inst_mem_in_wire[272]), .B(inst_mem_in_wire[304]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1043 ) );
  MUX \Inst_Mem/U1058  ( .A(inst_mem_in_wire[336]), .B(inst_mem_in_wire[368]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1042 ) );
  MUX \Inst_Mem/U1057  ( .A(\Inst_Mem/n1040 ), .B(\Inst_Mem/n1039 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1041 ) );
  MUX \Inst_Mem/U1056  ( .A(inst_mem_in_wire[400]), .B(inst_mem_in_wire[432]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1040 ) );
  MUX \Inst_Mem/U1055  ( .A(inst_mem_in_wire[464]), .B(inst_mem_in_wire[496]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1039 ) );
  MUX \Inst_Mem/U1054  ( .A(\Inst_Mem/n1037 ), .B(\Inst_Mem/n1030 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1038 ) );
  MUX \Inst_Mem/U1053  ( .A(\Inst_Mem/n1036 ), .B(\Inst_Mem/n1033 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1037 ) );
  MUX \Inst_Mem/U1052  ( .A(\Inst_Mem/n1035 ), .B(\Inst_Mem/n1034 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1036 ) );
  MUX \Inst_Mem/U1051  ( .A(inst_mem_in_wire[528]), .B(inst_mem_in_wire[560]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1035 ) );
  MUX \Inst_Mem/U1050  ( .A(inst_mem_in_wire[592]), .B(inst_mem_in_wire[624]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1034 ) );
  MUX \Inst_Mem/U1049  ( .A(\Inst_Mem/n1032 ), .B(\Inst_Mem/n1031 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1033 ) );
  MUX \Inst_Mem/U1048  ( .A(inst_mem_in_wire[656]), .B(inst_mem_in_wire[688]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1032 ) );
  MUX \Inst_Mem/U1047  ( .A(inst_mem_in_wire[720]), .B(inst_mem_in_wire[752]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1031 ) );
  MUX \Inst_Mem/U1046  ( .A(\Inst_Mem/n1029 ), .B(\Inst_Mem/n1026 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1030 ) );
  MUX \Inst_Mem/U1045  ( .A(\Inst_Mem/n1028 ), .B(\Inst_Mem/n1027 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1029 ) );
  MUX \Inst_Mem/U1044  ( .A(inst_mem_in_wire[784]), .B(inst_mem_in_wire[816]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1028 ) );
  MUX \Inst_Mem/U1043  ( .A(inst_mem_in_wire[848]), .B(inst_mem_in_wire[880]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1027 ) );
  MUX \Inst_Mem/U1042  ( .A(\Inst_Mem/n1025 ), .B(\Inst_Mem/n1024 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1026 ) );
  MUX \Inst_Mem/U1041  ( .A(inst_mem_in_wire[912]), .B(inst_mem_in_wire[944]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1025 ) );
  MUX \Inst_Mem/U1040  ( .A(inst_mem_in_wire[976]), .B(inst_mem_in_wire[1008]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1024 ) );
  MUX \Inst_Mem/U1039  ( .A(\Inst_Mem/n1022 ), .B(\Inst_Mem/n1007 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n1023 ) );
  MUX \Inst_Mem/U1038  ( .A(\Inst_Mem/n1021 ), .B(\Inst_Mem/n1014 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1022 ) );
  MUX \Inst_Mem/U1037  ( .A(\Inst_Mem/n1020 ), .B(\Inst_Mem/n1017 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1021 ) );
  MUX \Inst_Mem/U1036  ( .A(\Inst_Mem/n1019 ), .B(\Inst_Mem/n1018 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1020 ) );
  MUX \Inst_Mem/U1035  ( .A(inst_mem_in_wire[1040]), .B(inst_mem_in_wire[1072]), .S(pc_current[2]), .Z(\Inst_Mem/n1019 ) );
  MUX \Inst_Mem/U1034  ( .A(inst_mem_in_wire[1104]), .B(inst_mem_in_wire[1136]), .S(pc_current[2]), .Z(\Inst_Mem/n1018 ) );
  MUX \Inst_Mem/U1033  ( .A(\Inst_Mem/n1016 ), .B(\Inst_Mem/n1015 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1017 ) );
  MUX \Inst_Mem/U1032  ( .A(inst_mem_in_wire[1168]), .B(inst_mem_in_wire[1200]), .S(pc_current[2]), .Z(\Inst_Mem/n1016 ) );
  MUX \Inst_Mem/U1031  ( .A(inst_mem_in_wire[1232]), .B(inst_mem_in_wire[1264]), .S(pc_current[2]), .Z(\Inst_Mem/n1015 ) );
  MUX \Inst_Mem/U1030  ( .A(\Inst_Mem/n1013 ), .B(\Inst_Mem/n1010 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1014 ) );
  MUX \Inst_Mem/U1029  ( .A(\Inst_Mem/n1012 ), .B(\Inst_Mem/n1011 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1013 ) );
  MUX \Inst_Mem/U1028  ( .A(inst_mem_in_wire[1296]), .B(inst_mem_in_wire[1328]), .S(pc_current[2]), .Z(\Inst_Mem/n1012 ) );
  MUX \Inst_Mem/U1027  ( .A(inst_mem_in_wire[1360]), .B(inst_mem_in_wire[1392]), .S(pc_current[2]), .Z(\Inst_Mem/n1011 ) );
  MUX \Inst_Mem/U1026  ( .A(\Inst_Mem/n1009 ), .B(\Inst_Mem/n1008 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1010 ) );
  MUX \Inst_Mem/U1025  ( .A(inst_mem_in_wire[1424]), .B(inst_mem_in_wire[1456]), .S(pc_current[2]), .Z(\Inst_Mem/n1009 ) );
  MUX \Inst_Mem/U1024  ( .A(inst_mem_in_wire[1488]), .B(inst_mem_in_wire[1520]), .S(pc_current[2]), .Z(\Inst_Mem/n1008 ) );
  MUX \Inst_Mem/U1023  ( .A(\Inst_Mem/n1006 ), .B(\Inst_Mem/n999 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n1007 ) );
  MUX \Inst_Mem/U1022  ( .A(\Inst_Mem/n1005 ), .B(\Inst_Mem/n1002 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n1006 ) );
  MUX \Inst_Mem/U1021  ( .A(\Inst_Mem/n1004 ), .B(\Inst_Mem/n1003 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1005 ) );
  MUX \Inst_Mem/U1020  ( .A(inst_mem_in_wire[1552]), .B(inst_mem_in_wire[1584]), .S(pc_current[2]), .Z(\Inst_Mem/n1004 ) );
  MUX \Inst_Mem/U1019  ( .A(inst_mem_in_wire[1616]), .B(inst_mem_in_wire[1648]), .S(pc_current[2]), .Z(\Inst_Mem/n1003 ) );
  MUX \Inst_Mem/U1018  ( .A(\Inst_Mem/n1001 ), .B(\Inst_Mem/n1000 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n1002 ) );
  MUX \Inst_Mem/U1017  ( .A(inst_mem_in_wire[1680]), .B(inst_mem_in_wire[1712]), .S(pc_current[2]), .Z(\Inst_Mem/n1001 ) );
  MUX \Inst_Mem/U1016  ( .A(inst_mem_in_wire[1744]), .B(inst_mem_in_wire[1776]), .S(pc_current[2]), .Z(\Inst_Mem/n1000 ) );
  MUX \Inst_Mem/U1015  ( .A(\Inst_Mem/n998 ), .B(\Inst_Mem/n995 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n999 ) );
  MUX \Inst_Mem/U1014  ( .A(\Inst_Mem/n997 ), .B(\Inst_Mem/n996 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n998 ) );
  MUX \Inst_Mem/U1013  ( .A(inst_mem_in_wire[1808]), .B(inst_mem_in_wire[1840]), .S(pc_current[2]), .Z(\Inst_Mem/n997 ) );
  MUX \Inst_Mem/U1012  ( .A(inst_mem_in_wire[1872]), .B(inst_mem_in_wire[1904]), .S(pc_current[2]), .Z(\Inst_Mem/n996 ) );
  MUX \Inst_Mem/U1011  ( .A(\Inst_Mem/n994 ), .B(\Inst_Mem/n993 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n995 ) );
  MUX \Inst_Mem/U1010  ( .A(inst_mem_in_wire[1936]), .B(inst_mem_in_wire[1968]), .S(pc_current[2]), .Z(\Inst_Mem/n994 ) );
  MUX \Inst_Mem/U1009  ( .A(inst_mem_in_wire[2000]), .B(inst_mem_in_wire[2032]), .S(pc_current[2]), .Z(\Inst_Mem/n993 ) );
  MUX \Inst_Mem/U1008  ( .A(\Inst_Mem/n992 ), .B(\Inst_Mem/n961 ), .S(
        pc_current[7]), .Z(imm[15]) );
  MUX \Inst_Mem/U1007  ( .A(\Inst_Mem/n991 ), .B(\Inst_Mem/n976 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n992 ) );
  MUX \Inst_Mem/U1006  ( .A(\Inst_Mem/n990 ), .B(\Inst_Mem/n983 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n991 ) );
  MUX \Inst_Mem/U1005  ( .A(\Inst_Mem/n989 ), .B(\Inst_Mem/n986 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n990 ) );
  MUX \Inst_Mem/U1004  ( .A(\Inst_Mem/n988 ), .B(\Inst_Mem/n987 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n989 ) );
  MUX \Inst_Mem/U1003  ( .A(inst_mem_in_wire[15]), .B(inst_mem_in_wire[47]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n988 ) );
  MUX \Inst_Mem/U1002  ( .A(inst_mem_in_wire[79]), .B(inst_mem_in_wire[111]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n987 ) );
  MUX \Inst_Mem/U1001  ( .A(\Inst_Mem/n985 ), .B(\Inst_Mem/n984 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n986 ) );
  MUX \Inst_Mem/U1000  ( .A(inst_mem_in_wire[143]), .B(inst_mem_in_wire[175]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n985 ) );
  MUX \Inst_Mem/U999  ( .A(inst_mem_in_wire[207]), .B(inst_mem_in_wire[239]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n984 ) );
  MUX \Inst_Mem/U998  ( .A(\Inst_Mem/n982 ), .B(\Inst_Mem/n979 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n983 ) );
  MUX \Inst_Mem/U997  ( .A(\Inst_Mem/n981 ), .B(\Inst_Mem/n980 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n982 ) );
  MUX \Inst_Mem/U996  ( .A(inst_mem_in_wire[271]), .B(inst_mem_in_wire[303]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n981 ) );
  MUX \Inst_Mem/U995  ( .A(inst_mem_in_wire[335]), .B(inst_mem_in_wire[367]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n980 ) );
  MUX \Inst_Mem/U994  ( .A(\Inst_Mem/n978 ), .B(\Inst_Mem/n977 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n979 ) );
  MUX \Inst_Mem/U993  ( .A(inst_mem_in_wire[399]), .B(inst_mem_in_wire[431]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n978 ) );
  MUX \Inst_Mem/U992  ( .A(inst_mem_in_wire[463]), .B(inst_mem_in_wire[495]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n977 ) );
  MUX \Inst_Mem/U991  ( .A(\Inst_Mem/n975 ), .B(\Inst_Mem/n968 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n976 ) );
  MUX \Inst_Mem/U990  ( .A(\Inst_Mem/n974 ), .B(\Inst_Mem/n971 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n975 ) );
  MUX \Inst_Mem/U989  ( .A(\Inst_Mem/n973 ), .B(\Inst_Mem/n972 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n974 ) );
  MUX \Inst_Mem/U988  ( .A(inst_mem_in_wire[527]), .B(inst_mem_in_wire[559]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n973 ) );
  MUX \Inst_Mem/U987  ( .A(inst_mem_in_wire[591]), .B(inst_mem_in_wire[623]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n972 ) );
  MUX \Inst_Mem/U986  ( .A(\Inst_Mem/n970 ), .B(\Inst_Mem/n969 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n971 ) );
  MUX \Inst_Mem/U985  ( .A(inst_mem_in_wire[655]), .B(inst_mem_in_wire[687]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n970 ) );
  MUX \Inst_Mem/U984  ( .A(inst_mem_in_wire[719]), .B(inst_mem_in_wire[751]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n969 ) );
  MUX \Inst_Mem/U983  ( .A(\Inst_Mem/n967 ), .B(\Inst_Mem/n964 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n968 ) );
  MUX \Inst_Mem/U982  ( .A(\Inst_Mem/n966 ), .B(\Inst_Mem/n965 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n967 ) );
  MUX \Inst_Mem/U981  ( .A(inst_mem_in_wire[783]), .B(inst_mem_in_wire[815]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n966 ) );
  MUX \Inst_Mem/U980  ( .A(inst_mem_in_wire[847]), .B(inst_mem_in_wire[879]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n965 ) );
  MUX \Inst_Mem/U979  ( .A(\Inst_Mem/n963 ), .B(\Inst_Mem/n962 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n964 ) );
  MUX \Inst_Mem/U978  ( .A(inst_mem_in_wire[911]), .B(inst_mem_in_wire[943]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n963 ) );
  MUX \Inst_Mem/U977  ( .A(inst_mem_in_wire[975]), .B(inst_mem_in_wire[1007]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n962 ) );
  MUX \Inst_Mem/U976  ( .A(\Inst_Mem/n960 ), .B(\Inst_Mem/n945 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n961 ) );
  MUX \Inst_Mem/U975  ( .A(\Inst_Mem/n959 ), .B(\Inst_Mem/n952 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n960 ) );
  MUX \Inst_Mem/U974  ( .A(\Inst_Mem/n958 ), .B(\Inst_Mem/n955 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n959 ) );
  MUX \Inst_Mem/U973  ( .A(\Inst_Mem/n957 ), .B(\Inst_Mem/n956 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n958 ) );
  MUX \Inst_Mem/U972  ( .A(inst_mem_in_wire[1039]), .B(inst_mem_in_wire[1071]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n957 ) );
  MUX \Inst_Mem/U971  ( .A(inst_mem_in_wire[1103]), .B(inst_mem_in_wire[1135]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n956 ) );
  MUX \Inst_Mem/U970  ( .A(\Inst_Mem/n954 ), .B(\Inst_Mem/n953 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n955 ) );
  MUX \Inst_Mem/U969  ( .A(inst_mem_in_wire[1167]), .B(inst_mem_in_wire[1199]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n954 ) );
  MUX \Inst_Mem/U968  ( .A(inst_mem_in_wire[1231]), .B(inst_mem_in_wire[1263]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n953 ) );
  MUX \Inst_Mem/U967  ( .A(\Inst_Mem/n951 ), .B(\Inst_Mem/n948 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n952 ) );
  MUX \Inst_Mem/U966  ( .A(\Inst_Mem/n950 ), .B(\Inst_Mem/n949 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n951 ) );
  MUX \Inst_Mem/U965  ( .A(inst_mem_in_wire[1295]), .B(inst_mem_in_wire[1327]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n950 ) );
  MUX \Inst_Mem/U964  ( .A(inst_mem_in_wire[1359]), .B(inst_mem_in_wire[1391]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n949 ) );
  MUX \Inst_Mem/U963  ( .A(\Inst_Mem/n947 ), .B(\Inst_Mem/n946 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n948 ) );
  MUX \Inst_Mem/U962  ( .A(inst_mem_in_wire[1423]), .B(inst_mem_in_wire[1455]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n947 ) );
  MUX \Inst_Mem/U961  ( .A(inst_mem_in_wire[1487]), .B(inst_mem_in_wire[1519]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n946 ) );
  MUX \Inst_Mem/U960  ( .A(\Inst_Mem/n944 ), .B(\Inst_Mem/n937 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n945 ) );
  MUX \Inst_Mem/U959  ( .A(\Inst_Mem/n943 ), .B(\Inst_Mem/n940 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n944 ) );
  MUX \Inst_Mem/U958  ( .A(\Inst_Mem/n942 ), .B(\Inst_Mem/n941 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n943 ) );
  MUX \Inst_Mem/U957  ( .A(inst_mem_in_wire[1551]), .B(inst_mem_in_wire[1583]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n942 ) );
  MUX \Inst_Mem/U956  ( .A(inst_mem_in_wire[1615]), .B(inst_mem_in_wire[1647]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n941 ) );
  MUX \Inst_Mem/U955  ( .A(\Inst_Mem/n939 ), .B(\Inst_Mem/n938 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n940 ) );
  MUX \Inst_Mem/U954  ( .A(inst_mem_in_wire[1679]), .B(inst_mem_in_wire[1711]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n939 ) );
  MUX \Inst_Mem/U953  ( .A(inst_mem_in_wire[1743]), .B(inst_mem_in_wire[1775]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n938 ) );
  MUX \Inst_Mem/U952  ( .A(\Inst_Mem/n936 ), .B(\Inst_Mem/n933 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n937 ) );
  MUX \Inst_Mem/U951  ( .A(\Inst_Mem/n935 ), .B(\Inst_Mem/n934 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n936 ) );
  MUX \Inst_Mem/U950  ( .A(inst_mem_in_wire[1807]), .B(inst_mem_in_wire[1839]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n935 ) );
  MUX \Inst_Mem/U949  ( .A(inst_mem_in_wire[1871]), .B(inst_mem_in_wire[1903]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n934 ) );
  MUX \Inst_Mem/U948  ( .A(\Inst_Mem/n932 ), .B(\Inst_Mem/n931 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n933 ) );
  MUX \Inst_Mem/U947  ( .A(inst_mem_in_wire[1935]), .B(inst_mem_in_wire[1967]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n932 ) );
  MUX \Inst_Mem/U946  ( .A(inst_mem_in_wire[1999]), .B(inst_mem_in_wire[2031]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n931 ) );
  MUX \Inst_Mem/U945  ( .A(\Inst_Mem/n930 ), .B(\Inst_Mem/n899 ), .S(
        pc_current[7]), .Z(imm[14]) );
  MUX \Inst_Mem/U944  ( .A(\Inst_Mem/n929 ), .B(\Inst_Mem/n914 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n930 ) );
  MUX \Inst_Mem/U943  ( .A(\Inst_Mem/n928 ), .B(\Inst_Mem/n921 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n929 ) );
  MUX \Inst_Mem/U942  ( .A(\Inst_Mem/n927 ), .B(\Inst_Mem/n924 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n928 ) );
  MUX \Inst_Mem/U941  ( .A(\Inst_Mem/n926 ), .B(\Inst_Mem/n925 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n927 ) );
  MUX \Inst_Mem/U940  ( .A(inst_mem_in_wire[14]), .B(inst_mem_in_wire[46]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n926 ) );
  MUX \Inst_Mem/U939  ( .A(inst_mem_in_wire[78]), .B(inst_mem_in_wire[110]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n925 ) );
  MUX \Inst_Mem/U938  ( .A(\Inst_Mem/n923 ), .B(\Inst_Mem/n922 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n924 ) );
  MUX \Inst_Mem/U937  ( .A(inst_mem_in_wire[142]), .B(inst_mem_in_wire[174]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n923 ) );
  MUX \Inst_Mem/U936  ( .A(inst_mem_in_wire[206]), .B(inst_mem_in_wire[238]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n922 ) );
  MUX \Inst_Mem/U935  ( .A(\Inst_Mem/n920 ), .B(\Inst_Mem/n917 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n921 ) );
  MUX \Inst_Mem/U934  ( .A(\Inst_Mem/n919 ), .B(\Inst_Mem/n918 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n920 ) );
  MUX \Inst_Mem/U933  ( .A(inst_mem_in_wire[270]), .B(inst_mem_in_wire[302]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n919 ) );
  MUX \Inst_Mem/U932  ( .A(inst_mem_in_wire[334]), .B(inst_mem_in_wire[366]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n918 ) );
  MUX \Inst_Mem/U931  ( .A(\Inst_Mem/n916 ), .B(\Inst_Mem/n915 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n917 ) );
  MUX \Inst_Mem/U930  ( .A(inst_mem_in_wire[398]), .B(inst_mem_in_wire[430]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n916 ) );
  MUX \Inst_Mem/U929  ( .A(inst_mem_in_wire[462]), .B(inst_mem_in_wire[494]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n915 ) );
  MUX \Inst_Mem/U928  ( .A(\Inst_Mem/n913 ), .B(\Inst_Mem/n906 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n914 ) );
  MUX \Inst_Mem/U927  ( .A(\Inst_Mem/n912 ), .B(\Inst_Mem/n909 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n913 ) );
  MUX \Inst_Mem/U926  ( .A(\Inst_Mem/n911 ), .B(\Inst_Mem/n910 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n912 ) );
  MUX \Inst_Mem/U925  ( .A(inst_mem_in_wire[526]), .B(inst_mem_in_wire[558]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n911 ) );
  MUX \Inst_Mem/U924  ( .A(inst_mem_in_wire[590]), .B(inst_mem_in_wire[622]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n910 ) );
  MUX \Inst_Mem/U923  ( .A(\Inst_Mem/n908 ), .B(\Inst_Mem/n907 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n909 ) );
  MUX \Inst_Mem/U922  ( .A(inst_mem_in_wire[654]), .B(inst_mem_in_wire[686]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n908 ) );
  MUX \Inst_Mem/U921  ( .A(inst_mem_in_wire[718]), .B(inst_mem_in_wire[750]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n907 ) );
  MUX \Inst_Mem/U920  ( .A(\Inst_Mem/n905 ), .B(\Inst_Mem/n902 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n906 ) );
  MUX \Inst_Mem/U919  ( .A(\Inst_Mem/n904 ), .B(\Inst_Mem/n903 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n905 ) );
  MUX \Inst_Mem/U918  ( .A(inst_mem_in_wire[782]), .B(inst_mem_in_wire[814]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n904 ) );
  MUX \Inst_Mem/U917  ( .A(inst_mem_in_wire[846]), .B(inst_mem_in_wire[878]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n903 ) );
  MUX \Inst_Mem/U916  ( .A(\Inst_Mem/n901 ), .B(\Inst_Mem/n900 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n902 ) );
  MUX \Inst_Mem/U915  ( .A(inst_mem_in_wire[910]), .B(inst_mem_in_wire[942]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n901 ) );
  MUX \Inst_Mem/U914  ( .A(inst_mem_in_wire[974]), .B(inst_mem_in_wire[1006]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n900 ) );
  MUX \Inst_Mem/U913  ( .A(\Inst_Mem/n898 ), .B(\Inst_Mem/n883 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n899 ) );
  MUX \Inst_Mem/U912  ( .A(\Inst_Mem/n897 ), .B(\Inst_Mem/n890 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n898 ) );
  MUX \Inst_Mem/U911  ( .A(\Inst_Mem/n896 ), .B(\Inst_Mem/n893 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n897 ) );
  MUX \Inst_Mem/U910  ( .A(\Inst_Mem/n895 ), .B(\Inst_Mem/n894 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n896 ) );
  MUX \Inst_Mem/U909  ( .A(inst_mem_in_wire[1038]), .B(inst_mem_in_wire[1070]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n895 ) );
  MUX \Inst_Mem/U908  ( .A(inst_mem_in_wire[1102]), .B(inst_mem_in_wire[1134]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n894 ) );
  MUX \Inst_Mem/U907  ( .A(\Inst_Mem/n892 ), .B(\Inst_Mem/n891 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n893 ) );
  MUX \Inst_Mem/U906  ( .A(inst_mem_in_wire[1166]), .B(inst_mem_in_wire[1198]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n892 ) );
  MUX \Inst_Mem/U905  ( .A(inst_mem_in_wire[1230]), .B(inst_mem_in_wire[1262]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n891 ) );
  MUX \Inst_Mem/U904  ( .A(\Inst_Mem/n889 ), .B(\Inst_Mem/n886 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n890 ) );
  MUX \Inst_Mem/U903  ( .A(\Inst_Mem/n888 ), .B(\Inst_Mem/n887 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n889 ) );
  MUX \Inst_Mem/U902  ( .A(inst_mem_in_wire[1294]), .B(inst_mem_in_wire[1326]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n888 ) );
  MUX \Inst_Mem/U901  ( .A(inst_mem_in_wire[1358]), .B(inst_mem_in_wire[1390]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n887 ) );
  MUX \Inst_Mem/U900  ( .A(\Inst_Mem/n885 ), .B(\Inst_Mem/n884 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n886 ) );
  MUX \Inst_Mem/U899  ( .A(inst_mem_in_wire[1422]), .B(inst_mem_in_wire[1454]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n885 ) );
  MUX \Inst_Mem/U898  ( .A(inst_mem_in_wire[1486]), .B(inst_mem_in_wire[1518]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n884 ) );
  MUX \Inst_Mem/U897  ( .A(\Inst_Mem/n882 ), .B(\Inst_Mem/n875 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n883 ) );
  MUX \Inst_Mem/U896  ( .A(\Inst_Mem/n881 ), .B(\Inst_Mem/n878 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n882 ) );
  MUX \Inst_Mem/U895  ( .A(\Inst_Mem/n880 ), .B(\Inst_Mem/n879 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n881 ) );
  MUX \Inst_Mem/U894  ( .A(inst_mem_in_wire[1550]), .B(inst_mem_in_wire[1582]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n880 ) );
  MUX \Inst_Mem/U893  ( .A(inst_mem_in_wire[1614]), .B(inst_mem_in_wire[1646]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n879 ) );
  MUX \Inst_Mem/U892  ( .A(\Inst_Mem/n877 ), .B(\Inst_Mem/n876 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n878 ) );
  MUX \Inst_Mem/U891  ( .A(inst_mem_in_wire[1678]), .B(inst_mem_in_wire[1710]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n877 ) );
  MUX \Inst_Mem/U890  ( .A(inst_mem_in_wire[1742]), .B(inst_mem_in_wire[1774]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n876 ) );
  MUX \Inst_Mem/U889  ( .A(\Inst_Mem/n874 ), .B(\Inst_Mem/n871 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n875 ) );
  MUX \Inst_Mem/U888  ( .A(\Inst_Mem/n873 ), .B(\Inst_Mem/n872 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n874 ) );
  MUX \Inst_Mem/U887  ( .A(inst_mem_in_wire[1806]), .B(inst_mem_in_wire[1838]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n873 ) );
  MUX \Inst_Mem/U886  ( .A(inst_mem_in_wire[1870]), .B(inst_mem_in_wire[1902]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n872 ) );
  MUX \Inst_Mem/U885  ( .A(\Inst_Mem/n870 ), .B(\Inst_Mem/n869 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n871 ) );
  MUX \Inst_Mem/U884  ( .A(inst_mem_in_wire[1934]), .B(inst_mem_in_wire[1966]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n870 ) );
  MUX \Inst_Mem/U883  ( .A(inst_mem_in_wire[1998]), .B(inst_mem_in_wire[2030]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n869 ) );
  MUX \Inst_Mem/U882  ( .A(\Inst_Mem/n868 ), .B(\Inst_Mem/n837 ), .S(
        pc_current[7]), .Z(imm[13]) );
  MUX \Inst_Mem/U881  ( .A(\Inst_Mem/n867 ), .B(\Inst_Mem/n852 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n868 ) );
  MUX \Inst_Mem/U880  ( .A(\Inst_Mem/n866 ), .B(\Inst_Mem/n859 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n867 ) );
  MUX \Inst_Mem/U879  ( .A(\Inst_Mem/n865 ), .B(\Inst_Mem/n862 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n866 ) );
  MUX \Inst_Mem/U878  ( .A(\Inst_Mem/n864 ), .B(\Inst_Mem/n863 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n865 ) );
  MUX \Inst_Mem/U877  ( .A(inst_mem_in_wire[13]), .B(inst_mem_in_wire[45]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n864 ) );
  MUX \Inst_Mem/U876  ( .A(inst_mem_in_wire[77]), .B(inst_mem_in_wire[109]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n863 ) );
  MUX \Inst_Mem/U875  ( .A(\Inst_Mem/n861 ), .B(\Inst_Mem/n860 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n862 ) );
  MUX \Inst_Mem/U874  ( .A(inst_mem_in_wire[141]), .B(inst_mem_in_wire[173]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n861 ) );
  MUX \Inst_Mem/U873  ( .A(inst_mem_in_wire[205]), .B(inst_mem_in_wire[237]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n860 ) );
  MUX \Inst_Mem/U872  ( .A(\Inst_Mem/n858 ), .B(\Inst_Mem/n855 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n859 ) );
  MUX \Inst_Mem/U871  ( .A(\Inst_Mem/n857 ), .B(\Inst_Mem/n856 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n858 ) );
  MUX \Inst_Mem/U870  ( .A(inst_mem_in_wire[269]), .B(inst_mem_in_wire[301]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n857 ) );
  MUX \Inst_Mem/U869  ( .A(inst_mem_in_wire[333]), .B(inst_mem_in_wire[365]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n856 ) );
  MUX \Inst_Mem/U868  ( .A(\Inst_Mem/n854 ), .B(\Inst_Mem/n853 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n855 ) );
  MUX \Inst_Mem/U867  ( .A(inst_mem_in_wire[397]), .B(inst_mem_in_wire[429]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n854 ) );
  MUX \Inst_Mem/U866  ( .A(inst_mem_in_wire[461]), .B(inst_mem_in_wire[493]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n853 ) );
  MUX \Inst_Mem/U865  ( .A(\Inst_Mem/n851 ), .B(\Inst_Mem/n844 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n852 ) );
  MUX \Inst_Mem/U864  ( .A(\Inst_Mem/n850 ), .B(\Inst_Mem/n847 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n851 ) );
  MUX \Inst_Mem/U863  ( .A(\Inst_Mem/n849 ), .B(\Inst_Mem/n848 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n850 ) );
  MUX \Inst_Mem/U862  ( .A(inst_mem_in_wire[525]), .B(inst_mem_in_wire[557]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n849 ) );
  MUX \Inst_Mem/U861  ( .A(inst_mem_in_wire[589]), .B(inst_mem_in_wire[621]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n848 ) );
  MUX \Inst_Mem/U860  ( .A(\Inst_Mem/n846 ), .B(\Inst_Mem/n845 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n847 ) );
  MUX \Inst_Mem/U859  ( .A(inst_mem_in_wire[653]), .B(inst_mem_in_wire[685]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n846 ) );
  MUX \Inst_Mem/U858  ( .A(inst_mem_in_wire[717]), .B(inst_mem_in_wire[749]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n845 ) );
  MUX \Inst_Mem/U857  ( .A(\Inst_Mem/n843 ), .B(\Inst_Mem/n840 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n844 ) );
  MUX \Inst_Mem/U856  ( .A(\Inst_Mem/n842 ), .B(\Inst_Mem/n841 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n843 ) );
  MUX \Inst_Mem/U855  ( .A(inst_mem_in_wire[781]), .B(inst_mem_in_wire[813]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n842 ) );
  MUX \Inst_Mem/U854  ( .A(inst_mem_in_wire[845]), .B(inst_mem_in_wire[877]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n841 ) );
  MUX \Inst_Mem/U853  ( .A(\Inst_Mem/n839 ), .B(\Inst_Mem/n838 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n840 ) );
  MUX \Inst_Mem/U852  ( .A(inst_mem_in_wire[909]), .B(inst_mem_in_wire[941]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n839 ) );
  MUX \Inst_Mem/U851  ( .A(inst_mem_in_wire[973]), .B(inst_mem_in_wire[1005]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n838 ) );
  MUX \Inst_Mem/U850  ( .A(\Inst_Mem/n836 ), .B(\Inst_Mem/n821 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n837 ) );
  MUX \Inst_Mem/U849  ( .A(\Inst_Mem/n835 ), .B(\Inst_Mem/n828 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n836 ) );
  MUX \Inst_Mem/U848  ( .A(\Inst_Mem/n834 ), .B(\Inst_Mem/n831 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n835 ) );
  MUX \Inst_Mem/U847  ( .A(\Inst_Mem/n833 ), .B(\Inst_Mem/n832 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n834 ) );
  MUX \Inst_Mem/U846  ( .A(inst_mem_in_wire[1037]), .B(inst_mem_in_wire[1069]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n833 ) );
  MUX \Inst_Mem/U845  ( .A(inst_mem_in_wire[1101]), .B(inst_mem_in_wire[1133]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n832 ) );
  MUX \Inst_Mem/U844  ( .A(\Inst_Mem/n830 ), .B(\Inst_Mem/n829 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n831 ) );
  MUX \Inst_Mem/U843  ( .A(inst_mem_in_wire[1165]), .B(inst_mem_in_wire[1197]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n830 ) );
  MUX \Inst_Mem/U842  ( .A(inst_mem_in_wire[1229]), .B(inst_mem_in_wire[1261]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n829 ) );
  MUX \Inst_Mem/U841  ( .A(\Inst_Mem/n827 ), .B(\Inst_Mem/n824 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n828 ) );
  MUX \Inst_Mem/U840  ( .A(\Inst_Mem/n826 ), .B(\Inst_Mem/n825 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n827 ) );
  MUX \Inst_Mem/U839  ( .A(inst_mem_in_wire[1293]), .B(inst_mem_in_wire[1325]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n826 ) );
  MUX \Inst_Mem/U838  ( .A(inst_mem_in_wire[1357]), .B(inst_mem_in_wire[1389]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n825 ) );
  MUX \Inst_Mem/U837  ( .A(\Inst_Mem/n823 ), .B(\Inst_Mem/n822 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n824 ) );
  MUX \Inst_Mem/U836  ( .A(inst_mem_in_wire[1421]), .B(inst_mem_in_wire[1453]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n823 ) );
  MUX \Inst_Mem/U835  ( .A(inst_mem_in_wire[1485]), .B(inst_mem_in_wire[1517]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n822 ) );
  MUX \Inst_Mem/U834  ( .A(\Inst_Mem/n820 ), .B(\Inst_Mem/n813 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n821 ) );
  MUX \Inst_Mem/U833  ( .A(\Inst_Mem/n819 ), .B(\Inst_Mem/n816 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n820 ) );
  MUX \Inst_Mem/U832  ( .A(\Inst_Mem/n818 ), .B(\Inst_Mem/n817 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n819 ) );
  MUX \Inst_Mem/U831  ( .A(inst_mem_in_wire[1549]), .B(inst_mem_in_wire[1581]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n818 ) );
  MUX \Inst_Mem/U830  ( .A(inst_mem_in_wire[1613]), .B(inst_mem_in_wire[1645]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n817 ) );
  MUX \Inst_Mem/U829  ( .A(\Inst_Mem/n815 ), .B(\Inst_Mem/n814 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n816 ) );
  MUX \Inst_Mem/U828  ( .A(inst_mem_in_wire[1677]), .B(inst_mem_in_wire[1709]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n815 ) );
  MUX \Inst_Mem/U827  ( .A(inst_mem_in_wire[1741]), .B(inst_mem_in_wire[1773]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n814 ) );
  MUX \Inst_Mem/U826  ( .A(\Inst_Mem/n812 ), .B(\Inst_Mem/n809 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n813 ) );
  MUX \Inst_Mem/U825  ( .A(\Inst_Mem/n811 ), .B(\Inst_Mem/n810 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n812 ) );
  MUX \Inst_Mem/U824  ( .A(inst_mem_in_wire[1805]), .B(inst_mem_in_wire[1837]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n811 ) );
  MUX \Inst_Mem/U823  ( .A(inst_mem_in_wire[1869]), .B(inst_mem_in_wire[1901]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n810 ) );
  MUX \Inst_Mem/U822  ( .A(\Inst_Mem/n808 ), .B(\Inst_Mem/n807 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n809 ) );
  MUX \Inst_Mem/U821  ( .A(inst_mem_in_wire[1933]), .B(inst_mem_in_wire[1965]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n808 ) );
  MUX \Inst_Mem/U820  ( .A(inst_mem_in_wire[1997]), .B(inst_mem_in_wire[2029]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n807 ) );
  MUX \Inst_Mem/U819  ( .A(\Inst_Mem/n806 ), .B(\Inst_Mem/n775 ), .S(
        pc_current[7]), .Z(imm[12]) );
  MUX \Inst_Mem/U818  ( .A(\Inst_Mem/n805 ), .B(\Inst_Mem/n790 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n806 ) );
  MUX \Inst_Mem/U817  ( .A(\Inst_Mem/n804 ), .B(\Inst_Mem/n797 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n805 ) );
  MUX \Inst_Mem/U816  ( .A(\Inst_Mem/n803 ), .B(\Inst_Mem/n800 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n804 ) );
  MUX \Inst_Mem/U815  ( .A(\Inst_Mem/n802 ), .B(\Inst_Mem/n801 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n803 ) );
  MUX \Inst_Mem/U814  ( .A(inst_mem_in_wire[12]), .B(inst_mem_in_wire[44]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n802 ) );
  MUX \Inst_Mem/U813  ( .A(inst_mem_in_wire[76]), .B(inst_mem_in_wire[108]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n801 ) );
  MUX \Inst_Mem/U812  ( .A(\Inst_Mem/n799 ), .B(\Inst_Mem/n798 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n800 ) );
  MUX \Inst_Mem/U811  ( .A(inst_mem_in_wire[140]), .B(inst_mem_in_wire[172]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n799 ) );
  MUX \Inst_Mem/U810  ( .A(inst_mem_in_wire[204]), .B(inst_mem_in_wire[236]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n798 ) );
  MUX \Inst_Mem/U809  ( .A(\Inst_Mem/n796 ), .B(\Inst_Mem/n793 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n797 ) );
  MUX \Inst_Mem/U808  ( .A(\Inst_Mem/n795 ), .B(\Inst_Mem/n794 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n796 ) );
  MUX \Inst_Mem/U807  ( .A(inst_mem_in_wire[268]), .B(inst_mem_in_wire[300]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n795 ) );
  MUX \Inst_Mem/U806  ( .A(inst_mem_in_wire[332]), .B(inst_mem_in_wire[364]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n794 ) );
  MUX \Inst_Mem/U805  ( .A(\Inst_Mem/n792 ), .B(\Inst_Mem/n791 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n793 ) );
  MUX \Inst_Mem/U804  ( .A(inst_mem_in_wire[396]), .B(inst_mem_in_wire[428]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n792 ) );
  MUX \Inst_Mem/U803  ( .A(inst_mem_in_wire[460]), .B(inst_mem_in_wire[492]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n791 ) );
  MUX \Inst_Mem/U802  ( .A(\Inst_Mem/n789 ), .B(\Inst_Mem/n782 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n790 ) );
  MUX \Inst_Mem/U801  ( .A(\Inst_Mem/n788 ), .B(\Inst_Mem/n785 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n789 ) );
  MUX \Inst_Mem/U800  ( .A(\Inst_Mem/n787 ), .B(\Inst_Mem/n786 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n788 ) );
  MUX \Inst_Mem/U799  ( .A(inst_mem_in_wire[524]), .B(inst_mem_in_wire[556]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n787 ) );
  MUX \Inst_Mem/U798  ( .A(inst_mem_in_wire[588]), .B(inst_mem_in_wire[620]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n786 ) );
  MUX \Inst_Mem/U797  ( .A(\Inst_Mem/n784 ), .B(\Inst_Mem/n783 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n785 ) );
  MUX \Inst_Mem/U796  ( .A(inst_mem_in_wire[652]), .B(inst_mem_in_wire[684]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n784 ) );
  MUX \Inst_Mem/U795  ( .A(inst_mem_in_wire[716]), .B(inst_mem_in_wire[748]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n783 ) );
  MUX \Inst_Mem/U794  ( .A(\Inst_Mem/n781 ), .B(\Inst_Mem/n778 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n782 ) );
  MUX \Inst_Mem/U793  ( .A(\Inst_Mem/n780 ), .B(\Inst_Mem/n779 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n781 ) );
  MUX \Inst_Mem/U792  ( .A(inst_mem_in_wire[780]), .B(inst_mem_in_wire[812]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n780 ) );
  MUX \Inst_Mem/U791  ( .A(inst_mem_in_wire[844]), .B(inst_mem_in_wire[876]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n779 ) );
  MUX \Inst_Mem/U790  ( .A(\Inst_Mem/n777 ), .B(\Inst_Mem/n776 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n778 ) );
  MUX \Inst_Mem/U789  ( .A(inst_mem_in_wire[908]), .B(inst_mem_in_wire[940]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n777 ) );
  MUX \Inst_Mem/U788  ( .A(inst_mem_in_wire[972]), .B(inst_mem_in_wire[1004]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n776 ) );
  MUX \Inst_Mem/U787  ( .A(\Inst_Mem/n774 ), .B(\Inst_Mem/n759 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n775 ) );
  MUX \Inst_Mem/U786  ( .A(\Inst_Mem/n773 ), .B(\Inst_Mem/n766 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n774 ) );
  MUX \Inst_Mem/U785  ( .A(\Inst_Mem/n772 ), .B(\Inst_Mem/n769 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n773 ) );
  MUX \Inst_Mem/U784  ( .A(\Inst_Mem/n771 ), .B(\Inst_Mem/n770 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n772 ) );
  MUX \Inst_Mem/U783  ( .A(inst_mem_in_wire[1036]), .B(inst_mem_in_wire[1068]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n771 ) );
  MUX \Inst_Mem/U782  ( .A(inst_mem_in_wire[1100]), .B(inst_mem_in_wire[1132]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n770 ) );
  MUX \Inst_Mem/U781  ( .A(\Inst_Mem/n768 ), .B(\Inst_Mem/n767 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n769 ) );
  MUX \Inst_Mem/U780  ( .A(inst_mem_in_wire[1164]), .B(inst_mem_in_wire[1196]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n768 ) );
  MUX \Inst_Mem/U779  ( .A(inst_mem_in_wire[1228]), .B(inst_mem_in_wire[1260]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n767 ) );
  MUX \Inst_Mem/U778  ( .A(\Inst_Mem/n765 ), .B(\Inst_Mem/n762 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n766 ) );
  MUX \Inst_Mem/U777  ( .A(\Inst_Mem/n764 ), .B(\Inst_Mem/n763 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n765 ) );
  MUX \Inst_Mem/U776  ( .A(inst_mem_in_wire[1292]), .B(inst_mem_in_wire[1324]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n764 ) );
  MUX \Inst_Mem/U775  ( .A(inst_mem_in_wire[1356]), .B(inst_mem_in_wire[1388]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n763 ) );
  MUX \Inst_Mem/U774  ( .A(\Inst_Mem/n761 ), .B(\Inst_Mem/n760 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n762 ) );
  MUX \Inst_Mem/U773  ( .A(inst_mem_in_wire[1420]), .B(inst_mem_in_wire[1452]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n761 ) );
  MUX \Inst_Mem/U772  ( .A(inst_mem_in_wire[1484]), .B(inst_mem_in_wire[1516]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n760 ) );
  MUX \Inst_Mem/U771  ( .A(\Inst_Mem/n758 ), .B(\Inst_Mem/n751 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n759 ) );
  MUX \Inst_Mem/U770  ( .A(\Inst_Mem/n757 ), .B(\Inst_Mem/n754 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n758 ) );
  MUX \Inst_Mem/U769  ( .A(\Inst_Mem/n756 ), .B(\Inst_Mem/n755 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n757 ) );
  MUX \Inst_Mem/U768  ( .A(inst_mem_in_wire[1548]), .B(inst_mem_in_wire[1580]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n756 ) );
  MUX \Inst_Mem/U767  ( .A(inst_mem_in_wire[1612]), .B(inst_mem_in_wire[1644]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n755 ) );
  MUX \Inst_Mem/U766  ( .A(\Inst_Mem/n753 ), .B(\Inst_Mem/n752 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n754 ) );
  MUX \Inst_Mem/U765  ( .A(inst_mem_in_wire[1676]), .B(inst_mem_in_wire[1708]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n753 ) );
  MUX \Inst_Mem/U764  ( .A(inst_mem_in_wire[1740]), .B(inst_mem_in_wire[1772]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n752 ) );
  MUX \Inst_Mem/U763  ( .A(\Inst_Mem/n750 ), .B(\Inst_Mem/n747 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n751 ) );
  MUX \Inst_Mem/U762  ( .A(\Inst_Mem/n749 ), .B(\Inst_Mem/n748 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n750 ) );
  MUX \Inst_Mem/U761  ( .A(inst_mem_in_wire[1804]), .B(inst_mem_in_wire[1836]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n749 ) );
  MUX \Inst_Mem/U760  ( .A(inst_mem_in_wire[1868]), .B(inst_mem_in_wire[1900]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n748 ) );
  MUX \Inst_Mem/U759  ( .A(\Inst_Mem/n746 ), .B(\Inst_Mem/n745 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n747 ) );
  MUX \Inst_Mem/U758  ( .A(inst_mem_in_wire[1932]), .B(inst_mem_in_wire[1964]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n746 ) );
  MUX \Inst_Mem/U757  ( .A(inst_mem_in_wire[1996]), .B(inst_mem_in_wire[2028]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n745 ) );
  MUX \Inst_Mem/U756  ( .A(\Inst_Mem/n744 ), .B(\Inst_Mem/n713 ), .S(
        pc_current[7]), .Z(imm[11]) );
  MUX \Inst_Mem/U755  ( .A(\Inst_Mem/n743 ), .B(\Inst_Mem/n728 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n744 ) );
  MUX \Inst_Mem/U754  ( .A(\Inst_Mem/n742 ), .B(\Inst_Mem/n735 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n743 ) );
  MUX \Inst_Mem/U753  ( .A(\Inst_Mem/n741 ), .B(\Inst_Mem/n738 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n742 ) );
  MUX \Inst_Mem/U752  ( .A(\Inst_Mem/n740 ), .B(\Inst_Mem/n739 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n741 ) );
  MUX \Inst_Mem/U751  ( .A(inst_mem_in_wire[11]), .B(inst_mem_in_wire[43]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n740 ) );
  MUX \Inst_Mem/U750  ( .A(inst_mem_in_wire[75]), .B(inst_mem_in_wire[107]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n739 ) );
  MUX \Inst_Mem/U749  ( .A(\Inst_Mem/n737 ), .B(\Inst_Mem/n736 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n738 ) );
  MUX \Inst_Mem/U748  ( .A(inst_mem_in_wire[139]), .B(inst_mem_in_wire[171]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n737 ) );
  MUX \Inst_Mem/U747  ( .A(inst_mem_in_wire[203]), .B(inst_mem_in_wire[235]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n736 ) );
  MUX \Inst_Mem/U746  ( .A(\Inst_Mem/n734 ), .B(\Inst_Mem/n731 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n735 ) );
  MUX \Inst_Mem/U745  ( .A(\Inst_Mem/n733 ), .B(\Inst_Mem/n732 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n734 ) );
  MUX \Inst_Mem/U744  ( .A(inst_mem_in_wire[267]), .B(inst_mem_in_wire[299]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n733 ) );
  MUX \Inst_Mem/U743  ( .A(inst_mem_in_wire[331]), .B(inst_mem_in_wire[363]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n732 ) );
  MUX \Inst_Mem/U742  ( .A(\Inst_Mem/n730 ), .B(\Inst_Mem/n729 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n731 ) );
  MUX \Inst_Mem/U741  ( .A(inst_mem_in_wire[395]), .B(inst_mem_in_wire[427]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n730 ) );
  MUX \Inst_Mem/U740  ( .A(inst_mem_in_wire[459]), .B(inst_mem_in_wire[491]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n729 ) );
  MUX \Inst_Mem/U739  ( .A(\Inst_Mem/n727 ), .B(\Inst_Mem/n720 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n728 ) );
  MUX \Inst_Mem/U738  ( .A(\Inst_Mem/n726 ), .B(\Inst_Mem/n723 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n727 ) );
  MUX \Inst_Mem/U737  ( .A(\Inst_Mem/n725 ), .B(\Inst_Mem/n724 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n726 ) );
  MUX \Inst_Mem/U736  ( .A(inst_mem_in_wire[523]), .B(inst_mem_in_wire[555]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n725 ) );
  MUX \Inst_Mem/U735  ( .A(inst_mem_in_wire[587]), .B(inst_mem_in_wire[619]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n724 ) );
  MUX \Inst_Mem/U734  ( .A(\Inst_Mem/n722 ), .B(\Inst_Mem/n721 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n723 ) );
  MUX \Inst_Mem/U733  ( .A(inst_mem_in_wire[651]), .B(inst_mem_in_wire[683]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n722 ) );
  MUX \Inst_Mem/U732  ( .A(inst_mem_in_wire[715]), .B(inst_mem_in_wire[747]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n721 ) );
  MUX \Inst_Mem/U731  ( .A(\Inst_Mem/n719 ), .B(\Inst_Mem/n716 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n720 ) );
  MUX \Inst_Mem/U730  ( .A(\Inst_Mem/n718 ), .B(\Inst_Mem/n717 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n719 ) );
  MUX \Inst_Mem/U729  ( .A(inst_mem_in_wire[779]), .B(inst_mem_in_wire[811]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n718 ) );
  MUX \Inst_Mem/U728  ( .A(inst_mem_in_wire[843]), .B(inst_mem_in_wire[875]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n717 ) );
  MUX \Inst_Mem/U727  ( .A(\Inst_Mem/n715 ), .B(\Inst_Mem/n714 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n716 ) );
  MUX \Inst_Mem/U726  ( .A(inst_mem_in_wire[907]), .B(inst_mem_in_wire[939]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n715 ) );
  MUX \Inst_Mem/U725  ( .A(inst_mem_in_wire[971]), .B(inst_mem_in_wire[1003]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n714 ) );
  MUX \Inst_Mem/U724  ( .A(\Inst_Mem/n712 ), .B(\Inst_Mem/n697 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n713 ) );
  MUX \Inst_Mem/U723  ( .A(\Inst_Mem/n711 ), .B(\Inst_Mem/n704 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n712 ) );
  MUX \Inst_Mem/U722  ( .A(\Inst_Mem/n710 ), .B(\Inst_Mem/n707 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n711 ) );
  MUX \Inst_Mem/U721  ( .A(\Inst_Mem/n709 ), .B(\Inst_Mem/n708 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n710 ) );
  MUX \Inst_Mem/U720  ( .A(inst_mem_in_wire[1035]), .B(inst_mem_in_wire[1067]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n709 ) );
  MUX \Inst_Mem/U719  ( .A(inst_mem_in_wire[1099]), .B(inst_mem_in_wire[1131]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n708 ) );
  MUX \Inst_Mem/U718  ( .A(\Inst_Mem/n706 ), .B(\Inst_Mem/n705 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n707 ) );
  MUX \Inst_Mem/U717  ( .A(inst_mem_in_wire[1163]), .B(inst_mem_in_wire[1195]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n706 ) );
  MUX \Inst_Mem/U716  ( .A(inst_mem_in_wire[1227]), .B(inst_mem_in_wire[1259]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n705 ) );
  MUX \Inst_Mem/U715  ( .A(\Inst_Mem/n703 ), .B(\Inst_Mem/n700 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n704 ) );
  MUX \Inst_Mem/U714  ( .A(\Inst_Mem/n702 ), .B(\Inst_Mem/n701 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n703 ) );
  MUX \Inst_Mem/U713  ( .A(inst_mem_in_wire[1291]), .B(inst_mem_in_wire[1323]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n702 ) );
  MUX \Inst_Mem/U712  ( .A(inst_mem_in_wire[1355]), .B(inst_mem_in_wire[1387]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n701 ) );
  MUX \Inst_Mem/U711  ( .A(\Inst_Mem/n699 ), .B(\Inst_Mem/n698 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n700 ) );
  MUX \Inst_Mem/U710  ( .A(inst_mem_in_wire[1419]), .B(inst_mem_in_wire[1451]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n699 ) );
  MUX \Inst_Mem/U709  ( .A(inst_mem_in_wire[1483]), .B(inst_mem_in_wire[1515]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n698 ) );
  MUX \Inst_Mem/U708  ( .A(\Inst_Mem/n696 ), .B(\Inst_Mem/n689 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n697 ) );
  MUX \Inst_Mem/U707  ( .A(\Inst_Mem/n695 ), .B(\Inst_Mem/n692 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n696 ) );
  MUX \Inst_Mem/U706  ( .A(\Inst_Mem/n694 ), .B(\Inst_Mem/n693 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n695 ) );
  MUX \Inst_Mem/U705  ( .A(inst_mem_in_wire[1547]), .B(inst_mem_in_wire[1579]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n694 ) );
  MUX \Inst_Mem/U704  ( .A(inst_mem_in_wire[1611]), .B(inst_mem_in_wire[1643]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n693 ) );
  MUX \Inst_Mem/U703  ( .A(\Inst_Mem/n691 ), .B(\Inst_Mem/n690 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n692 ) );
  MUX \Inst_Mem/U702  ( .A(inst_mem_in_wire[1675]), .B(inst_mem_in_wire[1707]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n691 ) );
  MUX \Inst_Mem/U701  ( .A(inst_mem_in_wire[1739]), .B(inst_mem_in_wire[1771]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n690 ) );
  MUX \Inst_Mem/U700  ( .A(\Inst_Mem/n688 ), .B(\Inst_Mem/n685 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n689 ) );
  MUX \Inst_Mem/U699  ( .A(\Inst_Mem/n687 ), .B(\Inst_Mem/n686 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n688 ) );
  MUX \Inst_Mem/U698  ( .A(inst_mem_in_wire[1803]), .B(inst_mem_in_wire[1835]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n687 ) );
  MUX \Inst_Mem/U697  ( .A(inst_mem_in_wire[1867]), .B(inst_mem_in_wire[1899]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n686 ) );
  MUX \Inst_Mem/U696  ( .A(\Inst_Mem/n684 ), .B(\Inst_Mem/n683 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n685 ) );
  MUX \Inst_Mem/U695  ( .A(inst_mem_in_wire[1931]), .B(inst_mem_in_wire[1963]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n684 ) );
  MUX \Inst_Mem/U694  ( .A(inst_mem_in_wire[1995]), .B(inst_mem_in_wire[2027]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n683 ) );
  MUX \Inst_Mem/U693  ( .A(\Inst_Mem/n682 ), .B(\Inst_Mem/n651 ), .S(
        pc_current[7]), .Z(imm[10]) );
  MUX \Inst_Mem/U692  ( .A(\Inst_Mem/n681 ), .B(\Inst_Mem/n666 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n682 ) );
  MUX \Inst_Mem/U691  ( .A(\Inst_Mem/n680 ), .B(\Inst_Mem/n673 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n681 ) );
  MUX \Inst_Mem/U690  ( .A(\Inst_Mem/n679 ), .B(\Inst_Mem/n676 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n680 ) );
  MUX \Inst_Mem/U689  ( .A(\Inst_Mem/n678 ), .B(\Inst_Mem/n677 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n679 ) );
  MUX \Inst_Mem/U688  ( .A(inst_mem_in_wire[10]), .B(inst_mem_in_wire[42]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n678 ) );
  MUX \Inst_Mem/U687  ( .A(inst_mem_in_wire[74]), .B(inst_mem_in_wire[106]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n677 ) );
  MUX \Inst_Mem/U686  ( .A(\Inst_Mem/n675 ), .B(\Inst_Mem/n674 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n676 ) );
  MUX \Inst_Mem/U685  ( .A(inst_mem_in_wire[138]), .B(inst_mem_in_wire[170]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n675 ) );
  MUX \Inst_Mem/U684  ( .A(inst_mem_in_wire[202]), .B(inst_mem_in_wire[234]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n674 ) );
  MUX \Inst_Mem/U683  ( .A(\Inst_Mem/n672 ), .B(\Inst_Mem/n669 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n673 ) );
  MUX \Inst_Mem/U682  ( .A(\Inst_Mem/n671 ), .B(\Inst_Mem/n670 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n672 ) );
  MUX \Inst_Mem/U681  ( .A(inst_mem_in_wire[266]), .B(inst_mem_in_wire[298]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n671 ) );
  MUX \Inst_Mem/U680  ( .A(inst_mem_in_wire[330]), .B(inst_mem_in_wire[362]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n670 ) );
  MUX \Inst_Mem/U679  ( .A(\Inst_Mem/n668 ), .B(\Inst_Mem/n667 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n669 ) );
  MUX \Inst_Mem/U678  ( .A(inst_mem_in_wire[394]), .B(inst_mem_in_wire[426]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n668 ) );
  MUX \Inst_Mem/U677  ( .A(inst_mem_in_wire[458]), .B(inst_mem_in_wire[490]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n667 ) );
  MUX \Inst_Mem/U676  ( .A(\Inst_Mem/n665 ), .B(\Inst_Mem/n658 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n666 ) );
  MUX \Inst_Mem/U675  ( .A(\Inst_Mem/n664 ), .B(\Inst_Mem/n661 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n665 ) );
  MUX \Inst_Mem/U674  ( .A(\Inst_Mem/n663 ), .B(\Inst_Mem/n662 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n664 ) );
  MUX \Inst_Mem/U673  ( .A(inst_mem_in_wire[522]), .B(inst_mem_in_wire[554]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n663 ) );
  MUX \Inst_Mem/U672  ( .A(inst_mem_in_wire[586]), .B(inst_mem_in_wire[618]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n662 ) );
  MUX \Inst_Mem/U671  ( .A(\Inst_Mem/n660 ), .B(\Inst_Mem/n659 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n661 ) );
  MUX \Inst_Mem/U670  ( .A(inst_mem_in_wire[650]), .B(inst_mem_in_wire[682]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n660 ) );
  MUX \Inst_Mem/U669  ( .A(inst_mem_in_wire[714]), .B(inst_mem_in_wire[746]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n659 ) );
  MUX \Inst_Mem/U668  ( .A(\Inst_Mem/n657 ), .B(\Inst_Mem/n654 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n658 ) );
  MUX \Inst_Mem/U667  ( .A(\Inst_Mem/n656 ), .B(\Inst_Mem/n655 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n657 ) );
  MUX \Inst_Mem/U666  ( .A(inst_mem_in_wire[778]), .B(inst_mem_in_wire[810]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n656 ) );
  MUX \Inst_Mem/U665  ( .A(inst_mem_in_wire[842]), .B(inst_mem_in_wire[874]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n655 ) );
  MUX \Inst_Mem/U664  ( .A(\Inst_Mem/n653 ), .B(\Inst_Mem/n652 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n654 ) );
  MUX \Inst_Mem/U663  ( .A(inst_mem_in_wire[906]), .B(inst_mem_in_wire[938]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n653 ) );
  MUX \Inst_Mem/U662  ( .A(inst_mem_in_wire[970]), .B(inst_mem_in_wire[1002]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n652 ) );
  MUX \Inst_Mem/U661  ( .A(\Inst_Mem/n650 ), .B(\Inst_Mem/n635 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n651 ) );
  MUX \Inst_Mem/U660  ( .A(\Inst_Mem/n649 ), .B(\Inst_Mem/n642 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n650 ) );
  MUX \Inst_Mem/U659  ( .A(\Inst_Mem/n648 ), .B(\Inst_Mem/n645 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n649 ) );
  MUX \Inst_Mem/U658  ( .A(\Inst_Mem/n647 ), .B(\Inst_Mem/n646 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n648 ) );
  MUX \Inst_Mem/U657  ( .A(inst_mem_in_wire[1034]), .B(inst_mem_in_wire[1066]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n647 ) );
  MUX \Inst_Mem/U656  ( .A(inst_mem_in_wire[1098]), .B(inst_mem_in_wire[1130]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n646 ) );
  MUX \Inst_Mem/U655  ( .A(\Inst_Mem/n644 ), .B(\Inst_Mem/n643 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n645 ) );
  MUX \Inst_Mem/U654  ( .A(inst_mem_in_wire[1162]), .B(inst_mem_in_wire[1194]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n644 ) );
  MUX \Inst_Mem/U653  ( .A(inst_mem_in_wire[1226]), .B(inst_mem_in_wire[1258]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n643 ) );
  MUX \Inst_Mem/U652  ( .A(\Inst_Mem/n641 ), .B(\Inst_Mem/n638 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n642 ) );
  MUX \Inst_Mem/U651  ( .A(\Inst_Mem/n640 ), .B(\Inst_Mem/n639 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n641 ) );
  MUX \Inst_Mem/U650  ( .A(inst_mem_in_wire[1290]), .B(inst_mem_in_wire[1322]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n640 ) );
  MUX \Inst_Mem/U649  ( .A(inst_mem_in_wire[1354]), .B(inst_mem_in_wire[1386]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n639 ) );
  MUX \Inst_Mem/U648  ( .A(\Inst_Mem/n637 ), .B(\Inst_Mem/n636 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n638 ) );
  MUX \Inst_Mem/U647  ( .A(inst_mem_in_wire[1418]), .B(inst_mem_in_wire[1450]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n637 ) );
  MUX \Inst_Mem/U646  ( .A(inst_mem_in_wire[1482]), .B(inst_mem_in_wire[1514]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n636 ) );
  MUX \Inst_Mem/U645  ( .A(\Inst_Mem/n634 ), .B(\Inst_Mem/n627 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n635 ) );
  MUX \Inst_Mem/U644  ( .A(\Inst_Mem/n633 ), .B(\Inst_Mem/n630 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n634 ) );
  MUX \Inst_Mem/U643  ( .A(\Inst_Mem/n632 ), .B(\Inst_Mem/n631 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n633 ) );
  MUX \Inst_Mem/U642  ( .A(inst_mem_in_wire[1546]), .B(inst_mem_in_wire[1578]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n632 ) );
  MUX \Inst_Mem/U641  ( .A(inst_mem_in_wire[1610]), .B(inst_mem_in_wire[1642]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n631 ) );
  MUX \Inst_Mem/U640  ( .A(\Inst_Mem/n629 ), .B(\Inst_Mem/n628 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n630 ) );
  MUX \Inst_Mem/U639  ( .A(inst_mem_in_wire[1674]), .B(inst_mem_in_wire[1706]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n629 ) );
  MUX \Inst_Mem/U638  ( .A(inst_mem_in_wire[1738]), .B(inst_mem_in_wire[1770]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n628 ) );
  MUX \Inst_Mem/U637  ( .A(\Inst_Mem/n626 ), .B(\Inst_Mem/n623 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n627 ) );
  MUX \Inst_Mem/U636  ( .A(\Inst_Mem/n625 ), .B(\Inst_Mem/n624 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n626 ) );
  MUX \Inst_Mem/U635  ( .A(inst_mem_in_wire[1802]), .B(inst_mem_in_wire[1834]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n625 ) );
  MUX \Inst_Mem/U634  ( .A(inst_mem_in_wire[1866]), .B(inst_mem_in_wire[1898]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n624 ) );
  MUX \Inst_Mem/U633  ( .A(\Inst_Mem/n622 ), .B(\Inst_Mem/n621 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n623 ) );
  MUX \Inst_Mem/U632  ( .A(inst_mem_in_wire[1930]), .B(inst_mem_in_wire[1962]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n622 ) );
  MUX \Inst_Mem/U631  ( .A(inst_mem_in_wire[1994]), .B(inst_mem_in_wire[2026]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n621 ) );
  MUX \Inst_Mem/U630  ( .A(\Inst_Mem/n620 ), .B(\Inst_Mem/n589 ), .S(
        pc_current[7]), .Z(imm[9]) );
  MUX \Inst_Mem/U629  ( .A(\Inst_Mem/n619 ), .B(\Inst_Mem/n604 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n620 ) );
  MUX \Inst_Mem/U628  ( .A(\Inst_Mem/n618 ), .B(\Inst_Mem/n611 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n619 ) );
  MUX \Inst_Mem/U627  ( .A(\Inst_Mem/n617 ), .B(\Inst_Mem/n614 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n618 ) );
  MUX \Inst_Mem/U626  ( .A(\Inst_Mem/n616 ), .B(\Inst_Mem/n615 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n617 ) );
  MUX \Inst_Mem/U625  ( .A(inst_mem_in_wire[9]), .B(inst_mem_in_wire[41]), .S(
        pc_current[2]), .Z(\Inst_Mem/n616 ) );
  MUX \Inst_Mem/U624  ( .A(inst_mem_in_wire[73]), .B(inst_mem_in_wire[105]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n615 ) );
  MUX \Inst_Mem/U623  ( .A(\Inst_Mem/n613 ), .B(\Inst_Mem/n612 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n614 ) );
  MUX \Inst_Mem/U622  ( .A(inst_mem_in_wire[137]), .B(inst_mem_in_wire[169]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n613 ) );
  MUX \Inst_Mem/U621  ( .A(inst_mem_in_wire[201]), .B(inst_mem_in_wire[233]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n612 ) );
  MUX \Inst_Mem/U620  ( .A(\Inst_Mem/n610 ), .B(\Inst_Mem/n607 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n611 ) );
  MUX \Inst_Mem/U619  ( .A(\Inst_Mem/n609 ), .B(\Inst_Mem/n608 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n610 ) );
  MUX \Inst_Mem/U618  ( .A(inst_mem_in_wire[265]), .B(inst_mem_in_wire[297]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n609 ) );
  MUX \Inst_Mem/U617  ( .A(inst_mem_in_wire[329]), .B(inst_mem_in_wire[361]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n608 ) );
  MUX \Inst_Mem/U616  ( .A(\Inst_Mem/n606 ), .B(\Inst_Mem/n605 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n607 ) );
  MUX \Inst_Mem/U615  ( .A(inst_mem_in_wire[393]), .B(inst_mem_in_wire[425]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n606 ) );
  MUX \Inst_Mem/U614  ( .A(inst_mem_in_wire[457]), .B(inst_mem_in_wire[489]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n605 ) );
  MUX \Inst_Mem/U613  ( .A(\Inst_Mem/n603 ), .B(\Inst_Mem/n596 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n604 ) );
  MUX \Inst_Mem/U612  ( .A(\Inst_Mem/n602 ), .B(\Inst_Mem/n599 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n603 ) );
  MUX \Inst_Mem/U611  ( .A(\Inst_Mem/n601 ), .B(\Inst_Mem/n600 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n602 ) );
  MUX \Inst_Mem/U610  ( .A(inst_mem_in_wire[521]), .B(inst_mem_in_wire[553]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n601 ) );
  MUX \Inst_Mem/U609  ( .A(inst_mem_in_wire[585]), .B(inst_mem_in_wire[617]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n600 ) );
  MUX \Inst_Mem/U608  ( .A(\Inst_Mem/n598 ), .B(\Inst_Mem/n597 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n599 ) );
  MUX \Inst_Mem/U607  ( .A(inst_mem_in_wire[649]), .B(inst_mem_in_wire[681]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n598 ) );
  MUX \Inst_Mem/U606  ( .A(inst_mem_in_wire[713]), .B(inst_mem_in_wire[745]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n597 ) );
  MUX \Inst_Mem/U605  ( .A(\Inst_Mem/n595 ), .B(\Inst_Mem/n592 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n596 ) );
  MUX \Inst_Mem/U604  ( .A(\Inst_Mem/n594 ), .B(\Inst_Mem/n593 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n595 ) );
  MUX \Inst_Mem/U603  ( .A(inst_mem_in_wire[777]), .B(inst_mem_in_wire[809]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n594 ) );
  MUX \Inst_Mem/U602  ( .A(inst_mem_in_wire[841]), .B(inst_mem_in_wire[873]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n593 ) );
  MUX \Inst_Mem/U601  ( .A(\Inst_Mem/n591 ), .B(\Inst_Mem/n590 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n592 ) );
  MUX \Inst_Mem/U600  ( .A(inst_mem_in_wire[905]), .B(inst_mem_in_wire[937]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n591 ) );
  MUX \Inst_Mem/U599  ( .A(inst_mem_in_wire[969]), .B(inst_mem_in_wire[1001]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n590 ) );
  MUX \Inst_Mem/U598  ( .A(\Inst_Mem/n588 ), .B(\Inst_Mem/n573 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n589 ) );
  MUX \Inst_Mem/U597  ( .A(\Inst_Mem/n587 ), .B(\Inst_Mem/n580 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n588 ) );
  MUX \Inst_Mem/U596  ( .A(\Inst_Mem/n586 ), .B(\Inst_Mem/n583 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n587 ) );
  MUX \Inst_Mem/U595  ( .A(\Inst_Mem/n585 ), .B(\Inst_Mem/n584 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n586 ) );
  MUX \Inst_Mem/U594  ( .A(inst_mem_in_wire[1033]), .B(inst_mem_in_wire[1065]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n585 ) );
  MUX \Inst_Mem/U593  ( .A(inst_mem_in_wire[1097]), .B(inst_mem_in_wire[1129]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n584 ) );
  MUX \Inst_Mem/U592  ( .A(\Inst_Mem/n582 ), .B(\Inst_Mem/n581 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n583 ) );
  MUX \Inst_Mem/U591  ( .A(inst_mem_in_wire[1161]), .B(inst_mem_in_wire[1193]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n582 ) );
  MUX \Inst_Mem/U590  ( .A(inst_mem_in_wire[1225]), .B(inst_mem_in_wire[1257]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n581 ) );
  MUX \Inst_Mem/U589  ( .A(\Inst_Mem/n579 ), .B(\Inst_Mem/n576 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n580 ) );
  MUX \Inst_Mem/U588  ( .A(\Inst_Mem/n578 ), .B(\Inst_Mem/n577 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n579 ) );
  MUX \Inst_Mem/U587  ( .A(inst_mem_in_wire[1289]), .B(inst_mem_in_wire[1321]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n578 ) );
  MUX \Inst_Mem/U586  ( .A(inst_mem_in_wire[1353]), .B(inst_mem_in_wire[1385]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n577 ) );
  MUX \Inst_Mem/U585  ( .A(\Inst_Mem/n575 ), .B(\Inst_Mem/n574 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n576 ) );
  MUX \Inst_Mem/U584  ( .A(inst_mem_in_wire[1417]), .B(inst_mem_in_wire[1449]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n575 ) );
  MUX \Inst_Mem/U583  ( .A(inst_mem_in_wire[1481]), .B(inst_mem_in_wire[1513]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n574 ) );
  MUX \Inst_Mem/U582  ( .A(\Inst_Mem/n572 ), .B(\Inst_Mem/n565 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n573 ) );
  MUX \Inst_Mem/U581  ( .A(\Inst_Mem/n571 ), .B(\Inst_Mem/n568 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n572 ) );
  MUX \Inst_Mem/U580  ( .A(\Inst_Mem/n570 ), .B(\Inst_Mem/n569 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n571 ) );
  MUX \Inst_Mem/U579  ( .A(inst_mem_in_wire[1545]), .B(inst_mem_in_wire[1577]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n570 ) );
  MUX \Inst_Mem/U578  ( .A(inst_mem_in_wire[1609]), .B(inst_mem_in_wire[1641]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n569 ) );
  MUX \Inst_Mem/U577  ( .A(\Inst_Mem/n567 ), .B(\Inst_Mem/n566 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n568 ) );
  MUX \Inst_Mem/U576  ( .A(inst_mem_in_wire[1673]), .B(inst_mem_in_wire[1705]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n567 ) );
  MUX \Inst_Mem/U575  ( .A(inst_mem_in_wire[1737]), .B(inst_mem_in_wire[1769]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n566 ) );
  MUX \Inst_Mem/U574  ( .A(\Inst_Mem/n564 ), .B(\Inst_Mem/n561 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n565 ) );
  MUX \Inst_Mem/U573  ( .A(\Inst_Mem/n563 ), .B(\Inst_Mem/n562 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n564 ) );
  MUX \Inst_Mem/U572  ( .A(inst_mem_in_wire[1801]), .B(inst_mem_in_wire[1833]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n563 ) );
  MUX \Inst_Mem/U571  ( .A(inst_mem_in_wire[1865]), .B(inst_mem_in_wire[1897]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n562 ) );
  MUX \Inst_Mem/U570  ( .A(\Inst_Mem/n560 ), .B(\Inst_Mem/n559 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n561 ) );
  MUX \Inst_Mem/U569  ( .A(inst_mem_in_wire[1929]), .B(inst_mem_in_wire[1961]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n560 ) );
  MUX \Inst_Mem/U568  ( .A(inst_mem_in_wire[1993]), .B(inst_mem_in_wire[2025]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n559 ) );
  MUX \Inst_Mem/U567  ( .A(\Inst_Mem/n558 ), .B(\Inst_Mem/n527 ), .S(
        pc_current[7]), .Z(imm[8]) );
  MUX \Inst_Mem/U566  ( .A(\Inst_Mem/n557 ), .B(\Inst_Mem/n542 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n558 ) );
  MUX \Inst_Mem/U565  ( .A(\Inst_Mem/n556 ), .B(\Inst_Mem/n549 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n557 ) );
  MUX \Inst_Mem/U564  ( .A(\Inst_Mem/n555 ), .B(\Inst_Mem/n552 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n556 ) );
  MUX \Inst_Mem/U563  ( .A(\Inst_Mem/n554 ), .B(\Inst_Mem/n553 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n555 ) );
  MUX \Inst_Mem/U562  ( .A(inst_mem_in_wire[8]), .B(inst_mem_in_wire[40]), .S(
        pc_current[2]), .Z(\Inst_Mem/n554 ) );
  MUX \Inst_Mem/U561  ( .A(inst_mem_in_wire[72]), .B(inst_mem_in_wire[104]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n553 ) );
  MUX \Inst_Mem/U560  ( .A(\Inst_Mem/n551 ), .B(\Inst_Mem/n550 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n552 ) );
  MUX \Inst_Mem/U559  ( .A(inst_mem_in_wire[136]), .B(inst_mem_in_wire[168]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n551 ) );
  MUX \Inst_Mem/U558  ( .A(inst_mem_in_wire[200]), .B(inst_mem_in_wire[232]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n550 ) );
  MUX \Inst_Mem/U557  ( .A(\Inst_Mem/n548 ), .B(\Inst_Mem/n545 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n549 ) );
  MUX \Inst_Mem/U556  ( .A(\Inst_Mem/n547 ), .B(\Inst_Mem/n546 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n548 ) );
  MUX \Inst_Mem/U555  ( .A(inst_mem_in_wire[264]), .B(inst_mem_in_wire[296]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n547 ) );
  MUX \Inst_Mem/U554  ( .A(inst_mem_in_wire[328]), .B(inst_mem_in_wire[360]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n546 ) );
  MUX \Inst_Mem/U553  ( .A(\Inst_Mem/n544 ), .B(\Inst_Mem/n543 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n545 ) );
  MUX \Inst_Mem/U552  ( .A(inst_mem_in_wire[392]), .B(inst_mem_in_wire[424]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n544 ) );
  MUX \Inst_Mem/U551  ( .A(inst_mem_in_wire[456]), .B(inst_mem_in_wire[488]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n543 ) );
  MUX \Inst_Mem/U550  ( .A(\Inst_Mem/n541 ), .B(\Inst_Mem/n534 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n542 ) );
  MUX \Inst_Mem/U549  ( .A(\Inst_Mem/n540 ), .B(\Inst_Mem/n537 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n541 ) );
  MUX \Inst_Mem/U548  ( .A(\Inst_Mem/n539 ), .B(\Inst_Mem/n538 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n540 ) );
  MUX \Inst_Mem/U547  ( .A(inst_mem_in_wire[520]), .B(inst_mem_in_wire[552]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n539 ) );
  MUX \Inst_Mem/U546  ( .A(inst_mem_in_wire[584]), .B(inst_mem_in_wire[616]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n538 ) );
  MUX \Inst_Mem/U545  ( .A(\Inst_Mem/n536 ), .B(\Inst_Mem/n535 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n537 ) );
  MUX \Inst_Mem/U544  ( .A(inst_mem_in_wire[648]), .B(inst_mem_in_wire[680]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n536 ) );
  MUX \Inst_Mem/U543  ( .A(inst_mem_in_wire[712]), .B(inst_mem_in_wire[744]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n535 ) );
  MUX \Inst_Mem/U542  ( .A(\Inst_Mem/n533 ), .B(\Inst_Mem/n530 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n534 ) );
  MUX \Inst_Mem/U541  ( .A(\Inst_Mem/n532 ), .B(\Inst_Mem/n531 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n533 ) );
  MUX \Inst_Mem/U540  ( .A(inst_mem_in_wire[776]), .B(inst_mem_in_wire[808]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n532 ) );
  MUX \Inst_Mem/U539  ( .A(inst_mem_in_wire[840]), .B(inst_mem_in_wire[872]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n531 ) );
  MUX \Inst_Mem/U538  ( .A(\Inst_Mem/n529 ), .B(\Inst_Mem/n528 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n530 ) );
  MUX \Inst_Mem/U537  ( .A(inst_mem_in_wire[904]), .B(inst_mem_in_wire[936]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n529 ) );
  MUX \Inst_Mem/U536  ( .A(inst_mem_in_wire[968]), .B(inst_mem_in_wire[1000]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n528 ) );
  MUX \Inst_Mem/U535  ( .A(\Inst_Mem/n526 ), .B(\Inst_Mem/n511 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n527 ) );
  MUX \Inst_Mem/U534  ( .A(\Inst_Mem/n525 ), .B(\Inst_Mem/n518 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n526 ) );
  MUX \Inst_Mem/U533  ( .A(\Inst_Mem/n524 ), .B(\Inst_Mem/n521 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n525 ) );
  MUX \Inst_Mem/U532  ( .A(\Inst_Mem/n523 ), .B(\Inst_Mem/n522 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n524 ) );
  MUX \Inst_Mem/U531  ( .A(inst_mem_in_wire[1032]), .B(inst_mem_in_wire[1064]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n523 ) );
  MUX \Inst_Mem/U530  ( .A(inst_mem_in_wire[1096]), .B(inst_mem_in_wire[1128]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n522 ) );
  MUX \Inst_Mem/U529  ( .A(\Inst_Mem/n520 ), .B(\Inst_Mem/n519 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n521 ) );
  MUX \Inst_Mem/U528  ( .A(inst_mem_in_wire[1160]), .B(inst_mem_in_wire[1192]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n520 ) );
  MUX \Inst_Mem/U527  ( .A(inst_mem_in_wire[1224]), .B(inst_mem_in_wire[1256]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n519 ) );
  MUX \Inst_Mem/U526  ( .A(\Inst_Mem/n517 ), .B(\Inst_Mem/n514 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n518 ) );
  MUX \Inst_Mem/U525  ( .A(\Inst_Mem/n516 ), .B(\Inst_Mem/n515 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n517 ) );
  MUX \Inst_Mem/U524  ( .A(inst_mem_in_wire[1288]), .B(inst_mem_in_wire[1320]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n516 ) );
  MUX \Inst_Mem/U523  ( .A(inst_mem_in_wire[1352]), .B(inst_mem_in_wire[1384]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n515 ) );
  MUX \Inst_Mem/U522  ( .A(\Inst_Mem/n513 ), .B(\Inst_Mem/n512 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n514 ) );
  MUX \Inst_Mem/U521  ( .A(inst_mem_in_wire[1416]), .B(inst_mem_in_wire[1448]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n513 ) );
  MUX \Inst_Mem/U520  ( .A(inst_mem_in_wire[1480]), .B(inst_mem_in_wire[1512]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n512 ) );
  MUX \Inst_Mem/U519  ( .A(\Inst_Mem/n510 ), .B(\Inst_Mem/n503 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n511 ) );
  MUX \Inst_Mem/U518  ( .A(\Inst_Mem/n509 ), .B(\Inst_Mem/n506 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n510 ) );
  MUX \Inst_Mem/U517  ( .A(\Inst_Mem/n508 ), .B(\Inst_Mem/n507 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n509 ) );
  MUX \Inst_Mem/U516  ( .A(inst_mem_in_wire[1544]), .B(inst_mem_in_wire[1576]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n508 ) );
  MUX \Inst_Mem/U515  ( .A(inst_mem_in_wire[1608]), .B(inst_mem_in_wire[1640]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n507 ) );
  MUX \Inst_Mem/U514  ( .A(\Inst_Mem/n505 ), .B(\Inst_Mem/n504 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n506 ) );
  MUX \Inst_Mem/U513  ( .A(inst_mem_in_wire[1672]), .B(inst_mem_in_wire[1704]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n505 ) );
  MUX \Inst_Mem/U512  ( .A(inst_mem_in_wire[1736]), .B(inst_mem_in_wire[1768]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n504 ) );
  MUX \Inst_Mem/U511  ( .A(\Inst_Mem/n502 ), .B(\Inst_Mem/n499 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n503 ) );
  MUX \Inst_Mem/U510  ( .A(\Inst_Mem/n501 ), .B(\Inst_Mem/n500 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n502 ) );
  MUX \Inst_Mem/U509  ( .A(inst_mem_in_wire[1800]), .B(inst_mem_in_wire[1832]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n501 ) );
  MUX \Inst_Mem/U508  ( .A(inst_mem_in_wire[1864]), .B(inst_mem_in_wire[1896]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n500 ) );
  MUX \Inst_Mem/U507  ( .A(\Inst_Mem/n498 ), .B(\Inst_Mem/n497 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n499 ) );
  MUX \Inst_Mem/U506  ( .A(inst_mem_in_wire[1928]), .B(inst_mem_in_wire[1960]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n498 ) );
  MUX \Inst_Mem/U505  ( .A(inst_mem_in_wire[1992]), .B(inst_mem_in_wire[2024]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n497 ) );
  MUX \Inst_Mem/U504  ( .A(\Inst_Mem/n496 ), .B(\Inst_Mem/n465 ), .S(
        pc_current[7]), .Z(imm[7]) );
  MUX \Inst_Mem/U503  ( .A(\Inst_Mem/n495 ), .B(\Inst_Mem/n480 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n496 ) );
  MUX \Inst_Mem/U502  ( .A(\Inst_Mem/n494 ), .B(\Inst_Mem/n487 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n495 ) );
  MUX \Inst_Mem/U501  ( .A(\Inst_Mem/n493 ), .B(\Inst_Mem/n490 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n494 ) );
  MUX \Inst_Mem/U500  ( .A(\Inst_Mem/n492 ), .B(\Inst_Mem/n491 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n493 ) );
  MUX \Inst_Mem/U499  ( .A(inst_mem_in_wire[7]), .B(inst_mem_in_wire[39]), .S(
        pc_current[2]), .Z(\Inst_Mem/n492 ) );
  MUX \Inst_Mem/U498  ( .A(inst_mem_in_wire[71]), .B(inst_mem_in_wire[103]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n491 ) );
  MUX \Inst_Mem/U497  ( .A(\Inst_Mem/n489 ), .B(\Inst_Mem/n488 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n490 ) );
  MUX \Inst_Mem/U496  ( .A(inst_mem_in_wire[135]), .B(inst_mem_in_wire[167]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n489 ) );
  MUX \Inst_Mem/U495  ( .A(inst_mem_in_wire[199]), .B(inst_mem_in_wire[231]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n488 ) );
  MUX \Inst_Mem/U494  ( .A(\Inst_Mem/n486 ), .B(\Inst_Mem/n483 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n487 ) );
  MUX \Inst_Mem/U493  ( .A(\Inst_Mem/n485 ), .B(\Inst_Mem/n484 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n486 ) );
  MUX \Inst_Mem/U492  ( .A(inst_mem_in_wire[263]), .B(inst_mem_in_wire[295]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n485 ) );
  MUX \Inst_Mem/U491  ( .A(inst_mem_in_wire[327]), .B(inst_mem_in_wire[359]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n484 ) );
  MUX \Inst_Mem/U490  ( .A(\Inst_Mem/n482 ), .B(\Inst_Mem/n481 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n483 ) );
  MUX \Inst_Mem/U489  ( .A(inst_mem_in_wire[391]), .B(inst_mem_in_wire[423]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n482 ) );
  MUX \Inst_Mem/U488  ( .A(inst_mem_in_wire[455]), .B(inst_mem_in_wire[487]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n481 ) );
  MUX \Inst_Mem/U487  ( .A(\Inst_Mem/n479 ), .B(\Inst_Mem/n472 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n480 ) );
  MUX \Inst_Mem/U486  ( .A(\Inst_Mem/n478 ), .B(\Inst_Mem/n475 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n479 ) );
  MUX \Inst_Mem/U485  ( .A(\Inst_Mem/n477 ), .B(\Inst_Mem/n476 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n478 ) );
  MUX \Inst_Mem/U484  ( .A(inst_mem_in_wire[519]), .B(inst_mem_in_wire[551]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n477 ) );
  MUX \Inst_Mem/U483  ( .A(inst_mem_in_wire[583]), .B(inst_mem_in_wire[615]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n476 ) );
  MUX \Inst_Mem/U482  ( .A(\Inst_Mem/n474 ), .B(\Inst_Mem/n473 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n475 ) );
  MUX \Inst_Mem/U481  ( .A(inst_mem_in_wire[647]), .B(inst_mem_in_wire[679]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n474 ) );
  MUX \Inst_Mem/U480  ( .A(inst_mem_in_wire[711]), .B(inst_mem_in_wire[743]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n473 ) );
  MUX \Inst_Mem/U479  ( .A(\Inst_Mem/n471 ), .B(\Inst_Mem/n468 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n472 ) );
  MUX \Inst_Mem/U478  ( .A(\Inst_Mem/n470 ), .B(\Inst_Mem/n469 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n471 ) );
  MUX \Inst_Mem/U477  ( .A(inst_mem_in_wire[775]), .B(inst_mem_in_wire[807]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n470 ) );
  MUX \Inst_Mem/U476  ( .A(inst_mem_in_wire[839]), .B(inst_mem_in_wire[871]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n469 ) );
  MUX \Inst_Mem/U475  ( .A(\Inst_Mem/n467 ), .B(\Inst_Mem/n466 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n468 ) );
  MUX \Inst_Mem/U474  ( .A(inst_mem_in_wire[903]), .B(inst_mem_in_wire[935]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n467 ) );
  MUX \Inst_Mem/U473  ( .A(inst_mem_in_wire[967]), .B(inst_mem_in_wire[999]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n466 ) );
  MUX \Inst_Mem/U472  ( .A(\Inst_Mem/n464 ), .B(\Inst_Mem/n449 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n465 ) );
  MUX \Inst_Mem/U471  ( .A(\Inst_Mem/n463 ), .B(\Inst_Mem/n456 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n464 ) );
  MUX \Inst_Mem/U470  ( .A(\Inst_Mem/n462 ), .B(\Inst_Mem/n459 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n463 ) );
  MUX \Inst_Mem/U469  ( .A(\Inst_Mem/n461 ), .B(\Inst_Mem/n460 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n462 ) );
  MUX \Inst_Mem/U468  ( .A(inst_mem_in_wire[1031]), .B(inst_mem_in_wire[1063]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n461 ) );
  MUX \Inst_Mem/U467  ( .A(inst_mem_in_wire[1095]), .B(inst_mem_in_wire[1127]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n460 ) );
  MUX \Inst_Mem/U466  ( .A(\Inst_Mem/n458 ), .B(\Inst_Mem/n457 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n459 ) );
  MUX \Inst_Mem/U465  ( .A(inst_mem_in_wire[1159]), .B(inst_mem_in_wire[1191]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n458 ) );
  MUX \Inst_Mem/U464  ( .A(inst_mem_in_wire[1223]), .B(inst_mem_in_wire[1255]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n457 ) );
  MUX \Inst_Mem/U463  ( .A(\Inst_Mem/n455 ), .B(\Inst_Mem/n452 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n456 ) );
  MUX \Inst_Mem/U462  ( .A(\Inst_Mem/n454 ), .B(\Inst_Mem/n453 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n455 ) );
  MUX \Inst_Mem/U461  ( .A(inst_mem_in_wire[1287]), .B(inst_mem_in_wire[1319]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n454 ) );
  MUX \Inst_Mem/U460  ( .A(inst_mem_in_wire[1351]), .B(inst_mem_in_wire[1383]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n453 ) );
  MUX \Inst_Mem/U459  ( .A(\Inst_Mem/n451 ), .B(\Inst_Mem/n450 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n452 ) );
  MUX \Inst_Mem/U458  ( .A(inst_mem_in_wire[1415]), .B(inst_mem_in_wire[1447]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n451 ) );
  MUX \Inst_Mem/U457  ( .A(inst_mem_in_wire[1479]), .B(inst_mem_in_wire[1511]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n450 ) );
  MUX \Inst_Mem/U456  ( .A(\Inst_Mem/n448 ), .B(\Inst_Mem/n441 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n449 ) );
  MUX \Inst_Mem/U455  ( .A(\Inst_Mem/n447 ), .B(\Inst_Mem/n444 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n448 ) );
  MUX \Inst_Mem/U454  ( .A(\Inst_Mem/n446 ), .B(\Inst_Mem/n445 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n447 ) );
  MUX \Inst_Mem/U453  ( .A(inst_mem_in_wire[1543]), .B(inst_mem_in_wire[1575]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n446 ) );
  MUX \Inst_Mem/U452  ( .A(inst_mem_in_wire[1607]), .B(inst_mem_in_wire[1639]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n445 ) );
  MUX \Inst_Mem/U451  ( .A(\Inst_Mem/n443 ), .B(\Inst_Mem/n442 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n444 ) );
  MUX \Inst_Mem/U450  ( .A(inst_mem_in_wire[1671]), .B(inst_mem_in_wire[1703]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n443 ) );
  MUX \Inst_Mem/U449  ( .A(inst_mem_in_wire[1735]), .B(inst_mem_in_wire[1767]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n442 ) );
  MUX \Inst_Mem/U448  ( .A(\Inst_Mem/n440 ), .B(\Inst_Mem/n437 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n441 ) );
  MUX \Inst_Mem/U447  ( .A(\Inst_Mem/n439 ), .B(\Inst_Mem/n438 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n440 ) );
  MUX \Inst_Mem/U446  ( .A(inst_mem_in_wire[1799]), .B(inst_mem_in_wire[1831]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n439 ) );
  MUX \Inst_Mem/U445  ( .A(inst_mem_in_wire[1863]), .B(inst_mem_in_wire[1895]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n438 ) );
  MUX \Inst_Mem/U444  ( .A(\Inst_Mem/n436 ), .B(\Inst_Mem/n435 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n437 ) );
  MUX \Inst_Mem/U443  ( .A(inst_mem_in_wire[1927]), .B(inst_mem_in_wire[1959]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n436 ) );
  MUX \Inst_Mem/U442  ( .A(inst_mem_in_wire[1991]), .B(inst_mem_in_wire[2023]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n435 ) );
  MUX \Inst_Mem/U441  ( .A(\Inst_Mem/n434 ), .B(\Inst_Mem/n403 ), .S(
        pc_current[7]), .Z(imm[6]) );
  MUX \Inst_Mem/U440  ( .A(\Inst_Mem/n433 ), .B(\Inst_Mem/n418 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n434 ) );
  MUX \Inst_Mem/U439  ( .A(\Inst_Mem/n432 ), .B(\Inst_Mem/n425 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n433 ) );
  MUX \Inst_Mem/U438  ( .A(\Inst_Mem/n431 ), .B(\Inst_Mem/n428 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n432 ) );
  MUX \Inst_Mem/U437  ( .A(\Inst_Mem/n430 ), .B(\Inst_Mem/n429 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n431 ) );
  MUX \Inst_Mem/U436  ( .A(inst_mem_in_wire[6]), .B(inst_mem_in_wire[38]), .S(
        pc_current[2]), .Z(\Inst_Mem/n430 ) );
  MUX \Inst_Mem/U435  ( .A(inst_mem_in_wire[70]), .B(inst_mem_in_wire[102]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n429 ) );
  MUX \Inst_Mem/U434  ( .A(\Inst_Mem/n427 ), .B(\Inst_Mem/n426 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n428 ) );
  MUX \Inst_Mem/U433  ( .A(inst_mem_in_wire[134]), .B(inst_mem_in_wire[166]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n427 ) );
  MUX \Inst_Mem/U432  ( .A(inst_mem_in_wire[198]), .B(inst_mem_in_wire[230]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n426 ) );
  MUX \Inst_Mem/U431  ( .A(\Inst_Mem/n424 ), .B(\Inst_Mem/n421 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n425 ) );
  MUX \Inst_Mem/U430  ( .A(\Inst_Mem/n423 ), .B(\Inst_Mem/n422 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n424 ) );
  MUX \Inst_Mem/U429  ( .A(inst_mem_in_wire[262]), .B(inst_mem_in_wire[294]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n423 ) );
  MUX \Inst_Mem/U428  ( .A(inst_mem_in_wire[326]), .B(inst_mem_in_wire[358]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n422 ) );
  MUX \Inst_Mem/U427  ( .A(\Inst_Mem/n420 ), .B(\Inst_Mem/n419 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n421 ) );
  MUX \Inst_Mem/U426  ( .A(inst_mem_in_wire[390]), .B(inst_mem_in_wire[422]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n420 ) );
  MUX \Inst_Mem/U425  ( .A(inst_mem_in_wire[454]), .B(inst_mem_in_wire[486]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n419 ) );
  MUX \Inst_Mem/U424  ( .A(\Inst_Mem/n417 ), .B(\Inst_Mem/n410 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n418 ) );
  MUX \Inst_Mem/U423  ( .A(\Inst_Mem/n416 ), .B(\Inst_Mem/n413 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n417 ) );
  MUX \Inst_Mem/U422  ( .A(\Inst_Mem/n415 ), .B(\Inst_Mem/n414 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n416 ) );
  MUX \Inst_Mem/U421  ( .A(inst_mem_in_wire[518]), .B(inst_mem_in_wire[550]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n415 ) );
  MUX \Inst_Mem/U420  ( .A(inst_mem_in_wire[582]), .B(inst_mem_in_wire[614]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n414 ) );
  MUX \Inst_Mem/U419  ( .A(\Inst_Mem/n412 ), .B(\Inst_Mem/n411 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n413 ) );
  MUX \Inst_Mem/U418  ( .A(inst_mem_in_wire[646]), .B(inst_mem_in_wire[678]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n412 ) );
  MUX \Inst_Mem/U417  ( .A(inst_mem_in_wire[710]), .B(inst_mem_in_wire[742]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n411 ) );
  MUX \Inst_Mem/U416  ( .A(\Inst_Mem/n409 ), .B(\Inst_Mem/n406 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n410 ) );
  MUX \Inst_Mem/U415  ( .A(\Inst_Mem/n408 ), .B(\Inst_Mem/n407 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n409 ) );
  MUX \Inst_Mem/U414  ( .A(inst_mem_in_wire[774]), .B(inst_mem_in_wire[806]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n408 ) );
  MUX \Inst_Mem/U413  ( .A(inst_mem_in_wire[838]), .B(inst_mem_in_wire[870]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n407 ) );
  MUX \Inst_Mem/U412  ( .A(\Inst_Mem/n405 ), .B(\Inst_Mem/n404 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n406 ) );
  MUX \Inst_Mem/U411  ( .A(inst_mem_in_wire[902]), .B(inst_mem_in_wire[934]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n405 ) );
  MUX \Inst_Mem/U410  ( .A(inst_mem_in_wire[966]), .B(inst_mem_in_wire[998]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n404 ) );
  MUX \Inst_Mem/U409  ( .A(\Inst_Mem/n402 ), .B(\Inst_Mem/n387 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n403 ) );
  MUX \Inst_Mem/U408  ( .A(\Inst_Mem/n401 ), .B(\Inst_Mem/n394 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n402 ) );
  MUX \Inst_Mem/U407  ( .A(\Inst_Mem/n400 ), .B(\Inst_Mem/n397 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n401 ) );
  MUX \Inst_Mem/U406  ( .A(\Inst_Mem/n399 ), .B(\Inst_Mem/n398 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n400 ) );
  MUX \Inst_Mem/U405  ( .A(inst_mem_in_wire[1030]), .B(inst_mem_in_wire[1062]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n399 ) );
  MUX \Inst_Mem/U404  ( .A(inst_mem_in_wire[1094]), .B(inst_mem_in_wire[1126]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n398 ) );
  MUX \Inst_Mem/U403  ( .A(\Inst_Mem/n396 ), .B(\Inst_Mem/n395 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n397 ) );
  MUX \Inst_Mem/U402  ( .A(inst_mem_in_wire[1158]), .B(inst_mem_in_wire[1190]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n396 ) );
  MUX \Inst_Mem/U401  ( .A(inst_mem_in_wire[1222]), .B(inst_mem_in_wire[1254]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n395 ) );
  MUX \Inst_Mem/U400  ( .A(\Inst_Mem/n393 ), .B(\Inst_Mem/n390 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n394 ) );
  MUX \Inst_Mem/U399  ( .A(\Inst_Mem/n392 ), .B(\Inst_Mem/n391 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n393 ) );
  MUX \Inst_Mem/U398  ( .A(inst_mem_in_wire[1286]), .B(inst_mem_in_wire[1318]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n392 ) );
  MUX \Inst_Mem/U397  ( .A(inst_mem_in_wire[1350]), .B(inst_mem_in_wire[1382]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n391 ) );
  MUX \Inst_Mem/U396  ( .A(\Inst_Mem/n389 ), .B(\Inst_Mem/n388 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n390 ) );
  MUX \Inst_Mem/U395  ( .A(inst_mem_in_wire[1414]), .B(inst_mem_in_wire[1446]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n389 ) );
  MUX \Inst_Mem/U394  ( .A(inst_mem_in_wire[1478]), .B(inst_mem_in_wire[1510]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n388 ) );
  MUX \Inst_Mem/U393  ( .A(\Inst_Mem/n386 ), .B(\Inst_Mem/n379 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n387 ) );
  MUX \Inst_Mem/U392  ( .A(\Inst_Mem/n385 ), .B(\Inst_Mem/n382 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n386 ) );
  MUX \Inst_Mem/U391  ( .A(\Inst_Mem/n384 ), .B(\Inst_Mem/n383 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n385 ) );
  MUX \Inst_Mem/U390  ( .A(inst_mem_in_wire[1542]), .B(inst_mem_in_wire[1574]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n384 ) );
  MUX \Inst_Mem/U389  ( .A(inst_mem_in_wire[1606]), .B(inst_mem_in_wire[1638]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n383 ) );
  MUX \Inst_Mem/U388  ( .A(\Inst_Mem/n381 ), .B(\Inst_Mem/n380 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n382 ) );
  MUX \Inst_Mem/U387  ( .A(inst_mem_in_wire[1670]), .B(inst_mem_in_wire[1702]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n381 ) );
  MUX \Inst_Mem/U386  ( .A(inst_mem_in_wire[1734]), .B(inst_mem_in_wire[1766]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n380 ) );
  MUX \Inst_Mem/U385  ( .A(\Inst_Mem/n378 ), .B(\Inst_Mem/n375 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n379 ) );
  MUX \Inst_Mem/U384  ( .A(\Inst_Mem/n377 ), .B(\Inst_Mem/n376 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n378 ) );
  MUX \Inst_Mem/U383  ( .A(inst_mem_in_wire[1798]), .B(inst_mem_in_wire[1830]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n377 ) );
  MUX \Inst_Mem/U382  ( .A(inst_mem_in_wire[1862]), .B(inst_mem_in_wire[1894]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n376 ) );
  MUX \Inst_Mem/U381  ( .A(\Inst_Mem/n374 ), .B(\Inst_Mem/n373 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n375 ) );
  MUX \Inst_Mem/U380  ( .A(inst_mem_in_wire[1926]), .B(inst_mem_in_wire[1958]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n374 ) );
  MUX \Inst_Mem/U379  ( .A(inst_mem_in_wire[1990]), .B(inst_mem_in_wire[2022]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n373 ) );
  MUX \Inst_Mem/U378  ( .A(\Inst_Mem/n372 ), .B(\Inst_Mem/n341 ), .S(
        pc_current[7]), .Z(imm[5]) );
  MUX \Inst_Mem/U377  ( .A(\Inst_Mem/n371 ), .B(\Inst_Mem/n356 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n372 ) );
  MUX \Inst_Mem/U376  ( .A(\Inst_Mem/n370 ), .B(\Inst_Mem/n363 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n371 ) );
  MUX \Inst_Mem/U375  ( .A(\Inst_Mem/n369 ), .B(\Inst_Mem/n366 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n370 ) );
  MUX \Inst_Mem/U374  ( .A(\Inst_Mem/n368 ), .B(\Inst_Mem/n367 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n369 ) );
  MUX \Inst_Mem/U373  ( .A(inst_mem_in_wire[5]), .B(inst_mem_in_wire[37]), .S(
        pc_current[2]), .Z(\Inst_Mem/n368 ) );
  MUX \Inst_Mem/U372  ( .A(inst_mem_in_wire[69]), .B(inst_mem_in_wire[101]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n367 ) );
  MUX \Inst_Mem/U371  ( .A(\Inst_Mem/n365 ), .B(\Inst_Mem/n364 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n366 ) );
  MUX \Inst_Mem/U370  ( .A(inst_mem_in_wire[133]), .B(inst_mem_in_wire[165]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n365 ) );
  MUX \Inst_Mem/U369  ( .A(inst_mem_in_wire[197]), .B(inst_mem_in_wire[229]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n364 ) );
  MUX \Inst_Mem/U368  ( .A(\Inst_Mem/n362 ), .B(\Inst_Mem/n359 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n363 ) );
  MUX \Inst_Mem/U367  ( .A(\Inst_Mem/n361 ), .B(\Inst_Mem/n360 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n362 ) );
  MUX \Inst_Mem/U366  ( .A(inst_mem_in_wire[261]), .B(inst_mem_in_wire[293]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n361 ) );
  MUX \Inst_Mem/U365  ( .A(inst_mem_in_wire[325]), .B(inst_mem_in_wire[357]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n360 ) );
  MUX \Inst_Mem/U364  ( .A(\Inst_Mem/n358 ), .B(\Inst_Mem/n357 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n359 ) );
  MUX \Inst_Mem/U363  ( .A(inst_mem_in_wire[389]), .B(inst_mem_in_wire[421]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n358 ) );
  MUX \Inst_Mem/U362  ( .A(inst_mem_in_wire[453]), .B(inst_mem_in_wire[485]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n357 ) );
  MUX \Inst_Mem/U361  ( .A(\Inst_Mem/n355 ), .B(\Inst_Mem/n348 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n356 ) );
  MUX \Inst_Mem/U360  ( .A(\Inst_Mem/n354 ), .B(\Inst_Mem/n351 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n355 ) );
  MUX \Inst_Mem/U359  ( .A(\Inst_Mem/n353 ), .B(\Inst_Mem/n352 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n354 ) );
  MUX \Inst_Mem/U358  ( .A(inst_mem_in_wire[517]), .B(inst_mem_in_wire[549]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n353 ) );
  MUX \Inst_Mem/U357  ( .A(inst_mem_in_wire[581]), .B(inst_mem_in_wire[613]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n352 ) );
  MUX \Inst_Mem/U356  ( .A(\Inst_Mem/n350 ), .B(\Inst_Mem/n349 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n351 ) );
  MUX \Inst_Mem/U355  ( .A(inst_mem_in_wire[645]), .B(inst_mem_in_wire[677]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n350 ) );
  MUX \Inst_Mem/U354  ( .A(inst_mem_in_wire[709]), .B(inst_mem_in_wire[741]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n349 ) );
  MUX \Inst_Mem/U353  ( .A(\Inst_Mem/n347 ), .B(\Inst_Mem/n344 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n348 ) );
  MUX \Inst_Mem/U352  ( .A(\Inst_Mem/n346 ), .B(\Inst_Mem/n345 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n347 ) );
  MUX \Inst_Mem/U351  ( .A(inst_mem_in_wire[773]), .B(inst_mem_in_wire[805]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n346 ) );
  MUX \Inst_Mem/U350  ( .A(inst_mem_in_wire[837]), .B(inst_mem_in_wire[869]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n345 ) );
  MUX \Inst_Mem/U349  ( .A(\Inst_Mem/n343 ), .B(\Inst_Mem/n342 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n344 ) );
  MUX \Inst_Mem/U348  ( .A(inst_mem_in_wire[901]), .B(inst_mem_in_wire[933]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n343 ) );
  MUX \Inst_Mem/U347  ( .A(inst_mem_in_wire[965]), .B(inst_mem_in_wire[997]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n342 ) );
  MUX \Inst_Mem/U346  ( .A(\Inst_Mem/n340 ), .B(\Inst_Mem/n325 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n341 ) );
  MUX \Inst_Mem/U345  ( .A(\Inst_Mem/n339 ), .B(\Inst_Mem/n332 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n340 ) );
  MUX \Inst_Mem/U344  ( .A(\Inst_Mem/n338 ), .B(\Inst_Mem/n335 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n339 ) );
  MUX \Inst_Mem/U343  ( .A(\Inst_Mem/n337 ), .B(\Inst_Mem/n336 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n338 ) );
  MUX \Inst_Mem/U342  ( .A(inst_mem_in_wire[1029]), .B(inst_mem_in_wire[1061]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n337 ) );
  MUX \Inst_Mem/U341  ( .A(inst_mem_in_wire[1093]), .B(inst_mem_in_wire[1125]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n336 ) );
  MUX \Inst_Mem/U340  ( .A(\Inst_Mem/n334 ), .B(\Inst_Mem/n333 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n335 ) );
  MUX \Inst_Mem/U339  ( .A(inst_mem_in_wire[1157]), .B(inst_mem_in_wire[1189]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n334 ) );
  MUX \Inst_Mem/U338  ( .A(inst_mem_in_wire[1221]), .B(inst_mem_in_wire[1253]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n333 ) );
  MUX \Inst_Mem/U337  ( .A(\Inst_Mem/n331 ), .B(\Inst_Mem/n328 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n332 ) );
  MUX \Inst_Mem/U336  ( .A(\Inst_Mem/n330 ), .B(\Inst_Mem/n329 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n331 ) );
  MUX \Inst_Mem/U335  ( .A(inst_mem_in_wire[1285]), .B(inst_mem_in_wire[1317]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n330 ) );
  MUX \Inst_Mem/U334  ( .A(inst_mem_in_wire[1349]), .B(inst_mem_in_wire[1381]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n329 ) );
  MUX \Inst_Mem/U333  ( .A(\Inst_Mem/n327 ), .B(\Inst_Mem/n326 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n328 ) );
  MUX \Inst_Mem/U332  ( .A(inst_mem_in_wire[1413]), .B(inst_mem_in_wire[1445]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n327 ) );
  MUX \Inst_Mem/U331  ( .A(inst_mem_in_wire[1477]), .B(inst_mem_in_wire[1509]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n326 ) );
  MUX \Inst_Mem/U330  ( .A(\Inst_Mem/n324 ), .B(\Inst_Mem/n317 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n325 ) );
  MUX \Inst_Mem/U329  ( .A(\Inst_Mem/n323 ), .B(\Inst_Mem/n320 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n324 ) );
  MUX \Inst_Mem/U328  ( .A(\Inst_Mem/n322 ), .B(\Inst_Mem/n321 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n323 ) );
  MUX \Inst_Mem/U327  ( .A(inst_mem_in_wire[1541]), .B(inst_mem_in_wire[1573]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n322 ) );
  MUX \Inst_Mem/U326  ( .A(inst_mem_in_wire[1605]), .B(inst_mem_in_wire[1637]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n321 ) );
  MUX \Inst_Mem/U325  ( .A(\Inst_Mem/n319 ), .B(\Inst_Mem/n318 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n320 ) );
  MUX \Inst_Mem/U324  ( .A(inst_mem_in_wire[1669]), .B(inst_mem_in_wire[1701]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n319 ) );
  MUX \Inst_Mem/U323  ( .A(inst_mem_in_wire[1733]), .B(inst_mem_in_wire[1765]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n318 ) );
  MUX \Inst_Mem/U322  ( .A(\Inst_Mem/n316 ), .B(\Inst_Mem/n313 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n317 ) );
  MUX \Inst_Mem/U321  ( .A(\Inst_Mem/n315 ), .B(\Inst_Mem/n314 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n316 ) );
  MUX \Inst_Mem/U320  ( .A(inst_mem_in_wire[1797]), .B(inst_mem_in_wire[1829]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n315 ) );
  MUX \Inst_Mem/U319  ( .A(inst_mem_in_wire[1861]), .B(inst_mem_in_wire[1893]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n314 ) );
  MUX \Inst_Mem/U318  ( .A(\Inst_Mem/n312 ), .B(\Inst_Mem/n311 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n313 ) );
  MUX \Inst_Mem/U317  ( .A(inst_mem_in_wire[1925]), .B(inst_mem_in_wire[1957]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n312 ) );
  MUX \Inst_Mem/U316  ( .A(inst_mem_in_wire[1989]), .B(inst_mem_in_wire[2021]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n311 ) );
  MUX \Inst_Mem/U315  ( .A(\Inst_Mem/n310 ), .B(\Inst_Mem/n279 ), .S(
        pc_current[7]), .Z(imm[4]) );
  MUX \Inst_Mem/U314  ( .A(\Inst_Mem/n309 ), .B(\Inst_Mem/n294 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n310 ) );
  MUX \Inst_Mem/U313  ( .A(\Inst_Mem/n308 ), .B(\Inst_Mem/n301 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n309 ) );
  MUX \Inst_Mem/U312  ( .A(\Inst_Mem/n307 ), .B(\Inst_Mem/n304 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n308 ) );
  MUX \Inst_Mem/U311  ( .A(\Inst_Mem/n306 ), .B(\Inst_Mem/n305 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n307 ) );
  MUX \Inst_Mem/U310  ( .A(inst_mem_in_wire[4]), .B(inst_mem_in_wire[36]), .S(
        pc_current[2]), .Z(\Inst_Mem/n306 ) );
  MUX \Inst_Mem/U309  ( .A(inst_mem_in_wire[68]), .B(inst_mem_in_wire[100]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n305 ) );
  MUX \Inst_Mem/U308  ( .A(\Inst_Mem/n303 ), .B(\Inst_Mem/n302 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n304 ) );
  MUX \Inst_Mem/U307  ( .A(inst_mem_in_wire[132]), .B(inst_mem_in_wire[164]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n303 ) );
  MUX \Inst_Mem/U306  ( .A(inst_mem_in_wire[196]), .B(inst_mem_in_wire[228]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n302 ) );
  MUX \Inst_Mem/U305  ( .A(\Inst_Mem/n300 ), .B(\Inst_Mem/n297 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n301 ) );
  MUX \Inst_Mem/U304  ( .A(\Inst_Mem/n299 ), .B(\Inst_Mem/n298 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n300 ) );
  MUX \Inst_Mem/U303  ( .A(inst_mem_in_wire[260]), .B(inst_mem_in_wire[292]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n299 ) );
  MUX \Inst_Mem/U302  ( .A(inst_mem_in_wire[324]), .B(inst_mem_in_wire[356]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n298 ) );
  MUX \Inst_Mem/U301  ( .A(\Inst_Mem/n296 ), .B(\Inst_Mem/n295 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n297 ) );
  MUX \Inst_Mem/U300  ( .A(inst_mem_in_wire[388]), .B(inst_mem_in_wire[420]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n296 ) );
  MUX \Inst_Mem/U299  ( .A(inst_mem_in_wire[452]), .B(inst_mem_in_wire[484]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n295 ) );
  MUX \Inst_Mem/U298  ( .A(\Inst_Mem/n293 ), .B(\Inst_Mem/n286 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n294 ) );
  MUX \Inst_Mem/U297  ( .A(\Inst_Mem/n292 ), .B(\Inst_Mem/n289 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n293 ) );
  MUX \Inst_Mem/U296  ( .A(\Inst_Mem/n291 ), .B(\Inst_Mem/n290 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n292 ) );
  MUX \Inst_Mem/U295  ( .A(inst_mem_in_wire[516]), .B(inst_mem_in_wire[548]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n291 ) );
  MUX \Inst_Mem/U294  ( .A(inst_mem_in_wire[580]), .B(inst_mem_in_wire[612]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n290 ) );
  MUX \Inst_Mem/U293  ( .A(\Inst_Mem/n288 ), .B(\Inst_Mem/n287 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n289 ) );
  MUX \Inst_Mem/U292  ( .A(inst_mem_in_wire[644]), .B(inst_mem_in_wire[676]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n288 ) );
  MUX \Inst_Mem/U291  ( .A(inst_mem_in_wire[708]), .B(inst_mem_in_wire[740]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n287 ) );
  MUX \Inst_Mem/U290  ( .A(\Inst_Mem/n285 ), .B(\Inst_Mem/n282 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n286 ) );
  MUX \Inst_Mem/U289  ( .A(\Inst_Mem/n284 ), .B(\Inst_Mem/n283 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n285 ) );
  MUX \Inst_Mem/U288  ( .A(inst_mem_in_wire[772]), .B(inst_mem_in_wire[804]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n284 ) );
  MUX \Inst_Mem/U287  ( .A(inst_mem_in_wire[836]), .B(inst_mem_in_wire[868]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n283 ) );
  MUX \Inst_Mem/U286  ( .A(\Inst_Mem/n281 ), .B(\Inst_Mem/n280 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n282 ) );
  MUX \Inst_Mem/U285  ( .A(inst_mem_in_wire[900]), .B(inst_mem_in_wire[932]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n281 ) );
  MUX \Inst_Mem/U284  ( .A(inst_mem_in_wire[964]), .B(inst_mem_in_wire[996]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n280 ) );
  MUX \Inst_Mem/U283  ( .A(\Inst_Mem/n278 ), .B(\Inst_Mem/n263 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n279 ) );
  MUX \Inst_Mem/U282  ( .A(\Inst_Mem/n277 ), .B(\Inst_Mem/n270 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n278 ) );
  MUX \Inst_Mem/U281  ( .A(\Inst_Mem/n276 ), .B(\Inst_Mem/n273 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n277 ) );
  MUX \Inst_Mem/U280  ( .A(\Inst_Mem/n275 ), .B(\Inst_Mem/n274 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n276 ) );
  MUX \Inst_Mem/U279  ( .A(inst_mem_in_wire[1028]), .B(inst_mem_in_wire[1060]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n275 ) );
  MUX \Inst_Mem/U278  ( .A(inst_mem_in_wire[1092]), .B(inst_mem_in_wire[1124]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n274 ) );
  MUX \Inst_Mem/U277  ( .A(\Inst_Mem/n272 ), .B(\Inst_Mem/n271 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n273 ) );
  MUX \Inst_Mem/U276  ( .A(inst_mem_in_wire[1156]), .B(inst_mem_in_wire[1188]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n272 ) );
  MUX \Inst_Mem/U275  ( .A(inst_mem_in_wire[1220]), .B(inst_mem_in_wire[1252]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n271 ) );
  MUX \Inst_Mem/U274  ( .A(\Inst_Mem/n269 ), .B(\Inst_Mem/n266 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n270 ) );
  MUX \Inst_Mem/U273  ( .A(\Inst_Mem/n268 ), .B(\Inst_Mem/n267 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n269 ) );
  MUX \Inst_Mem/U272  ( .A(inst_mem_in_wire[1284]), .B(inst_mem_in_wire[1316]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n268 ) );
  MUX \Inst_Mem/U271  ( .A(inst_mem_in_wire[1348]), .B(inst_mem_in_wire[1380]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n267 ) );
  MUX \Inst_Mem/U270  ( .A(\Inst_Mem/n265 ), .B(\Inst_Mem/n264 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n266 ) );
  MUX \Inst_Mem/U269  ( .A(inst_mem_in_wire[1412]), .B(inst_mem_in_wire[1444]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n265 ) );
  MUX \Inst_Mem/U268  ( .A(inst_mem_in_wire[1476]), .B(inst_mem_in_wire[1508]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n264 ) );
  MUX \Inst_Mem/U267  ( .A(\Inst_Mem/n262 ), .B(\Inst_Mem/n255 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n263 ) );
  MUX \Inst_Mem/U266  ( .A(\Inst_Mem/n261 ), .B(\Inst_Mem/n258 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n262 ) );
  MUX \Inst_Mem/U265  ( .A(\Inst_Mem/n260 ), .B(\Inst_Mem/n259 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n261 ) );
  MUX \Inst_Mem/U264  ( .A(inst_mem_in_wire[1540]), .B(inst_mem_in_wire[1572]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n260 ) );
  MUX \Inst_Mem/U263  ( .A(inst_mem_in_wire[1604]), .B(inst_mem_in_wire[1636]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n259 ) );
  MUX \Inst_Mem/U262  ( .A(\Inst_Mem/n257 ), .B(\Inst_Mem/n256 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n258 ) );
  MUX \Inst_Mem/U261  ( .A(inst_mem_in_wire[1668]), .B(inst_mem_in_wire[1700]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n257 ) );
  MUX \Inst_Mem/U260  ( .A(inst_mem_in_wire[1732]), .B(inst_mem_in_wire[1764]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n256 ) );
  MUX \Inst_Mem/U259  ( .A(\Inst_Mem/n254 ), .B(\Inst_Mem/n251 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n255 ) );
  MUX \Inst_Mem/U258  ( .A(\Inst_Mem/n253 ), .B(\Inst_Mem/n252 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n254 ) );
  MUX \Inst_Mem/U257  ( .A(inst_mem_in_wire[1796]), .B(inst_mem_in_wire[1828]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n253 ) );
  MUX \Inst_Mem/U256  ( .A(inst_mem_in_wire[1860]), .B(inst_mem_in_wire[1892]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n252 ) );
  MUX \Inst_Mem/U255  ( .A(\Inst_Mem/n250 ), .B(\Inst_Mem/n249 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n251 ) );
  MUX \Inst_Mem/U254  ( .A(inst_mem_in_wire[1924]), .B(inst_mem_in_wire[1956]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n250 ) );
  MUX \Inst_Mem/U253  ( .A(inst_mem_in_wire[1988]), .B(inst_mem_in_wire[2020]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n249 ) );
  MUX \Inst_Mem/U252  ( .A(\Inst_Mem/n248 ), .B(\Inst_Mem/n217 ), .S(
        pc_current[7]), .Z(imm[3]) );
  MUX \Inst_Mem/U251  ( .A(\Inst_Mem/n247 ), .B(\Inst_Mem/n232 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n248 ) );
  MUX \Inst_Mem/U250  ( .A(\Inst_Mem/n246 ), .B(\Inst_Mem/n239 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n247 ) );
  MUX \Inst_Mem/U249  ( .A(\Inst_Mem/n245 ), .B(\Inst_Mem/n242 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n246 ) );
  MUX \Inst_Mem/U248  ( .A(\Inst_Mem/n244 ), .B(\Inst_Mem/n243 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n245 ) );
  MUX \Inst_Mem/U247  ( .A(inst_mem_in_wire[3]), .B(inst_mem_in_wire[35]), .S(
        pc_current[2]), .Z(\Inst_Mem/n244 ) );
  MUX \Inst_Mem/U246  ( .A(inst_mem_in_wire[67]), .B(inst_mem_in_wire[99]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n243 ) );
  MUX \Inst_Mem/U245  ( .A(\Inst_Mem/n241 ), .B(\Inst_Mem/n240 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n242 ) );
  MUX \Inst_Mem/U244  ( .A(inst_mem_in_wire[131]), .B(inst_mem_in_wire[163]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n241 ) );
  MUX \Inst_Mem/U243  ( .A(inst_mem_in_wire[195]), .B(inst_mem_in_wire[227]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n240 ) );
  MUX \Inst_Mem/U242  ( .A(\Inst_Mem/n238 ), .B(\Inst_Mem/n235 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n239 ) );
  MUX \Inst_Mem/U241  ( .A(\Inst_Mem/n237 ), .B(\Inst_Mem/n236 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n238 ) );
  MUX \Inst_Mem/U240  ( .A(inst_mem_in_wire[259]), .B(inst_mem_in_wire[291]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n237 ) );
  MUX \Inst_Mem/U239  ( .A(inst_mem_in_wire[323]), .B(inst_mem_in_wire[355]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n236 ) );
  MUX \Inst_Mem/U238  ( .A(\Inst_Mem/n234 ), .B(\Inst_Mem/n233 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n235 ) );
  MUX \Inst_Mem/U237  ( .A(inst_mem_in_wire[387]), .B(inst_mem_in_wire[419]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n234 ) );
  MUX \Inst_Mem/U236  ( .A(inst_mem_in_wire[451]), .B(inst_mem_in_wire[483]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n233 ) );
  MUX \Inst_Mem/U235  ( .A(\Inst_Mem/n231 ), .B(\Inst_Mem/n224 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n232 ) );
  MUX \Inst_Mem/U234  ( .A(\Inst_Mem/n230 ), .B(\Inst_Mem/n227 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n231 ) );
  MUX \Inst_Mem/U233  ( .A(\Inst_Mem/n229 ), .B(\Inst_Mem/n228 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n230 ) );
  MUX \Inst_Mem/U232  ( .A(inst_mem_in_wire[515]), .B(inst_mem_in_wire[547]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n229 ) );
  MUX \Inst_Mem/U231  ( .A(inst_mem_in_wire[579]), .B(inst_mem_in_wire[611]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n228 ) );
  MUX \Inst_Mem/U230  ( .A(\Inst_Mem/n226 ), .B(\Inst_Mem/n225 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n227 ) );
  MUX \Inst_Mem/U229  ( .A(inst_mem_in_wire[643]), .B(inst_mem_in_wire[675]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n226 ) );
  MUX \Inst_Mem/U228  ( .A(inst_mem_in_wire[707]), .B(inst_mem_in_wire[739]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n225 ) );
  MUX \Inst_Mem/U227  ( .A(\Inst_Mem/n223 ), .B(\Inst_Mem/n220 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n224 ) );
  MUX \Inst_Mem/U226  ( .A(\Inst_Mem/n222 ), .B(\Inst_Mem/n221 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n223 ) );
  MUX \Inst_Mem/U225  ( .A(inst_mem_in_wire[771]), .B(inst_mem_in_wire[803]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n222 ) );
  MUX \Inst_Mem/U224  ( .A(inst_mem_in_wire[835]), .B(inst_mem_in_wire[867]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n221 ) );
  MUX \Inst_Mem/U223  ( .A(\Inst_Mem/n219 ), .B(\Inst_Mem/n218 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n220 ) );
  MUX \Inst_Mem/U222  ( .A(inst_mem_in_wire[899]), .B(inst_mem_in_wire[931]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n219 ) );
  MUX \Inst_Mem/U221  ( .A(inst_mem_in_wire[963]), .B(inst_mem_in_wire[995]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n218 ) );
  MUX \Inst_Mem/U220  ( .A(\Inst_Mem/n216 ), .B(\Inst_Mem/n201 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n217 ) );
  MUX \Inst_Mem/U219  ( .A(\Inst_Mem/n215 ), .B(\Inst_Mem/n208 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n216 ) );
  MUX \Inst_Mem/U218  ( .A(\Inst_Mem/n214 ), .B(\Inst_Mem/n211 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n215 ) );
  MUX \Inst_Mem/U217  ( .A(\Inst_Mem/n213 ), .B(\Inst_Mem/n212 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n214 ) );
  MUX \Inst_Mem/U216  ( .A(inst_mem_in_wire[1027]), .B(inst_mem_in_wire[1059]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n213 ) );
  MUX \Inst_Mem/U215  ( .A(inst_mem_in_wire[1091]), .B(inst_mem_in_wire[1123]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n212 ) );
  MUX \Inst_Mem/U214  ( .A(\Inst_Mem/n210 ), .B(\Inst_Mem/n209 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n211 ) );
  MUX \Inst_Mem/U213  ( .A(inst_mem_in_wire[1155]), .B(inst_mem_in_wire[1187]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n210 ) );
  MUX \Inst_Mem/U212  ( .A(inst_mem_in_wire[1219]), .B(inst_mem_in_wire[1251]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n209 ) );
  MUX \Inst_Mem/U211  ( .A(\Inst_Mem/n207 ), .B(\Inst_Mem/n204 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n208 ) );
  MUX \Inst_Mem/U210  ( .A(\Inst_Mem/n206 ), .B(\Inst_Mem/n205 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n207 ) );
  MUX \Inst_Mem/U209  ( .A(inst_mem_in_wire[1283]), .B(inst_mem_in_wire[1315]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n206 ) );
  MUX \Inst_Mem/U208  ( .A(inst_mem_in_wire[1347]), .B(inst_mem_in_wire[1379]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n205 ) );
  MUX \Inst_Mem/U207  ( .A(\Inst_Mem/n203 ), .B(\Inst_Mem/n202 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n204 ) );
  MUX \Inst_Mem/U206  ( .A(inst_mem_in_wire[1411]), .B(inst_mem_in_wire[1443]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n203 ) );
  MUX \Inst_Mem/U205  ( .A(inst_mem_in_wire[1475]), .B(inst_mem_in_wire[1507]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n202 ) );
  MUX \Inst_Mem/U204  ( .A(\Inst_Mem/n200 ), .B(\Inst_Mem/n193 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n201 ) );
  MUX \Inst_Mem/U203  ( .A(\Inst_Mem/n199 ), .B(\Inst_Mem/n196 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n200 ) );
  MUX \Inst_Mem/U202  ( .A(\Inst_Mem/n198 ), .B(\Inst_Mem/n197 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n199 ) );
  MUX \Inst_Mem/U201  ( .A(inst_mem_in_wire[1539]), .B(inst_mem_in_wire[1571]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n198 ) );
  MUX \Inst_Mem/U200  ( .A(inst_mem_in_wire[1603]), .B(inst_mem_in_wire[1635]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n197 ) );
  MUX \Inst_Mem/U199  ( .A(\Inst_Mem/n195 ), .B(\Inst_Mem/n194 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n196 ) );
  MUX \Inst_Mem/U198  ( .A(inst_mem_in_wire[1667]), .B(inst_mem_in_wire[1699]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n195 ) );
  MUX \Inst_Mem/U197  ( .A(inst_mem_in_wire[1731]), .B(inst_mem_in_wire[1763]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n194 ) );
  MUX \Inst_Mem/U196  ( .A(\Inst_Mem/n192 ), .B(\Inst_Mem/n189 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n193 ) );
  MUX \Inst_Mem/U195  ( .A(\Inst_Mem/n191 ), .B(\Inst_Mem/n190 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n192 ) );
  MUX \Inst_Mem/U194  ( .A(inst_mem_in_wire[1795]), .B(inst_mem_in_wire[1827]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n191 ) );
  MUX \Inst_Mem/U193  ( .A(inst_mem_in_wire[1859]), .B(inst_mem_in_wire[1891]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n190 ) );
  MUX \Inst_Mem/U192  ( .A(\Inst_Mem/n188 ), .B(\Inst_Mem/n187 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n189 ) );
  MUX \Inst_Mem/U191  ( .A(inst_mem_in_wire[1923]), .B(inst_mem_in_wire[1955]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n188 ) );
  MUX \Inst_Mem/U190  ( .A(inst_mem_in_wire[1987]), .B(inst_mem_in_wire[2019]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n187 ) );
  MUX \Inst_Mem/U189  ( .A(\Inst_Mem/n186 ), .B(\Inst_Mem/n155 ), .S(
        pc_current[7]), .Z(imm[2]) );
  MUX \Inst_Mem/U188  ( .A(\Inst_Mem/n185 ), .B(\Inst_Mem/n170 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n186 ) );
  MUX \Inst_Mem/U187  ( .A(\Inst_Mem/n184 ), .B(\Inst_Mem/n177 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n185 ) );
  MUX \Inst_Mem/U186  ( .A(\Inst_Mem/n183 ), .B(\Inst_Mem/n180 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n184 ) );
  MUX \Inst_Mem/U185  ( .A(\Inst_Mem/n182 ), .B(\Inst_Mem/n181 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n183 ) );
  MUX \Inst_Mem/U184  ( .A(inst_mem_in_wire[2]), .B(inst_mem_in_wire[34]), .S(
        pc_current[2]), .Z(\Inst_Mem/n182 ) );
  MUX \Inst_Mem/U183  ( .A(inst_mem_in_wire[66]), .B(inst_mem_in_wire[98]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n181 ) );
  MUX \Inst_Mem/U182  ( .A(\Inst_Mem/n179 ), .B(\Inst_Mem/n178 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n180 ) );
  MUX \Inst_Mem/U181  ( .A(inst_mem_in_wire[130]), .B(inst_mem_in_wire[162]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n179 ) );
  MUX \Inst_Mem/U180  ( .A(inst_mem_in_wire[194]), .B(inst_mem_in_wire[226]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n178 ) );
  MUX \Inst_Mem/U179  ( .A(\Inst_Mem/n176 ), .B(\Inst_Mem/n173 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n177 ) );
  MUX \Inst_Mem/U178  ( .A(\Inst_Mem/n175 ), .B(\Inst_Mem/n174 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n176 ) );
  MUX \Inst_Mem/U177  ( .A(inst_mem_in_wire[258]), .B(inst_mem_in_wire[290]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n175 ) );
  MUX \Inst_Mem/U176  ( .A(inst_mem_in_wire[322]), .B(inst_mem_in_wire[354]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n174 ) );
  MUX \Inst_Mem/U175  ( .A(\Inst_Mem/n172 ), .B(\Inst_Mem/n171 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n173 ) );
  MUX \Inst_Mem/U174  ( .A(inst_mem_in_wire[386]), .B(inst_mem_in_wire[418]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n172 ) );
  MUX \Inst_Mem/U173  ( .A(inst_mem_in_wire[450]), .B(inst_mem_in_wire[482]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n171 ) );
  MUX \Inst_Mem/U172  ( .A(\Inst_Mem/n169 ), .B(\Inst_Mem/n162 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n170 ) );
  MUX \Inst_Mem/U171  ( .A(\Inst_Mem/n168 ), .B(\Inst_Mem/n165 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n169 ) );
  MUX \Inst_Mem/U170  ( .A(\Inst_Mem/n167 ), .B(\Inst_Mem/n166 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n168 ) );
  MUX \Inst_Mem/U169  ( .A(inst_mem_in_wire[514]), .B(inst_mem_in_wire[546]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n167 ) );
  MUX \Inst_Mem/U168  ( .A(inst_mem_in_wire[578]), .B(inst_mem_in_wire[610]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n166 ) );
  MUX \Inst_Mem/U167  ( .A(\Inst_Mem/n164 ), .B(\Inst_Mem/n163 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n165 ) );
  MUX \Inst_Mem/U166  ( .A(inst_mem_in_wire[642]), .B(inst_mem_in_wire[674]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n164 ) );
  MUX \Inst_Mem/U165  ( .A(inst_mem_in_wire[706]), .B(inst_mem_in_wire[738]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n163 ) );
  MUX \Inst_Mem/U164  ( .A(\Inst_Mem/n161 ), .B(\Inst_Mem/n158 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n162 ) );
  MUX \Inst_Mem/U163  ( .A(\Inst_Mem/n160 ), .B(\Inst_Mem/n159 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n161 ) );
  MUX \Inst_Mem/U162  ( .A(inst_mem_in_wire[770]), .B(inst_mem_in_wire[802]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n160 ) );
  MUX \Inst_Mem/U161  ( .A(inst_mem_in_wire[834]), .B(inst_mem_in_wire[866]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n159 ) );
  MUX \Inst_Mem/U160  ( .A(\Inst_Mem/n157 ), .B(\Inst_Mem/n156 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n158 ) );
  MUX \Inst_Mem/U159  ( .A(inst_mem_in_wire[898]), .B(inst_mem_in_wire[930]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n157 ) );
  MUX \Inst_Mem/U158  ( .A(inst_mem_in_wire[962]), .B(inst_mem_in_wire[994]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n156 ) );
  MUX \Inst_Mem/U157  ( .A(\Inst_Mem/n154 ), .B(\Inst_Mem/n139 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n155 ) );
  MUX \Inst_Mem/U156  ( .A(\Inst_Mem/n153 ), .B(\Inst_Mem/n146 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n154 ) );
  MUX \Inst_Mem/U155  ( .A(\Inst_Mem/n152 ), .B(\Inst_Mem/n149 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n153 ) );
  MUX \Inst_Mem/U154  ( .A(\Inst_Mem/n151 ), .B(\Inst_Mem/n150 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n152 ) );
  MUX \Inst_Mem/U153  ( .A(inst_mem_in_wire[1026]), .B(inst_mem_in_wire[1058]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n151 ) );
  MUX \Inst_Mem/U152  ( .A(inst_mem_in_wire[1090]), .B(inst_mem_in_wire[1122]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n150 ) );
  MUX \Inst_Mem/U151  ( .A(\Inst_Mem/n148 ), .B(\Inst_Mem/n147 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n149 ) );
  MUX \Inst_Mem/U150  ( .A(inst_mem_in_wire[1154]), .B(inst_mem_in_wire[1186]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n148 ) );
  MUX \Inst_Mem/U149  ( .A(inst_mem_in_wire[1218]), .B(inst_mem_in_wire[1250]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n147 ) );
  MUX \Inst_Mem/U148  ( .A(\Inst_Mem/n145 ), .B(\Inst_Mem/n142 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n146 ) );
  MUX \Inst_Mem/U147  ( .A(\Inst_Mem/n144 ), .B(\Inst_Mem/n143 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n145 ) );
  MUX \Inst_Mem/U146  ( .A(inst_mem_in_wire[1282]), .B(inst_mem_in_wire[1314]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n144 ) );
  MUX \Inst_Mem/U145  ( .A(inst_mem_in_wire[1346]), .B(inst_mem_in_wire[1378]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n143 ) );
  MUX \Inst_Mem/U144  ( .A(\Inst_Mem/n141 ), .B(\Inst_Mem/n140 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n142 ) );
  MUX \Inst_Mem/U143  ( .A(inst_mem_in_wire[1410]), .B(inst_mem_in_wire[1442]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n141 ) );
  MUX \Inst_Mem/U142  ( .A(inst_mem_in_wire[1474]), .B(inst_mem_in_wire[1506]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n140 ) );
  MUX \Inst_Mem/U141  ( .A(\Inst_Mem/n138 ), .B(\Inst_Mem/n131 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n139 ) );
  MUX \Inst_Mem/U140  ( .A(\Inst_Mem/n137 ), .B(\Inst_Mem/n134 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n138 ) );
  MUX \Inst_Mem/U139  ( .A(\Inst_Mem/n136 ), .B(\Inst_Mem/n135 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n137 ) );
  MUX \Inst_Mem/U138  ( .A(inst_mem_in_wire[1538]), .B(inst_mem_in_wire[1570]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n136 ) );
  MUX \Inst_Mem/U137  ( .A(inst_mem_in_wire[1602]), .B(inst_mem_in_wire[1634]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n135 ) );
  MUX \Inst_Mem/U136  ( .A(\Inst_Mem/n133 ), .B(\Inst_Mem/n132 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n134 ) );
  MUX \Inst_Mem/U135  ( .A(inst_mem_in_wire[1666]), .B(inst_mem_in_wire[1698]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n133 ) );
  MUX \Inst_Mem/U134  ( .A(inst_mem_in_wire[1730]), .B(inst_mem_in_wire[1762]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n132 ) );
  MUX \Inst_Mem/U133  ( .A(\Inst_Mem/n130 ), .B(\Inst_Mem/n127 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n131 ) );
  MUX \Inst_Mem/U132  ( .A(\Inst_Mem/n129 ), .B(\Inst_Mem/n128 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n130 ) );
  MUX \Inst_Mem/U131  ( .A(inst_mem_in_wire[1794]), .B(inst_mem_in_wire[1826]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n129 ) );
  MUX \Inst_Mem/U130  ( .A(inst_mem_in_wire[1858]), .B(inst_mem_in_wire[1890]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n128 ) );
  MUX \Inst_Mem/U129  ( .A(\Inst_Mem/n126 ), .B(\Inst_Mem/n125 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n127 ) );
  MUX \Inst_Mem/U128  ( .A(inst_mem_in_wire[1922]), .B(inst_mem_in_wire[1954]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n126 ) );
  MUX \Inst_Mem/U127  ( .A(inst_mem_in_wire[1986]), .B(inst_mem_in_wire[2018]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n125 ) );
  MUX \Inst_Mem/U126  ( .A(\Inst_Mem/n124 ), .B(\Inst_Mem/n93 ), .S(
        pc_current[7]), .Z(imm[1]) );
  MUX \Inst_Mem/U125  ( .A(\Inst_Mem/n123 ), .B(\Inst_Mem/n108 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n124 ) );
  MUX \Inst_Mem/U124  ( .A(\Inst_Mem/n122 ), .B(\Inst_Mem/n115 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n123 ) );
  MUX \Inst_Mem/U123  ( .A(\Inst_Mem/n121 ), .B(\Inst_Mem/n118 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n122 ) );
  MUX \Inst_Mem/U122  ( .A(\Inst_Mem/n120 ), .B(\Inst_Mem/n119 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n121 ) );
  MUX \Inst_Mem/U121  ( .A(inst_mem_in_wire[1]), .B(inst_mem_in_wire[33]), .S(
        pc_current[2]), .Z(\Inst_Mem/n120 ) );
  MUX \Inst_Mem/U120  ( .A(inst_mem_in_wire[65]), .B(inst_mem_in_wire[97]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n119 ) );
  MUX \Inst_Mem/U119  ( .A(\Inst_Mem/n117 ), .B(\Inst_Mem/n116 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n118 ) );
  MUX \Inst_Mem/U118  ( .A(inst_mem_in_wire[129]), .B(inst_mem_in_wire[161]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n117 ) );
  MUX \Inst_Mem/U117  ( .A(inst_mem_in_wire[193]), .B(inst_mem_in_wire[225]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n116 ) );
  MUX \Inst_Mem/U116  ( .A(\Inst_Mem/n114 ), .B(\Inst_Mem/n111 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n115 ) );
  MUX \Inst_Mem/U115  ( .A(\Inst_Mem/n113 ), .B(\Inst_Mem/n112 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n114 ) );
  MUX \Inst_Mem/U114  ( .A(inst_mem_in_wire[257]), .B(inst_mem_in_wire[289]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n113 ) );
  MUX \Inst_Mem/U113  ( .A(inst_mem_in_wire[321]), .B(inst_mem_in_wire[353]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n112 ) );
  MUX \Inst_Mem/U112  ( .A(\Inst_Mem/n110 ), .B(\Inst_Mem/n109 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n111 ) );
  MUX \Inst_Mem/U111  ( .A(inst_mem_in_wire[385]), .B(inst_mem_in_wire[417]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n110 ) );
  MUX \Inst_Mem/U110  ( .A(inst_mem_in_wire[449]), .B(inst_mem_in_wire[481]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n109 ) );
  MUX \Inst_Mem/U109  ( .A(\Inst_Mem/n107 ), .B(\Inst_Mem/n100 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n108 ) );
  MUX \Inst_Mem/U108  ( .A(\Inst_Mem/n106 ), .B(\Inst_Mem/n103 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n107 ) );
  MUX \Inst_Mem/U107  ( .A(\Inst_Mem/n105 ), .B(\Inst_Mem/n104 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n106 ) );
  MUX \Inst_Mem/U106  ( .A(inst_mem_in_wire[513]), .B(inst_mem_in_wire[545]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n105 ) );
  MUX \Inst_Mem/U105  ( .A(inst_mem_in_wire[577]), .B(inst_mem_in_wire[609]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n104 ) );
  MUX \Inst_Mem/U104  ( .A(\Inst_Mem/n102 ), .B(\Inst_Mem/n101 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n103 ) );
  MUX \Inst_Mem/U103  ( .A(inst_mem_in_wire[641]), .B(inst_mem_in_wire[673]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n102 ) );
  MUX \Inst_Mem/U102  ( .A(inst_mem_in_wire[705]), .B(inst_mem_in_wire[737]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n101 ) );
  MUX \Inst_Mem/U101  ( .A(\Inst_Mem/n99 ), .B(\Inst_Mem/n96 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n100 ) );
  MUX \Inst_Mem/U100  ( .A(\Inst_Mem/n98 ), .B(\Inst_Mem/n97 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n99 ) );
  MUX \Inst_Mem/U99  ( .A(inst_mem_in_wire[769]), .B(inst_mem_in_wire[801]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n98 ) );
  MUX \Inst_Mem/U98  ( .A(inst_mem_in_wire[833]), .B(inst_mem_in_wire[865]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n97 ) );
  MUX \Inst_Mem/U97  ( .A(\Inst_Mem/n95 ), .B(\Inst_Mem/n94 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n96 ) );
  MUX \Inst_Mem/U96  ( .A(inst_mem_in_wire[897]), .B(inst_mem_in_wire[929]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n95 ) );
  MUX \Inst_Mem/U95  ( .A(inst_mem_in_wire[961]), .B(inst_mem_in_wire[993]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n94 ) );
  MUX \Inst_Mem/U94  ( .A(\Inst_Mem/n92 ), .B(\Inst_Mem/n77 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n93 ) );
  MUX \Inst_Mem/U93  ( .A(\Inst_Mem/n91 ), .B(\Inst_Mem/n84 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n92 ) );
  MUX \Inst_Mem/U92  ( .A(\Inst_Mem/n90 ), .B(\Inst_Mem/n87 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n91 ) );
  MUX \Inst_Mem/U91  ( .A(\Inst_Mem/n89 ), .B(\Inst_Mem/n88 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n90 ) );
  MUX \Inst_Mem/U90  ( .A(inst_mem_in_wire[1025]), .B(inst_mem_in_wire[1057]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n89 ) );
  MUX \Inst_Mem/U89  ( .A(inst_mem_in_wire[1089]), .B(inst_mem_in_wire[1121]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n88 ) );
  MUX \Inst_Mem/U88  ( .A(\Inst_Mem/n86 ), .B(\Inst_Mem/n85 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n87 ) );
  MUX \Inst_Mem/U87  ( .A(inst_mem_in_wire[1153]), .B(inst_mem_in_wire[1185]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n86 ) );
  MUX \Inst_Mem/U86  ( .A(inst_mem_in_wire[1217]), .B(inst_mem_in_wire[1249]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n85 ) );
  MUX \Inst_Mem/U85  ( .A(\Inst_Mem/n83 ), .B(\Inst_Mem/n80 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n84 ) );
  MUX \Inst_Mem/U84  ( .A(\Inst_Mem/n82 ), .B(\Inst_Mem/n81 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n83 ) );
  MUX \Inst_Mem/U83  ( .A(inst_mem_in_wire[1281]), .B(inst_mem_in_wire[1313]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n82 ) );
  MUX \Inst_Mem/U82  ( .A(inst_mem_in_wire[1345]), .B(inst_mem_in_wire[1377]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n81 ) );
  MUX \Inst_Mem/U81  ( .A(\Inst_Mem/n79 ), .B(\Inst_Mem/n78 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n80 ) );
  MUX \Inst_Mem/U80  ( .A(inst_mem_in_wire[1409]), .B(inst_mem_in_wire[1441]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n79 ) );
  MUX \Inst_Mem/U79  ( .A(inst_mem_in_wire[1473]), .B(inst_mem_in_wire[1505]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n78 ) );
  MUX \Inst_Mem/U78  ( .A(\Inst_Mem/n76 ), .B(\Inst_Mem/n69 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n77 ) );
  MUX \Inst_Mem/U77  ( .A(\Inst_Mem/n75 ), .B(\Inst_Mem/n72 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n76 ) );
  MUX \Inst_Mem/U76  ( .A(\Inst_Mem/n74 ), .B(\Inst_Mem/n73 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n75 ) );
  MUX \Inst_Mem/U75  ( .A(inst_mem_in_wire[1537]), .B(inst_mem_in_wire[1569]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n74 ) );
  MUX \Inst_Mem/U74  ( .A(inst_mem_in_wire[1601]), .B(inst_mem_in_wire[1633]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n73 ) );
  MUX \Inst_Mem/U73  ( .A(\Inst_Mem/n71 ), .B(\Inst_Mem/n70 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n72 ) );
  MUX \Inst_Mem/U72  ( .A(inst_mem_in_wire[1665]), .B(inst_mem_in_wire[1697]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n71 ) );
  MUX \Inst_Mem/U71  ( .A(inst_mem_in_wire[1729]), .B(inst_mem_in_wire[1761]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n70 ) );
  MUX \Inst_Mem/U70  ( .A(\Inst_Mem/n68 ), .B(\Inst_Mem/n65 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n69 ) );
  MUX \Inst_Mem/U69  ( .A(\Inst_Mem/n67 ), .B(\Inst_Mem/n66 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n68 ) );
  MUX \Inst_Mem/U68  ( .A(inst_mem_in_wire[1793]), .B(inst_mem_in_wire[1825]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n67 ) );
  MUX \Inst_Mem/U67  ( .A(inst_mem_in_wire[1857]), .B(inst_mem_in_wire[1889]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n66 ) );
  MUX \Inst_Mem/U66  ( .A(\Inst_Mem/n64 ), .B(\Inst_Mem/n63 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n65 ) );
  MUX \Inst_Mem/U65  ( .A(inst_mem_in_wire[1921]), .B(inst_mem_in_wire[1953]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n64 ) );
  MUX \Inst_Mem/U64  ( .A(inst_mem_in_wire[1985]), .B(inst_mem_in_wire[2017]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n63 ) );
  MUX \Inst_Mem/U63  ( .A(\Inst_Mem/n62 ), .B(\Inst_Mem/n31 ), .S(
        pc_current[7]), .Z(imm[0]) );
  MUX \Inst_Mem/U62  ( .A(\Inst_Mem/n61 ), .B(\Inst_Mem/n46 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n62 ) );
  MUX \Inst_Mem/U61  ( .A(\Inst_Mem/n60 ), .B(\Inst_Mem/n53 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n61 ) );
  MUX \Inst_Mem/U60  ( .A(\Inst_Mem/n59 ), .B(\Inst_Mem/n56 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n60 ) );
  MUX \Inst_Mem/U59  ( .A(\Inst_Mem/n58 ), .B(\Inst_Mem/n57 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n59 ) );
  MUX \Inst_Mem/U58  ( .A(inst_mem_in_wire[0]), .B(inst_mem_in_wire[32]), .S(
        pc_current[2]), .Z(\Inst_Mem/n58 ) );
  MUX \Inst_Mem/U57  ( .A(inst_mem_in_wire[64]), .B(inst_mem_in_wire[96]), .S(
        pc_current[2]), .Z(\Inst_Mem/n57 ) );
  MUX \Inst_Mem/U56  ( .A(\Inst_Mem/n55 ), .B(\Inst_Mem/n54 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n56 ) );
  MUX \Inst_Mem/U55  ( .A(inst_mem_in_wire[128]), .B(inst_mem_in_wire[160]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n55 ) );
  MUX \Inst_Mem/U54  ( .A(inst_mem_in_wire[192]), .B(inst_mem_in_wire[224]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n54 ) );
  MUX \Inst_Mem/U53  ( .A(\Inst_Mem/n52 ), .B(\Inst_Mem/n49 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n53 ) );
  MUX \Inst_Mem/U52  ( .A(\Inst_Mem/n51 ), .B(\Inst_Mem/n50 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n52 ) );
  MUX \Inst_Mem/U51  ( .A(inst_mem_in_wire[256]), .B(inst_mem_in_wire[288]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n51 ) );
  MUX \Inst_Mem/U50  ( .A(inst_mem_in_wire[320]), .B(inst_mem_in_wire[352]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n50 ) );
  MUX \Inst_Mem/U49  ( .A(\Inst_Mem/n48 ), .B(\Inst_Mem/n47 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n49 ) );
  MUX \Inst_Mem/U48  ( .A(inst_mem_in_wire[384]), .B(inst_mem_in_wire[416]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n48 ) );
  MUX \Inst_Mem/U47  ( .A(inst_mem_in_wire[448]), .B(inst_mem_in_wire[480]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n47 ) );
  MUX \Inst_Mem/U46  ( .A(\Inst_Mem/n45 ), .B(\Inst_Mem/n38 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n46 ) );
  MUX \Inst_Mem/U45  ( .A(\Inst_Mem/n44 ), .B(\Inst_Mem/n41 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n45 ) );
  MUX \Inst_Mem/U44  ( .A(\Inst_Mem/n43 ), .B(\Inst_Mem/n42 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n44 ) );
  MUX \Inst_Mem/U43  ( .A(inst_mem_in_wire[512]), .B(inst_mem_in_wire[544]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n43 ) );
  MUX \Inst_Mem/U42  ( .A(inst_mem_in_wire[576]), .B(inst_mem_in_wire[608]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n42 ) );
  MUX \Inst_Mem/U41  ( .A(\Inst_Mem/n40 ), .B(\Inst_Mem/n39 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n41 ) );
  MUX \Inst_Mem/U40  ( .A(inst_mem_in_wire[640]), .B(inst_mem_in_wire[672]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n40 ) );
  MUX \Inst_Mem/U39  ( .A(inst_mem_in_wire[704]), .B(inst_mem_in_wire[736]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n39 ) );
  MUX \Inst_Mem/U38  ( .A(\Inst_Mem/n37 ), .B(\Inst_Mem/n34 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n38 ) );
  MUX \Inst_Mem/U37  ( .A(\Inst_Mem/n36 ), .B(\Inst_Mem/n35 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n37 ) );
  MUX \Inst_Mem/U36  ( .A(inst_mem_in_wire[768]), .B(inst_mem_in_wire[800]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n36 ) );
  MUX \Inst_Mem/U35  ( .A(inst_mem_in_wire[832]), .B(inst_mem_in_wire[864]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n35 ) );
  MUX \Inst_Mem/U34  ( .A(\Inst_Mem/n33 ), .B(\Inst_Mem/n32 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n34 ) );
  MUX \Inst_Mem/U33  ( .A(inst_mem_in_wire[896]), .B(inst_mem_in_wire[928]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n33 ) );
  MUX \Inst_Mem/U32  ( .A(inst_mem_in_wire[960]), .B(inst_mem_in_wire[992]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n32 ) );
  MUX \Inst_Mem/U31  ( .A(\Inst_Mem/n30 ), .B(\Inst_Mem/n15 ), .S(
        pc_current[6]), .Z(\Inst_Mem/n31 ) );
  MUX \Inst_Mem/U30  ( .A(\Inst_Mem/n29 ), .B(\Inst_Mem/n22 ), .S(
        pc_current[5]), .Z(\Inst_Mem/n30 ) );
  MUX \Inst_Mem/U29  ( .A(\Inst_Mem/n28 ), .B(\Inst_Mem/n25 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n29 ) );
  MUX \Inst_Mem/U28  ( .A(\Inst_Mem/n27 ), .B(\Inst_Mem/n26 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n28 ) );
  MUX \Inst_Mem/U27  ( .A(inst_mem_in_wire[1024]), .B(inst_mem_in_wire[1056]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n27 ) );
  MUX \Inst_Mem/U26  ( .A(inst_mem_in_wire[1088]), .B(inst_mem_in_wire[1120]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n26 ) );
  MUX \Inst_Mem/U25  ( .A(\Inst_Mem/n24 ), .B(\Inst_Mem/n23 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n25 ) );
  MUX \Inst_Mem/U24  ( .A(inst_mem_in_wire[1152]), .B(inst_mem_in_wire[1184]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n24 ) );
  MUX \Inst_Mem/U23  ( .A(inst_mem_in_wire[1216]), .B(inst_mem_in_wire[1248]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n23 ) );
  MUX \Inst_Mem/U22  ( .A(\Inst_Mem/n21 ), .B(\Inst_Mem/n18 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n22 ) );
  MUX \Inst_Mem/U21  ( .A(\Inst_Mem/n20 ), .B(\Inst_Mem/n19 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n21 ) );
  MUX \Inst_Mem/U20  ( .A(inst_mem_in_wire[1280]), .B(inst_mem_in_wire[1312]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n20 ) );
  MUX \Inst_Mem/U19  ( .A(inst_mem_in_wire[1344]), .B(inst_mem_in_wire[1376]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n19 ) );
  MUX \Inst_Mem/U18  ( .A(\Inst_Mem/n17 ), .B(\Inst_Mem/n16 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n18 ) );
  MUX \Inst_Mem/U17  ( .A(inst_mem_in_wire[1408]), .B(inst_mem_in_wire[1440]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n17 ) );
  MUX \Inst_Mem/U16  ( .A(inst_mem_in_wire[1472]), .B(inst_mem_in_wire[1504]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n16 ) );
  MUX \Inst_Mem/U15  ( .A(\Inst_Mem/n14 ), .B(\Inst_Mem/n7 ), .S(pc_current[5]), .Z(\Inst_Mem/n15 ) );
  MUX \Inst_Mem/U14  ( .A(\Inst_Mem/n13 ), .B(\Inst_Mem/n10 ), .S(
        pc_current[4]), .Z(\Inst_Mem/n14 ) );
  MUX \Inst_Mem/U13  ( .A(\Inst_Mem/n12 ), .B(\Inst_Mem/n11 ), .S(
        pc_current[3]), .Z(\Inst_Mem/n13 ) );
  MUX \Inst_Mem/U12  ( .A(inst_mem_in_wire[1536]), .B(inst_mem_in_wire[1568]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n12 ) );
  MUX \Inst_Mem/U11  ( .A(inst_mem_in_wire[1600]), .B(inst_mem_in_wire[1632]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n11 ) );
  MUX \Inst_Mem/U10  ( .A(\Inst_Mem/n9 ), .B(\Inst_Mem/n8 ), .S(pc_current[3]), 
        .Z(\Inst_Mem/n10 ) );
  MUX \Inst_Mem/U9  ( .A(inst_mem_in_wire[1664]), .B(inst_mem_in_wire[1696]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n9 ) );
  MUX \Inst_Mem/U8  ( .A(inst_mem_in_wire[1728]), .B(inst_mem_in_wire[1760]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n8 ) );
  MUX \Inst_Mem/U7  ( .A(\Inst_Mem/n6 ), .B(\Inst_Mem/n3 ), .S(pc_current[4]), 
        .Z(\Inst_Mem/n7 ) );
  MUX \Inst_Mem/U6  ( .A(\Inst_Mem/n5 ), .B(\Inst_Mem/n4 ), .S(pc_current[3]), 
        .Z(\Inst_Mem/n6 ) );
  MUX \Inst_Mem/U5  ( .A(inst_mem_in_wire[1792]), .B(inst_mem_in_wire[1824]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n5 ) );
  MUX \Inst_Mem/U4  ( .A(inst_mem_in_wire[1856]), .B(inst_mem_in_wire[1888]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n4 ) );
  MUX \Inst_Mem/U3  ( .A(\Inst_Mem/n2 ), .B(\Inst_Mem/n1 ), .S(pc_current[3]), 
        .Z(\Inst_Mem/n3 ) );
  MUX \Inst_Mem/U2  ( .A(inst_mem_in_wire[1920]), .B(inst_mem_in_wire[1952]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n2 ) );
  MUX \Inst_Mem/U1  ( .A(inst_mem_in_wire[1984]), .B(inst_mem_in_wire[2016]), 
        .S(pc_current[2]), .Z(\Inst_Mem/n1 ) );
  MUX \Data_Mem/U8280  ( .A(\Data_Mem/n8247 ), .B(\Data_Mem/n8216 ), .S(N24), 
        .Z(c_memory[31]) );
  MUX \Data_Mem/U8279  ( .A(\Data_Mem/n8246 ), .B(\Data_Mem/n8231 ), .S(N25), 
        .Z(\Data_Mem/n8247 ) );
  MUX \Data_Mem/U8278  ( .A(\Data_Mem/n8245 ), .B(\Data_Mem/n8238 ), .S(N26), 
        .Z(\Data_Mem/n8246 ) );
  MUX \Data_Mem/U8277  ( .A(\Data_Mem/n8244 ), .B(\Data_Mem/n8241 ), .S(N27), 
        .Z(\Data_Mem/n8245 ) );
  MUX \Data_Mem/U8276  ( .A(\Data_Mem/n8243 ), .B(\Data_Mem/n8242 ), .S(N28), 
        .Z(\Data_Mem/n8244 ) );
  MUX \Data_Mem/U8275  ( .A(data_mem_out_wire[31]), .B(data_mem_out_wire[63]), 
        .S(N29), .Z(\Data_Mem/n8243 ) );
  MUX \Data_Mem/U8274  ( .A(data_mem_out_wire[95]), .B(data_mem_out_wire[127]), 
        .S(N29), .Z(\Data_Mem/n8242 ) );
  MUX \Data_Mem/U8273  ( .A(\Data_Mem/n8240 ), .B(\Data_Mem/n8239 ), .S(N28), 
        .Z(\Data_Mem/n8241 ) );
  MUX \Data_Mem/U8272  ( .A(data_mem_out_wire[159]), .B(data_mem_out_wire[191]), .S(N29), .Z(\Data_Mem/n8240 ) );
  MUX \Data_Mem/U8271  ( .A(data_mem_out_wire[223]), .B(data_mem_out_wire[255]), .S(N29), .Z(\Data_Mem/n8239 ) );
  MUX \Data_Mem/U8270  ( .A(\Data_Mem/n8237 ), .B(\Data_Mem/n8234 ), .S(N27), 
        .Z(\Data_Mem/n8238 ) );
  MUX \Data_Mem/U8269  ( .A(\Data_Mem/n8236 ), .B(\Data_Mem/n8235 ), .S(N28), 
        .Z(\Data_Mem/n8237 ) );
  MUX \Data_Mem/U8268  ( .A(data_mem_out_wire[287]), .B(data_mem_out_wire[319]), .S(N29), .Z(\Data_Mem/n8236 ) );
  MUX \Data_Mem/U8267  ( .A(data_mem_out_wire[351]), .B(data_mem_out_wire[383]), .S(N29), .Z(\Data_Mem/n8235 ) );
  MUX \Data_Mem/U8266  ( .A(\Data_Mem/n8233 ), .B(\Data_Mem/n8232 ), .S(N28), 
        .Z(\Data_Mem/n8234 ) );
  MUX \Data_Mem/U8265  ( .A(data_mem_out_wire[415]), .B(data_mem_out_wire[447]), .S(N29), .Z(\Data_Mem/n8233 ) );
  MUX \Data_Mem/U8264  ( .A(data_mem_out_wire[479]), .B(data_mem_out_wire[511]), .S(N29), .Z(\Data_Mem/n8232 ) );
  MUX \Data_Mem/U8263  ( .A(\Data_Mem/n8230 ), .B(\Data_Mem/n8223 ), .S(N26), 
        .Z(\Data_Mem/n8231 ) );
  MUX \Data_Mem/U8262  ( .A(\Data_Mem/n8229 ), .B(\Data_Mem/n8226 ), .S(N27), 
        .Z(\Data_Mem/n8230 ) );
  MUX \Data_Mem/U8261  ( .A(\Data_Mem/n8228 ), .B(\Data_Mem/n8227 ), .S(N28), 
        .Z(\Data_Mem/n8229 ) );
  MUX \Data_Mem/U8260  ( .A(data_mem_out_wire[543]), .B(data_mem_out_wire[575]), .S(N29), .Z(\Data_Mem/n8228 ) );
  MUX \Data_Mem/U8259  ( .A(data_mem_out_wire[607]), .B(data_mem_out_wire[639]), .S(N29), .Z(\Data_Mem/n8227 ) );
  MUX \Data_Mem/U8258  ( .A(\Data_Mem/n8225 ), .B(\Data_Mem/n8224 ), .S(N28), 
        .Z(\Data_Mem/n8226 ) );
  MUX \Data_Mem/U8257  ( .A(data_mem_out_wire[671]), .B(data_mem_out_wire[703]), .S(N29), .Z(\Data_Mem/n8225 ) );
  MUX \Data_Mem/U8256  ( .A(data_mem_out_wire[735]), .B(data_mem_out_wire[767]), .S(N29), .Z(\Data_Mem/n8224 ) );
  MUX \Data_Mem/U8255  ( .A(\Data_Mem/n8222 ), .B(\Data_Mem/n8219 ), .S(N27), 
        .Z(\Data_Mem/n8223 ) );
  MUX \Data_Mem/U8254  ( .A(\Data_Mem/n8221 ), .B(\Data_Mem/n8220 ), .S(N28), 
        .Z(\Data_Mem/n8222 ) );
  MUX \Data_Mem/U8253  ( .A(data_mem_out_wire[799]), .B(data_mem_out_wire[831]), .S(N29), .Z(\Data_Mem/n8221 ) );
  MUX \Data_Mem/U8252  ( .A(data_mem_out_wire[863]), .B(data_mem_out_wire[895]), .S(N29), .Z(\Data_Mem/n8220 ) );
  MUX \Data_Mem/U8251  ( .A(\Data_Mem/n8218 ), .B(\Data_Mem/n8217 ), .S(N28), 
        .Z(\Data_Mem/n8219 ) );
  MUX \Data_Mem/U8250  ( .A(data_mem_out_wire[927]), .B(data_mem_out_wire[959]), .S(N29), .Z(\Data_Mem/n8218 ) );
  MUX \Data_Mem/U8249  ( .A(data_mem_out_wire[991]), .B(
        data_mem_out_wire[1023]), .S(N29), .Z(\Data_Mem/n8217 ) );
  MUX \Data_Mem/U8248  ( .A(\Data_Mem/n8215 ), .B(\Data_Mem/n8200 ), .S(N25), 
        .Z(\Data_Mem/n8216 ) );
  MUX \Data_Mem/U8247  ( .A(\Data_Mem/n8214 ), .B(\Data_Mem/n8207 ), .S(N26), 
        .Z(\Data_Mem/n8215 ) );
  MUX \Data_Mem/U8246  ( .A(\Data_Mem/n8213 ), .B(\Data_Mem/n8210 ), .S(N27), 
        .Z(\Data_Mem/n8214 ) );
  MUX \Data_Mem/U8245  ( .A(\Data_Mem/n8212 ), .B(\Data_Mem/n8211 ), .S(N28), 
        .Z(\Data_Mem/n8213 ) );
  MUX \Data_Mem/U8244  ( .A(data_mem_out_wire[1055]), .B(
        data_mem_out_wire[1087]), .S(N29), .Z(\Data_Mem/n8212 ) );
  MUX \Data_Mem/U8243  ( .A(data_mem_out_wire[1119]), .B(
        data_mem_out_wire[1151]), .S(N29), .Z(\Data_Mem/n8211 ) );
  MUX \Data_Mem/U8242  ( .A(\Data_Mem/n8209 ), .B(\Data_Mem/n8208 ), .S(N28), 
        .Z(\Data_Mem/n8210 ) );
  MUX \Data_Mem/U8241  ( .A(data_mem_out_wire[1183]), .B(
        data_mem_out_wire[1215]), .S(N29), .Z(\Data_Mem/n8209 ) );
  MUX \Data_Mem/U8240  ( .A(data_mem_out_wire[1247]), .B(
        data_mem_out_wire[1279]), .S(N29), .Z(\Data_Mem/n8208 ) );
  MUX \Data_Mem/U8239  ( .A(\Data_Mem/n8206 ), .B(\Data_Mem/n8203 ), .S(N27), 
        .Z(\Data_Mem/n8207 ) );
  MUX \Data_Mem/U8238  ( .A(\Data_Mem/n8205 ), .B(\Data_Mem/n8204 ), .S(N28), 
        .Z(\Data_Mem/n8206 ) );
  MUX \Data_Mem/U8237  ( .A(data_mem_out_wire[1311]), .B(
        data_mem_out_wire[1343]), .S(N29), .Z(\Data_Mem/n8205 ) );
  MUX \Data_Mem/U8236  ( .A(data_mem_out_wire[1375]), .B(
        data_mem_out_wire[1407]), .S(N29), .Z(\Data_Mem/n8204 ) );
  MUX \Data_Mem/U8235  ( .A(\Data_Mem/n8202 ), .B(\Data_Mem/n8201 ), .S(N28), 
        .Z(\Data_Mem/n8203 ) );
  MUX \Data_Mem/U8234  ( .A(data_mem_out_wire[1439]), .B(
        data_mem_out_wire[1471]), .S(N29), .Z(\Data_Mem/n8202 ) );
  MUX \Data_Mem/U8233  ( .A(data_mem_out_wire[1503]), .B(
        data_mem_out_wire[1535]), .S(N29), .Z(\Data_Mem/n8201 ) );
  MUX \Data_Mem/U8232  ( .A(\Data_Mem/n8199 ), .B(\Data_Mem/n8192 ), .S(N26), 
        .Z(\Data_Mem/n8200 ) );
  MUX \Data_Mem/U8231  ( .A(\Data_Mem/n8198 ), .B(\Data_Mem/n8195 ), .S(N27), 
        .Z(\Data_Mem/n8199 ) );
  MUX \Data_Mem/U8230  ( .A(\Data_Mem/n8197 ), .B(\Data_Mem/n8196 ), .S(N28), 
        .Z(\Data_Mem/n8198 ) );
  MUX \Data_Mem/U8229  ( .A(data_mem_out_wire[1567]), .B(
        data_mem_out_wire[1599]), .S(N29), .Z(\Data_Mem/n8197 ) );
  MUX \Data_Mem/U8228  ( .A(data_mem_out_wire[1631]), .B(
        data_mem_out_wire[1663]), .S(N29), .Z(\Data_Mem/n8196 ) );
  MUX \Data_Mem/U8227  ( .A(\Data_Mem/n8194 ), .B(\Data_Mem/n8193 ), .S(N28), 
        .Z(\Data_Mem/n8195 ) );
  MUX \Data_Mem/U8226  ( .A(data_mem_out_wire[1695]), .B(
        data_mem_out_wire[1727]), .S(N29), .Z(\Data_Mem/n8194 ) );
  MUX \Data_Mem/U8225  ( .A(data_mem_out_wire[1759]), .B(
        data_mem_out_wire[1791]), .S(N29), .Z(\Data_Mem/n8193 ) );
  MUX \Data_Mem/U8224  ( .A(\Data_Mem/n8191 ), .B(\Data_Mem/n8188 ), .S(N27), 
        .Z(\Data_Mem/n8192 ) );
  MUX \Data_Mem/U8223  ( .A(\Data_Mem/n8190 ), .B(\Data_Mem/n8189 ), .S(N28), 
        .Z(\Data_Mem/n8191 ) );
  MUX \Data_Mem/U8222  ( .A(data_mem_out_wire[1823]), .B(
        data_mem_out_wire[1855]), .S(N29), .Z(\Data_Mem/n8190 ) );
  MUX \Data_Mem/U8221  ( .A(data_mem_out_wire[1887]), .B(
        data_mem_out_wire[1919]), .S(N29), .Z(\Data_Mem/n8189 ) );
  MUX \Data_Mem/U8220  ( .A(\Data_Mem/n8187 ), .B(\Data_Mem/n8186 ), .S(N28), 
        .Z(\Data_Mem/n8188 ) );
  MUX \Data_Mem/U8219  ( .A(data_mem_out_wire[1951]), .B(
        data_mem_out_wire[1983]), .S(N29), .Z(\Data_Mem/n8187 ) );
  MUX \Data_Mem/U8218  ( .A(data_mem_out_wire[2015]), .B(
        data_mem_out_wire[2047]), .S(N29), .Z(\Data_Mem/n8186 ) );
  MUX \Data_Mem/U8217  ( .A(\Data_Mem/n8185 ), .B(\Data_Mem/n8154 ), .S(N24), 
        .Z(c_memory[30]) );
  MUX \Data_Mem/U8216  ( .A(\Data_Mem/n8184 ), .B(\Data_Mem/n8169 ), .S(N25), 
        .Z(\Data_Mem/n8185 ) );
  MUX \Data_Mem/U8215  ( .A(\Data_Mem/n8183 ), .B(\Data_Mem/n8176 ), .S(N26), 
        .Z(\Data_Mem/n8184 ) );
  MUX \Data_Mem/U8214  ( .A(\Data_Mem/n8182 ), .B(\Data_Mem/n8179 ), .S(N27), 
        .Z(\Data_Mem/n8183 ) );
  MUX \Data_Mem/U8213  ( .A(\Data_Mem/n8181 ), .B(\Data_Mem/n8180 ), .S(N28), 
        .Z(\Data_Mem/n8182 ) );
  MUX \Data_Mem/U8212  ( .A(data_mem_out_wire[30]), .B(data_mem_out_wire[62]), 
        .S(N29), .Z(\Data_Mem/n8181 ) );
  MUX \Data_Mem/U8211  ( .A(data_mem_out_wire[94]), .B(data_mem_out_wire[126]), 
        .S(N29), .Z(\Data_Mem/n8180 ) );
  MUX \Data_Mem/U8210  ( .A(\Data_Mem/n8178 ), .B(\Data_Mem/n8177 ), .S(N28), 
        .Z(\Data_Mem/n8179 ) );
  MUX \Data_Mem/U8209  ( .A(data_mem_out_wire[158]), .B(data_mem_out_wire[190]), .S(N29), .Z(\Data_Mem/n8178 ) );
  MUX \Data_Mem/U8208  ( .A(data_mem_out_wire[222]), .B(data_mem_out_wire[254]), .S(N29), .Z(\Data_Mem/n8177 ) );
  MUX \Data_Mem/U8207  ( .A(\Data_Mem/n8175 ), .B(\Data_Mem/n8172 ), .S(N27), 
        .Z(\Data_Mem/n8176 ) );
  MUX \Data_Mem/U8206  ( .A(\Data_Mem/n8174 ), .B(\Data_Mem/n8173 ), .S(N28), 
        .Z(\Data_Mem/n8175 ) );
  MUX \Data_Mem/U8205  ( .A(data_mem_out_wire[286]), .B(data_mem_out_wire[318]), .S(N29), .Z(\Data_Mem/n8174 ) );
  MUX \Data_Mem/U8204  ( .A(data_mem_out_wire[350]), .B(data_mem_out_wire[382]), .S(N29), .Z(\Data_Mem/n8173 ) );
  MUX \Data_Mem/U8203  ( .A(\Data_Mem/n8171 ), .B(\Data_Mem/n8170 ), .S(N28), 
        .Z(\Data_Mem/n8172 ) );
  MUX \Data_Mem/U8202  ( .A(data_mem_out_wire[414]), .B(data_mem_out_wire[446]), .S(N29), .Z(\Data_Mem/n8171 ) );
  MUX \Data_Mem/U8201  ( .A(data_mem_out_wire[478]), .B(data_mem_out_wire[510]), .S(N29), .Z(\Data_Mem/n8170 ) );
  MUX \Data_Mem/U8200  ( .A(\Data_Mem/n8168 ), .B(\Data_Mem/n8161 ), .S(N26), 
        .Z(\Data_Mem/n8169 ) );
  MUX \Data_Mem/U8199  ( .A(\Data_Mem/n8167 ), .B(\Data_Mem/n8164 ), .S(N27), 
        .Z(\Data_Mem/n8168 ) );
  MUX \Data_Mem/U8198  ( .A(\Data_Mem/n8166 ), .B(\Data_Mem/n8165 ), .S(N28), 
        .Z(\Data_Mem/n8167 ) );
  MUX \Data_Mem/U8197  ( .A(data_mem_out_wire[542]), .B(data_mem_out_wire[574]), .S(N29), .Z(\Data_Mem/n8166 ) );
  MUX \Data_Mem/U8196  ( .A(data_mem_out_wire[606]), .B(data_mem_out_wire[638]), .S(N29), .Z(\Data_Mem/n8165 ) );
  MUX \Data_Mem/U8195  ( .A(\Data_Mem/n8163 ), .B(\Data_Mem/n8162 ), .S(N28), 
        .Z(\Data_Mem/n8164 ) );
  MUX \Data_Mem/U8194  ( .A(data_mem_out_wire[670]), .B(data_mem_out_wire[702]), .S(N29), .Z(\Data_Mem/n8163 ) );
  MUX \Data_Mem/U8193  ( .A(data_mem_out_wire[734]), .B(data_mem_out_wire[766]), .S(N29), .Z(\Data_Mem/n8162 ) );
  MUX \Data_Mem/U8192  ( .A(\Data_Mem/n8160 ), .B(\Data_Mem/n8157 ), .S(N27), 
        .Z(\Data_Mem/n8161 ) );
  MUX \Data_Mem/U8191  ( .A(\Data_Mem/n8159 ), .B(\Data_Mem/n8158 ), .S(N28), 
        .Z(\Data_Mem/n8160 ) );
  MUX \Data_Mem/U8190  ( .A(data_mem_out_wire[798]), .B(data_mem_out_wire[830]), .S(N29), .Z(\Data_Mem/n8159 ) );
  MUX \Data_Mem/U8189  ( .A(data_mem_out_wire[862]), .B(data_mem_out_wire[894]), .S(N29), .Z(\Data_Mem/n8158 ) );
  MUX \Data_Mem/U8188  ( .A(\Data_Mem/n8156 ), .B(\Data_Mem/n8155 ), .S(N28), 
        .Z(\Data_Mem/n8157 ) );
  MUX \Data_Mem/U8187  ( .A(data_mem_out_wire[926]), .B(data_mem_out_wire[958]), .S(N29), .Z(\Data_Mem/n8156 ) );
  MUX \Data_Mem/U8186  ( .A(data_mem_out_wire[990]), .B(
        data_mem_out_wire[1022]), .S(N29), .Z(\Data_Mem/n8155 ) );
  MUX \Data_Mem/U8185  ( .A(\Data_Mem/n8153 ), .B(\Data_Mem/n8138 ), .S(N25), 
        .Z(\Data_Mem/n8154 ) );
  MUX \Data_Mem/U8184  ( .A(\Data_Mem/n8152 ), .B(\Data_Mem/n8145 ), .S(N26), 
        .Z(\Data_Mem/n8153 ) );
  MUX \Data_Mem/U8183  ( .A(\Data_Mem/n8151 ), .B(\Data_Mem/n8148 ), .S(N27), 
        .Z(\Data_Mem/n8152 ) );
  MUX \Data_Mem/U8182  ( .A(\Data_Mem/n8150 ), .B(\Data_Mem/n8149 ), .S(N28), 
        .Z(\Data_Mem/n8151 ) );
  MUX \Data_Mem/U8181  ( .A(data_mem_out_wire[1054]), .B(
        data_mem_out_wire[1086]), .S(N29), .Z(\Data_Mem/n8150 ) );
  MUX \Data_Mem/U8180  ( .A(data_mem_out_wire[1118]), .B(
        data_mem_out_wire[1150]), .S(N29), .Z(\Data_Mem/n8149 ) );
  MUX \Data_Mem/U8179  ( .A(\Data_Mem/n8147 ), .B(\Data_Mem/n8146 ), .S(N28), 
        .Z(\Data_Mem/n8148 ) );
  MUX \Data_Mem/U8178  ( .A(data_mem_out_wire[1182]), .B(
        data_mem_out_wire[1214]), .S(N29), .Z(\Data_Mem/n8147 ) );
  MUX \Data_Mem/U8177  ( .A(data_mem_out_wire[1246]), .B(
        data_mem_out_wire[1278]), .S(N29), .Z(\Data_Mem/n8146 ) );
  MUX \Data_Mem/U8176  ( .A(\Data_Mem/n8144 ), .B(\Data_Mem/n8141 ), .S(N27), 
        .Z(\Data_Mem/n8145 ) );
  MUX \Data_Mem/U8175  ( .A(\Data_Mem/n8143 ), .B(\Data_Mem/n8142 ), .S(N28), 
        .Z(\Data_Mem/n8144 ) );
  MUX \Data_Mem/U8174  ( .A(data_mem_out_wire[1310]), .B(
        data_mem_out_wire[1342]), .S(N29), .Z(\Data_Mem/n8143 ) );
  MUX \Data_Mem/U8173  ( .A(data_mem_out_wire[1374]), .B(
        data_mem_out_wire[1406]), .S(N29), .Z(\Data_Mem/n8142 ) );
  MUX \Data_Mem/U8172  ( .A(\Data_Mem/n8140 ), .B(\Data_Mem/n8139 ), .S(N28), 
        .Z(\Data_Mem/n8141 ) );
  MUX \Data_Mem/U8171  ( .A(data_mem_out_wire[1438]), .B(
        data_mem_out_wire[1470]), .S(N29), .Z(\Data_Mem/n8140 ) );
  MUX \Data_Mem/U8170  ( .A(data_mem_out_wire[1502]), .B(
        data_mem_out_wire[1534]), .S(N29), .Z(\Data_Mem/n8139 ) );
  MUX \Data_Mem/U8169  ( .A(\Data_Mem/n8137 ), .B(\Data_Mem/n8130 ), .S(N26), 
        .Z(\Data_Mem/n8138 ) );
  MUX \Data_Mem/U8168  ( .A(\Data_Mem/n8136 ), .B(\Data_Mem/n8133 ), .S(N27), 
        .Z(\Data_Mem/n8137 ) );
  MUX \Data_Mem/U8167  ( .A(\Data_Mem/n8135 ), .B(\Data_Mem/n8134 ), .S(N28), 
        .Z(\Data_Mem/n8136 ) );
  MUX \Data_Mem/U8166  ( .A(data_mem_out_wire[1566]), .B(
        data_mem_out_wire[1598]), .S(N29), .Z(\Data_Mem/n8135 ) );
  MUX \Data_Mem/U8165  ( .A(data_mem_out_wire[1630]), .B(
        data_mem_out_wire[1662]), .S(N29), .Z(\Data_Mem/n8134 ) );
  MUX \Data_Mem/U8164  ( .A(\Data_Mem/n8132 ), .B(\Data_Mem/n8131 ), .S(N28), 
        .Z(\Data_Mem/n8133 ) );
  MUX \Data_Mem/U8163  ( .A(data_mem_out_wire[1694]), .B(
        data_mem_out_wire[1726]), .S(N29), .Z(\Data_Mem/n8132 ) );
  MUX \Data_Mem/U8162  ( .A(data_mem_out_wire[1758]), .B(
        data_mem_out_wire[1790]), .S(N29), .Z(\Data_Mem/n8131 ) );
  MUX \Data_Mem/U8161  ( .A(\Data_Mem/n8129 ), .B(\Data_Mem/n8126 ), .S(N27), 
        .Z(\Data_Mem/n8130 ) );
  MUX \Data_Mem/U8160  ( .A(\Data_Mem/n8128 ), .B(\Data_Mem/n8127 ), .S(N28), 
        .Z(\Data_Mem/n8129 ) );
  MUX \Data_Mem/U8159  ( .A(data_mem_out_wire[1822]), .B(
        data_mem_out_wire[1854]), .S(N29), .Z(\Data_Mem/n8128 ) );
  MUX \Data_Mem/U8158  ( .A(data_mem_out_wire[1886]), .B(
        data_mem_out_wire[1918]), .S(N29), .Z(\Data_Mem/n8127 ) );
  MUX \Data_Mem/U8157  ( .A(\Data_Mem/n8125 ), .B(\Data_Mem/n8124 ), .S(N28), 
        .Z(\Data_Mem/n8126 ) );
  MUX \Data_Mem/U8156  ( .A(data_mem_out_wire[1950]), .B(
        data_mem_out_wire[1982]), .S(N29), .Z(\Data_Mem/n8125 ) );
  MUX \Data_Mem/U8155  ( .A(data_mem_out_wire[2014]), .B(
        data_mem_out_wire[2046]), .S(N29), .Z(\Data_Mem/n8124 ) );
  MUX \Data_Mem/U8154  ( .A(\Data_Mem/n8123 ), .B(\Data_Mem/n8092 ), .S(N24), 
        .Z(c_memory[29]) );
  MUX \Data_Mem/U8153  ( .A(\Data_Mem/n8122 ), .B(\Data_Mem/n8107 ), .S(N25), 
        .Z(\Data_Mem/n8123 ) );
  MUX \Data_Mem/U8152  ( .A(\Data_Mem/n8121 ), .B(\Data_Mem/n8114 ), .S(N26), 
        .Z(\Data_Mem/n8122 ) );
  MUX \Data_Mem/U8151  ( .A(\Data_Mem/n8120 ), .B(\Data_Mem/n8117 ), .S(N27), 
        .Z(\Data_Mem/n8121 ) );
  MUX \Data_Mem/U8150  ( .A(\Data_Mem/n8119 ), .B(\Data_Mem/n8118 ), .S(N28), 
        .Z(\Data_Mem/n8120 ) );
  MUX \Data_Mem/U8149  ( .A(data_mem_out_wire[29]), .B(data_mem_out_wire[61]), 
        .S(N29), .Z(\Data_Mem/n8119 ) );
  MUX \Data_Mem/U8148  ( .A(data_mem_out_wire[93]), .B(data_mem_out_wire[125]), 
        .S(N29), .Z(\Data_Mem/n8118 ) );
  MUX \Data_Mem/U8147  ( .A(\Data_Mem/n8116 ), .B(\Data_Mem/n8115 ), .S(N28), 
        .Z(\Data_Mem/n8117 ) );
  MUX \Data_Mem/U8146  ( .A(data_mem_out_wire[157]), .B(data_mem_out_wire[189]), .S(N29), .Z(\Data_Mem/n8116 ) );
  MUX \Data_Mem/U8145  ( .A(data_mem_out_wire[221]), .B(data_mem_out_wire[253]), .S(N29), .Z(\Data_Mem/n8115 ) );
  MUX \Data_Mem/U8144  ( .A(\Data_Mem/n8113 ), .B(\Data_Mem/n8110 ), .S(N27), 
        .Z(\Data_Mem/n8114 ) );
  MUX \Data_Mem/U8143  ( .A(\Data_Mem/n8112 ), .B(\Data_Mem/n8111 ), .S(N28), 
        .Z(\Data_Mem/n8113 ) );
  MUX \Data_Mem/U8142  ( .A(data_mem_out_wire[285]), .B(data_mem_out_wire[317]), .S(N29), .Z(\Data_Mem/n8112 ) );
  MUX \Data_Mem/U8141  ( .A(data_mem_out_wire[349]), .B(data_mem_out_wire[381]), .S(N29), .Z(\Data_Mem/n8111 ) );
  MUX \Data_Mem/U8140  ( .A(\Data_Mem/n8109 ), .B(\Data_Mem/n8108 ), .S(N28), 
        .Z(\Data_Mem/n8110 ) );
  MUX \Data_Mem/U8139  ( .A(data_mem_out_wire[413]), .B(data_mem_out_wire[445]), .S(N29), .Z(\Data_Mem/n8109 ) );
  MUX \Data_Mem/U8138  ( .A(data_mem_out_wire[477]), .B(data_mem_out_wire[509]), .S(N29), .Z(\Data_Mem/n8108 ) );
  MUX \Data_Mem/U8137  ( .A(\Data_Mem/n8106 ), .B(\Data_Mem/n8099 ), .S(N26), 
        .Z(\Data_Mem/n8107 ) );
  MUX \Data_Mem/U8136  ( .A(\Data_Mem/n8105 ), .B(\Data_Mem/n8102 ), .S(N27), 
        .Z(\Data_Mem/n8106 ) );
  MUX \Data_Mem/U8135  ( .A(\Data_Mem/n8104 ), .B(\Data_Mem/n8103 ), .S(N28), 
        .Z(\Data_Mem/n8105 ) );
  MUX \Data_Mem/U8134  ( .A(data_mem_out_wire[541]), .B(data_mem_out_wire[573]), .S(N29), .Z(\Data_Mem/n8104 ) );
  MUX \Data_Mem/U8133  ( .A(data_mem_out_wire[605]), .B(data_mem_out_wire[637]), .S(N29), .Z(\Data_Mem/n8103 ) );
  MUX \Data_Mem/U8132  ( .A(\Data_Mem/n8101 ), .B(\Data_Mem/n8100 ), .S(N28), 
        .Z(\Data_Mem/n8102 ) );
  MUX \Data_Mem/U8131  ( .A(data_mem_out_wire[669]), .B(data_mem_out_wire[701]), .S(N29), .Z(\Data_Mem/n8101 ) );
  MUX \Data_Mem/U8130  ( .A(data_mem_out_wire[733]), .B(data_mem_out_wire[765]), .S(N29), .Z(\Data_Mem/n8100 ) );
  MUX \Data_Mem/U8129  ( .A(\Data_Mem/n8098 ), .B(\Data_Mem/n8095 ), .S(N27), 
        .Z(\Data_Mem/n8099 ) );
  MUX \Data_Mem/U8128  ( .A(\Data_Mem/n8097 ), .B(\Data_Mem/n8096 ), .S(N28), 
        .Z(\Data_Mem/n8098 ) );
  MUX \Data_Mem/U8127  ( .A(data_mem_out_wire[797]), .B(data_mem_out_wire[829]), .S(N29), .Z(\Data_Mem/n8097 ) );
  MUX \Data_Mem/U8126  ( .A(data_mem_out_wire[861]), .B(data_mem_out_wire[893]), .S(N29), .Z(\Data_Mem/n8096 ) );
  MUX \Data_Mem/U8125  ( .A(\Data_Mem/n8094 ), .B(\Data_Mem/n8093 ), .S(N28), 
        .Z(\Data_Mem/n8095 ) );
  MUX \Data_Mem/U8124  ( .A(data_mem_out_wire[925]), .B(data_mem_out_wire[957]), .S(N29), .Z(\Data_Mem/n8094 ) );
  MUX \Data_Mem/U8123  ( .A(data_mem_out_wire[989]), .B(
        data_mem_out_wire[1021]), .S(N29), .Z(\Data_Mem/n8093 ) );
  MUX \Data_Mem/U8122  ( .A(\Data_Mem/n8091 ), .B(\Data_Mem/n8076 ), .S(N25), 
        .Z(\Data_Mem/n8092 ) );
  MUX \Data_Mem/U8121  ( .A(\Data_Mem/n8090 ), .B(\Data_Mem/n8083 ), .S(N26), 
        .Z(\Data_Mem/n8091 ) );
  MUX \Data_Mem/U8120  ( .A(\Data_Mem/n8089 ), .B(\Data_Mem/n8086 ), .S(N27), 
        .Z(\Data_Mem/n8090 ) );
  MUX \Data_Mem/U8119  ( .A(\Data_Mem/n8088 ), .B(\Data_Mem/n8087 ), .S(N28), 
        .Z(\Data_Mem/n8089 ) );
  MUX \Data_Mem/U8118  ( .A(data_mem_out_wire[1053]), .B(
        data_mem_out_wire[1085]), .S(N29), .Z(\Data_Mem/n8088 ) );
  MUX \Data_Mem/U8117  ( .A(data_mem_out_wire[1117]), .B(
        data_mem_out_wire[1149]), .S(N29), .Z(\Data_Mem/n8087 ) );
  MUX \Data_Mem/U8116  ( .A(\Data_Mem/n8085 ), .B(\Data_Mem/n8084 ), .S(N28), 
        .Z(\Data_Mem/n8086 ) );
  MUX \Data_Mem/U8115  ( .A(data_mem_out_wire[1181]), .B(
        data_mem_out_wire[1213]), .S(N29), .Z(\Data_Mem/n8085 ) );
  MUX \Data_Mem/U8114  ( .A(data_mem_out_wire[1245]), .B(
        data_mem_out_wire[1277]), .S(N29), .Z(\Data_Mem/n8084 ) );
  MUX \Data_Mem/U8113  ( .A(\Data_Mem/n8082 ), .B(\Data_Mem/n8079 ), .S(N27), 
        .Z(\Data_Mem/n8083 ) );
  MUX \Data_Mem/U8112  ( .A(\Data_Mem/n8081 ), .B(\Data_Mem/n8080 ), .S(N28), 
        .Z(\Data_Mem/n8082 ) );
  MUX \Data_Mem/U8111  ( .A(data_mem_out_wire[1309]), .B(
        data_mem_out_wire[1341]), .S(N29), .Z(\Data_Mem/n8081 ) );
  MUX \Data_Mem/U8110  ( .A(data_mem_out_wire[1373]), .B(
        data_mem_out_wire[1405]), .S(N29), .Z(\Data_Mem/n8080 ) );
  MUX \Data_Mem/U8109  ( .A(\Data_Mem/n8078 ), .B(\Data_Mem/n8077 ), .S(N28), 
        .Z(\Data_Mem/n8079 ) );
  MUX \Data_Mem/U8108  ( .A(data_mem_out_wire[1437]), .B(
        data_mem_out_wire[1469]), .S(N29), .Z(\Data_Mem/n8078 ) );
  MUX \Data_Mem/U8107  ( .A(data_mem_out_wire[1501]), .B(
        data_mem_out_wire[1533]), .S(N29), .Z(\Data_Mem/n8077 ) );
  MUX \Data_Mem/U8106  ( .A(\Data_Mem/n8075 ), .B(\Data_Mem/n8068 ), .S(N26), 
        .Z(\Data_Mem/n8076 ) );
  MUX \Data_Mem/U8105  ( .A(\Data_Mem/n8074 ), .B(\Data_Mem/n8071 ), .S(N27), 
        .Z(\Data_Mem/n8075 ) );
  MUX \Data_Mem/U8104  ( .A(\Data_Mem/n8073 ), .B(\Data_Mem/n8072 ), .S(N28), 
        .Z(\Data_Mem/n8074 ) );
  MUX \Data_Mem/U8103  ( .A(data_mem_out_wire[1565]), .B(
        data_mem_out_wire[1597]), .S(N29), .Z(\Data_Mem/n8073 ) );
  MUX \Data_Mem/U8102  ( .A(data_mem_out_wire[1629]), .B(
        data_mem_out_wire[1661]), .S(N29), .Z(\Data_Mem/n8072 ) );
  MUX \Data_Mem/U8101  ( .A(\Data_Mem/n8070 ), .B(\Data_Mem/n8069 ), .S(N28), 
        .Z(\Data_Mem/n8071 ) );
  MUX \Data_Mem/U8100  ( .A(data_mem_out_wire[1693]), .B(
        data_mem_out_wire[1725]), .S(N29), .Z(\Data_Mem/n8070 ) );
  MUX \Data_Mem/U8099  ( .A(data_mem_out_wire[1757]), .B(
        data_mem_out_wire[1789]), .S(N29), .Z(\Data_Mem/n8069 ) );
  MUX \Data_Mem/U8098  ( .A(\Data_Mem/n8067 ), .B(\Data_Mem/n8064 ), .S(N27), 
        .Z(\Data_Mem/n8068 ) );
  MUX \Data_Mem/U8097  ( .A(\Data_Mem/n8066 ), .B(\Data_Mem/n8065 ), .S(N28), 
        .Z(\Data_Mem/n8067 ) );
  MUX \Data_Mem/U8096  ( .A(data_mem_out_wire[1821]), .B(
        data_mem_out_wire[1853]), .S(N29), .Z(\Data_Mem/n8066 ) );
  MUX \Data_Mem/U8095  ( .A(data_mem_out_wire[1885]), .B(
        data_mem_out_wire[1917]), .S(N29), .Z(\Data_Mem/n8065 ) );
  MUX \Data_Mem/U8094  ( .A(\Data_Mem/n8063 ), .B(\Data_Mem/n8062 ), .S(N28), 
        .Z(\Data_Mem/n8064 ) );
  MUX \Data_Mem/U8093  ( .A(data_mem_out_wire[1949]), .B(
        data_mem_out_wire[1981]), .S(N29), .Z(\Data_Mem/n8063 ) );
  MUX \Data_Mem/U8092  ( .A(data_mem_out_wire[2013]), .B(
        data_mem_out_wire[2045]), .S(N29), .Z(\Data_Mem/n8062 ) );
  MUX \Data_Mem/U8091  ( .A(\Data_Mem/n8061 ), .B(\Data_Mem/n8030 ), .S(N24), 
        .Z(c_memory[28]) );
  MUX \Data_Mem/U8090  ( .A(\Data_Mem/n8060 ), .B(\Data_Mem/n8045 ), .S(N25), 
        .Z(\Data_Mem/n8061 ) );
  MUX \Data_Mem/U8089  ( .A(\Data_Mem/n8059 ), .B(\Data_Mem/n8052 ), .S(N26), 
        .Z(\Data_Mem/n8060 ) );
  MUX \Data_Mem/U8088  ( .A(\Data_Mem/n8058 ), .B(\Data_Mem/n8055 ), .S(N27), 
        .Z(\Data_Mem/n8059 ) );
  MUX \Data_Mem/U8087  ( .A(\Data_Mem/n8057 ), .B(\Data_Mem/n8056 ), .S(N28), 
        .Z(\Data_Mem/n8058 ) );
  MUX \Data_Mem/U8086  ( .A(data_mem_out_wire[28]), .B(data_mem_out_wire[60]), 
        .S(N29), .Z(\Data_Mem/n8057 ) );
  MUX \Data_Mem/U8085  ( .A(data_mem_out_wire[92]), .B(data_mem_out_wire[124]), 
        .S(N29), .Z(\Data_Mem/n8056 ) );
  MUX \Data_Mem/U8084  ( .A(\Data_Mem/n8054 ), .B(\Data_Mem/n8053 ), .S(N28), 
        .Z(\Data_Mem/n8055 ) );
  MUX \Data_Mem/U8083  ( .A(data_mem_out_wire[156]), .B(data_mem_out_wire[188]), .S(N29), .Z(\Data_Mem/n8054 ) );
  MUX \Data_Mem/U8082  ( .A(data_mem_out_wire[220]), .B(data_mem_out_wire[252]), .S(N29), .Z(\Data_Mem/n8053 ) );
  MUX \Data_Mem/U8081  ( .A(\Data_Mem/n8051 ), .B(\Data_Mem/n8048 ), .S(N27), 
        .Z(\Data_Mem/n8052 ) );
  MUX \Data_Mem/U8080  ( .A(\Data_Mem/n8050 ), .B(\Data_Mem/n8049 ), .S(N28), 
        .Z(\Data_Mem/n8051 ) );
  MUX \Data_Mem/U8079  ( .A(data_mem_out_wire[284]), .B(data_mem_out_wire[316]), .S(N29), .Z(\Data_Mem/n8050 ) );
  MUX \Data_Mem/U8078  ( .A(data_mem_out_wire[348]), .B(data_mem_out_wire[380]), .S(N29), .Z(\Data_Mem/n8049 ) );
  MUX \Data_Mem/U8077  ( .A(\Data_Mem/n8047 ), .B(\Data_Mem/n8046 ), .S(N28), 
        .Z(\Data_Mem/n8048 ) );
  MUX \Data_Mem/U8076  ( .A(data_mem_out_wire[412]), .B(data_mem_out_wire[444]), .S(N29), .Z(\Data_Mem/n8047 ) );
  MUX \Data_Mem/U8075  ( .A(data_mem_out_wire[476]), .B(data_mem_out_wire[508]), .S(N29), .Z(\Data_Mem/n8046 ) );
  MUX \Data_Mem/U8074  ( .A(\Data_Mem/n8044 ), .B(\Data_Mem/n8037 ), .S(N26), 
        .Z(\Data_Mem/n8045 ) );
  MUX \Data_Mem/U8073  ( .A(\Data_Mem/n8043 ), .B(\Data_Mem/n8040 ), .S(N27), 
        .Z(\Data_Mem/n8044 ) );
  MUX \Data_Mem/U8072  ( .A(\Data_Mem/n8042 ), .B(\Data_Mem/n8041 ), .S(N28), 
        .Z(\Data_Mem/n8043 ) );
  MUX \Data_Mem/U8071  ( .A(data_mem_out_wire[540]), .B(data_mem_out_wire[572]), .S(N29), .Z(\Data_Mem/n8042 ) );
  MUX \Data_Mem/U8070  ( .A(data_mem_out_wire[604]), .B(data_mem_out_wire[636]), .S(N29), .Z(\Data_Mem/n8041 ) );
  MUX \Data_Mem/U8069  ( .A(\Data_Mem/n8039 ), .B(\Data_Mem/n8038 ), .S(N28), 
        .Z(\Data_Mem/n8040 ) );
  MUX \Data_Mem/U8068  ( .A(data_mem_out_wire[668]), .B(data_mem_out_wire[700]), .S(N29), .Z(\Data_Mem/n8039 ) );
  MUX \Data_Mem/U8067  ( .A(data_mem_out_wire[732]), .B(data_mem_out_wire[764]), .S(N29), .Z(\Data_Mem/n8038 ) );
  MUX \Data_Mem/U8066  ( .A(\Data_Mem/n8036 ), .B(\Data_Mem/n8033 ), .S(N27), 
        .Z(\Data_Mem/n8037 ) );
  MUX \Data_Mem/U8065  ( .A(\Data_Mem/n8035 ), .B(\Data_Mem/n8034 ), .S(N28), 
        .Z(\Data_Mem/n8036 ) );
  MUX \Data_Mem/U8064  ( .A(data_mem_out_wire[796]), .B(data_mem_out_wire[828]), .S(N29), .Z(\Data_Mem/n8035 ) );
  MUX \Data_Mem/U8063  ( .A(data_mem_out_wire[860]), .B(data_mem_out_wire[892]), .S(N29), .Z(\Data_Mem/n8034 ) );
  MUX \Data_Mem/U8062  ( .A(\Data_Mem/n8032 ), .B(\Data_Mem/n8031 ), .S(N28), 
        .Z(\Data_Mem/n8033 ) );
  MUX \Data_Mem/U8061  ( .A(data_mem_out_wire[924]), .B(data_mem_out_wire[956]), .S(N29), .Z(\Data_Mem/n8032 ) );
  MUX \Data_Mem/U8060  ( .A(data_mem_out_wire[988]), .B(
        data_mem_out_wire[1020]), .S(N29), .Z(\Data_Mem/n8031 ) );
  MUX \Data_Mem/U8059  ( .A(\Data_Mem/n8029 ), .B(\Data_Mem/n8014 ), .S(N25), 
        .Z(\Data_Mem/n8030 ) );
  MUX \Data_Mem/U8058  ( .A(\Data_Mem/n8028 ), .B(\Data_Mem/n8021 ), .S(N26), 
        .Z(\Data_Mem/n8029 ) );
  MUX \Data_Mem/U8057  ( .A(\Data_Mem/n8027 ), .B(\Data_Mem/n8024 ), .S(N27), 
        .Z(\Data_Mem/n8028 ) );
  MUX \Data_Mem/U8056  ( .A(\Data_Mem/n8026 ), .B(\Data_Mem/n8025 ), .S(N28), 
        .Z(\Data_Mem/n8027 ) );
  MUX \Data_Mem/U8055  ( .A(data_mem_out_wire[1052]), .B(
        data_mem_out_wire[1084]), .S(N29), .Z(\Data_Mem/n8026 ) );
  MUX \Data_Mem/U8054  ( .A(data_mem_out_wire[1116]), .B(
        data_mem_out_wire[1148]), .S(N29), .Z(\Data_Mem/n8025 ) );
  MUX \Data_Mem/U8053  ( .A(\Data_Mem/n8023 ), .B(\Data_Mem/n8022 ), .S(N28), 
        .Z(\Data_Mem/n8024 ) );
  MUX \Data_Mem/U8052  ( .A(data_mem_out_wire[1180]), .B(
        data_mem_out_wire[1212]), .S(N29), .Z(\Data_Mem/n8023 ) );
  MUX \Data_Mem/U8051  ( .A(data_mem_out_wire[1244]), .B(
        data_mem_out_wire[1276]), .S(N29), .Z(\Data_Mem/n8022 ) );
  MUX \Data_Mem/U8050  ( .A(\Data_Mem/n8020 ), .B(\Data_Mem/n8017 ), .S(N27), 
        .Z(\Data_Mem/n8021 ) );
  MUX \Data_Mem/U8049  ( .A(\Data_Mem/n8019 ), .B(\Data_Mem/n8018 ), .S(N28), 
        .Z(\Data_Mem/n8020 ) );
  MUX \Data_Mem/U8048  ( .A(data_mem_out_wire[1308]), .B(
        data_mem_out_wire[1340]), .S(N29), .Z(\Data_Mem/n8019 ) );
  MUX \Data_Mem/U8047  ( .A(data_mem_out_wire[1372]), .B(
        data_mem_out_wire[1404]), .S(N29), .Z(\Data_Mem/n8018 ) );
  MUX \Data_Mem/U8046  ( .A(\Data_Mem/n8016 ), .B(\Data_Mem/n8015 ), .S(N28), 
        .Z(\Data_Mem/n8017 ) );
  MUX \Data_Mem/U8045  ( .A(data_mem_out_wire[1436]), .B(
        data_mem_out_wire[1468]), .S(N29), .Z(\Data_Mem/n8016 ) );
  MUX \Data_Mem/U8044  ( .A(data_mem_out_wire[1500]), .B(
        data_mem_out_wire[1532]), .S(N29), .Z(\Data_Mem/n8015 ) );
  MUX \Data_Mem/U8043  ( .A(\Data_Mem/n8013 ), .B(\Data_Mem/n8006 ), .S(N26), 
        .Z(\Data_Mem/n8014 ) );
  MUX \Data_Mem/U8042  ( .A(\Data_Mem/n8012 ), .B(\Data_Mem/n8009 ), .S(N27), 
        .Z(\Data_Mem/n8013 ) );
  MUX \Data_Mem/U8041  ( .A(\Data_Mem/n8011 ), .B(\Data_Mem/n8010 ), .S(N28), 
        .Z(\Data_Mem/n8012 ) );
  MUX \Data_Mem/U8040  ( .A(data_mem_out_wire[1564]), .B(
        data_mem_out_wire[1596]), .S(N29), .Z(\Data_Mem/n8011 ) );
  MUX \Data_Mem/U8039  ( .A(data_mem_out_wire[1628]), .B(
        data_mem_out_wire[1660]), .S(N29), .Z(\Data_Mem/n8010 ) );
  MUX \Data_Mem/U8038  ( .A(\Data_Mem/n8008 ), .B(\Data_Mem/n8007 ), .S(N28), 
        .Z(\Data_Mem/n8009 ) );
  MUX \Data_Mem/U8037  ( .A(data_mem_out_wire[1692]), .B(
        data_mem_out_wire[1724]), .S(N29), .Z(\Data_Mem/n8008 ) );
  MUX \Data_Mem/U8036  ( .A(data_mem_out_wire[1756]), .B(
        data_mem_out_wire[1788]), .S(N29), .Z(\Data_Mem/n8007 ) );
  MUX \Data_Mem/U8035  ( .A(\Data_Mem/n8005 ), .B(\Data_Mem/n8002 ), .S(N27), 
        .Z(\Data_Mem/n8006 ) );
  MUX \Data_Mem/U8034  ( .A(\Data_Mem/n8004 ), .B(\Data_Mem/n8003 ), .S(N28), 
        .Z(\Data_Mem/n8005 ) );
  MUX \Data_Mem/U8033  ( .A(data_mem_out_wire[1820]), .B(
        data_mem_out_wire[1852]), .S(N29), .Z(\Data_Mem/n8004 ) );
  MUX \Data_Mem/U8032  ( .A(data_mem_out_wire[1884]), .B(
        data_mem_out_wire[1916]), .S(N29), .Z(\Data_Mem/n8003 ) );
  MUX \Data_Mem/U8031  ( .A(\Data_Mem/n8001 ), .B(\Data_Mem/n8000 ), .S(N28), 
        .Z(\Data_Mem/n8002 ) );
  MUX \Data_Mem/U8030  ( .A(data_mem_out_wire[1948]), .B(
        data_mem_out_wire[1980]), .S(N29), .Z(\Data_Mem/n8001 ) );
  MUX \Data_Mem/U8029  ( .A(data_mem_out_wire[2012]), .B(
        data_mem_out_wire[2044]), .S(N29), .Z(\Data_Mem/n8000 ) );
  MUX \Data_Mem/U8028  ( .A(\Data_Mem/n7999 ), .B(\Data_Mem/n7968 ), .S(N24), 
        .Z(c_memory[27]) );
  MUX \Data_Mem/U8027  ( .A(\Data_Mem/n7998 ), .B(\Data_Mem/n7983 ), .S(N25), 
        .Z(\Data_Mem/n7999 ) );
  MUX \Data_Mem/U8026  ( .A(\Data_Mem/n7997 ), .B(\Data_Mem/n7990 ), .S(N26), 
        .Z(\Data_Mem/n7998 ) );
  MUX \Data_Mem/U8025  ( .A(\Data_Mem/n7996 ), .B(\Data_Mem/n7993 ), .S(N27), 
        .Z(\Data_Mem/n7997 ) );
  MUX \Data_Mem/U8024  ( .A(\Data_Mem/n7995 ), .B(\Data_Mem/n7994 ), .S(N28), 
        .Z(\Data_Mem/n7996 ) );
  MUX \Data_Mem/U8023  ( .A(data_mem_out_wire[27]), .B(data_mem_out_wire[59]), 
        .S(N29), .Z(\Data_Mem/n7995 ) );
  MUX \Data_Mem/U8022  ( .A(data_mem_out_wire[91]), .B(data_mem_out_wire[123]), 
        .S(N29), .Z(\Data_Mem/n7994 ) );
  MUX \Data_Mem/U8021  ( .A(\Data_Mem/n7992 ), .B(\Data_Mem/n7991 ), .S(N28), 
        .Z(\Data_Mem/n7993 ) );
  MUX \Data_Mem/U8020  ( .A(data_mem_out_wire[155]), .B(data_mem_out_wire[187]), .S(N29), .Z(\Data_Mem/n7992 ) );
  MUX \Data_Mem/U8019  ( .A(data_mem_out_wire[219]), .B(data_mem_out_wire[251]), .S(N29), .Z(\Data_Mem/n7991 ) );
  MUX \Data_Mem/U8018  ( .A(\Data_Mem/n7989 ), .B(\Data_Mem/n7986 ), .S(N27), 
        .Z(\Data_Mem/n7990 ) );
  MUX \Data_Mem/U8017  ( .A(\Data_Mem/n7988 ), .B(\Data_Mem/n7987 ), .S(N28), 
        .Z(\Data_Mem/n7989 ) );
  MUX \Data_Mem/U8016  ( .A(data_mem_out_wire[283]), .B(data_mem_out_wire[315]), .S(N29), .Z(\Data_Mem/n7988 ) );
  MUX \Data_Mem/U8015  ( .A(data_mem_out_wire[347]), .B(data_mem_out_wire[379]), .S(N29), .Z(\Data_Mem/n7987 ) );
  MUX \Data_Mem/U8014  ( .A(\Data_Mem/n7985 ), .B(\Data_Mem/n7984 ), .S(N28), 
        .Z(\Data_Mem/n7986 ) );
  MUX \Data_Mem/U8013  ( .A(data_mem_out_wire[411]), .B(data_mem_out_wire[443]), .S(N29), .Z(\Data_Mem/n7985 ) );
  MUX \Data_Mem/U8012  ( .A(data_mem_out_wire[475]), .B(data_mem_out_wire[507]), .S(N29), .Z(\Data_Mem/n7984 ) );
  MUX \Data_Mem/U8011  ( .A(\Data_Mem/n7982 ), .B(\Data_Mem/n7975 ), .S(N26), 
        .Z(\Data_Mem/n7983 ) );
  MUX \Data_Mem/U8010  ( .A(\Data_Mem/n7981 ), .B(\Data_Mem/n7978 ), .S(N27), 
        .Z(\Data_Mem/n7982 ) );
  MUX \Data_Mem/U8009  ( .A(\Data_Mem/n7980 ), .B(\Data_Mem/n7979 ), .S(N28), 
        .Z(\Data_Mem/n7981 ) );
  MUX \Data_Mem/U8008  ( .A(data_mem_out_wire[539]), .B(data_mem_out_wire[571]), .S(N29), .Z(\Data_Mem/n7980 ) );
  MUX \Data_Mem/U8007  ( .A(data_mem_out_wire[603]), .B(data_mem_out_wire[635]), .S(N29), .Z(\Data_Mem/n7979 ) );
  MUX \Data_Mem/U8006  ( .A(\Data_Mem/n7977 ), .B(\Data_Mem/n7976 ), .S(N28), 
        .Z(\Data_Mem/n7978 ) );
  MUX \Data_Mem/U8005  ( .A(data_mem_out_wire[667]), .B(data_mem_out_wire[699]), .S(N29), .Z(\Data_Mem/n7977 ) );
  MUX \Data_Mem/U8004  ( .A(data_mem_out_wire[731]), .B(data_mem_out_wire[763]), .S(N29), .Z(\Data_Mem/n7976 ) );
  MUX \Data_Mem/U8003  ( .A(\Data_Mem/n7974 ), .B(\Data_Mem/n7971 ), .S(N27), 
        .Z(\Data_Mem/n7975 ) );
  MUX \Data_Mem/U8002  ( .A(\Data_Mem/n7973 ), .B(\Data_Mem/n7972 ), .S(N28), 
        .Z(\Data_Mem/n7974 ) );
  MUX \Data_Mem/U8001  ( .A(data_mem_out_wire[795]), .B(data_mem_out_wire[827]), .S(N29), .Z(\Data_Mem/n7973 ) );
  MUX \Data_Mem/U8000  ( .A(data_mem_out_wire[859]), .B(data_mem_out_wire[891]), .S(N29), .Z(\Data_Mem/n7972 ) );
  MUX \Data_Mem/U7999  ( .A(\Data_Mem/n7970 ), .B(\Data_Mem/n7969 ), .S(N28), 
        .Z(\Data_Mem/n7971 ) );
  MUX \Data_Mem/U7998  ( .A(data_mem_out_wire[923]), .B(data_mem_out_wire[955]), .S(N29), .Z(\Data_Mem/n7970 ) );
  MUX \Data_Mem/U7997  ( .A(data_mem_out_wire[987]), .B(
        data_mem_out_wire[1019]), .S(N29), .Z(\Data_Mem/n7969 ) );
  MUX \Data_Mem/U7996  ( .A(\Data_Mem/n7967 ), .B(\Data_Mem/n7952 ), .S(N25), 
        .Z(\Data_Mem/n7968 ) );
  MUX \Data_Mem/U7995  ( .A(\Data_Mem/n7966 ), .B(\Data_Mem/n7959 ), .S(N26), 
        .Z(\Data_Mem/n7967 ) );
  MUX \Data_Mem/U7994  ( .A(\Data_Mem/n7965 ), .B(\Data_Mem/n7962 ), .S(N27), 
        .Z(\Data_Mem/n7966 ) );
  MUX \Data_Mem/U7993  ( .A(\Data_Mem/n7964 ), .B(\Data_Mem/n7963 ), .S(N28), 
        .Z(\Data_Mem/n7965 ) );
  MUX \Data_Mem/U7992  ( .A(data_mem_out_wire[1051]), .B(
        data_mem_out_wire[1083]), .S(N29), .Z(\Data_Mem/n7964 ) );
  MUX \Data_Mem/U7991  ( .A(data_mem_out_wire[1115]), .B(
        data_mem_out_wire[1147]), .S(N29), .Z(\Data_Mem/n7963 ) );
  MUX \Data_Mem/U7990  ( .A(\Data_Mem/n7961 ), .B(\Data_Mem/n7960 ), .S(N28), 
        .Z(\Data_Mem/n7962 ) );
  MUX \Data_Mem/U7989  ( .A(data_mem_out_wire[1179]), .B(
        data_mem_out_wire[1211]), .S(N29), .Z(\Data_Mem/n7961 ) );
  MUX \Data_Mem/U7988  ( .A(data_mem_out_wire[1243]), .B(
        data_mem_out_wire[1275]), .S(N29), .Z(\Data_Mem/n7960 ) );
  MUX \Data_Mem/U7987  ( .A(\Data_Mem/n7958 ), .B(\Data_Mem/n7955 ), .S(N27), 
        .Z(\Data_Mem/n7959 ) );
  MUX \Data_Mem/U7986  ( .A(\Data_Mem/n7957 ), .B(\Data_Mem/n7956 ), .S(N28), 
        .Z(\Data_Mem/n7958 ) );
  MUX \Data_Mem/U7985  ( .A(data_mem_out_wire[1307]), .B(
        data_mem_out_wire[1339]), .S(N29), .Z(\Data_Mem/n7957 ) );
  MUX \Data_Mem/U7984  ( .A(data_mem_out_wire[1371]), .B(
        data_mem_out_wire[1403]), .S(N29), .Z(\Data_Mem/n7956 ) );
  MUX \Data_Mem/U7983  ( .A(\Data_Mem/n7954 ), .B(\Data_Mem/n7953 ), .S(N28), 
        .Z(\Data_Mem/n7955 ) );
  MUX \Data_Mem/U7982  ( .A(data_mem_out_wire[1435]), .B(
        data_mem_out_wire[1467]), .S(N29), .Z(\Data_Mem/n7954 ) );
  MUX \Data_Mem/U7981  ( .A(data_mem_out_wire[1499]), .B(
        data_mem_out_wire[1531]), .S(N29), .Z(\Data_Mem/n7953 ) );
  MUX \Data_Mem/U7980  ( .A(\Data_Mem/n7951 ), .B(\Data_Mem/n7944 ), .S(N26), 
        .Z(\Data_Mem/n7952 ) );
  MUX \Data_Mem/U7979  ( .A(\Data_Mem/n7950 ), .B(\Data_Mem/n7947 ), .S(N27), 
        .Z(\Data_Mem/n7951 ) );
  MUX \Data_Mem/U7978  ( .A(\Data_Mem/n7949 ), .B(\Data_Mem/n7948 ), .S(N28), 
        .Z(\Data_Mem/n7950 ) );
  MUX \Data_Mem/U7977  ( .A(data_mem_out_wire[1563]), .B(
        data_mem_out_wire[1595]), .S(N29), .Z(\Data_Mem/n7949 ) );
  MUX \Data_Mem/U7976  ( .A(data_mem_out_wire[1627]), .B(
        data_mem_out_wire[1659]), .S(N29), .Z(\Data_Mem/n7948 ) );
  MUX \Data_Mem/U7975  ( .A(\Data_Mem/n7946 ), .B(\Data_Mem/n7945 ), .S(N28), 
        .Z(\Data_Mem/n7947 ) );
  MUX \Data_Mem/U7974  ( .A(data_mem_out_wire[1691]), .B(
        data_mem_out_wire[1723]), .S(N29), .Z(\Data_Mem/n7946 ) );
  MUX \Data_Mem/U7973  ( .A(data_mem_out_wire[1755]), .B(
        data_mem_out_wire[1787]), .S(N29), .Z(\Data_Mem/n7945 ) );
  MUX \Data_Mem/U7972  ( .A(\Data_Mem/n7943 ), .B(\Data_Mem/n7940 ), .S(N27), 
        .Z(\Data_Mem/n7944 ) );
  MUX \Data_Mem/U7971  ( .A(\Data_Mem/n7942 ), .B(\Data_Mem/n7941 ), .S(N28), 
        .Z(\Data_Mem/n7943 ) );
  MUX \Data_Mem/U7970  ( .A(data_mem_out_wire[1819]), .B(
        data_mem_out_wire[1851]), .S(N29), .Z(\Data_Mem/n7942 ) );
  MUX \Data_Mem/U7969  ( .A(data_mem_out_wire[1883]), .B(
        data_mem_out_wire[1915]), .S(N29), .Z(\Data_Mem/n7941 ) );
  MUX \Data_Mem/U7968  ( .A(\Data_Mem/n7939 ), .B(\Data_Mem/n7938 ), .S(N28), 
        .Z(\Data_Mem/n7940 ) );
  MUX \Data_Mem/U7967  ( .A(data_mem_out_wire[1947]), .B(
        data_mem_out_wire[1979]), .S(N29), .Z(\Data_Mem/n7939 ) );
  MUX \Data_Mem/U7966  ( .A(data_mem_out_wire[2011]), .B(
        data_mem_out_wire[2043]), .S(N29), .Z(\Data_Mem/n7938 ) );
  MUX \Data_Mem/U7965  ( .A(\Data_Mem/n7937 ), .B(\Data_Mem/n7906 ), .S(N24), 
        .Z(c_memory[26]) );
  MUX \Data_Mem/U7964  ( .A(\Data_Mem/n7936 ), .B(\Data_Mem/n7921 ), .S(N25), 
        .Z(\Data_Mem/n7937 ) );
  MUX \Data_Mem/U7963  ( .A(\Data_Mem/n7935 ), .B(\Data_Mem/n7928 ), .S(N26), 
        .Z(\Data_Mem/n7936 ) );
  MUX \Data_Mem/U7962  ( .A(\Data_Mem/n7934 ), .B(\Data_Mem/n7931 ), .S(N27), 
        .Z(\Data_Mem/n7935 ) );
  MUX \Data_Mem/U7961  ( .A(\Data_Mem/n7933 ), .B(\Data_Mem/n7932 ), .S(N28), 
        .Z(\Data_Mem/n7934 ) );
  MUX \Data_Mem/U7960  ( .A(data_mem_out_wire[26]), .B(data_mem_out_wire[58]), 
        .S(N29), .Z(\Data_Mem/n7933 ) );
  MUX \Data_Mem/U7959  ( .A(data_mem_out_wire[90]), .B(data_mem_out_wire[122]), 
        .S(N29), .Z(\Data_Mem/n7932 ) );
  MUX \Data_Mem/U7958  ( .A(\Data_Mem/n7930 ), .B(\Data_Mem/n7929 ), .S(N28), 
        .Z(\Data_Mem/n7931 ) );
  MUX \Data_Mem/U7957  ( .A(data_mem_out_wire[154]), .B(data_mem_out_wire[186]), .S(N29), .Z(\Data_Mem/n7930 ) );
  MUX \Data_Mem/U7956  ( .A(data_mem_out_wire[218]), .B(data_mem_out_wire[250]), .S(N29), .Z(\Data_Mem/n7929 ) );
  MUX \Data_Mem/U7955  ( .A(\Data_Mem/n7927 ), .B(\Data_Mem/n7924 ), .S(N27), 
        .Z(\Data_Mem/n7928 ) );
  MUX \Data_Mem/U7954  ( .A(\Data_Mem/n7926 ), .B(\Data_Mem/n7925 ), .S(N28), 
        .Z(\Data_Mem/n7927 ) );
  MUX \Data_Mem/U7953  ( .A(data_mem_out_wire[282]), .B(data_mem_out_wire[314]), .S(N29), .Z(\Data_Mem/n7926 ) );
  MUX \Data_Mem/U7952  ( .A(data_mem_out_wire[346]), .B(data_mem_out_wire[378]), .S(N29), .Z(\Data_Mem/n7925 ) );
  MUX \Data_Mem/U7951  ( .A(\Data_Mem/n7923 ), .B(\Data_Mem/n7922 ), .S(N28), 
        .Z(\Data_Mem/n7924 ) );
  MUX \Data_Mem/U7950  ( .A(data_mem_out_wire[410]), .B(data_mem_out_wire[442]), .S(N29), .Z(\Data_Mem/n7923 ) );
  MUX \Data_Mem/U7949  ( .A(data_mem_out_wire[474]), .B(data_mem_out_wire[506]), .S(N29), .Z(\Data_Mem/n7922 ) );
  MUX \Data_Mem/U7948  ( .A(\Data_Mem/n7920 ), .B(\Data_Mem/n7913 ), .S(N26), 
        .Z(\Data_Mem/n7921 ) );
  MUX \Data_Mem/U7947  ( .A(\Data_Mem/n7919 ), .B(\Data_Mem/n7916 ), .S(N27), 
        .Z(\Data_Mem/n7920 ) );
  MUX \Data_Mem/U7946  ( .A(\Data_Mem/n7918 ), .B(\Data_Mem/n7917 ), .S(N28), 
        .Z(\Data_Mem/n7919 ) );
  MUX \Data_Mem/U7945  ( .A(data_mem_out_wire[538]), .B(data_mem_out_wire[570]), .S(N29), .Z(\Data_Mem/n7918 ) );
  MUX \Data_Mem/U7944  ( .A(data_mem_out_wire[602]), .B(data_mem_out_wire[634]), .S(N29), .Z(\Data_Mem/n7917 ) );
  MUX \Data_Mem/U7943  ( .A(\Data_Mem/n7915 ), .B(\Data_Mem/n7914 ), .S(N28), 
        .Z(\Data_Mem/n7916 ) );
  MUX \Data_Mem/U7942  ( .A(data_mem_out_wire[666]), .B(data_mem_out_wire[698]), .S(N29), .Z(\Data_Mem/n7915 ) );
  MUX \Data_Mem/U7941  ( .A(data_mem_out_wire[730]), .B(data_mem_out_wire[762]), .S(N29), .Z(\Data_Mem/n7914 ) );
  MUX \Data_Mem/U7940  ( .A(\Data_Mem/n7912 ), .B(\Data_Mem/n7909 ), .S(N27), 
        .Z(\Data_Mem/n7913 ) );
  MUX \Data_Mem/U7939  ( .A(\Data_Mem/n7911 ), .B(\Data_Mem/n7910 ), .S(N28), 
        .Z(\Data_Mem/n7912 ) );
  MUX \Data_Mem/U7938  ( .A(data_mem_out_wire[794]), .B(data_mem_out_wire[826]), .S(N29), .Z(\Data_Mem/n7911 ) );
  MUX \Data_Mem/U7937  ( .A(data_mem_out_wire[858]), .B(data_mem_out_wire[890]), .S(N29), .Z(\Data_Mem/n7910 ) );
  MUX \Data_Mem/U7936  ( .A(\Data_Mem/n7908 ), .B(\Data_Mem/n7907 ), .S(N28), 
        .Z(\Data_Mem/n7909 ) );
  MUX \Data_Mem/U7935  ( .A(data_mem_out_wire[922]), .B(data_mem_out_wire[954]), .S(N29), .Z(\Data_Mem/n7908 ) );
  MUX \Data_Mem/U7934  ( .A(data_mem_out_wire[986]), .B(
        data_mem_out_wire[1018]), .S(N29), .Z(\Data_Mem/n7907 ) );
  MUX \Data_Mem/U7933  ( .A(\Data_Mem/n7905 ), .B(\Data_Mem/n7890 ), .S(N25), 
        .Z(\Data_Mem/n7906 ) );
  MUX \Data_Mem/U7932  ( .A(\Data_Mem/n7904 ), .B(\Data_Mem/n7897 ), .S(N26), 
        .Z(\Data_Mem/n7905 ) );
  MUX \Data_Mem/U7931  ( .A(\Data_Mem/n7903 ), .B(\Data_Mem/n7900 ), .S(N27), 
        .Z(\Data_Mem/n7904 ) );
  MUX \Data_Mem/U7930  ( .A(\Data_Mem/n7902 ), .B(\Data_Mem/n7901 ), .S(N28), 
        .Z(\Data_Mem/n7903 ) );
  MUX \Data_Mem/U7929  ( .A(data_mem_out_wire[1050]), .B(
        data_mem_out_wire[1082]), .S(N29), .Z(\Data_Mem/n7902 ) );
  MUX \Data_Mem/U7928  ( .A(data_mem_out_wire[1114]), .B(
        data_mem_out_wire[1146]), .S(N29), .Z(\Data_Mem/n7901 ) );
  MUX \Data_Mem/U7927  ( .A(\Data_Mem/n7899 ), .B(\Data_Mem/n7898 ), .S(N28), 
        .Z(\Data_Mem/n7900 ) );
  MUX \Data_Mem/U7926  ( .A(data_mem_out_wire[1178]), .B(
        data_mem_out_wire[1210]), .S(N29), .Z(\Data_Mem/n7899 ) );
  MUX \Data_Mem/U7925  ( .A(data_mem_out_wire[1242]), .B(
        data_mem_out_wire[1274]), .S(N29), .Z(\Data_Mem/n7898 ) );
  MUX \Data_Mem/U7924  ( .A(\Data_Mem/n7896 ), .B(\Data_Mem/n7893 ), .S(N27), 
        .Z(\Data_Mem/n7897 ) );
  MUX \Data_Mem/U7923  ( .A(\Data_Mem/n7895 ), .B(\Data_Mem/n7894 ), .S(N28), 
        .Z(\Data_Mem/n7896 ) );
  MUX \Data_Mem/U7922  ( .A(data_mem_out_wire[1306]), .B(
        data_mem_out_wire[1338]), .S(N29), .Z(\Data_Mem/n7895 ) );
  MUX \Data_Mem/U7921  ( .A(data_mem_out_wire[1370]), .B(
        data_mem_out_wire[1402]), .S(N29), .Z(\Data_Mem/n7894 ) );
  MUX \Data_Mem/U7920  ( .A(\Data_Mem/n7892 ), .B(\Data_Mem/n7891 ), .S(N28), 
        .Z(\Data_Mem/n7893 ) );
  MUX \Data_Mem/U7919  ( .A(data_mem_out_wire[1434]), .B(
        data_mem_out_wire[1466]), .S(N29), .Z(\Data_Mem/n7892 ) );
  MUX \Data_Mem/U7918  ( .A(data_mem_out_wire[1498]), .B(
        data_mem_out_wire[1530]), .S(N29), .Z(\Data_Mem/n7891 ) );
  MUX \Data_Mem/U7917  ( .A(\Data_Mem/n7889 ), .B(\Data_Mem/n7882 ), .S(N26), 
        .Z(\Data_Mem/n7890 ) );
  MUX \Data_Mem/U7916  ( .A(\Data_Mem/n7888 ), .B(\Data_Mem/n7885 ), .S(N27), 
        .Z(\Data_Mem/n7889 ) );
  MUX \Data_Mem/U7915  ( .A(\Data_Mem/n7887 ), .B(\Data_Mem/n7886 ), .S(N28), 
        .Z(\Data_Mem/n7888 ) );
  MUX \Data_Mem/U7914  ( .A(data_mem_out_wire[1562]), .B(
        data_mem_out_wire[1594]), .S(N29), .Z(\Data_Mem/n7887 ) );
  MUX \Data_Mem/U7913  ( .A(data_mem_out_wire[1626]), .B(
        data_mem_out_wire[1658]), .S(N29), .Z(\Data_Mem/n7886 ) );
  MUX \Data_Mem/U7912  ( .A(\Data_Mem/n7884 ), .B(\Data_Mem/n7883 ), .S(N28), 
        .Z(\Data_Mem/n7885 ) );
  MUX \Data_Mem/U7911  ( .A(data_mem_out_wire[1690]), .B(
        data_mem_out_wire[1722]), .S(N29), .Z(\Data_Mem/n7884 ) );
  MUX \Data_Mem/U7910  ( .A(data_mem_out_wire[1754]), .B(
        data_mem_out_wire[1786]), .S(N29), .Z(\Data_Mem/n7883 ) );
  MUX \Data_Mem/U7909  ( .A(\Data_Mem/n7881 ), .B(\Data_Mem/n7878 ), .S(N27), 
        .Z(\Data_Mem/n7882 ) );
  MUX \Data_Mem/U7908  ( .A(\Data_Mem/n7880 ), .B(\Data_Mem/n7879 ), .S(N28), 
        .Z(\Data_Mem/n7881 ) );
  MUX \Data_Mem/U7907  ( .A(data_mem_out_wire[1818]), .B(
        data_mem_out_wire[1850]), .S(N29), .Z(\Data_Mem/n7880 ) );
  MUX \Data_Mem/U7906  ( .A(data_mem_out_wire[1882]), .B(
        data_mem_out_wire[1914]), .S(N29), .Z(\Data_Mem/n7879 ) );
  MUX \Data_Mem/U7905  ( .A(\Data_Mem/n7877 ), .B(\Data_Mem/n7876 ), .S(N28), 
        .Z(\Data_Mem/n7878 ) );
  MUX \Data_Mem/U7904  ( .A(data_mem_out_wire[1946]), .B(
        data_mem_out_wire[1978]), .S(N29), .Z(\Data_Mem/n7877 ) );
  MUX \Data_Mem/U7903  ( .A(data_mem_out_wire[2010]), .B(
        data_mem_out_wire[2042]), .S(N29), .Z(\Data_Mem/n7876 ) );
  MUX \Data_Mem/U7902  ( .A(\Data_Mem/n7875 ), .B(\Data_Mem/n7844 ), .S(N24), 
        .Z(c_memory[25]) );
  MUX \Data_Mem/U7901  ( .A(\Data_Mem/n7874 ), .B(\Data_Mem/n7859 ), .S(N25), 
        .Z(\Data_Mem/n7875 ) );
  MUX \Data_Mem/U7900  ( .A(\Data_Mem/n7873 ), .B(\Data_Mem/n7866 ), .S(N26), 
        .Z(\Data_Mem/n7874 ) );
  MUX \Data_Mem/U7899  ( .A(\Data_Mem/n7872 ), .B(\Data_Mem/n7869 ), .S(N27), 
        .Z(\Data_Mem/n7873 ) );
  MUX \Data_Mem/U7898  ( .A(\Data_Mem/n7871 ), .B(\Data_Mem/n7870 ), .S(N28), 
        .Z(\Data_Mem/n7872 ) );
  MUX \Data_Mem/U7897  ( .A(data_mem_out_wire[25]), .B(data_mem_out_wire[57]), 
        .S(N29), .Z(\Data_Mem/n7871 ) );
  MUX \Data_Mem/U7896  ( .A(data_mem_out_wire[89]), .B(data_mem_out_wire[121]), 
        .S(N29), .Z(\Data_Mem/n7870 ) );
  MUX \Data_Mem/U7895  ( .A(\Data_Mem/n7868 ), .B(\Data_Mem/n7867 ), .S(N28), 
        .Z(\Data_Mem/n7869 ) );
  MUX \Data_Mem/U7894  ( .A(data_mem_out_wire[153]), .B(data_mem_out_wire[185]), .S(N29), .Z(\Data_Mem/n7868 ) );
  MUX \Data_Mem/U7893  ( .A(data_mem_out_wire[217]), .B(data_mem_out_wire[249]), .S(N29), .Z(\Data_Mem/n7867 ) );
  MUX \Data_Mem/U7892  ( .A(\Data_Mem/n7865 ), .B(\Data_Mem/n7862 ), .S(N27), 
        .Z(\Data_Mem/n7866 ) );
  MUX \Data_Mem/U7891  ( .A(\Data_Mem/n7864 ), .B(\Data_Mem/n7863 ), .S(N28), 
        .Z(\Data_Mem/n7865 ) );
  MUX \Data_Mem/U7890  ( .A(data_mem_out_wire[281]), .B(data_mem_out_wire[313]), .S(N29), .Z(\Data_Mem/n7864 ) );
  MUX \Data_Mem/U7889  ( .A(data_mem_out_wire[345]), .B(data_mem_out_wire[377]), .S(N29), .Z(\Data_Mem/n7863 ) );
  MUX \Data_Mem/U7888  ( .A(\Data_Mem/n7861 ), .B(\Data_Mem/n7860 ), .S(N28), 
        .Z(\Data_Mem/n7862 ) );
  MUX \Data_Mem/U7887  ( .A(data_mem_out_wire[409]), .B(data_mem_out_wire[441]), .S(N29), .Z(\Data_Mem/n7861 ) );
  MUX \Data_Mem/U7886  ( .A(data_mem_out_wire[473]), .B(data_mem_out_wire[505]), .S(N29), .Z(\Data_Mem/n7860 ) );
  MUX \Data_Mem/U7885  ( .A(\Data_Mem/n7858 ), .B(\Data_Mem/n7851 ), .S(N26), 
        .Z(\Data_Mem/n7859 ) );
  MUX \Data_Mem/U7884  ( .A(\Data_Mem/n7857 ), .B(\Data_Mem/n7854 ), .S(N27), 
        .Z(\Data_Mem/n7858 ) );
  MUX \Data_Mem/U7883  ( .A(\Data_Mem/n7856 ), .B(\Data_Mem/n7855 ), .S(N28), 
        .Z(\Data_Mem/n7857 ) );
  MUX \Data_Mem/U7882  ( .A(data_mem_out_wire[537]), .B(data_mem_out_wire[569]), .S(N29), .Z(\Data_Mem/n7856 ) );
  MUX \Data_Mem/U7881  ( .A(data_mem_out_wire[601]), .B(data_mem_out_wire[633]), .S(N29), .Z(\Data_Mem/n7855 ) );
  MUX \Data_Mem/U7880  ( .A(\Data_Mem/n7853 ), .B(\Data_Mem/n7852 ), .S(N28), 
        .Z(\Data_Mem/n7854 ) );
  MUX \Data_Mem/U7879  ( .A(data_mem_out_wire[665]), .B(data_mem_out_wire[697]), .S(N29), .Z(\Data_Mem/n7853 ) );
  MUX \Data_Mem/U7878  ( .A(data_mem_out_wire[729]), .B(data_mem_out_wire[761]), .S(N29), .Z(\Data_Mem/n7852 ) );
  MUX \Data_Mem/U7877  ( .A(\Data_Mem/n7850 ), .B(\Data_Mem/n7847 ), .S(N27), 
        .Z(\Data_Mem/n7851 ) );
  MUX \Data_Mem/U7876  ( .A(\Data_Mem/n7849 ), .B(\Data_Mem/n7848 ), .S(N28), 
        .Z(\Data_Mem/n7850 ) );
  MUX \Data_Mem/U7875  ( .A(data_mem_out_wire[793]), .B(data_mem_out_wire[825]), .S(N29), .Z(\Data_Mem/n7849 ) );
  MUX \Data_Mem/U7874  ( .A(data_mem_out_wire[857]), .B(data_mem_out_wire[889]), .S(N29), .Z(\Data_Mem/n7848 ) );
  MUX \Data_Mem/U7873  ( .A(\Data_Mem/n7846 ), .B(\Data_Mem/n7845 ), .S(N28), 
        .Z(\Data_Mem/n7847 ) );
  MUX \Data_Mem/U7872  ( .A(data_mem_out_wire[921]), .B(data_mem_out_wire[953]), .S(N29), .Z(\Data_Mem/n7846 ) );
  MUX \Data_Mem/U7871  ( .A(data_mem_out_wire[985]), .B(
        data_mem_out_wire[1017]), .S(N29), .Z(\Data_Mem/n7845 ) );
  MUX \Data_Mem/U7870  ( .A(\Data_Mem/n7843 ), .B(\Data_Mem/n7828 ), .S(N25), 
        .Z(\Data_Mem/n7844 ) );
  MUX \Data_Mem/U7869  ( .A(\Data_Mem/n7842 ), .B(\Data_Mem/n7835 ), .S(N26), 
        .Z(\Data_Mem/n7843 ) );
  MUX \Data_Mem/U7868  ( .A(\Data_Mem/n7841 ), .B(\Data_Mem/n7838 ), .S(N27), 
        .Z(\Data_Mem/n7842 ) );
  MUX \Data_Mem/U7867  ( .A(\Data_Mem/n7840 ), .B(\Data_Mem/n7839 ), .S(N28), 
        .Z(\Data_Mem/n7841 ) );
  MUX \Data_Mem/U7866  ( .A(data_mem_out_wire[1049]), .B(
        data_mem_out_wire[1081]), .S(N29), .Z(\Data_Mem/n7840 ) );
  MUX \Data_Mem/U7865  ( .A(data_mem_out_wire[1113]), .B(
        data_mem_out_wire[1145]), .S(N29), .Z(\Data_Mem/n7839 ) );
  MUX \Data_Mem/U7864  ( .A(\Data_Mem/n7837 ), .B(\Data_Mem/n7836 ), .S(N28), 
        .Z(\Data_Mem/n7838 ) );
  MUX \Data_Mem/U7863  ( .A(data_mem_out_wire[1177]), .B(
        data_mem_out_wire[1209]), .S(N29), .Z(\Data_Mem/n7837 ) );
  MUX \Data_Mem/U7862  ( .A(data_mem_out_wire[1241]), .B(
        data_mem_out_wire[1273]), .S(N29), .Z(\Data_Mem/n7836 ) );
  MUX \Data_Mem/U7861  ( .A(\Data_Mem/n7834 ), .B(\Data_Mem/n7831 ), .S(N27), 
        .Z(\Data_Mem/n7835 ) );
  MUX \Data_Mem/U7860  ( .A(\Data_Mem/n7833 ), .B(\Data_Mem/n7832 ), .S(N28), 
        .Z(\Data_Mem/n7834 ) );
  MUX \Data_Mem/U7859  ( .A(data_mem_out_wire[1305]), .B(
        data_mem_out_wire[1337]), .S(N29), .Z(\Data_Mem/n7833 ) );
  MUX \Data_Mem/U7858  ( .A(data_mem_out_wire[1369]), .B(
        data_mem_out_wire[1401]), .S(N29), .Z(\Data_Mem/n7832 ) );
  MUX \Data_Mem/U7857  ( .A(\Data_Mem/n7830 ), .B(\Data_Mem/n7829 ), .S(N28), 
        .Z(\Data_Mem/n7831 ) );
  MUX \Data_Mem/U7856  ( .A(data_mem_out_wire[1433]), .B(
        data_mem_out_wire[1465]), .S(N29), .Z(\Data_Mem/n7830 ) );
  MUX \Data_Mem/U7855  ( .A(data_mem_out_wire[1497]), .B(
        data_mem_out_wire[1529]), .S(N29), .Z(\Data_Mem/n7829 ) );
  MUX \Data_Mem/U7854  ( .A(\Data_Mem/n7827 ), .B(\Data_Mem/n7820 ), .S(N26), 
        .Z(\Data_Mem/n7828 ) );
  MUX \Data_Mem/U7853  ( .A(\Data_Mem/n7826 ), .B(\Data_Mem/n7823 ), .S(N27), 
        .Z(\Data_Mem/n7827 ) );
  MUX \Data_Mem/U7852  ( .A(\Data_Mem/n7825 ), .B(\Data_Mem/n7824 ), .S(N28), 
        .Z(\Data_Mem/n7826 ) );
  MUX \Data_Mem/U7851  ( .A(data_mem_out_wire[1561]), .B(
        data_mem_out_wire[1593]), .S(N29), .Z(\Data_Mem/n7825 ) );
  MUX \Data_Mem/U7850  ( .A(data_mem_out_wire[1625]), .B(
        data_mem_out_wire[1657]), .S(N29), .Z(\Data_Mem/n7824 ) );
  MUX \Data_Mem/U7849  ( .A(\Data_Mem/n7822 ), .B(\Data_Mem/n7821 ), .S(N28), 
        .Z(\Data_Mem/n7823 ) );
  MUX \Data_Mem/U7848  ( .A(data_mem_out_wire[1689]), .B(
        data_mem_out_wire[1721]), .S(N29), .Z(\Data_Mem/n7822 ) );
  MUX \Data_Mem/U7847  ( .A(data_mem_out_wire[1753]), .B(
        data_mem_out_wire[1785]), .S(N29), .Z(\Data_Mem/n7821 ) );
  MUX \Data_Mem/U7846  ( .A(\Data_Mem/n7819 ), .B(\Data_Mem/n7816 ), .S(N27), 
        .Z(\Data_Mem/n7820 ) );
  MUX \Data_Mem/U7845  ( .A(\Data_Mem/n7818 ), .B(\Data_Mem/n7817 ), .S(N28), 
        .Z(\Data_Mem/n7819 ) );
  MUX \Data_Mem/U7844  ( .A(data_mem_out_wire[1817]), .B(
        data_mem_out_wire[1849]), .S(N29), .Z(\Data_Mem/n7818 ) );
  MUX \Data_Mem/U7843  ( .A(data_mem_out_wire[1881]), .B(
        data_mem_out_wire[1913]), .S(N29), .Z(\Data_Mem/n7817 ) );
  MUX \Data_Mem/U7842  ( .A(\Data_Mem/n7815 ), .B(\Data_Mem/n7814 ), .S(N28), 
        .Z(\Data_Mem/n7816 ) );
  MUX \Data_Mem/U7841  ( .A(data_mem_out_wire[1945]), .B(
        data_mem_out_wire[1977]), .S(N29), .Z(\Data_Mem/n7815 ) );
  MUX \Data_Mem/U7840  ( .A(data_mem_out_wire[2009]), .B(
        data_mem_out_wire[2041]), .S(N29), .Z(\Data_Mem/n7814 ) );
  MUX \Data_Mem/U7839  ( .A(\Data_Mem/n7813 ), .B(\Data_Mem/n7782 ), .S(N24), 
        .Z(c_memory[24]) );
  MUX \Data_Mem/U7838  ( .A(\Data_Mem/n7812 ), .B(\Data_Mem/n7797 ), .S(N25), 
        .Z(\Data_Mem/n7813 ) );
  MUX \Data_Mem/U7837  ( .A(\Data_Mem/n7811 ), .B(\Data_Mem/n7804 ), .S(N26), 
        .Z(\Data_Mem/n7812 ) );
  MUX \Data_Mem/U7836  ( .A(\Data_Mem/n7810 ), .B(\Data_Mem/n7807 ), .S(N27), 
        .Z(\Data_Mem/n7811 ) );
  MUX \Data_Mem/U7835  ( .A(\Data_Mem/n7809 ), .B(\Data_Mem/n7808 ), .S(N28), 
        .Z(\Data_Mem/n7810 ) );
  MUX \Data_Mem/U7834  ( .A(data_mem_out_wire[24]), .B(data_mem_out_wire[56]), 
        .S(N29), .Z(\Data_Mem/n7809 ) );
  MUX \Data_Mem/U7833  ( .A(data_mem_out_wire[88]), .B(data_mem_out_wire[120]), 
        .S(N29), .Z(\Data_Mem/n7808 ) );
  MUX \Data_Mem/U7832  ( .A(\Data_Mem/n7806 ), .B(\Data_Mem/n7805 ), .S(N28), 
        .Z(\Data_Mem/n7807 ) );
  MUX \Data_Mem/U7831  ( .A(data_mem_out_wire[152]), .B(data_mem_out_wire[184]), .S(N29), .Z(\Data_Mem/n7806 ) );
  MUX \Data_Mem/U7830  ( .A(data_mem_out_wire[216]), .B(data_mem_out_wire[248]), .S(N29), .Z(\Data_Mem/n7805 ) );
  MUX \Data_Mem/U7829  ( .A(\Data_Mem/n7803 ), .B(\Data_Mem/n7800 ), .S(N27), 
        .Z(\Data_Mem/n7804 ) );
  MUX \Data_Mem/U7828  ( .A(\Data_Mem/n7802 ), .B(\Data_Mem/n7801 ), .S(N28), 
        .Z(\Data_Mem/n7803 ) );
  MUX \Data_Mem/U7827  ( .A(data_mem_out_wire[280]), .B(data_mem_out_wire[312]), .S(N29), .Z(\Data_Mem/n7802 ) );
  MUX \Data_Mem/U7826  ( .A(data_mem_out_wire[344]), .B(data_mem_out_wire[376]), .S(N29), .Z(\Data_Mem/n7801 ) );
  MUX \Data_Mem/U7825  ( .A(\Data_Mem/n7799 ), .B(\Data_Mem/n7798 ), .S(N28), 
        .Z(\Data_Mem/n7800 ) );
  MUX \Data_Mem/U7824  ( .A(data_mem_out_wire[408]), .B(data_mem_out_wire[440]), .S(N29), .Z(\Data_Mem/n7799 ) );
  MUX \Data_Mem/U7823  ( .A(data_mem_out_wire[472]), .B(data_mem_out_wire[504]), .S(N29), .Z(\Data_Mem/n7798 ) );
  MUX \Data_Mem/U7822  ( .A(\Data_Mem/n7796 ), .B(\Data_Mem/n7789 ), .S(N26), 
        .Z(\Data_Mem/n7797 ) );
  MUX \Data_Mem/U7821  ( .A(\Data_Mem/n7795 ), .B(\Data_Mem/n7792 ), .S(N27), 
        .Z(\Data_Mem/n7796 ) );
  MUX \Data_Mem/U7820  ( .A(\Data_Mem/n7794 ), .B(\Data_Mem/n7793 ), .S(N28), 
        .Z(\Data_Mem/n7795 ) );
  MUX \Data_Mem/U7819  ( .A(data_mem_out_wire[536]), .B(data_mem_out_wire[568]), .S(N29), .Z(\Data_Mem/n7794 ) );
  MUX \Data_Mem/U7818  ( .A(data_mem_out_wire[600]), .B(data_mem_out_wire[632]), .S(N29), .Z(\Data_Mem/n7793 ) );
  MUX \Data_Mem/U7817  ( .A(\Data_Mem/n7791 ), .B(\Data_Mem/n7790 ), .S(N28), 
        .Z(\Data_Mem/n7792 ) );
  MUX \Data_Mem/U7816  ( .A(data_mem_out_wire[664]), .B(data_mem_out_wire[696]), .S(N29), .Z(\Data_Mem/n7791 ) );
  MUX \Data_Mem/U7815  ( .A(data_mem_out_wire[728]), .B(data_mem_out_wire[760]), .S(N29), .Z(\Data_Mem/n7790 ) );
  MUX \Data_Mem/U7814  ( .A(\Data_Mem/n7788 ), .B(\Data_Mem/n7785 ), .S(N27), 
        .Z(\Data_Mem/n7789 ) );
  MUX \Data_Mem/U7813  ( .A(\Data_Mem/n7787 ), .B(\Data_Mem/n7786 ), .S(N28), 
        .Z(\Data_Mem/n7788 ) );
  MUX \Data_Mem/U7812  ( .A(data_mem_out_wire[792]), .B(data_mem_out_wire[824]), .S(N29), .Z(\Data_Mem/n7787 ) );
  MUX \Data_Mem/U7811  ( .A(data_mem_out_wire[856]), .B(data_mem_out_wire[888]), .S(N29), .Z(\Data_Mem/n7786 ) );
  MUX \Data_Mem/U7810  ( .A(\Data_Mem/n7784 ), .B(\Data_Mem/n7783 ), .S(N28), 
        .Z(\Data_Mem/n7785 ) );
  MUX \Data_Mem/U7809  ( .A(data_mem_out_wire[920]), .B(data_mem_out_wire[952]), .S(N29), .Z(\Data_Mem/n7784 ) );
  MUX \Data_Mem/U7808  ( .A(data_mem_out_wire[984]), .B(
        data_mem_out_wire[1016]), .S(N29), .Z(\Data_Mem/n7783 ) );
  MUX \Data_Mem/U7807  ( .A(\Data_Mem/n7781 ), .B(\Data_Mem/n7766 ), .S(N25), 
        .Z(\Data_Mem/n7782 ) );
  MUX \Data_Mem/U7806  ( .A(\Data_Mem/n7780 ), .B(\Data_Mem/n7773 ), .S(N26), 
        .Z(\Data_Mem/n7781 ) );
  MUX \Data_Mem/U7805  ( .A(\Data_Mem/n7779 ), .B(\Data_Mem/n7776 ), .S(N27), 
        .Z(\Data_Mem/n7780 ) );
  MUX \Data_Mem/U7804  ( .A(\Data_Mem/n7778 ), .B(\Data_Mem/n7777 ), .S(N28), 
        .Z(\Data_Mem/n7779 ) );
  MUX \Data_Mem/U7803  ( .A(data_mem_out_wire[1048]), .B(
        data_mem_out_wire[1080]), .S(N29), .Z(\Data_Mem/n7778 ) );
  MUX \Data_Mem/U7802  ( .A(data_mem_out_wire[1112]), .B(
        data_mem_out_wire[1144]), .S(N29), .Z(\Data_Mem/n7777 ) );
  MUX \Data_Mem/U7801  ( .A(\Data_Mem/n7775 ), .B(\Data_Mem/n7774 ), .S(N28), 
        .Z(\Data_Mem/n7776 ) );
  MUX \Data_Mem/U7800  ( .A(data_mem_out_wire[1176]), .B(
        data_mem_out_wire[1208]), .S(N29), .Z(\Data_Mem/n7775 ) );
  MUX \Data_Mem/U7799  ( .A(data_mem_out_wire[1240]), .B(
        data_mem_out_wire[1272]), .S(N29), .Z(\Data_Mem/n7774 ) );
  MUX \Data_Mem/U7798  ( .A(\Data_Mem/n7772 ), .B(\Data_Mem/n7769 ), .S(N27), 
        .Z(\Data_Mem/n7773 ) );
  MUX \Data_Mem/U7797  ( .A(\Data_Mem/n7771 ), .B(\Data_Mem/n7770 ), .S(N28), 
        .Z(\Data_Mem/n7772 ) );
  MUX \Data_Mem/U7796  ( .A(data_mem_out_wire[1304]), .B(
        data_mem_out_wire[1336]), .S(N29), .Z(\Data_Mem/n7771 ) );
  MUX \Data_Mem/U7795  ( .A(data_mem_out_wire[1368]), .B(
        data_mem_out_wire[1400]), .S(N29), .Z(\Data_Mem/n7770 ) );
  MUX \Data_Mem/U7794  ( .A(\Data_Mem/n7768 ), .B(\Data_Mem/n7767 ), .S(N28), 
        .Z(\Data_Mem/n7769 ) );
  MUX \Data_Mem/U7793  ( .A(data_mem_out_wire[1432]), .B(
        data_mem_out_wire[1464]), .S(N29), .Z(\Data_Mem/n7768 ) );
  MUX \Data_Mem/U7792  ( .A(data_mem_out_wire[1496]), .B(
        data_mem_out_wire[1528]), .S(N29), .Z(\Data_Mem/n7767 ) );
  MUX \Data_Mem/U7791  ( .A(\Data_Mem/n7765 ), .B(\Data_Mem/n7758 ), .S(N26), 
        .Z(\Data_Mem/n7766 ) );
  MUX \Data_Mem/U7790  ( .A(\Data_Mem/n7764 ), .B(\Data_Mem/n7761 ), .S(N27), 
        .Z(\Data_Mem/n7765 ) );
  MUX \Data_Mem/U7789  ( .A(\Data_Mem/n7763 ), .B(\Data_Mem/n7762 ), .S(N28), 
        .Z(\Data_Mem/n7764 ) );
  MUX \Data_Mem/U7788  ( .A(data_mem_out_wire[1560]), .B(
        data_mem_out_wire[1592]), .S(N29), .Z(\Data_Mem/n7763 ) );
  MUX \Data_Mem/U7787  ( .A(data_mem_out_wire[1624]), .B(
        data_mem_out_wire[1656]), .S(N29), .Z(\Data_Mem/n7762 ) );
  MUX \Data_Mem/U7786  ( .A(\Data_Mem/n7760 ), .B(\Data_Mem/n7759 ), .S(N28), 
        .Z(\Data_Mem/n7761 ) );
  MUX \Data_Mem/U7785  ( .A(data_mem_out_wire[1688]), .B(
        data_mem_out_wire[1720]), .S(N29), .Z(\Data_Mem/n7760 ) );
  MUX \Data_Mem/U7784  ( .A(data_mem_out_wire[1752]), .B(
        data_mem_out_wire[1784]), .S(N29), .Z(\Data_Mem/n7759 ) );
  MUX \Data_Mem/U7783  ( .A(\Data_Mem/n7757 ), .B(\Data_Mem/n7754 ), .S(N27), 
        .Z(\Data_Mem/n7758 ) );
  MUX \Data_Mem/U7782  ( .A(\Data_Mem/n7756 ), .B(\Data_Mem/n7755 ), .S(N28), 
        .Z(\Data_Mem/n7757 ) );
  MUX \Data_Mem/U7781  ( .A(data_mem_out_wire[1816]), .B(
        data_mem_out_wire[1848]), .S(N29), .Z(\Data_Mem/n7756 ) );
  MUX \Data_Mem/U7780  ( .A(data_mem_out_wire[1880]), .B(
        data_mem_out_wire[1912]), .S(N29), .Z(\Data_Mem/n7755 ) );
  MUX \Data_Mem/U7779  ( .A(\Data_Mem/n7753 ), .B(\Data_Mem/n7752 ), .S(N28), 
        .Z(\Data_Mem/n7754 ) );
  MUX \Data_Mem/U7778  ( .A(data_mem_out_wire[1944]), .B(
        data_mem_out_wire[1976]), .S(N29), .Z(\Data_Mem/n7753 ) );
  MUX \Data_Mem/U7777  ( .A(data_mem_out_wire[2008]), .B(
        data_mem_out_wire[2040]), .S(N29), .Z(\Data_Mem/n7752 ) );
  MUX \Data_Mem/U7776  ( .A(\Data_Mem/n7751 ), .B(\Data_Mem/n7720 ), .S(N24), 
        .Z(c_memory[23]) );
  MUX \Data_Mem/U7775  ( .A(\Data_Mem/n7750 ), .B(\Data_Mem/n7735 ), .S(N25), 
        .Z(\Data_Mem/n7751 ) );
  MUX \Data_Mem/U7774  ( .A(\Data_Mem/n7749 ), .B(\Data_Mem/n7742 ), .S(N26), 
        .Z(\Data_Mem/n7750 ) );
  MUX \Data_Mem/U7773  ( .A(\Data_Mem/n7748 ), .B(\Data_Mem/n7745 ), .S(N27), 
        .Z(\Data_Mem/n7749 ) );
  MUX \Data_Mem/U7772  ( .A(\Data_Mem/n7747 ), .B(\Data_Mem/n7746 ), .S(N28), 
        .Z(\Data_Mem/n7748 ) );
  MUX \Data_Mem/U7771  ( .A(data_mem_out_wire[23]), .B(data_mem_out_wire[55]), 
        .S(N29), .Z(\Data_Mem/n7747 ) );
  MUX \Data_Mem/U7770  ( .A(data_mem_out_wire[87]), .B(data_mem_out_wire[119]), 
        .S(N29), .Z(\Data_Mem/n7746 ) );
  MUX \Data_Mem/U7769  ( .A(\Data_Mem/n7744 ), .B(\Data_Mem/n7743 ), .S(N28), 
        .Z(\Data_Mem/n7745 ) );
  MUX \Data_Mem/U7768  ( .A(data_mem_out_wire[151]), .B(data_mem_out_wire[183]), .S(N29), .Z(\Data_Mem/n7744 ) );
  MUX \Data_Mem/U7767  ( .A(data_mem_out_wire[215]), .B(data_mem_out_wire[247]), .S(N29), .Z(\Data_Mem/n7743 ) );
  MUX \Data_Mem/U7766  ( .A(\Data_Mem/n7741 ), .B(\Data_Mem/n7738 ), .S(N27), 
        .Z(\Data_Mem/n7742 ) );
  MUX \Data_Mem/U7765  ( .A(\Data_Mem/n7740 ), .B(\Data_Mem/n7739 ), .S(N28), 
        .Z(\Data_Mem/n7741 ) );
  MUX \Data_Mem/U7764  ( .A(data_mem_out_wire[279]), .B(data_mem_out_wire[311]), .S(N29), .Z(\Data_Mem/n7740 ) );
  MUX \Data_Mem/U7763  ( .A(data_mem_out_wire[343]), .B(data_mem_out_wire[375]), .S(N29), .Z(\Data_Mem/n7739 ) );
  MUX \Data_Mem/U7762  ( .A(\Data_Mem/n7737 ), .B(\Data_Mem/n7736 ), .S(N28), 
        .Z(\Data_Mem/n7738 ) );
  MUX \Data_Mem/U7761  ( .A(data_mem_out_wire[407]), .B(data_mem_out_wire[439]), .S(N29), .Z(\Data_Mem/n7737 ) );
  MUX \Data_Mem/U7760  ( .A(data_mem_out_wire[471]), .B(data_mem_out_wire[503]), .S(N29), .Z(\Data_Mem/n7736 ) );
  MUX \Data_Mem/U7759  ( .A(\Data_Mem/n7734 ), .B(\Data_Mem/n7727 ), .S(N26), 
        .Z(\Data_Mem/n7735 ) );
  MUX \Data_Mem/U7758  ( .A(\Data_Mem/n7733 ), .B(\Data_Mem/n7730 ), .S(N27), 
        .Z(\Data_Mem/n7734 ) );
  MUX \Data_Mem/U7757  ( .A(\Data_Mem/n7732 ), .B(\Data_Mem/n7731 ), .S(N28), 
        .Z(\Data_Mem/n7733 ) );
  MUX \Data_Mem/U7756  ( .A(data_mem_out_wire[535]), .B(data_mem_out_wire[567]), .S(N29), .Z(\Data_Mem/n7732 ) );
  MUX \Data_Mem/U7755  ( .A(data_mem_out_wire[599]), .B(data_mem_out_wire[631]), .S(N29), .Z(\Data_Mem/n7731 ) );
  MUX \Data_Mem/U7754  ( .A(\Data_Mem/n7729 ), .B(\Data_Mem/n7728 ), .S(N28), 
        .Z(\Data_Mem/n7730 ) );
  MUX \Data_Mem/U7753  ( .A(data_mem_out_wire[663]), .B(data_mem_out_wire[695]), .S(N29), .Z(\Data_Mem/n7729 ) );
  MUX \Data_Mem/U7752  ( .A(data_mem_out_wire[727]), .B(data_mem_out_wire[759]), .S(N29), .Z(\Data_Mem/n7728 ) );
  MUX \Data_Mem/U7751  ( .A(\Data_Mem/n7726 ), .B(\Data_Mem/n7723 ), .S(N27), 
        .Z(\Data_Mem/n7727 ) );
  MUX \Data_Mem/U7750  ( .A(\Data_Mem/n7725 ), .B(\Data_Mem/n7724 ), .S(N28), 
        .Z(\Data_Mem/n7726 ) );
  MUX \Data_Mem/U7749  ( .A(data_mem_out_wire[791]), .B(data_mem_out_wire[823]), .S(N29), .Z(\Data_Mem/n7725 ) );
  MUX \Data_Mem/U7748  ( .A(data_mem_out_wire[855]), .B(data_mem_out_wire[887]), .S(N29), .Z(\Data_Mem/n7724 ) );
  MUX \Data_Mem/U7747  ( .A(\Data_Mem/n7722 ), .B(\Data_Mem/n7721 ), .S(N28), 
        .Z(\Data_Mem/n7723 ) );
  MUX \Data_Mem/U7746  ( .A(data_mem_out_wire[919]), .B(data_mem_out_wire[951]), .S(N29), .Z(\Data_Mem/n7722 ) );
  MUX \Data_Mem/U7745  ( .A(data_mem_out_wire[983]), .B(
        data_mem_out_wire[1015]), .S(N29), .Z(\Data_Mem/n7721 ) );
  MUX \Data_Mem/U7744  ( .A(\Data_Mem/n7719 ), .B(\Data_Mem/n7704 ), .S(N25), 
        .Z(\Data_Mem/n7720 ) );
  MUX \Data_Mem/U7743  ( .A(\Data_Mem/n7718 ), .B(\Data_Mem/n7711 ), .S(N26), 
        .Z(\Data_Mem/n7719 ) );
  MUX \Data_Mem/U7742  ( .A(\Data_Mem/n7717 ), .B(\Data_Mem/n7714 ), .S(N27), 
        .Z(\Data_Mem/n7718 ) );
  MUX \Data_Mem/U7741  ( .A(\Data_Mem/n7716 ), .B(\Data_Mem/n7715 ), .S(N28), 
        .Z(\Data_Mem/n7717 ) );
  MUX \Data_Mem/U7740  ( .A(data_mem_out_wire[1047]), .B(
        data_mem_out_wire[1079]), .S(N29), .Z(\Data_Mem/n7716 ) );
  MUX \Data_Mem/U7739  ( .A(data_mem_out_wire[1111]), .B(
        data_mem_out_wire[1143]), .S(N29), .Z(\Data_Mem/n7715 ) );
  MUX \Data_Mem/U7738  ( .A(\Data_Mem/n7713 ), .B(\Data_Mem/n7712 ), .S(N28), 
        .Z(\Data_Mem/n7714 ) );
  MUX \Data_Mem/U7737  ( .A(data_mem_out_wire[1175]), .B(
        data_mem_out_wire[1207]), .S(N29), .Z(\Data_Mem/n7713 ) );
  MUX \Data_Mem/U7736  ( .A(data_mem_out_wire[1239]), .B(
        data_mem_out_wire[1271]), .S(N29), .Z(\Data_Mem/n7712 ) );
  MUX \Data_Mem/U7735  ( .A(\Data_Mem/n7710 ), .B(\Data_Mem/n7707 ), .S(N27), 
        .Z(\Data_Mem/n7711 ) );
  MUX \Data_Mem/U7734  ( .A(\Data_Mem/n7709 ), .B(\Data_Mem/n7708 ), .S(N28), 
        .Z(\Data_Mem/n7710 ) );
  MUX \Data_Mem/U7733  ( .A(data_mem_out_wire[1303]), .B(
        data_mem_out_wire[1335]), .S(N29), .Z(\Data_Mem/n7709 ) );
  MUX \Data_Mem/U7732  ( .A(data_mem_out_wire[1367]), .B(
        data_mem_out_wire[1399]), .S(N29), .Z(\Data_Mem/n7708 ) );
  MUX \Data_Mem/U7731  ( .A(\Data_Mem/n7706 ), .B(\Data_Mem/n7705 ), .S(N28), 
        .Z(\Data_Mem/n7707 ) );
  MUX \Data_Mem/U7730  ( .A(data_mem_out_wire[1431]), .B(
        data_mem_out_wire[1463]), .S(N29), .Z(\Data_Mem/n7706 ) );
  MUX \Data_Mem/U7729  ( .A(data_mem_out_wire[1495]), .B(
        data_mem_out_wire[1527]), .S(N29), .Z(\Data_Mem/n7705 ) );
  MUX \Data_Mem/U7728  ( .A(\Data_Mem/n7703 ), .B(\Data_Mem/n7696 ), .S(N26), 
        .Z(\Data_Mem/n7704 ) );
  MUX \Data_Mem/U7727  ( .A(\Data_Mem/n7702 ), .B(\Data_Mem/n7699 ), .S(N27), 
        .Z(\Data_Mem/n7703 ) );
  MUX \Data_Mem/U7726  ( .A(\Data_Mem/n7701 ), .B(\Data_Mem/n7700 ), .S(N28), 
        .Z(\Data_Mem/n7702 ) );
  MUX \Data_Mem/U7725  ( .A(data_mem_out_wire[1559]), .B(
        data_mem_out_wire[1591]), .S(N29), .Z(\Data_Mem/n7701 ) );
  MUX \Data_Mem/U7724  ( .A(data_mem_out_wire[1623]), .B(
        data_mem_out_wire[1655]), .S(N29), .Z(\Data_Mem/n7700 ) );
  MUX \Data_Mem/U7723  ( .A(\Data_Mem/n7698 ), .B(\Data_Mem/n7697 ), .S(N28), 
        .Z(\Data_Mem/n7699 ) );
  MUX \Data_Mem/U7722  ( .A(data_mem_out_wire[1687]), .B(
        data_mem_out_wire[1719]), .S(N29), .Z(\Data_Mem/n7698 ) );
  MUX \Data_Mem/U7721  ( .A(data_mem_out_wire[1751]), .B(
        data_mem_out_wire[1783]), .S(N29), .Z(\Data_Mem/n7697 ) );
  MUX \Data_Mem/U7720  ( .A(\Data_Mem/n7695 ), .B(\Data_Mem/n7692 ), .S(N27), 
        .Z(\Data_Mem/n7696 ) );
  MUX \Data_Mem/U7719  ( .A(\Data_Mem/n7694 ), .B(\Data_Mem/n7693 ), .S(N28), 
        .Z(\Data_Mem/n7695 ) );
  MUX \Data_Mem/U7718  ( .A(data_mem_out_wire[1815]), .B(
        data_mem_out_wire[1847]), .S(N29), .Z(\Data_Mem/n7694 ) );
  MUX \Data_Mem/U7717  ( .A(data_mem_out_wire[1879]), .B(
        data_mem_out_wire[1911]), .S(N29), .Z(\Data_Mem/n7693 ) );
  MUX \Data_Mem/U7716  ( .A(\Data_Mem/n7691 ), .B(\Data_Mem/n7690 ), .S(N28), 
        .Z(\Data_Mem/n7692 ) );
  MUX \Data_Mem/U7715  ( .A(data_mem_out_wire[1943]), .B(
        data_mem_out_wire[1975]), .S(N29), .Z(\Data_Mem/n7691 ) );
  MUX \Data_Mem/U7714  ( .A(data_mem_out_wire[2007]), .B(
        data_mem_out_wire[2039]), .S(N29), .Z(\Data_Mem/n7690 ) );
  MUX \Data_Mem/U7713  ( .A(\Data_Mem/n7689 ), .B(\Data_Mem/n7658 ), .S(N24), 
        .Z(c_memory[22]) );
  MUX \Data_Mem/U7712  ( .A(\Data_Mem/n7688 ), .B(\Data_Mem/n7673 ), .S(N25), 
        .Z(\Data_Mem/n7689 ) );
  MUX \Data_Mem/U7711  ( .A(\Data_Mem/n7687 ), .B(\Data_Mem/n7680 ), .S(N26), 
        .Z(\Data_Mem/n7688 ) );
  MUX \Data_Mem/U7710  ( .A(\Data_Mem/n7686 ), .B(\Data_Mem/n7683 ), .S(N27), 
        .Z(\Data_Mem/n7687 ) );
  MUX \Data_Mem/U7709  ( .A(\Data_Mem/n7685 ), .B(\Data_Mem/n7684 ), .S(N28), 
        .Z(\Data_Mem/n7686 ) );
  MUX \Data_Mem/U7708  ( .A(data_mem_out_wire[22]), .B(data_mem_out_wire[54]), 
        .S(N29), .Z(\Data_Mem/n7685 ) );
  MUX \Data_Mem/U7707  ( .A(data_mem_out_wire[86]), .B(data_mem_out_wire[118]), 
        .S(N29), .Z(\Data_Mem/n7684 ) );
  MUX \Data_Mem/U7706  ( .A(\Data_Mem/n7682 ), .B(\Data_Mem/n7681 ), .S(N28), 
        .Z(\Data_Mem/n7683 ) );
  MUX \Data_Mem/U7705  ( .A(data_mem_out_wire[150]), .B(data_mem_out_wire[182]), .S(N29), .Z(\Data_Mem/n7682 ) );
  MUX \Data_Mem/U7704  ( .A(data_mem_out_wire[214]), .B(data_mem_out_wire[246]), .S(N29), .Z(\Data_Mem/n7681 ) );
  MUX \Data_Mem/U7703  ( .A(\Data_Mem/n7679 ), .B(\Data_Mem/n7676 ), .S(N27), 
        .Z(\Data_Mem/n7680 ) );
  MUX \Data_Mem/U7702  ( .A(\Data_Mem/n7678 ), .B(\Data_Mem/n7677 ), .S(N28), 
        .Z(\Data_Mem/n7679 ) );
  MUX \Data_Mem/U7701  ( .A(data_mem_out_wire[278]), .B(data_mem_out_wire[310]), .S(N29), .Z(\Data_Mem/n7678 ) );
  MUX \Data_Mem/U7700  ( .A(data_mem_out_wire[342]), .B(data_mem_out_wire[374]), .S(N29), .Z(\Data_Mem/n7677 ) );
  MUX \Data_Mem/U7699  ( .A(\Data_Mem/n7675 ), .B(\Data_Mem/n7674 ), .S(N28), 
        .Z(\Data_Mem/n7676 ) );
  MUX \Data_Mem/U7698  ( .A(data_mem_out_wire[406]), .B(data_mem_out_wire[438]), .S(N29), .Z(\Data_Mem/n7675 ) );
  MUX \Data_Mem/U7697  ( .A(data_mem_out_wire[470]), .B(data_mem_out_wire[502]), .S(N29), .Z(\Data_Mem/n7674 ) );
  MUX \Data_Mem/U7696  ( .A(\Data_Mem/n7672 ), .B(\Data_Mem/n7665 ), .S(N26), 
        .Z(\Data_Mem/n7673 ) );
  MUX \Data_Mem/U7695  ( .A(\Data_Mem/n7671 ), .B(\Data_Mem/n7668 ), .S(N27), 
        .Z(\Data_Mem/n7672 ) );
  MUX \Data_Mem/U7694  ( .A(\Data_Mem/n7670 ), .B(\Data_Mem/n7669 ), .S(N28), 
        .Z(\Data_Mem/n7671 ) );
  MUX \Data_Mem/U7693  ( .A(data_mem_out_wire[534]), .B(data_mem_out_wire[566]), .S(N29), .Z(\Data_Mem/n7670 ) );
  MUX \Data_Mem/U7692  ( .A(data_mem_out_wire[598]), .B(data_mem_out_wire[630]), .S(N29), .Z(\Data_Mem/n7669 ) );
  MUX \Data_Mem/U7691  ( .A(\Data_Mem/n7667 ), .B(\Data_Mem/n7666 ), .S(N28), 
        .Z(\Data_Mem/n7668 ) );
  MUX \Data_Mem/U7690  ( .A(data_mem_out_wire[662]), .B(data_mem_out_wire[694]), .S(N29), .Z(\Data_Mem/n7667 ) );
  MUX \Data_Mem/U7689  ( .A(data_mem_out_wire[726]), .B(data_mem_out_wire[758]), .S(N29), .Z(\Data_Mem/n7666 ) );
  MUX \Data_Mem/U7688  ( .A(\Data_Mem/n7664 ), .B(\Data_Mem/n7661 ), .S(N27), 
        .Z(\Data_Mem/n7665 ) );
  MUX \Data_Mem/U7687  ( .A(\Data_Mem/n7663 ), .B(\Data_Mem/n7662 ), .S(N28), 
        .Z(\Data_Mem/n7664 ) );
  MUX \Data_Mem/U7686  ( .A(data_mem_out_wire[790]), .B(data_mem_out_wire[822]), .S(N29), .Z(\Data_Mem/n7663 ) );
  MUX \Data_Mem/U7685  ( .A(data_mem_out_wire[854]), .B(data_mem_out_wire[886]), .S(N29), .Z(\Data_Mem/n7662 ) );
  MUX \Data_Mem/U7684  ( .A(\Data_Mem/n7660 ), .B(\Data_Mem/n7659 ), .S(N28), 
        .Z(\Data_Mem/n7661 ) );
  MUX \Data_Mem/U7683  ( .A(data_mem_out_wire[918]), .B(data_mem_out_wire[950]), .S(N29), .Z(\Data_Mem/n7660 ) );
  MUX \Data_Mem/U7682  ( .A(data_mem_out_wire[982]), .B(
        data_mem_out_wire[1014]), .S(N29), .Z(\Data_Mem/n7659 ) );
  MUX \Data_Mem/U7681  ( .A(\Data_Mem/n7657 ), .B(\Data_Mem/n7642 ), .S(N25), 
        .Z(\Data_Mem/n7658 ) );
  MUX \Data_Mem/U7680  ( .A(\Data_Mem/n7656 ), .B(\Data_Mem/n7649 ), .S(N26), 
        .Z(\Data_Mem/n7657 ) );
  MUX \Data_Mem/U7679  ( .A(\Data_Mem/n7655 ), .B(\Data_Mem/n7652 ), .S(N27), 
        .Z(\Data_Mem/n7656 ) );
  MUX \Data_Mem/U7678  ( .A(\Data_Mem/n7654 ), .B(\Data_Mem/n7653 ), .S(N28), 
        .Z(\Data_Mem/n7655 ) );
  MUX \Data_Mem/U7677  ( .A(data_mem_out_wire[1046]), .B(
        data_mem_out_wire[1078]), .S(N29), .Z(\Data_Mem/n7654 ) );
  MUX \Data_Mem/U7676  ( .A(data_mem_out_wire[1110]), .B(
        data_mem_out_wire[1142]), .S(N29), .Z(\Data_Mem/n7653 ) );
  MUX \Data_Mem/U7675  ( .A(\Data_Mem/n7651 ), .B(\Data_Mem/n7650 ), .S(N28), 
        .Z(\Data_Mem/n7652 ) );
  MUX \Data_Mem/U7674  ( .A(data_mem_out_wire[1174]), .B(
        data_mem_out_wire[1206]), .S(N29), .Z(\Data_Mem/n7651 ) );
  MUX \Data_Mem/U7673  ( .A(data_mem_out_wire[1238]), .B(
        data_mem_out_wire[1270]), .S(N29), .Z(\Data_Mem/n7650 ) );
  MUX \Data_Mem/U7672  ( .A(\Data_Mem/n7648 ), .B(\Data_Mem/n7645 ), .S(N27), 
        .Z(\Data_Mem/n7649 ) );
  MUX \Data_Mem/U7671  ( .A(\Data_Mem/n7647 ), .B(\Data_Mem/n7646 ), .S(N28), 
        .Z(\Data_Mem/n7648 ) );
  MUX \Data_Mem/U7670  ( .A(data_mem_out_wire[1302]), .B(
        data_mem_out_wire[1334]), .S(N29), .Z(\Data_Mem/n7647 ) );
  MUX \Data_Mem/U7669  ( .A(data_mem_out_wire[1366]), .B(
        data_mem_out_wire[1398]), .S(N29), .Z(\Data_Mem/n7646 ) );
  MUX \Data_Mem/U7668  ( .A(\Data_Mem/n7644 ), .B(\Data_Mem/n7643 ), .S(N28), 
        .Z(\Data_Mem/n7645 ) );
  MUX \Data_Mem/U7667  ( .A(data_mem_out_wire[1430]), .B(
        data_mem_out_wire[1462]), .S(N29), .Z(\Data_Mem/n7644 ) );
  MUX \Data_Mem/U7666  ( .A(data_mem_out_wire[1494]), .B(
        data_mem_out_wire[1526]), .S(N29), .Z(\Data_Mem/n7643 ) );
  MUX \Data_Mem/U7665  ( .A(\Data_Mem/n7641 ), .B(\Data_Mem/n7634 ), .S(N26), 
        .Z(\Data_Mem/n7642 ) );
  MUX \Data_Mem/U7664  ( .A(\Data_Mem/n7640 ), .B(\Data_Mem/n7637 ), .S(N27), 
        .Z(\Data_Mem/n7641 ) );
  MUX \Data_Mem/U7663  ( .A(\Data_Mem/n7639 ), .B(\Data_Mem/n7638 ), .S(N28), 
        .Z(\Data_Mem/n7640 ) );
  MUX \Data_Mem/U7662  ( .A(data_mem_out_wire[1558]), .B(
        data_mem_out_wire[1590]), .S(N29), .Z(\Data_Mem/n7639 ) );
  MUX \Data_Mem/U7661  ( .A(data_mem_out_wire[1622]), .B(
        data_mem_out_wire[1654]), .S(N29), .Z(\Data_Mem/n7638 ) );
  MUX \Data_Mem/U7660  ( .A(\Data_Mem/n7636 ), .B(\Data_Mem/n7635 ), .S(N28), 
        .Z(\Data_Mem/n7637 ) );
  MUX \Data_Mem/U7659  ( .A(data_mem_out_wire[1686]), .B(
        data_mem_out_wire[1718]), .S(N29), .Z(\Data_Mem/n7636 ) );
  MUX \Data_Mem/U7658  ( .A(data_mem_out_wire[1750]), .B(
        data_mem_out_wire[1782]), .S(N29), .Z(\Data_Mem/n7635 ) );
  MUX \Data_Mem/U7657  ( .A(\Data_Mem/n7633 ), .B(\Data_Mem/n7630 ), .S(N27), 
        .Z(\Data_Mem/n7634 ) );
  MUX \Data_Mem/U7656  ( .A(\Data_Mem/n7632 ), .B(\Data_Mem/n7631 ), .S(N28), 
        .Z(\Data_Mem/n7633 ) );
  MUX \Data_Mem/U7655  ( .A(data_mem_out_wire[1814]), .B(
        data_mem_out_wire[1846]), .S(N29), .Z(\Data_Mem/n7632 ) );
  MUX \Data_Mem/U7654  ( .A(data_mem_out_wire[1878]), .B(
        data_mem_out_wire[1910]), .S(N29), .Z(\Data_Mem/n7631 ) );
  MUX \Data_Mem/U7653  ( .A(\Data_Mem/n7629 ), .B(\Data_Mem/n7628 ), .S(N28), 
        .Z(\Data_Mem/n7630 ) );
  MUX \Data_Mem/U7652  ( .A(data_mem_out_wire[1942]), .B(
        data_mem_out_wire[1974]), .S(N29), .Z(\Data_Mem/n7629 ) );
  MUX \Data_Mem/U7651  ( .A(data_mem_out_wire[2006]), .B(
        data_mem_out_wire[2038]), .S(N29), .Z(\Data_Mem/n7628 ) );
  MUX \Data_Mem/U7650  ( .A(\Data_Mem/n7627 ), .B(\Data_Mem/n7596 ), .S(N24), 
        .Z(c_memory[21]) );
  MUX \Data_Mem/U7649  ( .A(\Data_Mem/n7626 ), .B(\Data_Mem/n7611 ), .S(N25), 
        .Z(\Data_Mem/n7627 ) );
  MUX \Data_Mem/U7648  ( .A(\Data_Mem/n7625 ), .B(\Data_Mem/n7618 ), .S(N26), 
        .Z(\Data_Mem/n7626 ) );
  MUX \Data_Mem/U7647  ( .A(\Data_Mem/n7624 ), .B(\Data_Mem/n7621 ), .S(N27), 
        .Z(\Data_Mem/n7625 ) );
  MUX \Data_Mem/U7646  ( .A(\Data_Mem/n7623 ), .B(\Data_Mem/n7622 ), .S(N28), 
        .Z(\Data_Mem/n7624 ) );
  MUX \Data_Mem/U7645  ( .A(data_mem_out_wire[21]), .B(data_mem_out_wire[53]), 
        .S(N29), .Z(\Data_Mem/n7623 ) );
  MUX \Data_Mem/U7644  ( .A(data_mem_out_wire[85]), .B(data_mem_out_wire[117]), 
        .S(N29), .Z(\Data_Mem/n7622 ) );
  MUX \Data_Mem/U7643  ( .A(\Data_Mem/n7620 ), .B(\Data_Mem/n7619 ), .S(N28), 
        .Z(\Data_Mem/n7621 ) );
  MUX \Data_Mem/U7642  ( .A(data_mem_out_wire[149]), .B(data_mem_out_wire[181]), .S(N29), .Z(\Data_Mem/n7620 ) );
  MUX \Data_Mem/U7641  ( .A(data_mem_out_wire[213]), .B(data_mem_out_wire[245]), .S(N29), .Z(\Data_Mem/n7619 ) );
  MUX \Data_Mem/U7640  ( .A(\Data_Mem/n7617 ), .B(\Data_Mem/n7614 ), .S(N27), 
        .Z(\Data_Mem/n7618 ) );
  MUX \Data_Mem/U7639  ( .A(\Data_Mem/n7616 ), .B(\Data_Mem/n7615 ), .S(N28), 
        .Z(\Data_Mem/n7617 ) );
  MUX \Data_Mem/U7638  ( .A(data_mem_out_wire[277]), .B(data_mem_out_wire[309]), .S(N29), .Z(\Data_Mem/n7616 ) );
  MUX \Data_Mem/U7637  ( .A(data_mem_out_wire[341]), .B(data_mem_out_wire[373]), .S(N29), .Z(\Data_Mem/n7615 ) );
  MUX \Data_Mem/U7636  ( .A(\Data_Mem/n7613 ), .B(\Data_Mem/n7612 ), .S(N28), 
        .Z(\Data_Mem/n7614 ) );
  MUX \Data_Mem/U7635  ( .A(data_mem_out_wire[405]), .B(data_mem_out_wire[437]), .S(N29), .Z(\Data_Mem/n7613 ) );
  MUX \Data_Mem/U7634  ( .A(data_mem_out_wire[469]), .B(data_mem_out_wire[501]), .S(N29), .Z(\Data_Mem/n7612 ) );
  MUX \Data_Mem/U7633  ( .A(\Data_Mem/n7610 ), .B(\Data_Mem/n7603 ), .S(N26), 
        .Z(\Data_Mem/n7611 ) );
  MUX \Data_Mem/U7632  ( .A(\Data_Mem/n7609 ), .B(\Data_Mem/n7606 ), .S(N27), 
        .Z(\Data_Mem/n7610 ) );
  MUX \Data_Mem/U7631  ( .A(\Data_Mem/n7608 ), .B(\Data_Mem/n7607 ), .S(N28), 
        .Z(\Data_Mem/n7609 ) );
  MUX \Data_Mem/U7630  ( .A(data_mem_out_wire[533]), .B(data_mem_out_wire[565]), .S(N29), .Z(\Data_Mem/n7608 ) );
  MUX \Data_Mem/U7629  ( .A(data_mem_out_wire[597]), .B(data_mem_out_wire[629]), .S(N29), .Z(\Data_Mem/n7607 ) );
  MUX \Data_Mem/U7628  ( .A(\Data_Mem/n7605 ), .B(\Data_Mem/n7604 ), .S(N28), 
        .Z(\Data_Mem/n7606 ) );
  MUX \Data_Mem/U7627  ( .A(data_mem_out_wire[661]), .B(data_mem_out_wire[693]), .S(N29), .Z(\Data_Mem/n7605 ) );
  MUX \Data_Mem/U7626  ( .A(data_mem_out_wire[725]), .B(data_mem_out_wire[757]), .S(N29), .Z(\Data_Mem/n7604 ) );
  MUX \Data_Mem/U7625  ( .A(\Data_Mem/n7602 ), .B(\Data_Mem/n7599 ), .S(N27), 
        .Z(\Data_Mem/n7603 ) );
  MUX \Data_Mem/U7624  ( .A(\Data_Mem/n7601 ), .B(\Data_Mem/n7600 ), .S(N28), 
        .Z(\Data_Mem/n7602 ) );
  MUX \Data_Mem/U7623  ( .A(data_mem_out_wire[789]), .B(data_mem_out_wire[821]), .S(N29), .Z(\Data_Mem/n7601 ) );
  MUX \Data_Mem/U7622  ( .A(data_mem_out_wire[853]), .B(data_mem_out_wire[885]), .S(N29), .Z(\Data_Mem/n7600 ) );
  MUX \Data_Mem/U7621  ( .A(\Data_Mem/n7598 ), .B(\Data_Mem/n7597 ), .S(N28), 
        .Z(\Data_Mem/n7599 ) );
  MUX \Data_Mem/U7620  ( .A(data_mem_out_wire[917]), .B(data_mem_out_wire[949]), .S(N29), .Z(\Data_Mem/n7598 ) );
  MUX \Data_Mem/U7619  ( .A(data_mem_out_wire[981]), .B(
        data_mem_out_wire[1013]), .S(N29), .Z(\Data_Mem/n7597 ) );
  MUX \Data_Mem/U7618  ( .A(\Data_Mem/n7595 ), .B(\Data_Mem/n7580 ), .S(N25), 
        .Z(\Data_Mem/n7596 ) );
  MUX \Data_Mem/U7617  ( .A(\Data_Mem/n7594 ), .B(\Data_Mem/n7587 ), .S(N26), 
        .Z(\Data_Mem/n7595 ) );
  MUX \Data_Mem/U7616  ( .A(\Data_Mem/n7593 ), .B(\Data_Mem/n7590 ), .S(N27), 
        .Z(\Data_Mem/n7594 ) );
  MUX \Data_Mem/U7615  ( .A(\Data_Mem/n7592 ), .B(\Data_Mem/n7591 ), .S(N28), 
        .Z(\Data_Mem/n7593 ) );
  MUX \Data_Mem/U7614  ( .A(data_mem_out_wire[1045]), .B(
        data_mem_out_wire[1077]), .S(N29), .Z(\Data_Mem/n7592 ) );
  MUX \Data_Mem/U7613  ( .A(data_mem_out_wire[1109]), .B(
        data_mem_out_wire[1141]), .S(N29), .Z(\Data_Mem/n7591 ) );
  MUX \Data_Mem/U7612  ( .A(\Data_Mem/n7589 ), .B(\Data_Mem/n7588 ), .S(N28), 
        .Z(\Data_Mem/n7590 ) );
  MUX \Data_Mem/U7611  ( .A(data_mem_out_wire[1173]), .B(
        data_mem_out_wire[1205]), .S(N29), .Z(\Data_Mem/n7589 ) );
  MUX \Data_Mem/U7610  ( .A(data_mem_out_wire[1237]), .B(
        data_mem_out_wire[1269]), .S(N29), .Z(\Data_Mem/n7588 ) );
  MUX \Data_Mem/U7609  ( .A(\Data_Mem/n7586 ), .B(\Data_Mem/n7583 ), .S(N27), 
        .Z(\Data_Mem/n7587 ) );
  MUX \Data_Mem/U7608  ( .A(\Data_Mem/n7585 ), .B(\Data_Mem/n7584 ), .S(N28), 
        .Z(\Data_Mem/n7586 ) );
  MUX \Data_Mem/U7607  ( .A(data_mem_out_wire[1301]), .B(
        data_mem_out_wire[1333]), .S(N29), .Z(\Data_Mem/n7585 ) );
  MUX \Data_Mem/U7606  ( .A(data_mem_out_wire[1365]), .B(
        data_mem_out_wire[1397]), .S(N29), .Z(\Data_Mem/n7584 ) );
  MUX \Data_Mem/U7605  ( .A(\Data_Mem/n7582 ), .B(\Data_Mem/n7581 ), .S(N28), 
        .Z(\Data_Mem/n7583 ) );
  MUX \Data_Mem/U7604  ( .A(data_mem_out_wire[1429]), .B(
        data_mem_out_wire[1461]), .S(N29), .Z(\Data_Mem/n7582 ) );
  MUX \Data_Mem/U7603  ( .A(data_mem_out_wire[1493]), .B(
        data_mem_out_wire[1525]), .S(N29), .Z(\Data_Mem/n7581 ) );
  MUX \Data_Mem/U7602  ( .A(\Data_Mem/n7579 ), .B(\Data_Mem/n7572 ), .S(N26), 
        .Z(\Data_Mem/n7580 ) );
  MUX \Data_Mem/U7601  ( .A(\Data_Mem/n7578 ), .B(\Data_Mem/n7575 ), .S(N27), 
        .Z(\Data_Mem/n7579 ) );
  MUX \Data_Mem/U7600  ( .A(\Data_Mem/n7577 ), .B(\Data_Mem/n7576 ), .S(N28), 
        .Z(\Data_Mem/n7578 ) );
  MUX \Data_Mem/U7599  ( .A(data_mem_out_wire[1557]), .B(
        data_mem_out_wire[1589]), .S(N29), .Z(\Data_Mem/n7577 ) );
  MUX \Data_Mem/U7598  ( .A(data_mem_out_wire[1621]), .B(
        data_mem_out_wire[1653]), .S(N29), .Z(\Data_Mem/n7576 ) );
  MUX \Data_Mem/U7597  ( .A(\Data_Mem/n7574 ), .B(\Data_Mem/n7573 ), .S(N28), 
        .Z(\Data_Mem/n7575 ) );
  MUX \Data_Mem/U7596  ( .A(data_mem_out_wire[1685]), .B(
        data_mem_out_wire[1717]), .S(N29), .Z(\Data_Mem/n7574 ) );
  MUX \Data_Mem/U7595  ( .A(data_mem_out_wire[1749]), .B(
        data_mem_out_wire[1781]), .S(N29), .Z(\Data_Mem/n7573 ) );
  MUX \Data_Mem/U7594  ( .A(\Data_Mem/n7571 ), .B(\Data_Mem/n7568 ), .S(N27), 
        .Z(\Data_Mem/n7572 ) );
  MUX \Data_Mem/U7593  ( .A(\Data_Mem/n7570 ), .B(\Data_Mem/n7569 ), .S(N28), 
        .Z(\Data_Mem/n7571 ) );
  MUX \Data_Mem/U7592  ( .A(data_mem_out_wire[1813]), .B(
        data_mem_out_wire[1845]), .S(N29), .Z(\Data_Mem/n7570 ) );
  MUX \Data_Mem/U7591  ( .A(data_mem_out_wire[1877]), .B(
        data_mem_out_wire[1909]), .S(N29), .Z(\Data_Mem/n7569 ) );
  MUX \Data_Mem/U7590  ( .A(\Data_Mem/n7567 ), .B(\Data_Mem/n7566 ), .S(N28), 
        .Z(\Data_Mem/n7568 ) );
  MUX \Data_Mem/U7589  ( .A(data_mem_out_wire[1941]), .B(
        data_mem_out_wire[1973]), .S(N29), .Z(\Data_Mem/n7567 ) );
  MUX \Data_Mem/U7588  ( .A(data_mem_out_wire[2005]), .B(
        data_mem_out_wire[2037]), .S(N29), .Z(\Data_Mem/n7566 ) );
  MUX \Data_Mem/U7587  ( .A(\Data_Mem/n7565 ), .B(\Data_Mem/n7534 ), .S(N24), 
        .Z(c_memory[20]) );
  MUX \Data_Mem/U7586  ( .A(\Data_Mem/n7564 ), .B(\Data_Mem/n7549 ), .S(N25), 
        .Z(\Data_Mem/n7565 ) );
  MUX \Data_Mem/U7585  ( .A(\Data_Mem/n7563 ), .B(\Data_Mem/n7556 ), .S(N26), 
        .Z(\Data_Mem/n7564 ) );
  MUX \Data_Mem/U7584  ( .A(\Data_Mem/n7562 ), .B(\Data_Mem/n7559 ), .S(N27), 
        .Z(\Data_Mem/n7563 ) );
  MUX \Data_Mem/U7583  ( .A(\Data_Mem/n7561 ), .B(\Data_Mem/n7560 ), .S(N28), 
        .Z(\Data_Mem/n7562 ) );
  MUX \Data_Mem/U7582  ( .A(data_mem_out_wire[20]), .B(data_mem_out_wire[52]), 
        .S(N29), .Z(\Data_Mem/n7561 ) );
  MUX \Data_Mem/U7581  ( .A(data_mem_out_wire[84]), .B(data_mem_out_wire[116]), 
        .S(N29), .Z(\Data_Mem/n7560 ) );
  MUX \Data_Mem/U7580  ( .A(\Data_Mem/n7558 ), .B(\Data_Mem/n7557 ), .S(N28), 
        .Z(\Data_Mem/n7559 ) );
  MUX \Data_Mem/U7579  ( .A(data_mem_out_wire[148]), .B(data_mem_out_wire[180]), .S(N29), .Z(\Data_Mem/n7558 ) );
  MUX \Data_Mem/U7578  ( .A(data_mem_out_wire[212]), .B(data_mem_out_wire[244]), .S(N29), .Z(\Data_Mem/n7557 ) );
  MUX \Data_Mem/U7577  ( .A(\Data_Mem/n7555 ), .B(\Data_Mem/n7552 ), .S(N27), 
        .Z(\Data_Mem/n7556 ) );
  MUX \Data_Mem/U7576  ( .A(\Data_Mem/n7554 ), .B(\Data_Mem/n7553 ), .S(N28), 
        .Z(\Data_Mem/n7555 ) );
  MUX \Data_Mem/U7575  ( .A(data_mem_out_wire[276]), .B(data_mem_out_wire[308]), .S(N29), .Z(\Data_Mem/n7554 ) );
  MUX \Data_Mem/U7574  ( .A(data_mem_out_wire[340]), .B(data_mem_out_wire[372]), .S(N29), .Z(\Data_Mem/n7553 ) );
  MUX \Data_Mem/U7573  ( .A(\Data_Mem/n7551 ), .B(\Data_Mem/n7550 ), .S(N28), 
        .Z(\Data_Mem/n7552 ) );
  MUX \Data_Mem/U7572  ( .A(data_mem_out_wire[404]), .B(data_mem_out_wire[436]), .S(N29), .Z(\Data_Mem/n7551 ) );
  MUX \Data_Mem/U7571  ( .A(data_mem_out_wire[468]), .B(data_mem_out_wire[500]), .S(N29), .Z(\Data_Mem/n7550 ) );
  MUX \Data_Mem/U7570  ( .A(\Data_Mem/n7548 ), .B(\Data_Mem/n7541 ), .S(N26), 
        .Z(\Data_Mem/n7549 ) );
  MUX \Data_Mem/U7569  ( .A(\Data_Mem/n7547 ), .B(\Data_Mem/n7544 ), .S(N27), 
        .Z(\Data_Mem/n7548 ) );
  MUX \Data_Mem/U7568  ( .A(\Data_Mem/n7546 ), .B(\Data_Mem/n7545 ), .S(N28), 
        .Z(\Data_Mem/n7547 ) );
  MUX \Data_Mem/U7567  ( .A(data_mem_out_wire[532]), .B(data_mem_out_wire[564]), .S(N29), .Z(\Data_Mem/n7546 ) );
  MUX \Data_Mem/U7566  ( .A(data_mem_out_wire[596]), .B(data_mem_out_wire[628]), .S(N29), .Z(\Data_Mem/n7545 ) );
  MUX \Data_Mem/U7565  ( .A(\Data_Mem/n7543 ), .B(\Data_Mem/n7542 ), .S(N28), 
        .Z(\Data_Mem/n7544 ) );
  MUX \Data_Mem/U7564  ( .A(data_mem_out_wire[660]), .B(data_mem_out_wire[692]), .S(N29), .Z(\Data_Mem/n7543 ) );
  MUX \Data_Mem/U7563  ( .A(data_mem_out_wire[724]), .B(data_mem_out_wire[756]), .S(N29), .Z(\Data_Mem/n7542 ) );
  MUX \Data_Mem/U7562  ( .A(\Data_Mem/n7540 ), .B(\Data_Mem/n7537 ), .S(N27), 
        .Z(\Data_Mem/n7541 ) );
  MUX \Data_Mem/U7561  ( .A(\Data_Mem/n7539 ), .B(\Data_Mem/n7538 ), .S(N28), 
        .Z(\Data_Mem/n7540 ) );
  MUX \Data_Mem/U7560  ( .A(data_mem_out_wire[788]), .B(data_mem_out_wire[820]), .S(N29), .Z(\Data_Mem/n7539 ) );
  MUX \Data_Mem/U7559  ( .A(data_mem_out_wire[852]), .B(data_mem_out_wire[884]), .S(N29), .Z(\Data_Mem/n7538 ) );
  MUX \Data_Mem/U7558  ( .A(\Data_Mem/n7536 ), .B(\Data_Mem/n7535 ), .S(N28), 
        .Z(\Data_Mem/n7537 ) );
  MUX \Data_Mem/U7557  ( .A(data_mem_out_wire[916]), .B(data_mem_out_wire[948]), .S(N29), .Z(\Data_Mem/n7536 ) );
  MUX \Data_Mem/U7556  ( .A(data_mem_out_wire[980]), .B(
        data_mem_out_wire[1012]), .S(N29), .Z(\Data_Mem/n7535 ) );
  MUX \Data_Mem/U7555  ( .A(\Data_Mem/n7533 ), .B(\Data_Mem/n7518 ), .S(N25), 
        .Z(\Data_Mem/n7534 ) );
  MUX \Data_Mem/U7554  ( .A(\Data_Mem/n7532 ), .B(\Data_Mem/n7525 ), .S(N26), 
        .Z(\Data_Mem/n7533 ) );
  MUX \Data_Mem/U7553  ( .A(\Data_Mem/n7531 ), .B(\Data_Mem/n7528 ), .S(N27), 
        .Z(\Data_Mem/n7532 ) );
  MUX \Data_Mem/U7552  ( .A(\Data_Mem/n7530 ), .B(\Data_Mem/n7529 ), .S(N28), 
        .Z(\Data_Mem/n7531 ) );
  MUX \Data_Mem/U7551  ( .A(data_mem_out_wire[1044]), .B(
        data_mem_out_wire[1076]), .S(N29), .Z(\Data_Mem/n7530 ) );
  MUX \Data_Mem/U7550  ( .A(data_mem_out_wire[1108]), .B(
        data_mem_out_wire[1140]), .S(N29), .Z(\Data_Mem/n7529 ) );
  MUX \Data_Mem/U7549  ( .A(\Data_Mem/n7527 ), .B(\Data_Mem/n7526 ), .S(N28), 
        .Z(\Data_Mem/n7528 ) );
  MUX \Data_Mem/U7548  ( .A(data_mem_out_wire[1172]), .B(
        data_mem_out_wire[1204]), .S(N29), .Z(\Data_Mem/n7527 ) );
  MUX \Data_Mem/U7547  ( .A(data_mem_out_wire[1236]), .B(
        data_mem_out_wire[1268]), .S(N29), .Z(\Data_Mem/n7526 ) );
  MUX \Data_Mem/U7546  ( .A(\Data_Mem/n7524 ), .B(\Data_Mem/n7521 ), .S(N27), 
        .Z(\Data_Mem/n7525 ) );
  MUX \Data_Mem/U7545  ( .A(\Data_Mem/n7523 ), .B(\Data_Mem/n7522 ), .S(N28), 
        .Z(\Data_Mem/n7524 ) );
  MUX \Data_Mem/U7544  ( .A(data_mem_out_wire[1300]), .B(
        data_mem_out_wire[1332]), .S(N29), .Z(\Data_Mem/n7523 ) );
  MUX \Data_Mem/U7543  ( .A(data_mem_out_wire[1364]), .B(
        data_mem_out_wire[1396]), .S(N29), .Z(\Data_Mem/n7522 ) );
  MUX \Data_Mem/U7542  ( .A(\Data_Mem/n7520 ), .B(\Data_Mem/n7519 ), .S(N28), 
        .Z(\Data_Mem/n7521 ) );
  MUX \Data_Mem/U7541  ( .A(data_mem_out_wire[1428]), .B(
        data_mem_out_wire[1460]), .S(N29), .Z(\Data_Mem/n7520 ) );
  MUX \Data_Mem/U7540  ( .A(data_mem_out_wire[1492]), .B(
        data_mem_out_wire[1524]), .S(N29), .Z(\Data_Mem/n7519 ) );
  MUX \Data_Mem/U7539  ( .A(\Data_Mem/n7517 ), .B(\Data_Mem/n7510 ), .S(N26), 
        .Z(\Data_Mem/n7518 ) );
  MUX \Data_Mem/U7538  ( .A(\Data_Mem/n7516 ), .B(\Data_Mem/n7513 ), .S(N27), 
        .Z(\Data_Mem/n7517 ) );
  MUX \Data_Mem/U7537  ( .A(\Data_Mem/n7515 ), .B(\Data_Mem/n7514 ), .S(N28), 
        .Z(\Data_Mem/n7516 ) );
  MUX \Data_Mem/U7536  ( .A(data_mem_out_wire[1556]), .B(
        data_mem_out_wire[1588]), .S(N29), .Z(\Data_Mem/n7515 ) );
  MUX \Data_Mem/U7535  ( .A(data_mem_out_wire[1620]), .B(
        data_mem_out_wire[1652]), .S(N29), .Z(\Data_Mem/n7514 ) );
  MUX \Data_Mem/U7534  ( .A(\Data_Mem/n7512 ), .B(\Data_Mem/n7511 ), .S(N28), 
        .Z(\Data_Mem/n7513 ) );
  MUX \Data_Mem/U7533  ( .A(data_mem_out_wire[1684]), .B(
        data_mem_out_wire[1716]), .S(N29), .Z(\Data_Mem/n7512 ) );
  MUX \Data_Mem/U7532  ( .A(data_mem_out_wire[1748]), .B(
        data_mem_out_wire[1780]), .S(N29), .Z(\Data_Mem/n7511 ) );
  MUX \Data_Mem/U7531  ( .A(\Data_Mem/n7509 ), .B(\Data_Mem/n7506 ), .S(N27), 
        .Z(\Data_Mem/n7510 ) );
  MUX \Data_Mem/U7530  ( .A(\Data_Mem/n7508 ), .B(\Data_Mem/n7507 ), .S(N28), 
        .Z(\Data_Mem/n7509 ) );
  MUX \Data_Mem/U7529  ( .A(data_mem_out_wire[1812]), .B(
        data_mem_out_wire[1844]), .S(N29), .Z(\Data_Mem/n7508 ) );
  MUX \Data_Mem/U7528  ( .A(data_mem_out_wire[1876]), .B(
        data_mem_out_wire[1908]), .S(N29), .Z(\Data_Mem/n7507 ) );
  MUX \Data_Mem/U7527  ( .A(\Data_Mem/n7505 ), .B(\Data_Mem/n7504 ), .S(N28), 
        .Z(\Data_Mem/n7506 ) );
  MUX \Data_Mem/U7526  ( .A(data_mem_out_wire[1940]), .B(
        data_mem_out_wire[1972]), .S(N29), .Z(\Data_Mem/n7505 ) );
  MUX \Data_Mem/U7525  ( .A(data_mem_out_wire[2004]), .B(
        data_mem_out_wire[2036]), .S(N29), .Z(\Data_Mem/n7504 ) );
  MUX \Data_Mem/U7524  ( .A(\Data_Mem/n7503 ), .B(\Data_Mem/n7472 ), .S(N24), 
        .Z(c_memory[19]) );
  MUX \Data_Mem/U7523  ( .A(\Data_Mem/n7502 ), .B(\Data_Mem/n7487 ), .S(N25), 
        .Z(\Data_Mem/n7503 ) );
  MUX \Data_Mem/U7522  ( .A(\Data_Mem/n7501 ), .B(\Data_Mem/n7494 ), .S(N26), 
        .Z(\Data_Mem/n7502 ) );
  MUX \Data_Mem/U7521  ( .A(\Data_Mem/n7500 ), .B(\Data_Mem/n7497 ), .S(N27), 
        .Z(\Data_Mem/n7501 ) );
  MUX \Data_Mem/U7520  ( .A(\Data_Mem/n7499 ), .B(\Data_Mem/n7498 ), .S(N28), 
        .Z(\Data_Mem/n7500 ) );
  MUX \Data_Mem/U7519  ( .A(data_mem_out_wire[19]), .B(data_mem_out_wire[51]), 
        .S(N29), .Z(\Data_Mem/n7499 ) );
  MUX \Data_Mem/U7518  ( .A(data_mem_out_wire[83]), .B(data_mem_out_wire[115]), 
        .S(N29), .Z(\Data_Mem/n7498 ) );
  MUX \Data_Mem/U7517  ( .A(\Data_Mem/n7496 ), .B(\Data_Mem/n7495 ), .S(N28), 
        .Z(\Data_Mem/n7497 ) );
  MUX \Data_Mem/U7516  ( .A(data_mem_out_wire[147]), .B(data_mem_out_wire[179]), .S(N29), .Z(\Data_Mem/n7496 ) );
  MUX \Data_Mem/U7515  ( .A(data_mem_out_wire[211]), .B(data_mem_out_wire[243]), .S(N29), .Z(\Data_Mem/n7495 ) );
  MUX \Data_Mem/U7514  ( .A(\Data_Mem/n7493 ), .B(\Data_Mem/n7490 ), .S(N27), 
        .Z(\Data_Mem/n7494 ) );
  MUX \Data_Mem/U7513  ( .A(\Data_Mem/n7492 ), .B(\Data_Mem/n7491 ), .S(N28), 
        .Z(\Data_Mem/n7493 ) );
  MUX \Data_Mem/U7512  ( .A(data_mem_out_wire[275]), .B(data_mem_out_wire[307]), .S(N29), .Z(\Data_Mem/n7492 ) );
  MUX \Data_Mem/U7511  ( .A(data_mem_out_wire[339]), .B(data_mem_out_wire[371]), .S(N29), .Z(\Data_Mem/n7491 ) );
  MUX \Data_Mem/U7510  ( .A(\Data_Mem/n7489 ), .B(\Data_Mem/n7488 ), .S(N28), 
        .Z(\Data_Mem/n7490 ) );
  MUX \Data_Mem/U7509  ( .A(data_mem_out_wire[403]), .B(data_mem_out_wire[435]), .S(N29), .Z(\Data_Mem/n7489 ) );
  MUX \Data_Mem/U7508  ( .A(data_mem_out_wire[467]), .B(data_mem_out_wire[499]), .S(N29), .Z(\Data_Mem/n7488 ) );
  MUX \Data_Mem/U7507  ( .A(\Data_Mem/n7486 ), .B(\Data_Mem/n7479 ), .S(N26), 
        .Z(\Data_Mem/n7487 ) );
  MUX \Data_Mem/U7506  ( .A(\Data_Mem/n7485 ), .B(\Data_Mem/n7482 ), .S(N27), 
        .Z(\Data_Mem/n7486 ) );
  MUX \Data_Mem/U7505  ( .A(\Data_Mem/n7484 ), .B(\Data_Mem/n7483 ), .S(N28), 
        .Z(\Data_Mem/n7485 ) );
  MUX \Data_Mem/U7504  ( .A(data_mem_out_wire[531]), .B(data_mem_out_wire[563]), .S(N29), .Z(\Data_Mem/n7484 ) );
  MUX \Data_Mem/U7503  ( .A(data_mem_out_wire[595]), .B(data_mem_out_wire[627]), .S(N29), .Z(\Data_Mem/n7483 ) );
  MUX \Data_Mem/U7502  ( .A(\Data_Mem/n7481 ), .B(\Data_Mem/n7480 ), .S(N28), 
        .Z(\Data_Mem/n7482 ) );
  MUX \Data_Mem/U7501  ( .A(data_mem_out_wire[659]), .B(data_mem_out_wire[691]), .S(N29), .Z(\Data_Mem/n7481 ) );
  MUX \Data_Mem/U7500  ( .A(data_mem_out_wire[723]), .B(data_mem_out_wire[755]), .S(N29), .Z(\Data_Mem/n7480 ) );
  MUX \Data_Mem/U7499  ( .A(\Data_Mem/n7478 ), .B(\Data_Mem/n7475 ), .S(N27), 
        .Z(\Data_Mem/n7479 ) );
  MUX \Data_Mem/U7498  ( .A(\Data_Mem/n7477 ), .B(\Data_Mem/n7476 ), .S(N28), 
        .Z(\Data_Mem/n7478 ) );
  MUX \Data_Mem/U7497  ( .A(data_mem_out_wire[787]), .B(data_mem_out_wire[819]), .S(N29), .Z(\Data_Mem/n7477 ) );
  MUX \Data_Mem/U7496  ( .A(data_mem_out_wire[851]), .B(data_mem_out_wire[883]), .S(N29), .Z(\Data_Mem/n7476 ) );
  MUX \Data_Mem/U7495  ( .A(\Data_Mem/n7474 ), .B(\Data_Mem/n7473 ), .S(N28), 
        .Z(\Data_Mem/n7475 ) );
  MUX \Data_Mem/U7494  ( .A(data_mem_out_wire[915]), .B(data_mem_out_wire[947]), .S(N29), .Z(\Data_Mem/n7474 ) );
  MUX \Data_Mem/U7493  ( .A(data_mem_out_wire[979]), .B(
        data_mem_out_wire[1011]), .S(N29), .Z(\Data_Mem/n7473 ) );
  MUX \Data_Mem/U7492  ( .A(\Data_Mem/n7471 ), .B(\Data_Mem/n7456 ), .S(N25), 
        .Z(\Data_Mem/n7472 ) );
  MUX \Data_Mem/U7491  ( .A(\Data_Mem/n7470 ), .B(\Data_Mem/n7463 ), .S(N26), 
        .Z(\Data_Mem/n7471 ) );
  MUX \Data_Mem/U7490  ( .A(\Data_Mem/n7469 ), .B(\Data_Mem/n7466 ), .S(N27), 
        .Z(\Data_Mem/n7470 ) );
  MUX \Data_Mem/U7489  ( .A(\Data_Mem/n7468 ), .B(\Data_Mem/n7467 ), .S(N28), 
        .Z(\Data_Mem/n7469 ) );
  MUX \Data_Mem/U7488  ( .A(data_mem_out_wire[1043]), .B(
        data_mem_out_wire[1075]), .S(N29), .Z(\Data_Mem/n7468 ) );
  MUX \Data_Mem/U7487  ( .A(data_mem_out_wire[1107]), .B(
        data_mem_out_wire[1139]), .S(N29), .Z(\Data_Mem/n7467 ) );
  MUX \Data_Mem/U7486  ( .A(\Data_Mem/n7465 ), .B(\Data_Mem/n7464 ), .S(N28), 
        .Z(\Data_Mem/n7466 ) );
  MUX \Data_Mem/U7485  ( .A(data_mem_out_wire[1171]), .B(
        data_mem_out_wire[1203]), .S(N29), .Z(\Data_Mem/n7465 ) );
  MUX \Data_Mem/U7484  ( .A(data_mem_out_wire[1235]), .B(
        data_mem_out_wire[1267]), .S(N29), .Z(\Data_Mem/n7464 ) );
  MUX \Data_Mem/U7483  ( .A(\Data_Mem/n7462 ), .B(\Data_Mem/n7459 ), .S(N27), 
        .Z(\Data_Mem/n7463 ) );
  MUX \Data_Mem/U7482  ( .A(\Data_Mem/n7461 ), .B(\Data_Mem/n7460 ), .S(N28), 
        .Z(\Data_Mem/n7462 ) );
  MUX \Data_Mem/U7481  ( .A(data_mem_out_wire[1299]), .B(
        data_mem_out_wire[1331]), .S(N29), .Z(\Data_Mem/n7461 ) );
  MUX \Data_Mem/U7480  ( .A(data_mem_out_wire[1363]), .B(
        data_mem_out_wire[1395]), .S(N29), .Z(\Data_Mem/n7460 ) );
  MUX \Data_Mem/U7479  ( .A(\Data_Mem/n7458 ), .B(\Data_Mem/n7457 ), .S(N28), 
        .Z(\Data_Mem/n7459 ) );
  MUX \Data_Mem/U7478  ( .A(data_mem_out_wire[1427]), .B(
        data_mem_out_wire[1459]), .S(N29), .Z(\Data_Mem/n7458 ) );
  MUX \Data_Mem/U7477  ( .A(data_mem_out_wire[1491]), .B(
        data_mem_out_wire[1523]), .S(N29), .Z(\Data_Mem/n7457 ) );
  MUX \Data_Mem/U7476  ( .A(\Data_Mem/n7455 ), .B(\Data_Mem/n7448 ), .S(N26), 
        .Z(\Data_Mem/n7456 ) );
  MUX \Data_Mem/U7475  ( .A(\Data_Mem/n7454 ), .B(\Data_Mem/n7451 ), .S(N27), 
        .Z(\Data_Mem/n7455 ) );
  MUX \Data_Mem/U7474  ( .A(\Data_Mem/n7453 ), .B(\Data_Mem/n7452 ), .S(N28), 
        .Z(\Data_Mem/n7454 ) );
  MUX \Data_Mem/U7473  ( .A(data_mem_out_wire[1555]), .B(
        data_mem_out_wire[1587]), .S(N29), .Z(\Data_Mem/n7453 ) );
  MUX \Data_Mem/U7472  ( .A(data_mem_out_wire[1619]), .B(
        data_mem_out_wire[1651]), .S(N29), .Z(\Data_Mem/n7452 ) );
  MUX \Data_Mem/U7471  ( .A(\Data_Mem/n7450 ), .B(\Data_Mem/n7449 ), .S(N28), 
        .Z(\Data_Mem/n7451 ) );
  MUX \Data_Mem/U7470  ( .A(data_mem_out_wire[1683]), .B(
        data_mem_out_wire[1715]), .S(N29), .Z(\Data_Mem/n7450 ) );
  MUX \Data_Mem/U7469  ( .A(data_mem_out_wire[1747]), .B(
        data_mem_out_wire[1779]), .S(N29), .Z(\Data_Mem/n7449 ) );
  MUX \Data_Mem/U7468  ( .A(\Data_Mem/n7447 ), .B(\Data_Mem/n7444 ), .S(N27), 
        .Z(\Data_Mem/n7448 ) );
  MUX \Data_Mem/U7467  ( .A(\Data_Mem/n7446 ), .B(\Data_Mem/n7445 ), .S(N28), 
        .Z(\Data_Mem/n7447 ) );
  MUX \Data_Mem/U7466  ( .A(data_mem_out_wire[1811]), .B(
        data_mem_out_wire[1843]), .S(N29), .Z(\Data_Mem/n7446 ) );
  MUX \Data_Mem/U7465  ( .A(data_mem_out_wire[1875]), .B(
        data_mem_out_wire[1907]), .S(N29), .Z(\Data_Mem/n7445 ) );
  MUX \Data_Mem/U7464  ( .A(\Data_Mem/n7443 ), .B(\Data_Mem/n7442 ), .S(N28), 
        .Z(\Data_Mem/n7444 ) );
  MUX \Data_Mem/U7463  ( .A(data_mem_out_wire[1939]), .B(
        data_mem_out_wire[1971]), .S(N29), .Z(\Data_Mem/n7443 ) );
  MUX \Data_Mem/U7462  ( .A(data_mem_out_wire[2003]), .B(
        data_mem_out_wire[2035]), .S(N29), .Z(\Data_Mem/n7442 ) );
  MUX \Data_Mem/U7461  ( .A(\Data_Mem/n7441 ), .B(\Data_Mem/n7410 ), .S(N24), 
        .Z(c_memory[18]) );
  MUX \Data_Mem/U7460  ( .A(\Data_Mem/n7440 ), .B(\Data_Mem/n7425 ), .S(N25), 
        .Z(\Data_Mem/n7441 ) );
  MUX \Data_Mem/U7459  ( .A(\Data_Mem/n7439 ), .B(\Data_Mem/n7432 ), .S(N26), 
        .Z(\Data_Mem/n7440 ) );
  MUX \Data_Mem/U7458  ( .A(\Data_Mem/n7438 ), .B(\Data_Mem/n7435 ), .S(N27), 
        .Z(\Data_Mem/n7439 ) );
  MUX \Data_Mem/U7457  ( .A(\Data_Mem/n7437 ), .B(\Data_Mem/n7436 ), .S(N28), 
        .Z(\Data_Mem/n7438 ) );
  MUX \Data_Mem/U7456  ( .A(data_mem_out_wire[18]), .B(data_mem_out_wire[50]), 
        .S(N29), .Z(\Data_Mem/n7437 ) );
  MUX \Data_Mem/U7455  ( .A(data_mem_out_wire[82]), .B(data_mem_out_wire[114]), 
        .S(N29), .Z(\Data_Mem/n7436 ) );
  MUX \Data_Mem/U7454  ( .A(\Data_Mem/n7434 ), .B(\Data_Mem/n7433 ), .S(N28), 
        .Z(\Data_Mem/n7435 ) );
  MUX \Data_Mem/U7453  ( .A(data_mem_out_wire[146]), .B(data_mem_out_wire[178]), .S(N29), .Z(\Data_Mem/n7434 ) );
  MUX \Data_Mem/U7452  ( .A(data_mem_out_wire[210]), .B(data_mem_out_wire[242]), .S(N29), .Z(\Data_Mem/n7433 ) );
  MUX \Data_Mem/U7451  ( .A(\Data_Mem/n7431 ), .B(\Data_Mem/n7428 ), .S(N27), 
        .Z(\Data_Mem/n7432 ) );
  MUX \Data_Mem/U7450  ( .A(\Data_Mem/n7430 ), .B(\Data_Mem/n7429 ), .S(N28), 
        .Z(\Data_Mem/n7431 ) );
  MUX \Data_Mem/U7449  ( .A(data_mem_out_wire[274]), .B(data_mem_out_wire[306]), .S(N29), .Z(\Data_Mem/n7430 ) );
  MUX \Data_Mem/U7448  ( .A(data_mem_out_wire[338]), .B(data_mem_out_wire[370]), .S(N29), .Z(\Data_Mem/n7429 ) );
  MUX \Data_Mem/U7447  ( .A(\Data_Mem/n7427 ), .B(\Data_Mem/n7426 ), .S(N28), 
        .Z(\Data_Mem/n7428 ) );
  MUX \Data_Mem/U7446  ( .A(data_mem_out_wire[402]), .B(data_mem_out_wire[434]), .S(N29), .Z(\Data_Mem/n7427 ) );
  MUX \Data_Mem/U7445  ( .A(data_mem_out_wire[466]), .B(data_mem_out_wire[498]), .S(N29), .Z(\Data_Mem/n7426 ) );
  MUX \Data_Mem/U7444  ( .A(\Data_Mem/n7424 ), .B(\Data_Mem/n7417 ), .S(N26), 
        .Z(\Data_Mem/n7425 ) );
  MUX \Data_Mem/U7443  ( .A(\Data_Mem/n7423 ), .B(\Data_Mem/n7420 ), .S(N27), 
        .Z(\Data_Mem/n7424 ) );
  MUX \Data_Mem/U7442  ( .A(\Data_Mem/n7422 ), .B(\Data_Mem/n7421 ), .S(N28), 
        .Z(\Data_Mem/n7423 ) );
  MUX \Data_Mem/U7441  ( .A(data_mem_out_wire[530]), .B(data_mem_out_wire[562]), .S(N29), .Z(\Data_Mem/n7422 ) );
  MUX \Data_Mem/U7440  ( .A(data_mem_out_wire[594]), .B(data_mem_out_wire[626]), .S(N29), .Z(\Data_Mem/n7421 ) );
  MUX \Data_Mem/U7439  ( .A(\Data_Mem/n7419 ), .B(\Data_Mem/n7418 ), .S(N28), 
        .Z(\Data_Mem/n7420 ) );
  MUX \Data_Mem/U7438  ( .A(data_mem_out_wire[658]), .B(data_mem_out_wire[690]), .S(N29), .Z(\Data_Mem/n7419 ) );
  MUX \Data_Mem/U7437  ( .A(data_mem_out_wire[722]), .B(data_mem_out_wire[754]), .S(N29), .Z(\Data_Mem/n7418 ) );
  MUX \Data_Mem/U7436  ( .A(\Data_Mem/n7416 ), .B(\Data_Mem/n7413 ), .S(N27), 
        .Z(\Data_Mem/n7417 ) );
  MUX \Data_Mem/U7435  ( .A(\Data_Mem/n7415 ), .B(\Data_Mem/n7414 ), .S(N28), 
        .Z(\Data_Mem/n7416 ) );
  MUX \Data_Mem/U7434  ( .A(data_mem_out_wire[786]), .B(data_mem_out_wire[818]), .S(N29), .Z(\Data_Mem/n7415 ) );
  MUX \Data_Mem/U7433  ( .A(data_mem_out_wire[850]), .B(data_mem_out_wire[882]), .S(N29), .Z(\Data_Mem/n7414 ) );
  MUX \Data_Mem/U7432  ( .A(\Data_Mem/n7412 ), .B(\Data_Mem/n7411 ), .S(N28), 
        .Z(\Data_Mem/n7413 ) );
  MUX \Data_Mem/U7431  ( .A(data_mem_out_wire[914]), .B(data_mem_out_wire[946]), .S(N29), .Z(\Data_Mem/n7412 ) );
  MUX \Data_Mem/U7430  ( .A(data_mem_out_wire[978]), .B(
        data_mem_out_wire[1010]), .S(N29), .Z(\Data_Mem/n7411 ) );
  MUX \Data_Mem/U7429  ( .A(\Data_Mem/n7409 ), .B(\Data_Mem/n7394 ), .S(N25), 
        .Z(\Data_Mem/n7410 ) );
  MUX \Data_Mem/U7428  ( .A(\Data_Mem/n7408 ), .B(\Data_Mem/n7401 ), .S(N26), 
        .Z(\Data_Mem/n7409 ) );
  MUX \Data_Mem/U7427  ( .A(\Data_Mem/n7407 ), .B(\Data_Mem/n7404 ), .S(N27), 
        .Z(\Data_Mem/n7408 ) );
  MUX \Data_Mem/U7426  ( .A(\Data_Mem/n7406 ), .B(\Data_Mem/n7405 ), .S(N28), 
        .Z(\Data_Mem/n7407 ) );
  MUX \Data_Mem/U7425  ( .A(data_mem_out_wire[1042]), .B(
        data_mem_out_wire[1074]), .S(N29), .Z(\Data_Mem/n7406 ) );
  MUX \Data_Mem/U7424  ( .A(data_mem_out_wire[1106]), .B(
        data_mem_out_wire[1138]), .S(N29), .Z(\Data_Mem/n7405 ) );
  MUX \Data_Mem/U7423  ( .A(\Data_Mem/n7403 ), .B(\Data_Mem/n7402 ), .S(N28), 
        .Z(\Data_Mem/n7404 ) );
  MUX \Data_Mem/U7422  ( .A(data_mem_out_wire[1170]), .B(
        data_mem_out_wire[1202]), .S(N29), .Z(\Data_Mem/n7403 ) );
  MUX \Data_Mem/U7421  ( .A(data_mem_out_wire[1234]), .B(
        data_mem_out_wire[1266]), .S(N29), .Z(\Data_Mem/n7402 ) );
  MUX \Data_Mem/U7420  ( .A(\Data_Mem/n7400 ), .B(\Data_Mem/n7397 ), .S(N27), 
        .Z(\Data_Mem/n7401 ) );
  MUX \Data_Mem/U7419  ( .A(\Data_Mem/n7399 ), .B(\Data_Mem/n7398 ), .S(N28), 
        .Z(\Data_Mem/n7400 ) );
  MUX \Data_Mem/U7418  ( .A(data_mem_out_wire[1298]), .B(
        data_mem_out_wire[1330]), .S(N29), .Z(\Data_Mem/n7399 ) );
  MUX \Data_Mem/U7417  ( .A(data_mem_out_wire[1362]), .B(
        data_mem_out_wire[1394]), .S(N29), .Z(\Data_Mem/n7398 ) );
  MUX \Data_Mem/U7416  ( .A(\Data_Mem/n7396 ), .B(\Data_Mem/n7395 ), .S(N28), 
        .Z(\Data_Mem/n7397 ) );
  MUX \Data_Mem/U7415  ( .A(data_mem_out_wire[1426]), .B(
        data_mem_out_wire[1458]), .S(N29), .Z(\Data_Mem/n7396 ) );
  MUX \Data_Mem/U7414  ( .A(data_mem_out_wire[1490]), .B(
        data_mem_out_wire[1522]), .S(N29), .Z(\Data_Mem/n7395 ) );
  MUX \Data_Mem/U7413  ( .A(\Data_Mem/n7393 ), .B(\Data_Mem/n7386 ), .S(N26), 
        .Z(\Data_Mem/n7394 ) );
  MUX \Data_Mem/U7412  ( .A(\Data_Mem/n7392 ), .B(\Data_Mem/n7389 ), .S(N27), 
        .Z(\Data_Mem/n7393 ) );
  MUX \Data_Mem/U7411  ( .A(\Data_Mem/n7391 ), .B(\Data_Mem/n7390 ), .S(N28), 
        .Z(\Data_Mem/n7392 ) );
  MUX \Data_Mem/U7410  ( .A(data_mem_out_wire[1554]), .B(
        data_mem_out_wire[1586]), .S(N29), .Z(\Data_Mem/n7391 ) );
  MUX \Data_Mem/U7409  ( .A(data_mem_out_wire[1618]), .B(
        data_mem_out_wire[1650]), .S(N29), .Z(\Data_Mem/n7390 ) );
  MUX \Data_Mem/U7408  ( .A(\Data_Mem/n7388 ), .B(\Data_Mem/n7387 ), .S(N28), 
        .Z(\Data_Mem/n7389 ) );
  MUX \Data_Mem/U7407  ( .A(data_mem_out_wire[1682]), .B(
        data_mem_out_wire[1714]), .S(N29), .Z(\Data_Mem/n7388 ) );
  MUX \Data_Mem/U7406  ( .A(data_mem_out_wire[1746]), .B(
        data_mem_out_wire[1778]), .S(N29), .Z(\Data_Mem/n7387 ) );
  MUX \Data_Mem/U7405  ( .A(\Data_Mem/n7385 ), .B(\Data_Mem/n7382 ), .S(N27), 
        .Z(\Data_Mem/n7386 ) );
  MUX \Data_Mem/U7404  ( .A(\Data_Mem/n7384 ), .B(\Data_Mem/n7383 ), .S(N28), 
        .Z(\Data_Mem/n7385 ) );
  MUX \Data_Mem/U7403  ( .A(data_mem_out_wire[1810]), .B(
        data_mem_out_wire[1842]), .S(N29), .Z(\Data_Mem/n7384 ) );
  MUX \Data_Mem/U7402  ( .A(data_mem_out_wire[1874]), .B(
        data_mem_out_wire[1906]), .S(N29), .Z(\Data_Mem/n7383 ) );
  MUX \Data_Mem/U7401  ( .A(\Data_Mem/n7381 ), .B(\Data_Mem/n7380 ), .S(N28), 
        .Z(\Data_Mem/n7382 ) );
  MUX \Data_Mem/U7400  ( .A(data_mem_out_wire[1938]), .B(
        data_mem_out_wire[1970]), .S(N29), .Z(\Data_Mem/n7381 ) );
  MUX \Data_Mem/U7399  ( .A(data_mem_out_wire[2002]), .B(
        data_mem_out_wire[2034]), .S(N29), .Z(\Data_Mem/n7380 ) );
  MUX \Data_Mem/U7398  ( .A(\Data_Mem/n7379 ), .B(\Data_Mem/n7348 ), .S(N24), 
        .Z(c_memory[17]) );
  MUX \Data_Mem/U7397  ( .A(\Data_Mem/n7378 ), .B(\Data_Mem/n7363 ), .S(N25), 
        .Z(\Data_Mem/n7379 ) );
  MUX \Data_Mem/U7396  ( .A(\Data_Mem/n7377 ), .B(\Data_Mem/n7370 ), .S(N26), 
        .Z(\Data_Mem/n7378 ) );
  MUX \Data_Mem/U7395  ( .A(\Data_Mem/n7376 ), .B(\Data_Mem/n7373 ), .S(N27), 
        .Z(\Data_Mem/n7377 ) );
  MUX \Data_Mem/U7394  ( .A(\Data_Mem/n7375 ), .B(\Data_Mem/n7374 ), .S(N28), 
        .Z(\Data_Mem/n7376 ) );
  MUX \Data_Mem/U7393  ( .A(data_mem_out_wire[17]), .B(data_mem_out_wire[49]), 
        .S(N29), .Z(\Data_Mem/n7375 ) );
  MUX \Data_Mem/U7392  ( .A(data_mem_out_wire[81]), .B(data_mem_out_wire[113]), 
        .S(N29), .Z(\Data_Mem/n7374 ) );
  MUX \Data_Mem/U7391  ( .A(\Data_Mem/n7372 ), .B(\Data_Mem/n7371 ), .S(N28), 
        .Z(\Data_Mem/n7373 ) );
  MUX \Data_Mem/U7390  ( .A(data_mem_out_wire[145]), .B(data_mem_out_wire[177]), .S(N29), .Z(\Data_Mem/n7372 ) );
  MUX \Data_Mem/U7389  ( .A(data_mem_out_wire[209]), .B(data_mem_out_wire[241]), .S(N29), .Z(\Data_Mem/n7371 ) );
  MUX \Data_Mem/U7388  ( .A(\Data_Mem/n7369 ), .B(\Data_Mem/n7366 ), .S(N27), 
        .Z(\Data_Mem/n7370 ) );
  MUX \Data_Mem/U7387  ( .A(\Data_Mem/n7368 ), .B(\Data_Mem/n7367 ), .S(N28), 
        .Z(\Data_Mem/n7369 ) );
  MUX \Data_Mem/U7386  ( .A(data_mem_out_wire[273]), .B(data_mem_out_wire[305]), .S(N29), .Z(\Data_Mem/n7368 ) );
  MUX \Data_Mem/U7385  ( .A(data_mem_out_wire[337]), .B(data_mem_out_wire[369]), .S(N29), .Z(\Data_Mem/n7367 ) );
  MUX \Data_Mem/U7384  ( .A(\Data_Mem/n7365 ), .B(\Data_Mem/n7364 ), .S(N28), 
        .Z(\Data_Mem/n7366 ) );
  MUX \Data_Mem/U7383  ( .A(data_mem_out_wire[401]), .B(data_mem_out_wire[433]), .S(N29), .Z(\Data_Mem/n7365 ) );
  MUX \Data_Mem/U7382  ( .A(data_mem_out_wire[465]), .B(data_mem_out_wire[497]), .S(N29), .Z(\Data_Mem/n7364 ) );
  MUX \Data_Mem/U7381  ( .A(\Data_Mem/n7362 ), .B(\Data_Mem/n7355 ), .S(N26), 
        .Z(\Data_Mem/n7363 ) );
  MUX \Data_Mem/U7380  ( .A(\Data_Mem/n7361 ), .B(\Data_Mem/n7358 ), .S(N27), 
        .Z(\Data_Mem/n7362 ) );
  MUX \Data_Mem/U7379  ( .A(\Data_Mem/n7360 ), .B(\Data_Mem/n7359 ), .S(N28), 
        .Z(\Data_Mem/n7361 ) );
  MUX \Data_Mem/U7378  ( .A(data_mem_out_wire[529]), .B(data_mem_out_wire[561]), .S(N29), .Z(\Data_Mem/n7360 ) );
  MUX \Data_Mem/U7377  ( .A(data_mem_out_wire[593]), .B(data_mem_out_wire[625]), .S(N29), .Z(\Data_Mem/n7359 ) );
  MUX \Data_Mem/U7376  ( .A(\Data_Mem/n7357 ), .B(\Data_Mem/n7356 ), .S(N28), 
        .Z(\Data_Mem/n7358 ) );
  MUX \Data_Mem/U7375  ( .A(data_mem_out_wire[657]), .B(data_mem_out_wire[689]), .S(N29), .Z(\Data_Mem/n7357 ) );
  MUX \Data_Mem/U7374  ( .A(data_mem_out_wire[721]), .B(data_mem_out_wire[753]), .S(N29), .Z(\Data_Mem/n7356 ) );
  MUX \Data_Mem/U7373  ( .A(\Data_Mem/n7354 ), .B(\Data_Mem/n7351 ), .S(N27), 
        .Z(\Data_Mem/n7355 ) );
  MUX \Data_Mem/U7372  ( .A(\Data_Mem/n7353 ), .B(\Data_Mem/n7352 ), .S(N28), 
        .Z(\Data_Mem/n7354 ) );
  MUX \Data_Mem/U7371  ( .A(data_mem_out_wire[785]), .B(data_mem_out_wire[817]), .S(N29), .Z(\Data_Mem/n7353 ) );
  MUX \Data_Mem/U7370  ( .A(data_mem_out_wire[849]), .B(data_mem_out_wire[881]), .S(N29), .Z(\Data_Mem/n7352 ) );
  MUX \Data_Mem/U7369  ( .A(\Data_Mem/n7350 ), .B(\Data_Mem/n7349 ), .S(N28), 
        .Z(\Data_Mem/n7351 ) );
  MUX \Data_Mem/U7368  ( .A(data_mem_out_wire[913]), .B(data_mem_out_wire[945]), .S(N29), .Z(\Data_Mem/n7350 ) );
  MUX \Data_Mem/U7367  ( .A(data_mem_out_wire[977]), .B(
        data_mem_out_wire[1009]), .S(N29), .Z(\Data_Mem/n7349 ) );
  MUX \Data_Mem/U7366  ( .A(\Data_Mem/n7347 ), .B(\Data_Mem/n7332 ), .S(N25), 
        .Z(\Data_Mem/n7348 ) );
  MUX \Data_Mem/U7365  ( .A(\Data_Mem/n7346 ), .B(\Data_Mem/n7339 ), .S(N26), 
        .Z(\Data_Mem/n7347 ) );
  MUX \Data_Mem/U7364  ( .A(\Data_Mem/n7345 ), .B(\Data_Mem/n7342 ), .S(N27), 
        .Z(\Data_Mem/n7346 ) );
  MUX \Data_Mem/U7363  ( .A(\Data_Mem/n7344 ), .B(\Data_Mem/n7343 ), .S(N28), 
        .Z(\Data_Mem/n7345 ) );
  MUX \Data_Mem/U7362  ( .A(data_mem_out_wire[1041]), .B(
        data_mem_out_wire[1073]), .S(N29), .Z(\Data_Mem/n7344 ) );
  MUX \Data_Mem/U7361  ( .A(data_mem_out_wire[1105]), .B(
        data_mem_out_wire[1137]), .S(N29), .Z(\Data_Mem/n7343 ) );
  MUX \Data_Mem/U7360  ( .A(\Data_Mem/n7341 ), .B(\Data_Mem/n7340 ), .S(N28), 
        .Z(\Data_Mem/n7342 ) );
  MUX \Data_Mem/U7359  ( .A(data_mem_out_wire[1169]), .B(
        data_mem_out_wire[1201]), .S(N29), .Z(\Data_Mem/n7341 ) );
  MUX \Data_Mem/U7358  ( .A(data_mem_out_wire[1233]), .B(
        data_mem_out_wire[1265]), .S(N29), .Z(\Data_Mem/n7340 ) );
  MUX \Data_Mem/U7357  ( .A(\Data_Mem/n7338 ), .B(\Data_Mem/n7335 ), .S(N27), 
        .Z(\Data_Mem/n7339 ) );
  MUX \Data_Mem/U7356  ( .A(\Data_Mem/n7337 ), .B(\Data_Mem/n7336 ), .S(N28), 
        .Z(\Data_Mem/n7338 ) );
  MUX \Data_Mem/U7355  ( .A(data_mem_out_wire[1297]), .B(
        data_mem_out_wire[1329]), .S(N29), .Z(\Data_Mem/n7337 ) );
  MUX \Data_Mem/U7354  ( .A(data_mem_out_wire[1361]), .B(
        data_mem_out_wire[1393]), .S(N29), .Z(\Data_Mem/n7336 ) );
  MUX \Data_Mem/U7353  ( .A(\Data_Mem/n7334 ), .B(\Data_Mem/n7333 ), .S(N28), 
        .Z(\Data_Mem/n7335 ) );
  MUX \Data_Mem/U7352  ( .A(data_mem_out_wire[1425]), .B(
        data_mem_out_wire[1457]), .S(N29), .Z(\Data_Mem/n7334 ) );
  MUX \Data_Mem/U7351  ( .A(data_mem_out_wire[1489]), .B(
        data_mem_out_wire[1521]), .S(N29), .Z(\Data_Mem/n7333 ) );
  MUX \Data_Mem/U7350  ( .A(\Data_Mem/n7331 ), .B(\Data_Mem/n7324 ), .S(N26), 
        .Z(\Data_Mem/n7332 ) );
  MUX \Data_Mem/U7349  ( .A(\Data_Mem/n7330 ), .B(\Data_Mem/n7327 ), .S(N27), 
        .Z(\Data_Mem/n7331 ) );
  MUX \Data_Mem/U7348  ( .A(\Data_Mem/n7329 ), .B(\Data_Mem/n7328 ), .S(N28), 
        .Z(\Data_Mem/n7330 ) );
  MUX \Data_Mem/U7347  ( .A(data_mem_out_wire[1553]), .B(
        data_mem_out_wire[1585]), .S(N29), .Z(\Data_Mem/n7329 ) );
  MUX \Data_Mem/U7346  ( .A(data_mem_out_wire[1617]), .B(
        data_mem_out_wire[1649]), .S(N29), .Z(\Data_Mem/n7328 ) );
  MUX \Data_Mem/U7345  ( .A(\Data_Mem/n7326 ), .B(\Data_Mem/n7325 ), .S(N28), 
        .Z(\Data_Mem/n7327 ) );
  MUX \Data_Mem/U7344  ( .A(data_mem_out_wire[1681]), .B(
        data_mem_out_wire[1713]), .S(N29), .Z(\Data_Mem/n7326 ) );
  MUX \Data_Mem/U7343  ( .A(data_mem_out_wire[1745]), .B(
        data_mem_out_wire[1777]), .S(N29), .Z(\Data_Mem/n7325 ) );
  MUX \Data_Mem/U7342  ( .A(\Data_Mem/n7323 ), .B(\Data_Mem/n7320 ), .S(N27), 
        .Z(\Data_Mem/n7324 ) );
  MUX \Data_Mem/U7341  ( .A(\Data_Mem/n7322 ), .B(\Data_Mem/n7321 ), .S(N28), 
        .Z(\Data_Mem/n7323 ) );
  MUX \Data_Mem/U7340  ( .A(data_mem_out_wire[1809]), .B(
        data_mem_out_wire[1841]), .S(N29), .Z(\Data_Mem/n7322 ) );
  MUX \Data_Mem/U7339  ( .A(data_mem_out_wire[1873]), .B(
        data_mem_out_wire[1905]), .S(N29), .Z(\Data_Mem/n7321 ) );
  MUX \Data_Mem/U7338  ( .A(\Data_Mem/n7319 ), .B(\Data_Mem/n7318 ), .S(N28), 
        .Z(\Data_Mem/n7320 ) );
  MUX \Data_Mem/U7337  ( .A(data_mem_out_wire[1937]), .B(
        data_mem_out_wire[1969]), .S(N29), .Z(\Data_Mem/n7319 ) );
  MUX \Data_Mem/U7336  ( .A(data_mem_out_wire[2001]), .B(
        data_mem_out_wire[2033]), .S(N29), .Z(\Data_Mem/n7318 ) );
  MUX \Data_Mem/U7335  ( .A(\Data_Mem/n7317 ), .B(\Data_Mem/n7286 ), .S(N24), 
        .Z(c_memory[16]) );
  MUX \Data_Mem/U7334  ( .A(\Data_Mem/n7316 ), .B(\Data_Mem/n7301 ), .S(N25), 
        .Z(\Data_Mem/n7317 ) );
  MUX \Data_Mem/U7333  ( .A(\Data_Mem/n7315 ), .B(\Data_Mem/n7308 ), .S(N26), 
        .Z(\Data_Mem/n7316 ) );
  MUX \Data_Mem/U7332  ( .A(\Data_Mem/n7314 ), .B(\Data_Mem/n7311 ), .S(N27), 
        .Z(\Data_Mem/n7315 ) );
  MUX \Data_Mem/U7331  ( .A(\Data_Mem/n7313 ), .B(\Data_Mem/n7312 ), .S(N28), 
        .Z(\Data_Mem/n7314 ) );
  MUX \Data_Mem/U7330  ( .A(data_mem_out_wire[16]), .B(data_mem_out_wire[48]), 
        .S(N29), .Z(\Data_Mem/n7313 ) );
  MUX \Data_Mem/U7329  ( .A(data_mem_out_wire[80]), .B(data_mem_out_wire[112]), 
        .S(N29), .Z(\Data_Mem/n7312 ) );
  MUX \Data_Mem/U7328  ( .A(\Data_Mem/n7310 ), .B(\Data_Mem/n7309 ), .S(N28), 
        .Z(\Data_Mem/n7311 ) );
  MUX \Data_Mem/U7327  ( .A(data_mem_out_wire[144]), .B(data_mem_out_wire[176]), .S(N29), .Z(\Data_Mem/n7310 ) );
  MUX \Data_Mem/U7326  ( .A(data_mem_out_wire[208]), .B(data_mem_out_wire[240]), .S(N29), .Z(\Data_Mem/n7309 ) );
  MUX \Data_Mem/U7325  ( .A(\Data_Mem/n7307 ), .B(\Data_Mem/n7304 ), .S(N27), 
        .Z(\Data_Mem/n7308 ) );
  MUX \Data_Mem/U7324  ( .A(\Data_Mem/n7306 ), .B(\Data_Mem/n7305 ), .S(N28), 
        .Z(\Data_Mem/n7307 ) );
  MUX \Data_Mem/U7323  ( .A(data_mem_out_wire[272]), .B(data_mem_out_wire[304]), .S(N29), .Z(\Data_Mem/n7306 ) );
  MUX \Data_Mem/U7322  ( .A(data_mem_out_wire[336]), .B(data_mem_out_wire[368]), .S(N29), .Z(\Data_Mem/n7305 ) );
  MUX \Data_Mem/U7321  ( .A(\Data_Mem/n7303 ), .B(\Data_Mem/n7302 ), .S(N28), 
        .Z(\Data_Mem/n7304 ) );
  MUX \Data_Mem/U7320  ( .A(data_mem_out_wire[400]), .B(data_mem_out_wire[432]), .S(N29), .Z(\Data_Mem/n7303 ) );
  MUX \Data_Mem/U7319  ( .A(data_mem_out_wire[464]), .B(data_mem_out_wire[496]), .S(N29), .Z(\Data_Mem/n7302 ) );
  MUX \Data_Mem/U7318  ( .A(\Data_Mem/n7300 ), .B(\Data_Mem/n7293 ), .S(N26), 
        .Z(\Data_Mem/n7301 ) );
  MUX \Data_Mem/U7317  ( .A(\Data_Mem/n7299 ), .B(\Data_Mem/n7296 ), .S(N27), 
        .Z(\Data_Mem/n7300 ) );
  MUX \Data_Mem/U7316  ( .A(\Data_Mem/n7298 ), .B(\Data_Mem/n7297 ), .S(N28), 
        .Z(\Data_Mem/n7299 ) );
  MUX \Data_Mem/U7315  ( .A(data_mem_out_wire[528]), .B(data_mem_out_wire[560]), .S(N29), .Z(\Data_Mem/n7298 ) );
  MUX \Data_Mem/U7314  ( .A(data_mem_out_wire[592]), .B(data_mem_out_wire[624]), .S(N29), .Z(\Data_Mem/n7297 ) );
  MUX \Data_Mem/U7313  ( .A(\Data_Mem/n7295 ), .B(\Data_Mem/n7294 ), .S(N28), 
        .Z(\Data_Mem/n7296 ) );
  MUX \Data_Mem/U7312  ( .A(data_mem_out_wire[656]), .B(data_mem_out_wire[688]), .S(N29), .Z(\Data_Mem/n7295 ) );
  MUX \Data_Mem/U7311  ( .A(data_mem_out_wire[720]), .B(data_mem_out_wire[752]), .S(N29), .Z(\Data_Mem/n7294 ) );
  MUX \Data_Mem/U7310  ( .A(\Data_Mem/n7292 ), .B(\Data_Mem/n7289 ), .S(N27), 
        .Z(\Data_Mem/n7293 ) );
  MUX \Data_Mem/U7309  ( .A(\Data_Mem/n7291 ), .B(\Data_Mem/n7290 ), .S(N28), 
        .Z(\Data_Mem/n7292 ) );
  MUX \Data_Mem/U7308  ( .A(data_mem_out_wire[784]), .B(data_mem_out_wire[816]), .S(N29), .Z(\Data_Mem/n7291 ) );
  MUX \Data_Mem/U7307  ( .A(data_mem_out_wire[848]), .B(data_mem_out_wire[880]), .S(N29), .Z(\Data_Mem/n7290 ) );
  MUX \Data_Mem/U7306  ( .A(\Data_Mem/n7288 ), .B(\Data_Mem/n7287 ), .S(N28), 
        .Z(\Data_Mem/n7289 ) );
  MUX \Data_Mem/U7305  ( .A(data_mem_out_wire[912]), .B(data_mem_out_wire[944]), .S(N29), .Z(\Data_Mem/n7288 ) );
  MUX \Data_Mem/U7304  ( .A(data_mem_out_wire[976]), .B(
        data_mem_out_wire[1008]), .S(N29), .Z(\Data_Mem/n7287 ) );
  MUX \Data_Mem/U7303  ( .A(\Data_Mem/n7285 ), .B(\Data_Mem/n7270 ), .S(N25), 
        .Z(\Data_Mem/n7286 ) );
  MUX \Data_Mem/U7302  ( .A(\Data_Mem/n7284 ), .B(\Data_Mem/n7277 ), .S(N26), 
        .Z(\Data_Mem/n7285 ) );
  MUX \Data_Mem/U7301  ( .A(\Data_Mem/n7283 ), .B(\Data_Mem/n7280 ), .S(N27), 
        .Z(\Data_Mem/n7284 ) );
  MUX \Data_Mem/U7300  ( .A(\Data_Mem/n7282 ), .B(\Data_Mem/n7281 ), .S(N28), 
        .Z(\Data_Mem/n7283 ) );
  MUX \Data_Mem/U7299  ( .A(data_mem_out_wire[1040]), .B(
        data_mem_out_wire[1072]), .S(N29), .Z(\Data_Mem/n7282 ) );
  MUX \Data_Mem/U7298  ( .A(data_mem_out_wire[1104]), .B(
        data_mem_out_wire[1136]), .S(N29), .Z(\Data_Mem/n7281 ) );
  MUX \Data_Mem/U7297  ( .A(\Data_Mem/n7279 ), .B(\Data_Mem/n7278 ), .S(N28), 
        .Z(\Data_Mem/n7280 ) );
  MUX \Data_Mem/U7296  ( .A(data_mem_out_wire[1168]), .B(
        data_mem_out_wire[1200]), .S(N29), .Z(\Data_Mem/n7279 ) );
  MUX \Data_Mem/U7295  ( .A(data_mem_out_wire[1232]), .B(
        data_mem_out_wire[1264]), .S(N29), .Z(\Data_Mem/n7278 ) );
  MUX \Data_Mem/U7294  ( .A(\Data_Mem/n7276 ), .B(\Data_Mem/n7273 ), .S(N27), 
        .Z(\Data_Mem/n7277 ) );
  MUX \Data_Mem/U7293  ( .A(\Data_Mem/n7275 ), .B(\Data_Mem/n7274 ), .S(N28), 
        .Z(\Data_Mem/n7276 ) );
  MUX \Data_Mem/U7292  ( .A(data_mem_out_wire[1296]), .B(
        data_mem_out_wire[1328]), .S(N29), .Z(\Data_Mem/n7275 ) );
  MUX \Data_Mem/U7291  ( .A(data_mem_out_wire[1360]), .B(
        data_mem_out_wire[1392]), .S(N29), .Z(\Data_Mem/n7274 ) );
  MUX \Data_Mem/U7290  ( .A(\Data_Mem/n7272 ), .B(\Data_Mem/n7271 ), .S(N28), 
        .Z(\Data_Mem/n7273 ) );
  MUX \Data_Mem/U7289  ( .A(data_mem_out_wire[1424]), .B(
        data_mem_out_wire[1456]), .S(N29), .Z(\Data_Mem/n7272 ) );
  MUX \Data_Mem/U7288  ( .A(data_mem_out_wire[1488]), .B(
        data_mem_out_wire[1520]), .S(N29), .Z(\Data_Mem/n7271 ) );
  MUX \Data_Mem/U7287  ( .A(\Data_Mem/n7269 ), .B(\Data_Mem/n7262 ), .S(N26), 
        .Z(\Data_Mem/n7270 ) );
  MUX \Data_Mem/U7286  ( .A(\Data_Mem/n7268 ), .B(\Data_Mem/n7265 ), .S(N27), 
        .Z(\Data_Mem/n7269 ) );
  MUX \Data_Mem/U7285  ( .A(\Data_Mem/n7267 ), .B(\Data_Mem/n7266 ), .S(N28), 
        .Z(\Data_Mem/n7268 ) );
  MUX \Data_Mem/U7284  ( .A(data_mem_out_wire[1552]), .B(
        data_mem_out_wire[1584]), .S(N29), .Z(\Data_Mem/n7267 ) );
  MUX \Data_Mem/U7283  ( .A(data_mem_out_wire[1616]), .B(
        data_mem_out_wire[1648]), .S(N29), .Z(\Data_Mem/n7266 ) );
  MUX \Data_Mem/U7282  ( .A(\Data_Mem/n7264 ), .B(\Data_Mem/n7263 ), .S(N28), 
        .Z(\Data_Mem/n7265 ) );
  MUX \Data_Mem/U7281  ( .A(data_mem_out_wire[1680]), .B(
        data_mem_out_wire[1712]), .S(N29), .Z(\Data_Mem/n7264 ) );
  MUX \Data_Mem/U7280  ( .A(data_mem_out_wire[1744]), .B(
        data_mem_out_wire[1776]), .S(N29), .Z(\Data_Mem/n7263 ) );
  MUX \Data_Mem/U7279  ( .A(\Data_Mem/n7261 ), .B(\Data_Mem/n7258 ), .S(N27), 
        .Z(\Data_Mem/n7262 ) );
  MUX \Data_Mem/U7278  ( .A(\Data_Mem/n7260 ), .B(\Data_Mem/n7259 ), .S(N28), 
        .Z(\Data_Mem/n7261 ) );
  MUX \Data_Mem/U7277  ( .A(data_mem_out_wire[1808]), .B(
        data_mem_out_wire[1840]), .S(N29), .Z(\Data_Mem/n7260 ) );
  MUX \Data_Mem/U7276  ( .A(data_mem_out_wire[1872]), .B(
        data_mem_out_wire[1904]), .S(N29), .Z(\Data_Mem/n7259 ) );
  MUX \Data_Mem/U7275  ( .A(\Data_Mem/n7257 ), .B(\Data_Mem/n7256 ), .S(N28), 
        .Z(\Data_Mem/n7258 ) );
  MUX \Data_Mem/U7274  ( .A(data_mem_out_wire[1936]), .B(
        data_mem_out_wire[1968]), .S(N29), .Z(\Data_Mem/n7257 ) );
  MUX \Data_Mem/U7273  ( .A(data_mem_out_wire[2000]), .B(
        data_mem_out_wire[2032]), .S(N29), .Z(\Data_Mem/n7256 ) );
  MUX \Data_Mem/U7272  ( .A(\Data_Mem/n7255 ), .B(\Data_Mem/n7224 ), .S(N24), 
        .Z(c_memory[15]) );
  MUX \Data_Mem/U7271  ( .A(\Data_Mem/n7254 ), .B(\Data_Mem/n7239 ), .S(N25), 
        .Z(\Data_Mem/n7255 ) );
  MUX \Data_Mem/U7270  ( .A(\Data_Mem/n7253 ), .B(\Data_Mem/n7246 ), .S(N26), 
        .Z(\Data_Mem/n7254 ) );
  MUX \Data_Mem/U7269  ( .A(\Data_Mem/n7252 ), .B(\Data_Mem/n7249 ), .S(N27), 
        .Z(\Data_Mem/n7253 ) );
  MUX \Data_Mem/U7268  ( .A(\Data_Mem/n7251 ), .B(\Data_Mem/n7250 ), .S(N28), 
        .Z(\Data_Mem/n7252 ) );
  MUX \Data_Mem/U7267  ( .A(data_mem_out_wire[15]), .B(data_mem_out_wire[47]), 
        .S(N29), .Z(\Data_Mem/n7251 ) );
  MUX \Data_Mem/U7266  ( .A(data_mem_out_wire[79]), .B(data_mem_out_wire[111]), 
        .S(N29), .Z(\Data_Mem/n7250 ) );
  MUX \Data_Mem/U7265  ( .A(\Data_Mem/n7248 ), .B(\Data_Mem/n7247 ), .S(N28), 
        .Z(\Data_Mem/n7249 ) );
  MUX \Data_Mem/U7264  ( .A(data_mem_out_wire[143]), .B(data_mem_out_wire[175]), .S(N29), .Z(\Data_Mem/n7248 ) );
  MUX \Data_Mem/U7263  ( .A(data_mem_out_wire[207]), .B(data_mem_out_wire[239]), .S(N29), .Z(\Data_Mem/n7247 ) );
  MUX \Data_Mem/U7262  ( .A(\Data_Mem/n7245 ), .B(\Data_Mem/n7242 ), .S(N27), 
        .Z(\Data_Mem/n7246 ) );
  MUX \Data_Mem/U7261  ( .A(\Data_Mem/n7244 ), .B(\Data_Mem/n7243 ), .S(N28), 
        .Z(\Data_Mem/n7245 ) );
  MUX \Data_Mem/U7260  ( .A(data_mem_out_wire[271]), .B(data_mem_out_wire[303]), .S(N29), .Z(\Data_Mem/n7244 ) );
  MUX \Data_Mem/U7259  ( .A(data_mem_out_wire[335]), .B(data_mem_out_wire[367]), .S(N29), .Z(\Data_Mem/n7243 ) );
  MUX \Data_Mem/U7258  ( .A(\Data_Mem/n7241 ), .B(\Data_Mem/n7240 ), .S(N28), 
        .Z(\Data_Mem/n7242 ) );
  MUX \Data_Mem/U7257  ( .A(data_mem_out_wire[399]), .B(data_mem_out_wire[431]), .S(N29), .Z(\Data_Mem/n7241 ) );
  MUX \Data_Mem/U7256  ( .A(data_mem_out_wire[463]), .B(data_mem_out_wire[495]), .S(N29), .Z(\Data_Mem/n7240 ) );
  MUX \Data_Mem/U7255  ( .A(\Data_Mem/n7238 ), .B(\Data_Mem/n7231 ), .S(N26), 
        .Z(\Data_Mem/n7239 ) );
  MUX \Data_Mem/U7254  ( .A(\Data_Mem/n7237 ), .B(\Data_Mem/n7234 ), .S(N27), 
        .Z(\Data_Mem/n7238 ) );
  MUX \Data_Mem/U7253  ( .A(\Data_Mem/n7236 ), .B(\Data_Mem/n7235 ), .S(N28), 
        .Z(\Data_Mem/n7237 ) );
  MUX \Data_Mem/U7252  ( .A(data_mem_out_wire[527]), .B(data_mem_out_wire[559]), .S(N29), .Z(\Data_Mem/n7236 ) );
  MUX \Data_Mem/U7251  ( .A(data_mem_out_wire[591]), .B(data_mem_out_wire[623]), .S(N29), .Z(\Data_Mem/n7235 ) );
  MUX \Data_Mem/U7250  ( .A(\Data_Mem/n7233 ), .B(\Data_Mem/n7232 ), .S(N28), 
        .Z(\Data_Mem/n7234 ) );
  MUX \Data_Mem/U7249  ( .A(data_mem_out_wire[655]), .B(data_mem_out_wire[687]), .S(N29), .Z(\Data_Mem/n7233 ) );
  MUX \Data_Mem/U7248  ( .A(data_mem_out_wire[719]), .B(data_mem_out_wire[751]), .S(N29), .Z(\Data_Mem/n7232 ) );
  MUX \Data_Mem/U7247  ( .A(\Data_Mem/n7230 ), .B(\Data_Mem/n7227 ), .S(N27), 
        .Z(\Data_Mem/n7231 ) );
  MUX \Data_Mem/U7246  ( .A(\Data_Mem/n7229 ), .B(\Data_Mem/n7228 ), .S(N28), 
        .Z(\Data_Mem/n7230 ) );
  MUX \Data_Mem/U7245  ( .A(data_mem_out_wire[783]), .B(data_mem_out_wire[815]), .S(N29), .Z(\Data_Mem/n7229 ) );
  MUX \Data_Mem/U7244  ( .A(data_mem_out_wire[847]), .B(data_mem_out_wire[879]), .S(N29), .Z(\Data_Mem/n7228 ) );
  MUX \Data_Mem/U7243  ( .A(\Data_Mem/n7226 ), .B(\Data_Mem/n7225 ), .S(N28), 
        .Z(\Data_Mem/n7227 ) );
  MUX \Data_Mem/U7242  ( .A(data_mem_out_wire[911]), .B(data_mem_out_wire[943]), .S(N29), .Z(\Data_Mem/n7226 ) );
  MUX \Data_Mem/U7241  ( .A(data_mem_out_wire[975]), .B(
        data_mem_out_wire[1007]), .S(N29), .Z(\Data_Mem/n7225 ) );
  MUX \Data_Mem/U7240  ( .A(\Data_Mem/n7223 ), .B(\Data_Mem/n7208 ), .S(N25), 
        .Z(\Data_Mem/n7224 ) );
  MUX \Data_Mem/U7239  ( .A(\Data_Mem/n7222 ), .B(\Data_Mem/n7215 ), .S(N26), 
        .Z(\Data_Mem/n7223 ) );
  MUX \Data_Mem/U7238  ( .A(\Data_Mem/n7221 ), .B(\Data_Mem/n7218 ), .S(N27), 
        .Z(\Data_Mem/n7222 ) );
  MUX \Data_Mem/U7237  ( .A(\Data_Mem/n7220 ), .B(\Data_Mem/n7219 ), .S(N28), 
        .Z(\Data_Mem/n7221 ) );
  MUX \Data_Mem/U7236  ( .A(data_mem_out_wire[1039]), .B(
        data_mem_out_wire[1071]), .S(N29), .Z(\Data_Mem/n7220 ) );
  MUX \Data_Mem/U7235  ( .A(data_mem_out_wire[1103]), .B(
        data_mem_out_wire[1135]), .S(N29), .Z(\Data_Mem/n7219 ) );
  MUX \Data_Mem/U7234  ( .A(\Data_Mem/n7217 ), .B(\Data_Mem/n7216 ), .S(N28), 
        .Z(\Data_Mem/n7218 ) );
  MUX \Data_Mem/U7233  ( .A(data_mem_out_wire[1167]), .B(
        data_mem_out_wire[1199]), .S(N29), .Z(\Data_Mem/n7217 ) );
  MUX \Data_Mem/U7232  ( .A(data_mem_out_wire[1231]), .B(
        data_mem_out_wire[1263]), .S(N29), .Z(\Data_Mem/n7216 ) );
  MUX \Data_Mem/U7231  ( .A(\Data_Mem/n7214 ), .B(\Data_Mem/n7211 ), .S(N27), 
        .Z(\Data_Mem/n7215 ) );
  MUX \Data_Mem/U7230  ( .A(\Data_Mem/n7213 ), .B(\Data_Mem/n7212 ), .S(N28), 
        .Z(\Data_Mem/n7214 ) );
  MUX \Data_Mem/U7229  ( .A(data_mem_out_wire[1295]), .B(
        data_mem_out_wire[1327]), .S(N29), .Z(\Data_Mem/n7213 ) );
  MUX \Data_Mem/U7228  ( .A(data_mem_out_wire[1359]), .B(
        data_mem_out_wire[1391]), .S(N29), .Z(\Data_Mem/n7212 ) );
  MUX \Data_Mem/U7227  ( .A(\Data_Mem/n7210 ), .B(\Data_Mem/n7209 ), .S(N28), 
        .Z(\Data_Mem/n7211 ) );
  MUX \Data_Mem/U7226  ( .A(data_mem_out_wire[1423]), .B(
        data_mem_out_wire[1455]), .S(N29), .Z(\Data_Mem/n7210 ) );
  MUX \Data_Mem/U7225  ( .A(data_mem_out_wire[1487]), .B(
        data_mem_out_wire[1519]), .S(N29), .Z(\Data_Mem/n7209 ) );
  MUX \Data_Mem/U7224  ( .A(\Data_Mem/n7207 ), .B(\Data_Mem/n7200 ), .S(N26), 
        .Z(\Data_Mem/n7208 ) );
  MUX \Data_Mem/U7223  ( .A(\Data_Mem/n7206 ), .B(\Data_Mem/n7203 ), .S(N27), 
        .Z(\Data_Mem/n7207 ) );
  MUX \Data_Mem/U7222  ( .A(\Data_Mem/n7205 ), .B(\Data_Mem/n7204 ), .S(N28), 
        .Z(\Data_Mem/n7206 ) );
  MUX \Data_Mem/U7221  ( .A(data_mem_out_wire[1551]), .B(
        data_mem_out_wire[1583]), .S(N29), .Z(\Data_Mem/n7205 ) );
  MUX \Data_Mem/U7220  ( .A(data_mem_out_wire[1615]), .B(
        data_mem_out_wire[1647]), .S(N29), .Z(\Data_Mem/n7204 ) );
  MUX \Data_Mem/U7219  ( .A(\Data_Mem/n7202 ), .B(\Data_Mem/n7201 ), .S(N28), 
        .Z(\Data_Mem/n7203 ) );
  MUX \Data_Mem/U7218  ( .A(data_mem_out_wire[1679]), .B(
        data_mem_out_wire[1711]), .S(N29), .Z(\Data_Mem/n7202 ) );
  MUX \Data_Mem/U7217  ( .A(data_mem_out_wire[1743]), .B(
        data_mem_out_wire[1775]), .S(N29), .Z(\Data_Mem/n7201 ) );
  MUX \Data_Mem/U7216  ( .A(\Data_Mem/n7199 ), .B(\Data_Mem/n7196 ), .S(N27), 
        .Z(\Data_Mem/n7200 ) );
  MUX \Data_Mem/U7215  ( .A(\Data_Mem/n7198 ), .B(\Data_Mem/n7197 ), .S(N28), 
        .Z(\Data_Mem/n7199 ) );
  MUX \Data_Mem/U7214  ( .A(data_mem_out_wire[1807]), .B(
        data_mem_out_wire[1839]), .S(N29), .Z(\Data_Mem/n7198 ) );
  MUX \Data_Mem/U7213  ( .A(data_mem_out_wire[1871]), .B(
        data_mem_out_wire[1903]), .S(N29), .Z(\Data_Mem/n7197 ) );
  MUX \Data_Mem/U7212  ( .A(\Data_Mem/n7195 ), .B(\Data_Mem/n7194 ), .S(N28), 
        .Z(\Data_Mem/n7196 ) );
  MUX \Data_Mem/U7211  ( .A(data_mem_out_wire[1935]), .B(
        data_mem_out_wire[1967]), .S(N29), .Z(\Data_Mem/n7195 ) );
  MUX \Data_Mem/U7210  ( .A(data_mem_out_wire[1999]), .B(
        data_mem_out_wire[2031]), .S(N29), .Z(\Data_Mem/n7194 ) );
  MUX \Data_Mem/U7209  ( .A(\Data_Mem/n7193 ), .B(\Data_Mem/n7162 ), .S(N24), 
        .Z(c_memory[14]) );
  MUX \Data_Mem/U7208  ( .A(\Data_Mem/n7192 ), .B(\Data_Mem/n7177 ), .S(N25), 
        .Z(\Data_Mem/n7193 ) );
  MUX \Data_Mem/U7207  ( .A(\Data_Mem/n7191 ), .B(\Data_Mem/n7184 ), .S(N26), 
        .Z(\Data_Mem/n7192 ) );
  MUX \Data_Mem/U7206  ( .A(\Data_Mem/n7190 ), .B(\Data_Mem/n7187 ), .S(N27), 
        .Z(\Data_Mem/n7191 ) );
  MUX \Data_Mem/U7205  ( .A(\Data_Mem/n7189 ), .B(\Data_Mem/n7188 ), .S(N28), 
        .Z(\Data_Mem/n7190 ) );
  MUX \Data_Mem/U7204  ( .A(data_mem_out_wire[14]), .B(data_mem_out_wire[46]), 
        .S(N29), .Z(\Data_Mem/n7189 ) );
  MUX \Data_Mem/U7203  ( .A(data_mem_out_wire[78]), .B(data_mem_out_wire[110]), 
        .S(N29), .Z(\Data_Mem/n7188 ) );
  MUX \Data_Mem/U7202  ( .A(\Data_Mem/n7186 ), .B(\Data_Mem/n7185 ), .S(N28), 
        .Z(\Data_Mem/n7187 ) );
  MUX \Data_Mem/U7201  ( .A(data_mem_out_wire[142]), .B(data_mem_out_wire[174]), .S(N29), .Z(\Data_Mem/n7186 ) );
  MUX \Data_Mem/U7200  ( .A(data_mem_out_wire[206]), .B(data_mem_out_wire[238]), .S(N29), .Z(\Data_Mem/n7185 ) );
  MUX \Data_Mem/U7199  ( .A(\Data_Mem/n7183 ), .B(\Data_Mem/n7180 ), .S(N27), 
        .Z(\Data_Mem/n7184 ) );
  MUX \Data_Mem/U7198  ( .A(\Data_Mem/n7182 ), .B(\Data_Mem/n7181 ), .S(N28), 
        .Z(\Data_Mem/n7183 ) );
  MUX \Data_Mem/U7197  ( .A(data_mem_out_wire[270]), .B(data_mem_out_wire[302]), .S(N29), .Z(\Data_Mem/n7182 ) );
  MUX \Data_Mem/U7196  ( .A(data_mem_out_wire[334]), .B(data_mem_out_wire[366]), .S(N29), .Z(\Data_Mem/n7181 ) );
  MUX \Data_Mem/U7195  ( .A(\Data_Mem/n7179 ), .B(\Data_Mem/n7178 ), .S(N28), 
        .Z(\Data_Mem/n7180 ) );
  MUX \Data_Mem/U7194  ( .A(data_mem_out_wire[398]), .B(data_mem_out_wire[430]), .S(N29), .Z(\Data_Mem/n7179 ) );
  MUX \Data_Mem/U7193  ( .A(data_mem_out_wire[462]), .B(data_mem_out_wire[494]), .S(N29), .Z(\Data_Mem/n7178 ) );
  MUX \Data_Mem/U7192  ( .A(\Data_Mem/n7176 ), .B(\Data_Mem/n7169 ), .S(N26), 
        .Z(\Data_Mem/n7177 ) );
  MUX \Data_Mem/U7191  ( .A(\Data_Mem/n7175 ), .B(\Data_Mem/n7172 ), .S(N27), 
        .Z(\Data_Mem/n7176 ) );
  MUX \Data_Mem/U7190  ( .A(\Data_Mem/n7174 ), .B(\Data_Mem/n7173 ), .S(N28), 
        .Z(\Data_Mem/n7175 ) );
  MUX \Data_Mem/U7189  ( .A(data_mem_out_wire[526]), .B(data_mem_out_wire[558]), .S(N29), .Z(\Data_Mem/n7174 ) );
  MUX \Data_Mem/U7188  ( .A(data_mem_out_wire[590]), .B(data_mem_out_wire[622]), .S(N29), .Z(\Data_Mem/n7173 ) );
  MUX \Data_Mem/U7187  ( .A(\Data_Mem/n7171 ), .B(\Data_Mem/n7170 ), .S(N28), 
        .Z(\Data_Mem/n7172 ) );
  MUX \Data_Mem/U7186  ( .A(data_mem_out_wire[654]), .B(data_mem_out_wire[686]), .S(N29), .Z(\Data_Mem/n7171 ) );
  MUX \Data_Mem/U7185  ( .A(data_mem_out_wire[718]), .B(data_mem_out_wire[750]), .S(N29), .Z(\Data_Mem/n7170 ) );
  MUX \Data_Mem/U7184  ( .A(\Data_Mem/n7168 ), .B(\Data_Mem/n7165 ), .S(N27), 
        .Z(\Data_Mem/n7169 ) );
  MUX \Data_Mem/U7183  ( .A(\Data_Mem/n7167 ), .B(\Data_Mem/n7166 ), .S(N28), 
        .Z(\Data_Mem/n7168 ) );
  MUX \Data_Mem/U7182  ( .A(data_mem_out_wire[782]), .B(data_mem_out_wire[814]), .S(N29), .Z(\Data_Mem/n7167 ) );
  MUX \Data_Mem/U7181  ( .A(data_mem_out_wire[846]), .B(data_mem_out_wire[878]), .S(N29), .Z(\Data_Mem/n7166 ) );
  MUX \Data_Mem/U7180  ( .A(\Data_Mem/n7164 ), .B(\Data_Mem/n7163 ), .S(N28), 
        .Z(\Data_Mem/n7165 ) );
  MUX \Data_Mem/U7179  ( .A(data_mem_out_wire[910]), .B(data_mem_out_wire[942]), .S(N29), .Z(\Data_Mem/n7164 ) );
  MUX \Data_Mem/U7178  ( .A(data_mem_out_wire[974]), .B(
        data_mem_out_wire[1006]), .S(N29), .Z(\Data_Mem/n7163 ) );
  MUX \Data_Mem/U7177  ( .A(\Data_Mem/n7161 ), .B(\Data_Mem/n7146 ), .S(N25), 
        .Z(\Data_Mem/n7162 ) );
  MUX \Data_Mem/U7176  ( .A(\Data_Mem/n7160 ), .B(\Data_Mem/n7153 ), .S(N26), 
        .Z(\Data_Mem/n7161 ) );
  MUX \Data_Mem/U7175  ( .A(\Data_Mem/n7159 ), .B(\Data_Mem/n7156 ), .S(N27), 
        .Z(\Data_Mem/n7160 ) );
  MUX \Data_Mem/U7174  ( .A(\Data_Mem/n7158 ), .B(\Data_Mem/n7157 ), .S(N28), 
        .Z(\Data_Mem/n7159 ) );
  MUX \Data_Mem/U7173  ( .A(data_mem_out_wire[1038]), .B(
        data_mem_out_wire[1070]), .S(N29), .Z(\Data_Mem/n7158 ) );
  MUX \Data_Mem/U7172  ( .A(data_mem_out_wire[1102]), .B(
        data_mem_out_wire[1134]), .S(N29), .Z(\Data_Mem/n7157 ) );
  MUX \Data_Mem/U7171  ( .A(\Data_Mem/n7155 ), .B(\Data_Mem/n7154 ), .S(N28), 
        .Z(\Data_Mem/n7156 ) );
  MUX \Data_Mem/U7170  ( .A(data_mem_out_wire[1166]), .B(
        data_mem_out_wire[1198]), .S(N29), .Z(\Data_Mem/n7155 ) );
  MUX \Data_Mem/U7169  ( .A(data_mem_out_wire[1230]), .B(
        data_mem_out_wire[1262]), .S(N29), .Z(\Data_Mem/n7154 ) );
  MUX \Data_Mem/U7168  ( .A(\Data_Mem/n7152 ), .B(\Data_Mem/n7149 ), .S(N27), 
        .Z(\Data_Mem/n7153 ) );
  MUX \Data_Mem/U7167  ( .A(\Data_Mem/n7151 ), .B(\Data_Mem/n7150 ), .S(N28), 
        .Z(\Data_Mem/n7152 ) );
  MUX \Data_Mem/U7166  ( .A(data_mem_out_wire[1294]), .B(
        data_mem_out_wire[1326]), .S(N29), .Z(\Data_Mem/n7151 ) );
  MUX \Data_Mem/U7165  ( .A(data_mem_out_wire[1358]), .B(
        data_mem_out_wire[1390]), .S(N29), .Z(\Data_Mem/n7150 ) );
  MUX \Data_Mem/U7164  ( .A(\Data_Mem/n7148 ), .B(\Data_Mem/n7147 ), .S(N28), 
        .Z(\Data_Mem/n7149 ) );
  MUX \Data_Mem/U7163  ( .A(data_mem_out_wire[1422]), .B(
        data_mem_out_wire[1454]), .S(N29), .Z(\Data_Mem/n7148 ) );
  MUX \Data_Mem/U7162  ( .A(data_mem_out_wire[1486]), .B(
        data_mem_out_wire[1518]), .S(N29), .Z(\Data_Mem/n7147 ) );
  MUX \Data_Mem/U7161  ( .A(\Data_Mem/n7145 ), .B(\Data_Mem/n7138 ), .S(N26), 
        .Z(\Data_Mem/n7146 ) );
  MUX \Data_Mem/U7160  ( .A(\Data_Mem/n7144 ), .B(\Data_Mem/n7141 ), .S(N27), 
        .Z(\Data_Mem/n7145 ) );
  MUX \Data_Mem/U7159  ( .A(\Data_Mem/n7143 ), .B(\Data_Mem/n7142 ), .S(N28), 
        .Z(\Data_Mem/n7144 ) );
  MUX \Data_Mem/U7158  ( .A(data_mem_out_wire[1550]), .B(
        data_mem_out_wire[1582]), .S(N29), .Z(\Data_Mem/n7143 ) );
  MUX \Data_Mem/U7157  ( .A(data_mem_out_wire[1614]), .B(
        data_mem_out_wire[1646]), .S(N29), .Z(\Data_Mem/n7142 ) );
  MUX \Data_Mem/U7156  ( .A(\Data_Mem/n7140 ), .B(\Data_Mem/n7139 ), .S(N28), 
        .Z(\Data_Mem/n7141 ) );
  MUX \Data_Mem/U7155  ( .A(data_mem_out_wire[1678]), .B(
        data_mem_out_wire[1710]), .S(N29), .Z(\Data_Mem/n7140 ) );
  MUX \Data_Mem/U7154  ( .A(data_mem_out_wire[1742]), .B(
        data_mem_out_wire[1774]), .S(N29), .Z(\Data_Mem/n7139 ) );
  MUX \Data_Mem/U7153  ( .A(\Data_Mem/n7137 ), .B(\Data_Mem/n7134 ), .S(N27), 
        .Z(\Data_Mem/n7138 ) );
  MUX \Data_Mem/U7152  ( .A(\Data_Mem/n7136 ), .B(\Data_Mem/n7135 ), .S(N28), 
        .Z(\Data_Mem/n7137 ) );
  MUX \Data_Mem/U7151  ( .A(data_mem_out_wire[1806]), .B(
        data_mem_out_wire[1838]), .S(N29), .Z(\Data_Mem/n7136 ) );
  MUX \Data_Mem/U7150  ( .A(data_mem_out_wire[1870]), .B(
        data_mem_out_wire[1902]), .S(N29), .Z(\Data_Mem/n7135 ) );
  MUX \Data_Mem/U7149  ( .A(\Data_Mem/n7133 ), .B(\Data_Mem/n7132 ), .S(N28), 
        .Z(\Data_Mem/n7134 ) );
  MUX \Data_Mem/U7148  ( .A(data_mem_out_wire[1934]), .B(
        data_mem_out_wire[1966]), .S(N29), .Z(\Data_Mem/n7133 ) );
  MUX \Data_Mem/U7147  ( .A(data_mem_out_wire[1998]), .B(
        data_mem_out_wire[2030]), .S(N29), .Z(\Data_Mem/n7132 ) );
  MUX \Data_Mem/U7146  ( .A(\Data_Mem/n7131 ), .B(\Data_Mem/n7100 ), .S(N24), 
        .Z(c_memory[13]) );
  MUX \Data_Mem/U7145  ( .A(\Data_Mem/n7130 ), .B(\Data_Mem/n7115 ), .S(N25), 
        .Z(\Data_Mem/n7131 ) );
  MUX \Data_Mem/U7144  ( .A(\Data_Mem/n7129 ), .B(\Data_Mem/n7122 ), .S(N26), 
        .Z(\Data_Mem/n7130 ) );
  MUX \Data_Mem/U7143  ( .A(\Data_Mem/n7128 ), .B(\Data_Mem/n7125 ), .S(N27), 
        .Z(\Data_Mem/n7129 ) );
  MUX \Data_Mem/U7142  ( .A(\Data_Mem/n7127 ), .B(\Data_Mem/n7126 ), .S(N28), 
        .Z(\Data_Mem/n7128 ) );
  MUX \Data_Mem/U7141  ( .A(data_mem_out_wire[13]), .B(data_mem_out_wire[45]), 
        .S(N29), .Z(\Data_Mem/n7127 ) );
  MUX \Data_Mem/U7140  ( .A(data_mem_out_wire[77]), .B(data_mem_out_wire[109]), 
        .S(N29), .Z(\Data_Mem/n7126 ) );
  MUX \Data_Mem/U7139  ( .A(\Data_Mem/n7124 ), .B(\Data_Mem/n7123 ), .S(N28), 
        .Z(\Data_Mem/n7125 ) );
  MUX \Data_Mem/U7138  ( .A(data_mem_out_wire[141]), .B(data_mem_out_wire[173]), .S(N29), .Z(\Data_Mem/n7124 ) );
  MUX \Data_Mem/U7137  ( .A(data_mem_out_wire[205]), .B(data_mem_out_wire[237]), .S(N29), .Z(\Data_Mem/n7123 ) );
  MUX \Data_Mem/U7136  ( .A(\Data_Mem/n7121 ), .B(\Data_Mem/n7118 ), .S(N27), 
        .Z(\Data_Mem/n7122 ) );
  MUX \Data_Mem/U7135  ( .A(\Data_Mem/n7120 ), .B(\Data_Mem/n7119 ), .S(N28), 
        .Z(\Data_Mem/n7121 ) );
  MUX \Data_Mem/U7134  ( .A(data_mem_out_wire[269]), .B(data_mem_out_wire[301]), .S(N29), .Z(\Data_Mem/n7120 ) );
  MUX \Data_Mem/U7133  ( .A(data_mem_out_wire[333]), .B(data_mem_out_wire[365]), .S(N29), .Z(\Data_Mem/n7119 ) );
  MUX \Data_Mem/U7132  ( .A(\Data_Mem/n7117 ), .B(\Data_Mem/n7116 ), .S(N28), 
        .Z(\Data_Mem/n7118 ) );
  MUX \Data_Mem/U7131  ( .A(data_mem_out_wire[397]), .B(data_mem_out_wire[429]), .S(N29), .Z(\Data_Mem/n7117 ) );
  MUX \Data_Mem/U7130  ( .A(data_mem_out_wire[461]), .B(data_mem_out_wire[493]), .S(N29), .Z(\Data_Mem/n7116 ) );
  MUX \Data_Mem/U7129  ( .A(\Data_Mem/n7114 ), .B(\Data_Mem/n7107 ), .S(N26), 
        .Z(\Data_Mem/n7115 ) );
  MUX \Data_Mem/U7128  ( .A(\Data_Mem/n7113 ), .B(\Data_Mem/n7110 ), .S(N27), 
        .Z(\Data_Mem/n7114 ) );
  MUX \Data_Mem/U7127  ( .A(\Data_Mem/n7112 ), .B(\Data_Mem/n7111 ), .S(N28), 
        .Z(\Data_Mem/n7113 ) );
  MUX \Data_Mem/U7126  ( .A(data_mem_out_wire[525]), .B(data_mem_out_wire[557]), .S(N29), .Z(\Data_Mem/n7112 ) );
  MUX \Data_Mem/U7125  ( .A(data_mem_out_wire[589]), .B(data_mem_out_wire[621]), .S(N29), .Z(\Data_Mem/n7111 ) );
  MUX \Data_Mem/U7124  ( .A(\Data_Mem/n7109 ), .B(\Data_Mem/n7108 ), .S(N28), 
        .Z(\Data_Mem/n7110 ) );
  MUX \Data_Mem/U7123  ( .A(data_mem_out_wire[653]), .B(data_mem_out_wire[685]), .S(N29), .Z(\Data_Mem/n7109 ) );
  MUX \Data_Mem/U7122  ( .A(data_mem_out_wire[717]), .B(data_mem_out_wire[749]), .S(N29), .Z(\Data_Mem/n7108 ) );
  MUX \Data_Mem/U7121  ( .A(\Data_Mem/n7106 ), .B(\Data_Mem/n7103 ), .S(N27), 
        .Z(\Data_Mem/n7107 ) );
  MUX \Data_Mem/U7120  ( .A(\Data_Mem/n7105 ), .B(\Data_Mem/n7104 ), .S(N28), 
        .Z(\Data_Mem/n7106 ) );
  MUX \Data_Mem/U7119  ( .A(data_mem_out_wire[781]), .B(data_mem_out_wire[813]), .S(N29), .Z(\Data_Mem/n7105 ) );
  MUX \Data_Mem/U7118  ( .A(data_mem_out_wire[845]), .B(data_mem_out_wire[877]), .S(N29), .Z(\Data_Mem/n7104 ) );
  MUX \Data_Mem/U7117  ( .A(\Data_Mem/n7102 ), .B(\Data_Mem/n7101 ), .S(N28), 
        .Z(\Data_Mem/n7103 ) );
  MUX \Data_Mem/U7116  ( .A(data_mem_out_wire[909]), .B(data_mem_out_wire[941]), .S(N29), .Z(\Data_Mem/n7102 ) );
  MUX \Data_Mem/U7115  ( .A(data_mem_out_wire[973]), .B(
        data_mem_out_wire[1005]), .S(N29), .Z(\Data_Mem/n7101 ) );
  MUX \Data_Mem/U7114  ( .A(\Data_Mem/n7099 ), .B(\Data_Mem/n7084 ), .S(N25), 
        .Z(\Data_Mem/n7100 ) );
  MUX \Data_Mem/U7113  ( .A(\Data_Mem/n7098 ), .B(\Data_Mem/n7091 ), .S(N26), 
        .Z(\Data_Mem/n7099 ) );
  MUX \Data_Mem/U7112  ( .A(\Data_Mem/n7097 ), .B(\Data_Mem/n7094 ), .S(N27), 
        .Z(\Data_Mem/n7098 ) );
  MUX \Data_Mem/U7111  ( .A(\Data_Mem/n7096 ), .B(\Data_Mem/n7095 ), .S(N28), 
        .Z(\Data_Mem/n7097 ) );
  MUX \Data_Mem/U7110  ( .A(data_mem_out_wire[1037]), .B(
        data_mem_out_wire[1069]), .S(N29), .Z(\Data_Mem/n7096 ) );
  MUX \Data_Mem/U7109  ( .A(data_mem_out_wire[1101]), .B(
        data_mem_out_wire[1133]), .S(N29), .Z(\Data_Mem/n7095 ) );
  MUX \Data_Mem/U7108  ( .A(\Data_Mem/n7093 ), .B(\Data_Mem/n7092 ), .S(N28), 
        .Z(\Data_Mem/n7094 ) );
  MUX \Data_Mem/U7107  ( .A(data_mem_out_wire[1165]), .B(
        data_mem_out_wire[1197]), .S(N29), .Z(\Data_Mem/n7093 ) );
  MUX \Data_Mem/U7106  ( .A(data_mem_out_wire[1229]), .B(
        data_mem_out_wire[1261]), .S(N29), .Z(\Data_Mem/n7092 ) );
  MUX \Data_Mem/U7105  ( .A(\Data_Mem/n7090 ), .B(\Data_Mem/n7087 ), .S(N27), 
        .Z(\Data_Mem/n7091 ) );
  MUX \Data_Mem/U7104  ( .A(\Data_Mem/n7089 ), .B(\Data_Mem/n7088 ), .S(N28), 
        .Z(\Data_Mem/n7090 ) );
  MUX \Data_Mem/U7103  ( .A(data_mem_out_wire[1293]), .B(
        data_mem_out_wire[1325]), .S(N29), .Z(\Data_Mem/n7089 ) );
  MUX \Data_Mem/U7102  ( .A(data_mem_out_wire[1357]), .B(
        data_mem_out_wire[1389]), .S(N29), .Z(\Data_Mem/n7088 ) );
  MUX \Data_Mem/U7101  ( .A(\Data_Mem/n7086 ), .B(\Data_Mem/n7085 ), .S(N28), 
        .Z(\Data_Mem/n7087 ) );
  MUX \Data_Mem/U7100  ( .A(data_mem_out_wire[1421]), .B(
        data_mem_out_wire[1453]), .S(N29), .Z(\Data_Mem/n7086 ) );
  MUX \Data_Mem/U7099  ( .A(data_mem_out_wire[1485]), .B(
        data_mem_out_wire[1517]), .S(N29), .Z(\Data_Mem/n7085 ) );
  MUX \Data_Mem/U7098  ( .A(\Data_Mem/n7083 ), .B(\Data_Mem/n7076 ), .S(N26), 
        .Z(\Data_Mem/n7084 ) );
  MUX \Data_Mem/U7097  ( .A(\Data_Mem/n7082 ), .B(\Data_Mem/n7079 ), .S(N27), 
        .Z(\Data_Mem/n7083 ) );
  MUX \Data_Mem/U7096  ( .A(\Data_Mem/n7081 ), .B(\Data_Mem/n7080 ), .S(N28), 
        .Z(\Data_Mem/n7082 ) );
  MUX \Data_Mem/U7095  ( .A(data_mem_out_wire[1549]), .B(
        data_mem_out_wire[1581]), .S(N29), .Z(\Data_Mem/n7081 ) );
  MUX \Data_Mem/U7094  ( .A(data_mem_out_wire[1613]), .B(
        data_mem_out_wire[1645]), .S(N29), .Z(\Data_Mem/n7080 ) );
  MUX \Data_Mem/U7093  ( .A(\Data_Mem/n7078 ), .B(\Data_Mem/n7077 ), .S(N28), 
        .Z(\Data_Mem/n7079 ) );
  MUX \Data_Mem/U7092  ( .A(data_mem_out_wire[1677]), .B(
        data_mem_out_wire[1709]), .S(N29), .Z(\Data_Mem/n7078 ) );
  MUX \Data_Mem/U7091  ( .A(data_mem_out_wire[1741]), .B(
        data_mem_out_wire[1773]), .S(N29), .Z(\Data_Mem/n7077 ) );
  MUX \Data_Mem/U7090  ( .A(\Data_Mem/n7075 ), .B(\Data_Mem/n7072 ), .S(N27), 
        .Z(\Data_Mem/n7076 ) );
  MUX \Data_Mem/U7089  ( .A(\Data_Mem/n7074 ), .B(\Data_Mem/n7073 ), .S(N28), 
        .Z(\Data_Mem/n7075 ) );
  MUX \Data_Mem/U7088  ( .A(data_mem_out_wire[1805]), .B(
        data_mem_out_wire[1837]), .S(N29), .Z(\Data_Mem/n7074 ) );
  MUX \Data_Mem/U7087  ( .A(data_mem_out_wire[1869]), .B(
        data_mem_out_wire[1901]), .S(N29), .Z(\Data_Mem/n7073 ) );
  MUX \Data_Mem/U7086  ( .A(\Data_Mem/n7071 ), .B(\Data_Mem/n7070 ), .S(N28), 
        .Z(\Data_Mem/n7072 ) );
  MUX \Data_Mem/U7085  ( .A(data_mem_out_wire[1933]), .B(
        data_mem_out_wire[1965]), .S(N29), .Z(\Data_Mem/n7071 ) );
  MUX \Data_Mem/U7084  ( .A(data_mem_out_wire[1997]), .B(
        data_mem_out_wire[2029]), .S(N29), .Z(\Data_Mem/n7070 ) );
  MUX \Data_Mem/U7083  ( .A(\Data_Mem/n7069 ), .B(\Data_Mem/n7038 ), .S(N24), 
        .Z(c_memory[12]) );
  MUX \Data_Mem/U7082  ( .A(\Data_Mem/n7068 ), .B(\Data_Mem/n7053 ), .S(N25), 
        .Z(\Data_Mem/n7069 ) );
  MUX \Data_Mem/U7081  ( .A(\Data_Mem/n7067 ), .B(\Data_Mem/n7060 ), .S(N26), 
        .Z(\Data_Mem/n7068 ) );
  MUX \Data_Mem/U7080  ( .A(\Data_Mem/n7066 ), .B(\Data_Mem/n7063 ), .S(N27), 
        .Z(\Data_Mem/n7067 ) );
  MUX \Data_Mem/U7079  ( .A(\Data_Mem/n7065 ), .B(\Data_Mem/n7064 ), .S(N28), 
        .Z(\Data_Mem/n7066 ) );
  MUX \Data_Mem/U7078  ( .A(data_mem_out_wire[12]), .B(data_mem_out_wire[44]), 
        .S(N29), .Z(\Data_Mem/n7065 ) );
  MUX \Data_Mem/U7077  ( .A(data_mem_out_wire[76]), .B(data_mem_out_wire[108]), 
        .S(N29), .Z(\Data_Mem/n7064 ) );
  MUX \Data_Mem/U7076  ( .A(\Data_Mem/n7062 ), .B(\Data_Mem/n7061 ), .S(N28), 
        .Z(\Data_Mem/n7063 ) );
  MUX \Data_Mem/U7075  ( .A(data_mem_out_wire[140]), .B(data_mem_out_wire[172]), .S(N29), .Z(\Data_Mem/n7062 ) );
  MUX \Data_Mem/U7074  ( .A(data_mem_out_wire[204]), .B(data_mem_out_wire[236]), .S(N29), .Z(\Data_Mem/n7061 ) );
  MUX \Data_Mem/U7073  ( .A(\Data_Mem/n7059 ), .B(\Data_Mem/n7056 ), .S(N27), 
        .Z(\Data_Mem/n7060 ) );
  MUX \Data_Mem/U7072  ( .A(\Data_Mem/n7058 ), .B(\Data_Mem/n7057 ), .S(N28), 
        .Z(\Data_Mem/n7059 ) );
  MUX \Data_Mem/U7071  ( .A(data_mem_out_wire[268]), .B(data_mem_out_wire[300]), .S(N29), .Z(\Data_Mem/n7058 ) );
  MUX \Data_Mem/U7070  ( .A(data_mem_out_wire[332]), .B(data_mem_out_wire[364]), .S(N29), .Z(\Data_Mem/n7057 ) );
  MUX \Data_Mem/U7069  ( .A(\Data_Mem/n7055 ), .B(\Data_Mem/n7054 ), .S(N28), 
        .Z(\Data_Mem/n7056 ) );
  MUX \Data_Mem/U7068  ( .A(data_mem_out_wire[396]), .B(data_mem_out_wire[428]), .S(N29), .Z(\Data_Mem/n7055 ) );
  MUX \Data_Mem/U7067  ( .A(data_mem_out_wire[460]), .B(data_mem_out_wire[492]), .S(N29), .Z(\Data_Mem/n7054 ) );
  MUX \Data_Mem/U7066  ( .A(\Data_Mem/n7052 ), .B(\Data_Mem/n7045 ), .S(N26), 
        .Z(\Data_Mem/n7053 ) );
  MUX \Data_Mem/U7065  ( .A(\Data_Mem/n7051 ), .B(\Data_Mem/n7048 ), .S(N27), 
        .Z(\Data_Mem/n7052 ) );
  MUX \Data_Mem/U7064  ( .A(\Data_Mem/n7050 ), .B(\Data_Mem/n7049 ), .S(N28), 
        .Z(\Data_Mem/n7051 ) );
  MUX \Data_Mem/U7063  ( .A(data_mem_out_wire[524]), .B(data_mem_out_wire[556]), .S(N29), .Z(\Data_Mem/n7050 ) );
  MUX \Data_Mem/U7062  ( .A(data_mem_out_wire[588]), .B(data_mem_out_wire[620]), .S(N29), .Z(\Data_Mem/n7049 ) );
  MUX \Data_Mem/U7061  ( .A(\Data_Mem/n7047 ), .B(\Data_Mem/n7046 ), .S(N28), 
        .Z(\Data_Mem/n7048 ) );
  MUX \Data_Mem/U7060  ( .A(data_mem_out_wire[652]), .B(data_mem_out_wire[684]), .S(N29), .Z(\Data_Mem/n7047 ) );
  MUX \Data_Mem/U7059  ( .A(data_mem_out_wire[716]), .B(data_mem_out_wire[748]), .S(N29), .Z(\Data_Mem/n7046 ) );
  MUX \Data_Mem/U7058  ( .A(\Data_Mem/n7044 ), .B(\Data_Mem/n7041 ), .S(N27), 
        .Z(\Data_Mem/n7045 ) );
  MUX \Data_Mem/U7057  ( .A(\Data_Mem/n7043 ), .B(\Data_Mem/n7042 ), .S(N28), 
        .Z(\Data_Mem/n7044 ) );
  MUX \Data_Mem/U7056  ( .A(data_mem_out_wire[780]), .B(data_mem_out_wire[812]), .S(N29), .Z(\Data_Mem/n7043 ) );
  MUX \Data_Mem/U7055  ( .A(data_mem_out_wire[844]), .B(data_mem_out_wire[876]), .S(N29), .Z(\Data_Mem/n7042 ) );
  MUX \Data_Mem/U7054  ( .A(\Data_Mem/n7040 ), .B(\Data_Mem/n7039 ), .S(N28), 
        .Z(\Data_Mem/n7041 ) );
  MUX \Data_Mem/U7053  ( .A(data_mem_out_wire[908]), .B(data_mem_out_wire[940]), .S(N29), .Z(\Data_Mem/n7040 ) );
  MUX \Data_Mem/U7052  ( .A(data_mem_out_wire[972]), .B(
        data_mem_out_wire[1004]), .S(N29), .Z(\Data_Mem/n7039 ) );
  MUX \Data_Mem/U7051  ( .A(\Data_Mem/n7037 ), .B(\Data_Mem/n7022 ), .S(N25), 
        .Z(\Data_Mem/n7038 ) );
  MUX \Data_Mem/U7050  ( .A(\Data_Mem/n7036 ), .B(\Data_Mem/n7029 ), .S(N26), 
        .Z(\Data_Mem/n7037 ) );
  MUX \Data_Mem/U7049  ( .A(\Data_Mem/n7035 ), .B(\Data_Mem/n7032 ), .S(N27), 
        .Z(\Data_Mem/n7036 ) );
  MUX \Data_Mem/U7048  ( .A(\Data_Mem/n7034 ), .B(\Data_Mem/n7033 ), .S(N28), 
        .Z(\Data_Mem/n7035 ) );
  MUX \Data_Mem/U7047  ( .A(data_mem_out_wire[1036]), .B(
        data_mem_out_wire[1068]), .S(N29), .Z(\Data_Mem/n7034 ) );
  MUX \Data_Mem/U7046  ( .A(data_mem_out_wire[1100]), .B(
        data_mem_out_wire[1132]), .S(N29), .Z(\Data_Mem/n7033 ) );
  MUX \Data_Mem/U7045  ( .A(\Data_Mem/n7031 ), .B(\Data_Mem/n7030 ), .S(N28), 
        .Z(\Data_Mem/n7032 ) );
  MUX \Data_Mem/U7044  ( .A(data_mem_out_wire[1164]), .B(
        data_mem_out_wire[1196]), .S(N29), .Z(\Data_Mem/n7031 ) );
  MUX \Data_Mem/U7043  ( .A(data_mem_out_wire[1228]), .B(
        data_mem_out_wire[1260]), .S(N29), .Z(\Data_Mem/n7030 ) );
  MUX \Data_Mem/U7042  ( .A(\Data_Mem/n7028 ), .B(\Data_Mem/n7025 ), .S(N27), 
        .Z(\Data_Mem/n7029 ) );
  MUX \Data_Mem/U7041  ( .A(\Data_Mem/n7027 ), .B(\Data_Mem/n7026 ), .S(N28), 
        .Z(\Data_Mem/n7028 ) );
  MUX \Data_Mem/U7040  ( .A(data_mem_out_wire[1292]), .B(
        data_mem_out_wire[1324]), .S(N29), .Z(\Data_Mem/n7027 ) );
  MUX \Data_Mem/U7039  ( .A(data_mem_out_wire[1356]), .B(
        data_mem_out_wire[1388]), .S(N29), .Z(\Data_Mem/n7026 ) );
  MUX \Data_Mem/U7038  ( .A(\Data_Mem/n7024 ), .B(\Data_Mem/n7023 ), .S(N28), 
        .Z(\Data_Mem/n7025 ) );
  MUX \Data_Mem/U7037  ( .A(data_mem_out_wire[1420]), .B(
        data_mem_out_wire[1452]), .S(N29), .Z(\Data_Mem/n7024 ) );
  MUX \Data_Mem/U7036  ( .A(data_mem_out_wire[1484]), .B(
        data_mem_out_wire[1516]), .S(N29), .Z(\Data_Mem/n7023 ) );
  MUX \Data_Mem/U7035  ( .A(\Data_Mem/n7021 ), .B(\Data_Mem/n7014 ), .S(N26), 
        .Z(\Data_Mem/n7022 ) );
  MUX \Data_Mem/U7034  ( .A(\Data_Mem/n7020 ), .B(\Data_Mem/n7017 ), .S(N27), 
        .Z(\Data_Mem/n7021 ) );
  MUX \Data_Mem/U7033  ( .A(\Data_Mem/n7019 ), .B(\Data_Mem/n7018 ), .S(N28), 
        .Z(\Data_Mem/n7020 ) );
  MUX \Data_Mem/U7032  ( .A(data_mem_out_wire[1548]), .B(
        data_mem_out_wire[1580]), .S(N29), .Z(\Data_Mem/n7019 ) );
  MUX \Data_Mem/U7031  ( .A(data_mem_out_wire[1612]), .B(
        data_mem_out_wire[1644]), .S(N29), .Z(\Data_Mem/n7018 ) );
  MUX \Data_Mem/U7030  ( .A(\Data_Mem/n7016 ), .B(\Data_Mem/n7015 ), .S(N28), 
        .Z(\Data_Mem/n7017 ) );
  MUX \Data_Mem/U7029  ( .A(data_mem_out_wire[1676]), .B(
        data_mem_out_wire[1708]), .S(N29), .Z(\Data_Mem/n7016 ) );
  MUX \Data_Mem/U7028  ( .A(data_mem_out_wire[1740]), .B(
        data_mem_out_wire[1772]), .S(N29), .Z(\Data_Mem/n7015 ) );
  MUX \Data_Mem/U7027  ( .A(\Data_Mem/n7013 ), .B(\Data_Mem/n7010 ), .S(N27), 
        .Z(\Data_Mem/n7014 ) );
  MUX \Data_Mem/U7026  ( .A(\Data_Mem/n7012 ), .B(\Data_Mem/n7011 ), .S(N28), 
        .Z(\Data_Mem/n7013 ) );
  MUX \Data_Mem/U7025  ( .A(data_mem_out_wire[1804]), .B(
        data_mem_out_wire[1836]), .S(N29), .Z(\Data_Mem/n7012 ) );
  MUX \Data_Mem/U7024  ( .A(data_mem_out_wire[1868]), .B(
        data_mem_out_wire[1900]), .S(N29), .Z(\Data_Mem/n7011 ) );
  MUX \Data_Mem/U7023  ( .A(\Data_Mem/n7009 ), .B(\Data_Mem/n7008 ), .S(N28), 
        .Z(\Data_Mem/n7010 ) );
  MUX \Data_Mem/U7022  ( .A(data_mem_out_wire[1932]), .B(
        data_mem_out_wire[1964]), .S(N29), .Z(\Data_Mem/n7009 ) );
  MUX \Data_Mem/U7021  ( .A(data_mem_out_wire[1996]), .B(
        data_mem_out_wire[2028]), .S(N29), .Z(\Data_Mem/n7008 ) );
  MUX \Data_Mem/U7020  ( .A(\Data_Mem/n7007 ), .B(\Data_Mem/n6976 ), .S(N24), 
        .Z(c_memory[11]) );
  MUX \Data_Mem/U7019  ( .A(\Data_Mem/n7006 ), .B(\Data_Mem/n6991 ), .S(N25), 
        .Z(\Data_Mem/n7007 ) );
  MUX \Data_Mem/U7018  ( .A(\Data_Mem/n7005 ), .B(\Data_Mem/n6998 ), .S(N26), 
        .Z(\Data_Mem/n7006 ) );
  MUX \Data_Mem/U7017  ( .A(\Data_Mem/n7004 ), .B(\Data_Mem/n7001 ), .S(N27), 
        .Z(\Data_Mem/n7005 ) );
  MUX \Data_Mem/U7016  ( .A(\Data_Mem/n7003 ), .B(\Data_Mem/n7002 ), .S(N28), 
        .Z(\Data_Mem/n7004 ) );
  MUX \Data_Mem/U7015  ( .A(data_mem_out_wire[11]), .B(data_mem_out_wire[43]), 
        .S(N29), .Z(\Data_Mem/n7003 ) );
  MUX \Data_Mem/U7014  ( .A(data_mem_out_wire[75]), .B(data_mem_out_wire[107]), 
        .S(N29), .Z(\Data_Mem/n7002 ) );
  MUX \Data_Mem/U7013  ( .A(\Data_Mem/n7000 ), .B(\Data_Mem/n6999 ), .S(N28), 
        .Z(\Data_Mem/n7001 ) );
  MUX \Data_Mem/U7012  ( .A(data_mem_out_wire[139]), .B(data_mem_out_wire[171]), .S(N29), .Z(\Data_Mem/n7000 ) );
  MUX \Data_Mem/U7011  ( .A(data_mem_out_wire[203]), .B(data_mem_out_wire[235]), .S(N29), .Z(\Data_Mem/n6999 ) );
  MUX \Data_Mem/U7010  ( .A(\Data_Mem/n6997 ), .B(\Data_Mem/n6994 ), .S(N27), 
        .Z(\Data_Mem/n6998 ) );
  MUX \Data_Mem/U7009  ( .A(\Data_Mem/n6996 ), .B(\Data_Mem/n6995 ), .S(N28), 
        .Z(\Data_Mem/n6997 ) );
  MUX \Data_Mem/U7008  ( .A(data_mem_out_wire[267]), .B(data_mem_out_wire[299]), .S(N29), .Z(\Data_Mem/n6996 ) );
  MUX \Data_Mem/U7007  ( .A(data_mem_out_wire[331]), .B(data_mem_out_wire[363]), .S(N29), .Z(\Data_Mem/n6995 ) );
  MUX \Data_Mem/U7006  ( .A(\Data_Mem/n6993 ), .B(\Data_Mem/n6992 ), .S(N28), 
        .Z(\Data_Mem/n6994 ) );
  MUX \Data_Mem/U7005  ( .A(data_mem_out_wire[395]), .B(data_mem_out_wire[427]), .S(N29), .Z(\Data_Mem/n6993 ) );
  MUX \Data_Mem/U7004  ( .A(data_mem_out_wire[459]), .B(data_mem_out_wire[491]), .S(N29), .Z(\Data_Mem/n6992 ) );
  MUX \Data_Mem/U7003  ( .A(\Data_Mem/n6990 ), .B(\Data_Mem/n6983 ), .S(N26), 
        .Z(\Data_Mem/n6991 ) );
  MUX \Data_Mem/U7002  ( .A(\Data_Mem/n6989 ), .B(\Data_Mem/n6986 ), .S(N27), 
        .Z(\Data_Mem/n6990 ) );
  MUX \Data_Mem/U7001  ( .A(\Data_Mem/n6988 ), .B(\Data_Mem/n6987 ), .S(N28), 
        .Z(\Data_Mem/n6989 ) );
  MUX \Data_Mem/U7000  ( .A(data_mem_out_wire[523]), .B(data_mem_out_wire[555]), .S(N29), .Z(\Data_Mem/n6988 ) );
  MUX \Data_Mem/U6999  ( .A(data_mem_out_wire[587]), .B(data_mem_out_wire[619]), .S(N29), .Z(\Data_Mem/n6987 ) );
  MUX \Data_Mem/U6998  ( .A(\Data_Mem/n6985 ), .B(\Data_Mem/n6984 ), .S(N28), 
        .Z(\Data_Mem/n6986 ) );
  MUX \Data_Mem/U6997  ( .A(data_mem_out_wire[651]), .B(data_mem_out_wire[683]), .S(N29), .Z(\Data_Mem/n6985 ) );
  MUX \Data_Mem/U6996  ( .A(data_mem_out_wire[715]), .B(data_mem_out_wire[747]), .S(N29), .Z(\Data_Mem/n6984 ) );
  MUX \Data_Mem/U6995  ( .A(\Data_Mem/n6982 ), .B(\Data_Mem/n6979 ), .S(N27), 
        .Z(\Data_Mem/n6983 ) );
  MUX \Data_Mem/U6994  ( .A(\Data_Mem/n6981 ), .B(\Data_Mem/n6980 ), .S(N28), 
        .Z(\Data_Mem/n6982 ) );
  MUX \Data_Mem/U6993  ( .A(data_mem_out_wire[779]), .B(data_mem_out_wire[811]), .S(N29), .Z(\Data_Mem/n6981 ) );
  MUX \Data_Mem/U6992  ( .A(data_mem_out_wire[843]), .B(data_mem_out_wire[875]), .S(N29), .Z(\Data_Mem/n6980 ) );
  MUX \Data_Mem/U6991  ( .A(\Data_Mem/n6978 ), .B(\Data_Mem/n6977 ), .S(N28), 
        .Z(\Data_Mem/n6979 ) );
  MUX \Data_Mem/U6990  ( .A(data_mem_out_wire[907]), .B(data_mem_out_wire[939]), .S(N29), .Z(\Data_Mem/n6978 ) );
  MUX \Data_Mem/U6989  ( .A(data_mem_out_wire[971]), .B(
        data_mem_out_wire[1003]), .S(N29), .Z(\Data_Mem/n6977 ) );
  MUX \Data_Mem/U6988  ( .A(\Data_Mem/n6975 ), .B(\Data_Mem/n6960 ), .S(N25), 
        .Z(\Data_Mem/n6976 ) );
  MUX \Data_Mem/U6987  ( .A(\Data_Mem/n6974 ), .B(\Data_Mem/n6967 ), .S(N26), 
        .Z(\Data_Mem/n6975 ) );
  MUX \Data_Mem/U6986  ( .A(\Data_Mem/n6973 ), .B(\Data_Mem/n6970 ), .S(N27), 
        .Z(\Data_Mem/n6974 ) );
  MUX \Data_Mem/U6985  ( .A(\Data_Mem/n6972 ), .B(\Data_Mem/n6971 ), .S(N28), 
        .Z(\Data_Mem/n6973 ) );
  MUX \Data_Mem/U6984  ( .A(data_mem_out_wire[1035]), .B(
        data_mem_out_wire[1067]), .S(N29), .Z(\Data_Mem/n6972 ) );
  MUX \Data_Mem/U6983  ( .A(data_mem_out_wire[1099]), .B(
        data_mem_out_wire[1131]), .S(N29), .Z(\Data_Mem/n6971 ) );
  MUX \Data_Mem/U6982  ( .A(\Data_Mem/n6969 ), .B(\Data_Mem/n6968 ), .S(N28), 
        .Z(\Data_Mem/n6970 ) );
  MUX \Data_Mem/U6981  ( .A(data_mem_out_wire[1163]), .B(
        data_mem_out_wire[1195]), .S(N29), .Z(\Data_Mem/n6969 ) );
  MUX \Data_Mem/U6980  ( .A(data_mem_out_wire[1227]), .B(
        data_mem_out_wire[1259]), .S(N29), .Z(\Data_Mem/n6968 ) );
  MUX \Data_Mem/U6979  ( .A(\Data_Mem/n6966 ), .B(\Data_Mem/n6963 ), .S(N27), 
        .Z(\Data_Mem/n6967 ) );
  MUX \Data_Mem/U6978  ( .A(\Data_Mem/n6965 ), .B(\Data_Mem/n6964 ), .S(N28), 
        .Z(\Data_Mem/n6966 ) );
  MUX \Data_Mem/U6977  ( .A(data_mem_out_wire[1291]), .B(
        data_mem_out_wire[1323]), .S(N29), .Z(\Data_Mem/n6965 ) );
  MUX \Data_Mem/U6976  ( .A(data_mem_out_wire[1355]), .B(
        data_mem_out_wire[1387]), .S(N29), .Z(\Data_Mem/n6964 ) );
  MUX \Data_Mem/U6975  ( .A(\Data_Mem/n6962 ), .B(\Data_Mem/n6961 ), .S(N28), 
        .Z(\Data_Mem/n6963 ) );
  MUX \Data_Mem/U6974  ( .A(data_mem_out_wire[1419]), .B(
        data_mem_out_wire[1451]), .S(N29), .Z(\Data_Mem/n6962 ) );
  MUX \Data_Mem/U6973  ( .A(data_mem_out_wire[1483]), .B(
        data_mem_out_wire[1515]), .S(N29), .Z(\Data_Mem/n6961 ) );
  MUX \Data_Mem/U6972  ( .A(\Data_Mem/n6959 ), .B(\Data_Mem/n6952 ), .S(N26), 
        .Z(\Data_Mem/n6960 ) );
  MUX \Data_Mem/U6971  ( .A(\Data_Mem/n6958 ), .B(\Data_Mem/n6955 ), .S(N27), 
        .Z(\Data_Mem/n6959 ) );
  MUX \Data_Mem/U6970  ( .A(\Data_Mem/n6957 ), .B(\Data_Mem/n6956 ), .S(N28), 
        .Z(\Data_Mem/n6958 ) );
  MUX \Data_Mem/U6969  ( .A(data_mem_out_wire[1547]), .B(
        data_mem_out_wire[1579]), .S(N29), .Z(\Data_Mem/n6957 ) );
  MUX \Data_Mem/U6968  ( .A(data_mem_out_wire[1611]), .B(
        data_mem_out_wire[1643]), .S(N29), .Z(\Data_Mem/n6956 ) );
  MUX \Data_Mem/U6967  ( .A(\Data_Mem/n6954 ), .B(\Data_Mem/n6953 ), .S(N28), 
        .Z(\Data_Mem/n6955 ) );
  MUX \Data_Mem/U6966  ( .A(data_mem_out_wire[1675]), .B(
        data_mem_out_wire[1707]), .S(N29), .Z(\Data_Mem/n6954 ) );
  MUX \Data_Mem/U6965  ( .A(data_mem_out_wire[1739]), .B(
        data_mem_out_wire[1771]), .S(N29), .Z(\Data_Mem/n6953 ) );
  MUX \Data_Mem/U6964  ( .A(\Data_Mem/n6951 ), .B(\Data_Mem/n6948 ), .S(N27), 
        .Z(\Data_Mem/n6952 ) );
  MUX \Data_Mem/U6963  ( .A(\Data_Mem/n6950 ), .B(\Data_Mem/n6949 ), .S(N28), 
        .Z(\Data_Mem/n6951 ) );
  MUX \Data_Mem/U6962  ( .A(data_mem_out_wire[1803]), .B(
        data_mem_out_wire[1835]), .S(N29), .Z(\Data_Mem/n6950 ) );
  MUX \Data_Mem/U6961  ( .A(data_mem_out_wire[1867]), .B(
        data_mem_out_wire[1899]), .S(N29), .Z(\Data_Mem/n6949 ) );
  MUX \Data_Mem/U6960  ( .A(\Data_Mem/n6947 ), .B(\Data_Mem/n6946 ), .S(N28), 
        .Z(\Data_Mem/n6948 ) );
  MUX \Data_Mem/U6959  ( .A(data_mem_out_wire[1931]), .B(
        data_mem_out_wire[1963]), .S(N29), .Z(\Data_Mem/n6947 ) );
  MUX \Data_Mem/U6958  ( .A(data_mem_out_wire[1995]), .B(
        data_mem_out_wire[2027]), .S(N29), .Z(\Data_Mem/n6946 ) );
  MUX \Data_Mem/U6957  ( .A(\Data_Mem/n6945 ), .B(\Data_Mem/n6914 ), .S(N24), 
        .Z(c_memory[10]) );
  MUX \Data_Mem/U6956  ( .A(\Data_Mem/n6944 ), .B(\Data_Mem/n6929 ), .S(N25), 
        .Z(\Data_Mem/n6945 ) );
  MUX \Data_Mem/U6955  ( .A(\Data_Mem/n6943 ), .B(\Data_Mem/n6936 ), .S(N26), 
        .Z(\Data_Mem/n6944 ) );
  MUX \Data_Mem/U6954  ( .A(\Data_Mem/n6942 ), .B(\Data_Mem/n6939 ), .S(N27), 
        .Z(\Data_Mem/n6943 ) );
  MUX \Data_Mem/U6953  ( .A(\Data_Mem/n6941 ), .B(\Data_Mem/n6940 ), .S(N28), 
        .Z(\Data_Mem/n6942 ) );
  MUX \Data_Mem/U6952  ( .A(data_mem_out_wire[10]), .B(data_mem_out_wire[42]), 
        .S(N29), .Z(\Data_Mem/n6941 ) );
  MUX \Data_Mem/U6951  ( .A(data_mem_out_wire[74]), .B(data_mem_out_wire[106]), 
        .S(N29), .Z(\Data_Mem/n6940 ) );
  MUX \Data_Mem/U6950  ( .A(\Data_Mem/n6938 ), .B(\Data_Mem/n6937 ), .S(N28), 
        .Z(\Data_Mem/n6939 ) );
  MUX \Data_Mem/U6949  ( .A(data_mem_out_wire[138]), .B(data_mem_out_wire[170]), .S(N29), .Z(\Data_Mem/n6938 ) );
  MUX \Data_Mem/U6948  ( .A(data_mem_out_wire[202]), .B(data_mem_out_wire[234]), .S(N29), .Z(\Data_Mem/n6937 ) );
  MUX \Data_Mem/U6947  ( .A(\Data_Mem/n6935 ), .B(\Data_Mem/n6932 ), .S(N27), 
        .Z(\Data_Mem/n6936 ) );
  MUX \Data_Mem/U6946  ( .A(\Data_Mem/n6934 ), .B(\Data_Mem/n6933 ), .S(N28), 
        .Z(\Data_Mem/n6935 ) );
  MUX \Data_Mem/U6945  ( .A(data_mem_out_wire[266]), .B(data_mem_out_wire[298]), .S(N29), .Z(\Data_Mem/n6934 ) );
  MUX \Data_Mem/U6944  ( .A(data_mem_out_wire[330]), .B(data_mem_out_wire[362]), .S(N29), .Z(\Data_Mem/n6933 ) );
  MUX \Data_Mem/U6943  ( .A(\Data_Mem/n6931 ), .B(\Data_Mem/n6930 ), .S(N28), 
        .Z(\Data_Mem/n6932 ) );
  MUX \Data_Mem/U6942  ( .A(data_mem_out_wire[394]), .B(data_mem_out_wire[426]), .S(N29), .Z(\Data_Mem/n6931 ) );
  MUX \Data_Mem/U6941  ( .A(data_mem_out_wire[458]), .B(data_mem_out_wire[490]), .S(N29), .Z(\Data_Mem/n6930 ) );
  MUX \Data_Mem/U6940  ( .A(\Data_Mem/n6928 ), .B(\Data_Mem/n6921 ), .S(N26), 
        .Z(\Data_Mem/n6929 ) );
  MUX \Data_Mem/U6939  ( .A(\Data_Mem/n6927 ), .B(\Data_Mem/n6924 ), .S(N27), 
        .Z(\Data_Mem/n6928 ) );
  MUX \Data_Mem/U6938  ( .A(\Data_Mem/n6926 ), .B(\Data_Mem/n6925 ), .S(N28), 
        .Z(\Data_Mem/n6927 ) );
  MUX \Data_Mem/U6937  ( .A(data_mem_out_wire[522]), .B(data_mem_out_wire[554]), .S(N29), .Z(\Data_Mem/n6926 ) );
  MUX \Data_Mem/U6936  ( .A(data_mem_out_wire[586]), .B(data_mem_out_wire[618]), .S(N29), .Z(\Data_Mem/n6925 ) );
  MUX \Data_Mem/U6935  ( .A(\Data_Mem/n6923 ), .B(\Data_Mem/n6922 ), .S(N28), 
        .Z(\Data_Mem/n6924 ) );
  MUX \Data_Mem/U6934  ( .A(data_mem_out_wire[650]), .B(data_mem_out_wire[682]), .S(N29), .Z(\Data_Mem/n6923 ) );
  MUX \Data_Mem/U6933  ( .A(data_mem_out_wire[714]), .B(data_mem_out_wire[746]), .S(N29), .Z(\Data_Mem/n6922 ) );
  MUX \Data_Mem/U6932  ( .A(\Data_Mem/n6920 ), .B(\Data_Mem/n6917 ), .S(N27), 
        .Z(\Data_Mem/n6921 ) );
  MUX \Data_Mem/U6931  ( .A(\Data_Mem/n6919 ), .B(\Data_Mem/n6918 ), .S(N28), 
        .Z(\Data_Mem/n6920 ) );
  MUX \Data_Mem/U6930  ( .A(data_mem_out_wire[778]), .B(data_mem_out_wire[810]), .S(N29), .Z(\Data_Mem/n6919 ) );
  MUX \Data_Mem/U6929  ( .A(data_mem_out_wire[842]), .B(data_mem_out_wire[874]), .S(N29), .Z(\Data_Mem/n6918 ) );
  MUX \Data_Mem/U6928  ( .A(\Data_Mem/n6916 ), .B(\Data_Mem/n6915 ), .S(N28), 
        .Z(\Data_Mem/n6917 ) );
  MUX \Data_Mem/U6927  ( .A(data_mem_out_wire[906]), .B(data_mem_out_wire[938]), .S(N29), .Z(\Data_Mem/n6916 ) );
  MUX \Data_Mem/U6926  ( .A(data_mem_out_wire[970]), .B(
        data_mem_out_wire[1002]), .S(N29), .Z(\Data_Mem/n6915 ) );
  MUX \Data_Mem/U6925  ( .A(\Data_Mem/n6913 ), .B(\Data_Mem/n6898 ), .S(N25), 
        .Z(\Data_Mem/n6914 ) );
  MUX \Data_Mem/U6924  ( .A(\Data_Mem/n6912 ), .B(\Data_Mem/n6905 ), .S(N26), 
        .Z(\Data_Mem/n6913 ) );
  MUX \Data_Mem/U6923  ( .A(\Data_Mem/n6911 ), .B(\Data_Mem/n6908 ), .S(N27), 
        .Z(\Data_Mem/n6912 ) );
  MUX \Data_Mem/U6922  ( .A(\Data_Mem/n6910 ), .B(\Data_Mem/n6909 ), .S(N28), 
        .Z(\Data_Mem/n6911 ) );
  MUX \Data_Mem/U6921  ( .A(data_mem_out_wire[1034]), .B(
        data_mem_out_wire[1066]), .S(N29), .Z(\Data_Mem/n6910 ) );
  MUX \Data_Mem/U6920  ( .A(data_mem_out_wire[1098]), .B(
        data_mem_out_wire[1130]), .S(N29), .Z(\Data_Mem/n6909 ) );
  MUX \Data_Mem/U6919  ( .A(\Data_Mem/n6907 ), .B(\Data_Mem/n6906 ), .S(N28), 
        .Z(\Data_Mem/n6908 ) );
  MUX \Data_Mem/U6918  ( .A(data_mem_out_wire[1162]), .B(
        data_mem_out_wire[1194]), .S(N29), .Z(\Data_Mem/n6907 ) );
  MUX \Data_Mem/U6917  ( .A(data_mem_out_wire[1226]), .B(
        data_mem_out_wire[1258]), .S(N29), .Z(\Data_Mem/n6906 ) );
  MUX \Data_Mem/U6916  ( .A(\Data_Mem/n6904 ), .B(\Data_Mem/n6901 ), .S(N27), 
        .Z(\Data_Mem/n6905 ) );
  MUX \Data_Mem/U6915  ( .A(\Data_Mem/n6903 ), .B(\Data_Mem/n6902 ), .S(N28), 
        .Z(\Data_Mem/n6904 ) );
  MUX \Data_Mem/U6914  ( .A(data_mem_out_wire[1290]), .B(
        data_mem_out_wire[1322]), .S(N29), .Z(\Data_Mem/n6903 ) );
  MUX \Data_Mem/U6913  ( .A(data_mem_out_wire[1354]), .B(
        data_mem_out_wire[1386]), .S(N29), .Z(\Data_Mem/n6902 ) );
  MUX \Data_Mem/U6912  ( .A(\Data_Mem/n6900 ), .B(\Data_Mem/n6899 ), .S(N28), 
        .Z(\Data_Mem/n6901 ) );
  MUX \Data_Mem/U6911  ( .A(data_mem_out_wire[1418]), .B(
        data_mem_out_wire[1450]), .S(N29), .Z(\Data_Mem/n6900 ) );
  MUX \Data_Mem/U6910  ( .A(data_mem_out_wire[1482]), .B(
        data_mem_out_wire[1514]), .S(N29), .Z(\Data_Mem/n6899 ) );
  MUX \Data_Mem/U6909  ( .A(\Data_Mem/n6897 ), .B(\Data_Mem/n6890 ), .S(N26), 
        .Z(\Data_Mem/n6898 ) );
  MUX \Data_Mem/U6908  ( .A(\Data_Mem/n6896 ), .B(\Data_Mem/n6893 ), .S(N27), 
        .Z(\Data_Mem/n6897 ) );
  MUX \Data_Mem/U6907  ( .A(\Data_Mem/n6895 ), .B(\Data_Mem/n6894 ), .S(N28), 
        .Z(\Data_Mem/n6896 ) );
  MUX \Data_Mem/U6906  ( .A(data_mem_out_wire[1546]), .B(
        data_mem_out_wire[1578]), .S(N29), .Z(\Data_Mem/n6895 ) );
  MUX \Data_Mem/U6905  ( .A(data_mem_out_wire[1610]), .B(
        data_mem_out_wire[1642]), .S(N29), .Z(\Data_Mem/n6894 ) );
  MUX \Data_Mem/U6904  ( .A(\Data_Mem/n6892 ), .B(\Data_Mem/n6891 ), .S(N28), 
        .Z(\Data_Mem/n6893 ) );
  MUX \Data_Mem/U6903  ( .A(data_mem_out_wire[1674]), .B(
        data_mem_out_wire[1706]), .S(N29), .Z(\Data_Mem/n6892 ) );
  MUX \Data_Mem/U6902  ( .A(data_mem_out_wire[1738]), .B(
        data_mem_out_wire[1770]), .S(N29), .Z(\Data_Mem/n6891 ) );
  MUX \Data_Mem/U6901  ( .A(\Data_Mem/n6889 ), .B(\Data_Mem/n6886 ), .S(N27), 
        .Z(\Data_Mem/n6890 ) );
  MUX \Data_Mem/U6900  ( .A(\Data_Mem/n6888 ), .B(\Data_Mem/n6887 ), .S(N28), 
        .Z(\Data_Mem/n6889 ) );
  MUX \Data_Mem/U6899  ( .A(data_mem_out_wire[1802]), .B(
        data_mem_out_wire[1834]), .S(N29), .Z(\Data_Mem/n6888 ) );
  MUX \Data_Mem/U6898  ( .A(data_mem_out_wire[1866]), .B(
        data_mem_out_wire[1898]), .S(N29), .Z(\Data_Mem/n6887 ) );
  MUX \Data_Mem/U6897  ( .A(\Data_Mem/n6885 ), .B(\Data_Mem/n6884 ), .S(N28), 
        .Z(\Data_Mem/n6886 ) );
  MUX \Data_Mem/U6896  ( .A(data_mem_out_wire[1930]), .B(
        data_mem_out_wire[1962]), .S(N29), .Z(\Data_Mem/n6885 ) );
  MUX \Data_Mem/U6895  ( .A(data_mem_out_wire[1994]), .B(
        data_mem_out_wire[2026]), .S(N29), .Z(\Data_Mem/n6884 ) );
  MUX \Data_Mem/U6894  ( .A(\Data_Mem/n6883 ), .B(\Data_Mem/n6852 ), .S(N24), 
        .Z(c_memory[9]) );
  MUX \Data_Mem/U6893  ( .A(\Data_Mem/n6882 ), .B(\Data_Mem/n6867 ), .S(N25), 
        .Z(\Data_Mem/n6883 ) );
  MUX \Data_Mem/U6892  ( .A(\Data_Mem/n6881 ), .B(\Data_Mem/n6874 ), .S(N26), 
        .Z(\Data_Mem/n6882 ) );
  MUX \Data_Mem/U6891  ( .A(\Data_Mem/n6880 ), .B(\Data_Mem/n6877 ), .S(N27), 
        .Z(\Data_Mem/n6881 ) );
  MUX \Data_Mem/U6890  ( .A(\Data_Mem/n6879 ), .B(\Data_Mem/n6878 ), .S(N28), 
        .Z(\Data_Mem/n6880 ) );
  MUX \Data_Mem/U6889  ( .A(data_mem_out_wire[9]), .B(data_mem_out_wire[41]), 
        .S(N29), .Z(\Data_Mem/n6879 ) );
  MUX \Data_Mem/U6888  ( .A(data_mem_out_wire[73]), .B(data_mem_out_wire[105]), 
        .S(N29), .Z(\Data_Mem/n6878 ) );
  MUX \Data_Mem/U6887  ( .A(\Data_Mem/n6876 ), .B(\Data_Mem/n6875 ), .S(N28), 
        .Z(\Data_Mem/n6877 ) );
  MUX \Data_Mem/U6886  ( .A(data_mem_out_wire[137]), .B(data_mem_out_wire[169]), .S(N29), .Z(\Data_Mem/n6876 ) );
  MUX \Data_Mem/U6885  ( .A(data_mem_out_wire[201]), .B(data_mem_out_wire[233]), .S(N29), .Z(\Data_Mem/n6875 ) );
  MUX \Data_Mem/U6884  ( .A(\Data_Mem/n6873 ), .B(\Data_Mem/n6870 ), .S(N27), 
        .Z(\Data_Mem/n6874 ) );
  MUX \Data_Mem/U6883  ( .A(\Data_Mem/n6872 ), .B(\Data_Mem/n6871 ), .S(N28), 
        .Z(\Data_Mem/n6873 ) );
  MUX \Data_Mem/U6882  ( .A(data_mem_out_wire[265]), .B(data_mem_out_wire[297]), .S(N29), .Z(\Data_Mem/n6872 ) );
  MUX \Data_Mem/U6881  ( .A(data_mem_out_wire[329]), .B(data_mem_out_wire[361]), .S(N29), .Z(\Data_Mem/n6871 ) );
  MUX \Data_Mem/U6880  ( .A(\Data_Mem/n6869 ), .B(\Data_Mem/n6868 ), .S(N28), 
        .Z(\Data_Mem/n6870 ) );
  MUX \Data_Mem/U6879  ( .A(data_mem_out_wire[393]), .B(data_mem_out_wire[425]), .S(N29), .Z(\Data_Mem/n6869 ) );
  MUX \Data_Mem/U6878  ( .A(data_mem_out_wire[457]), .B(data_mem_out_wire[489]), .S(N29), .Z(\Data_Mem/n6868 ) );
  MUX \Data_Mem/U6877  ( .A(\Data_Mem/n6866 ), .B(\Data_Mem/n6859 ), .S(N26), 
        .Z(\Data_Mem/n6867 ) );
  MUX \Data_Mem/U6876  ( .A(\Data_Mem/n6865 ), .B(\Data_Mem/n6862 ), .S(N27), 
        .Z(\Data_Mem/n6866 ) );
  MUX \Data_Mem/U6875  ( .A(\Data_Mem/n6864 ), .B(\Data_Mem/n6863 ), .S(N28), 
        .Z(\Data_Mem/n6865 ) );
  MUX \Data_Mem/U6874  ( .A(data_mem_out_wire[521]), .B(data_mem_out_wire[553]), .S(N29), .Z(\Data_Mem/n6864 ) );
  MUX \Data_Mem/U6873  ( .A(data_mem_out_wire[585]), .B(data_mem_out_wire[617]), .S(N29), .Z(\Data_Mem/n6863 ) );
  MUX \Data_Mem/U6872  ( .A(\Data_Mem/n6861 ), .B(\Data_Mem/n6860 ), .S(N28), 
        .Z(\Data_Mem/n6862 ) );
  MUX \Data_Mem/U6871  ( .A(data_mem_out_wire[649]), .B(data_mem_out_wire[681]), .S(N29), .Z(\Data_Mem/n6861 ) );
  MUX \Data_Mem/U6870  ( .A(data_mem_out_wire[713]), .B(data_mem_out_wire[745]), .S(N29), .Z(\Data_Mem/n6860 ) );
  MUX \Data_Mem/U6869  ( .A(\Data_Mem/n6858 ), .B(\Data_Mem/n6855 ), .S(N27), 
        .Z(\Data_Mem/n6859 ) );
  MUX \Data_Mem/U6868  ( .A(\Data_Mem/n6857 ), .B(\Data_Mem/n6856 ), .S(N28), 
        .Z(\Data_Mem/n6858 ) );
  MUX \Data_Mem/U6867  ( .A(data_mem_out_wire[777]), .B(data_mem_out_wire[809]), .S(N29), .Z(\Data_Mem/n6857 ) );
  MUX \Data_Mem/U6866  ( .A(data_mem_out_wire[841]), .B(data_mem_out_wire[873]), .S(N29), .Z(\Data_Mem/n6856 ) );
  MUX \Data_Mem/U6865  ( .A(\Data_Mem/n6854 ), .B(\Data_Mem/n6853 ), .S(N28), 
        .Z(\Data_Mem/n6855 ) );
  MUX \Data_Mem/U6864  ( .A(data_mem_out_wire[905]), .B(data_mem_out_wire[937]), .S(N29), .Z(\Data_Mem/n6854 ) );
  MUX \Data_Mem/U6863  ( .A(data_mem_out_wire[969]), .B(
        data_mem_out_wire[1001]), .S(N29), .Z(\Data_Mem/n6853 ) );
  MUX \Data_Mem/U6862  ( .A(\Data_Mem/n6851 ), .B(\Data_Mem/n6836 ), .S(N25), 
        .Z(\Data_Mem/n6852 ) );
  MUX \Data_Mem/U6861  ( .A(\Data_Mem/n6850 ), .B(\Data_Mem/n6843 ), .S(N26), 
        .Z(\Data_Mem/n6851 ) );
  MUX \Data_Mem/U6860  ( .A(\Data_Mem/n6849 ), .B(\Data_Mem/n6846 ), .S(N27), 
        .Z(\Data_Mem/n6850 ) );
  MUX \Data_Mem/U6859  ( .A(\Data_Mem/n6848 ), .B(\Data_Mem/n6847 ), .S(N28), 
        .Z(\Data_Mem/n6849 ) );
  MUX \Data_Mem/U6858  ( .A(data_mem_out_wire[1033]), .B(
        data_mem_out_wire[1065]), .S(N29), .Z(\Data_Mem/n6848 ) );
  MUX \Data_Mem/U6857  ( .A(data_mem_out_wire[1097]), .B(
        data_mem_out_wire[1129]), .S(N29), .Z(\Data_Mem/n6847 ) );
  MUX \Data_Mem/U6856  ( .A(\Data_Mem/n6845 ), .B(\Data_Mem/n6844 ), .S(N28), 
        .Z(\Data_Mem/n6846 ) );
  MUX \Data_Mem/U6855  ( .A(data_mem_out_wire[1161]), .B(
        data_mem_out_wire[1193]), .S(N29), .Z(\Data_Mem/n6845 ) );
  MUX \Data_Mem/U6854  ( .A(data_mem_out_wire[1225]), .B(
        data_mem_out_wire[1257]), .S(N29), .Z(\Data_Mem/n6844 ) );
  MUX \Data_Mem/U6853  ( .A(\Data_Mem/n6842 ), .B(\Data_Mem/n6839 ), .S(N27), 
        .Z(\Data_Mem/n6843 ) );
  MUX \Data_Mem/U6852  ( .A(\Data_Mem/n6841 ), .B(\Data_Mem/n6840 ), .S(N28), 
        .Z(\Data_Mem/n6842 ) );
  MUX \Data_Mem/U6851  ( .A(data_mem_out_wire[1289]), .B(
        data_mem_out_wire[1321]), .S(N29), .Z(\Data_Mem/n6841 ) );
  MUX \Data_Mem/U6850  ( .A(data_mem_out_wire[1353]), .B(
        data_mem_out_wire[1385]), .S(N29), .Z(\Data_Mem/n6840 ) );
  MUX \Data_Mem/U6849  ( .A(\Data_Mem/n6838 ), .B(\Data_Mem/n6837 ), .S(N28), 
        .Z(\Data_Mem/n6839 ) );
  MUX \Data_Mem/U6848  ( .A(data_mem_out_wire[1417]), .B(
        data_mem_out_wire[1449]), .S(N29), .Z(\Data_Mem/n6838 ) );
  MUX \Data_Mem/U6847  ( .A(data_mem_out_wire[1481]), .B(
        data_mem_out_wire[1513]), .S(N29), .Z(\Data_Mem/n6837 ) );
  MUX \Data_Mem/U6846  ( .A(\Data_Mem/n6835 ), .B(\Data_Mem/n6828 ), .S(N26), 
        .Z(\Data_Mem/n6836 ) );
  MUX \Data_Mem/U6845  ( .A(\Data_Mem/n6834 ), .B(\Data_Mem/n6831 ), .S(N27), 
        .Z(\Data_Mem/n6835 ) );
  MUX \Data_Mem/U6844  ( .A(\Data_Mem/n6833 ), .B(\Data_Mem/n6832 ), .S(N28), 
        .Z(\Data_Mem/n6834 ) );
  MUX \Data_Mem/U6843  ( .A(data_mem_out_wire[1545]), .B(
        data_mem_out_wire[1577]), .S(N29), .Z(\Data_Mem/n6833 ) );
  MUX \Data_Mem/U6842  ( .A(data_mem_out_wire[1609]), .B(
        data_mem_out_wire[1641]), .S(N29), .Z(\Data_Mem/n6832 ) );
  MUX \Data_Mem/U6841  ( .A(\Data_Mem/n6830 ), .B(\Data_Mem/n6829 ), .S(N28), 
        .Z(\Data_Mem/n6831 ) );
  MUX \Data_Mem/U6840  ( .A(data_mem_out_wire[1673]), .B(
        data_mem_out_wire[1705]), .S(N29), .Z(\Data_Mem/n6830 ) );
  MUX \Data_Mem/U6839  ( .A(data_mem_out_wire[1737]), .B(
        data_mem_out_wire[1769]), .S(N29), .Z(\Data_Mem/n6829 ) );
  MUX \Data_Mem/U6838  ( .A(\Data_Mem/n6827 ), .B(\Data_Mem/n6824 ), .S(N27), 
        .Z(\Data_Mem/n6828 ) );
  MUX \Data_Mem/U6837  ( .A(\Data_Mem/n6826 ), .B(\Data_Mem/n6825 ), .S(N28), 
        .Z(\Data_Mem/n6827 ) );
  MUX \Data_Mem/U6836  ( .A(data_mem_out_wire[1801]), .B(
        data_mem_out_wire[1833]), .S(N29), .Z(\Data_Mem/n6826 ) );
  MUX \Data_Mem/U6835  ( .A(data_mem_out_wire[1865]), .B(
        data_mem_out_wire[1897]), .S(N29), .Z(\Data_Mem/n6825 ) );
  MUX \Data_Mem/U6834  ( .A(\Data_Mem/n6823 ), .B(\Data_Mem/n6822 ), .S(N28), 
        .Z(\Data_Mem/n6824 ) );
  MUX \Data_Mem/U6833  ( .A(data_mem_out_wire[1929]), .B(
        data_mem_out_wire[1961]), .S(N29), .Z(\Data_Mem/n6823 ) );
  MUX \Data_Mem/U6832  ( .A(data_mem_out_wire[1993]), .B(
        data_mem_out_wire[2025]), .S(N29), .Z(\Data_Mem/n6822 ) );
  MUX \Data_Mem/U6831  ( .A(\Data_Mem/n6821 ), .B(\Data_Mem/n6790 ), .S(N24), 
        .Z(c_memory[8]) );
  MUX \Data_Mem/U6830  ( .A(\Data_Mem/n6820 ), .B(\Data_Mem/n6805 ), .S(N25), 
        .Z(\Data_Mem/n6821 ) );
  MUX \Data_Mem/U6829  ( .A(\Data_Mem/n6819 ), .B(\Data_Mem/n6812 ), .S(N26), 
        .Z(\Data_Mem/n6820 ) );
  MUX \Data_Mem/U6828  ( .A(\Data_Mem/n6818 ), .B(\Data_Mem/n6815 ), .S(N27), 
        .Z(\Data_Mem/n6819 ) );
  MUX \Data_Mem/U6827  ( .A(\Data_Mem/n6817 ), .B(\Data_Mem/n6816 ), .S(N28), 
        .Z(\Data_Mem/n6818 ) );
  MUX \Data_Mem/U6826  ( .A(data_mem_out_wire[8]), .B(data_mem_out_wire[40]), 
        .S(N29), .Z(\Data_Mem/n6817 ) );
  MUX \Data_Mem/U6825  ( .A(data_mem_out_wire[72]), .B(data_mem_out_wire[104]), 
        .S(N29), .Z(\Data_Mem/n6816 ) );
  MUX \Data_Mem/U6824  ( .A(\Data_Mem/n6814 ), .B(\Data_Mem/n6813 ), .S(N28), 
        .Z(\Data_Mem/n6815 ) );
  MUX \Data_Mem/U6823  ( .A(data_mem_out_wire[136]), .B(data_mem_out_wire[168]), .S(N29), .Z(\Data_Mem/n6814 ) );
  MUX \Data_Mem/U6822  ( .A(data_mem_out_wire[200]), .B(data_mem_out_wire[232]), .S(N29), .Z(\Data_Mem/n6813 ) );
  MUX \Data_Mem/U6821  ( .A(\Data_Mem/n6811 ), .B(\Data_Mem/n6808 ), .S(N27), 
        .Z(\Data_Mem/n6812 ) );
  MUX \Data_Mem/U6820  ( .A(\Data_Mem/n6810 ), .B(\Data_Mem/n6809 ), .S(N28), 
        .Z(\Data_Mem/n6811 ) );
  MUX \Data_Mem/U6819  ( .A(data_mem_out_wire[264]), .B(data_mem_out_wire[296]), .S(N29), .Z(\Data_Mem/n6810 ) );
  MUX \Data_Mem/U6818  ( .A(data_mem_out_wire[328]), .B(data_mem_out_wire[360]), .S(N29), .Z(\Data_Mem/n6809 ) );
  MUX \Data_Mem/U6817  ( .A(\Data_Mem/n6807 ), .B(\Data_Mem/n6806 ), .S(N28), 
        .Z(\Data_Mem/n6808 ) );
  MUX \Data_Mem/U6816  ( .A(data_mem_out_wire[392]), .B(data_mem_out_wire[424]), .S(N29), .Z(\Data_Mem/n6807 ) );
  MUX \Data_Mem/U6815  ( .A(data_mem_out_wire[456]), .B(data_mem_out_wire[488]), .S(N29), .Z(\Data_Mem/n6806 ) );
  MUX \Data_Mem/U6814  ( .A(\Data_Mem/n6804 ), .B(\Data_Mem/n6797 ), .S(N26), 
        .Z(\Data_Mem/n6805 ) );
  MUX \Data_Mem/U6813  ( .A(\Data_Mem/n6803 ), .B(\Data_Mem/n6800 ), .S(N27), 
        .Z(\Data_Mem/n6804 ) );
  MUX \Data_Mem/U6812  ( .A(\Data_Mem/n6802 ), .B(\Data_Mem/n6801 ), .S(N28), 
        .Z(\Data_Mem/n6803 ) );
  MUX \Data_Mem/U6811  ( .A(data_mem_out_wire[520]), .B(data_mem_out_wire[552]), .S(N29), .Z(\Data_Mem/n6802 ) );
  MUX \Data_Mem/U6810  ( .A(data_mem_out_wire[584]), .B(data_mem_out_wire[616]), .S(N29), .Z(\Data_Mem/n6801 ) );
  MUX \Data_Mem/U6809  ( .A(\Data_Mem/n6799 ), .B(\Data_Mem/n6798 ), .S(N28), 
        .Z(\Data_Mem/n6800 ) );
  MUX \Data_Mem/U6808  ( .A(data_mem_out_wire[648]), .B(data_mem_out_wire[680]), .S(N29), .Z(\Data_Mem/n6799 ) );
  MUX \Data_Mem/U6807  ( .A(data_mem_out_wire[712]), .B(data_mem_out_wire[744]), .S(N29), .Z(\Data_Mem/n6798 ) );
  MUX \Data_Mem/U6806  ( .A(\Data_Mem/n6796 ), .B(\Data_Mem/n6793 ), .S(N27), 
        .Z(\Data_Mem/n6797 ) );
  MUX \Data_Mem/U6805  ( .A(\Data_Mem/n6795 ), .B(\Data_Mem/n6794 ), .S(N28), 
        .Z(\Data_Mem/n6796 ) );
  MUX \Data_Mem/U6804  ( .A(data_mem_out_wire[776]), .B(data_mem_out_wire[808]), .S(N29), .Z(\Data_Mem/n6795 ) );
  MUX \Data_Mem/U6803  ( .A(data_mem_out_wire[840]), .B(data_mem_out_wire[872]), .S(N29), .Z(\Data_Mem/n6794 ) );
  MUX \Data_Mem/U6802  ( .A(\Data_Mem/n6792 ), .B(\Data_Mem/n6791 ), .S(N28), 
        .Z(\Data_Mem/n6793 ) );
  MUX \Data_Mem/U6801  ( .A(data_mem_out_wire[904]), .B(data_mem_out_wire[936]), .S(N29), .Z(\Data_Mem/n6792 ) );
  MUX \Data_Mem/U6800  ( .A(data_mem_out_wire[968]), .B(
        data_mem_out_wire[1000]), .S(N29), .Z(\Data_Mem/n6791 ) );
  MUX \Data_Mem/U6799  ( .A(\Data_Mem/n6789 ), .B(\Data_Mem/n6774 ), .S(N25), 
        .Z(\Data_Mem/n6790 ) );
  MUX \Data_Mem/U6798  ( .A(\Data_Mem/n6788 ), .B(\Data_Mem/n6781 ), .S(N26), 
        .Z(\Data_Mem/n6789 ) );
  MUX \Data_Mem/U6797  ( .A(\Data_Mem/n6787 ), .B(\Data_Mem/n6784 ), .S(N27), 
        .Z(\Data_Mem/n6788 ) );
  MUX \Data_Mem/U6796  ( .A(\Data_Mem/n6786 ), .B(\Data_Mem/n6785 ), .S(N28), 
        .Z(\Data_Mem/n6787 ) );
  MUX \Data_Mem/U6795  ( .A(data_mem_out_wire[1032]), .B(
        data_mem_out_wire[1064]), .S(N29), .Z(\Data_Mem/n6786 ) );
  MUX \Data_Mem/U6794  ( .A(data_mem_out_wire[1096]), .B(
        data_mem_out_wire[1128]), .S(N29), .Z(\Data_Mem/n6785 ) );
  MUX \Data_Mem/U6793  ( .A(\Data_Mem/n6783 ), .B(\Data_Mem/n6782 ), .S(N28), 
        .Z(\Data_Mem/n6784 ) );
  MUX \Data_Mem/U6792  ( .A(data_mem_out_wire[1160]), .B(
        data_mem_out_wire[1192]), .S(N29), .Z(\Data_Mem/n6783 ) );
  MUX \Data_Mem/U6791  ( .A(data_mem_out_wire[1224]), .B(
        data_mem_out_wire[1256]), .S(N29), .Z(\Data_Mem/n6782 ) );
  MUX \Data_Mem/U6790  ( .A(\Data_Mem/n6780 ), .B(\Data_Mem/n6777 ), .S(N27), 
        .Z(\Data_Mem/n6781 ) );
  MUX \Data_Mem/U6789  ( .A(\Data_Mem/n6779 ), .B(\Data_Mem/n6778 ), .S(N28), 
        .Z(\Data_Mem/n6780 ) );
  MUX \Data_Mem/U6788  ( .A(data_mem_out_wire[1288]), .B(
        data_mem_out_wire[1320]), .S(N29), .Z(\Data_Mem/n6779 ) );
  MUX \Data_Mem/U6787  ( .A(data_mem_out_wire[1352]), .B(
        data_mem_out_wire[1384]), .S(N29), .Z(\Data_Mem/n6778 ) );
  MUX \Data_Mem/U6786  ( .A(\Data_Mem/n6776 ), .B(\Data_Mem/n6775 ), .S(N28), 
        .Z(\Data_Mem/n6777 ) );
  MUX \Data_Mem/U6785  ( .A(data_mem_out_wire[1416]), .B(
        data_mem_out_wire[1448]), .S(N29), .Z(\Data_Mem/n6776 ) );
  MUX \Data_Mem/U6784  ( .A(data_mem_out_wire[1480]), .B(
        data_mem_out_wire[1512]), .S(N29), .Z(\Data_Mem/n6775 ) );
  MUX \Data_Mem/U6783  ( .A(\Data_Mem/n6773 ), .B(\Data_Mem/n6766 ), .S(N26), 
        .Z(\Data_Mem/n6774 ) );
  MUX \Data_Mem/U6782  ( .A(\Data_Mem/n6772 ), .B(\Data_Mem/n6769 ), .S(N27), 
        .Z(\Data_Mem/n6773 ) );
  MUX \Data_Mem/U6781  ( .A(\Data_Mem/n6771 ), .B(\Data_Mem/n6770 ), .S(N28), 
        .Z(\Data_Mem/n6772 ) );
  MUX \Data_Mem/U6780  ( .A(data_mem_out_wire[1544]), .B(
        data_mem_out_wire[1576]), .S(N29), .Z(\Data_Mem/n6771 ) );
  MUX \Data_Mem/U6779  ( .A(data_mem_out_wire[1608]), .B(
        data_mem_out_wire[1640]), .S(N29), .Z(\Data_Mem/n6770 ) );
  MUX \Data_Mem/U6778  ( .A(\Data_Mem/n6768 ), .B(\Data_Mem/n6767 ), .S(N28), 
        .Z(\Data_Mem/n6769 ) );
  MUX \Data_Mem/U6777  ( .A(data_mem_out_wire[1672]), .B(
        data_mem_out_wire[1704]), .S(N29), .Z(\Data_Mem/n6768 ) );
  MUX \Data_Mem/U6776  ( .A(data_mem_out_wire[1736]), .B(
        data_mem_out_wire[1768]), .S(N29), .Z(\Data_Mem/n6767 ) );
  MUX \Data_Mem/U6775  ( .A(\Data_Mem/n6765 ), .B(\Data_Mem/n6762 ), .S(N27), 
        .Z(\Data_Mem/n6766 ) );
  MUX \Data_Mem/U6774  ( .A(\Data_Mem/n6764 ), .B(\Data_Mem/n6763 ), .S(N28), 
        .Z(\Data_Mem/n6765 ) );
  MUX \Data_Mem/U6773  ( .A(data_mem_out_wire[1800]), .B(
        data_mem_out_wire[1832]), .S(N29), .Z(\Data_Mem/n6764 ) );
  MUX \Data_Mem/U6772  ( .A(data_mem_out_wire[1864]), .B(
        data_mem_out_wire[1896]), .S(N29), .Z(\Data_Mem/n6763 ) );
  MUX \Data_Mem/U6771  ( .A(\Data_Mem/n6761 ), .B(\Data_Mem/n6760 ), .S(N28), 
        .Z(\Data_Mem/n6762 ) );
  MUX \Data_Mem/U6770  ( .A(data_mem_out_wire[1928]), .B(
        data_mem_out_wire[1960]), .S(N29), .Z(\Data_Mem/n6761 ) );
  MUX \Data_Mem/U6769  ( .A(data_mem_out_wire[1992]), .B(
        data_mem_out_wire[2024]), .S(N29), .Z(\Data_Mem/n6760 ) );
  MUX \Data_Mem/U6768  ( .A(\Data_Mem/n6759 ), .B(\Data_Mem/n6728 ), .S(N24), 
        .Z(c_memory[7]) );
  MUX \Data_Mem/U6767  ( .A(\Data_Mem/n6758 ), .B(\Data_Mem/n6743 ), .S(N25), 
        .Z(\Data_Mem/n6759 ) );
  MUX \Data_Mem/U6766  ( .A(\Data_Mem/n6757 ), .B(\Data_Mem/n6750 ), .S(N26), 
        .Z(\Data_Mem/n6758 ) );
  MUX \Data_Mem/U6765  ( .A(\Data_Mem/n6756 ), .B(\Data_Mem/n6753 ), .S(N27), 
        .Z(\Data_Mem/n6757 ) );
  MUX \Data_Mem/U6764  ( .A(\Data_Mem/n6755 ), .B(\Data_Mem/n6754 ), .S(N28), 
        .Z(\Data_Mem/n6756 ) );
  MUX \Data_Mem/U6763  ( .A(data_mem_out_wire[7]), .B(data_mem_out_wire[39]), 
        .S(N29), .Z(\Data_Mem/n6755 ) );
  MUX \Data_Mem/U6762  ( .A(data_mem_out_wire[71]), .B(data_mem_out_wire[103]), 
        .S(N29), .Z(\Data_Mem/n6754 ) );
  MUX \Data_Mem/U6761  ( .A(\Data_Mem/n6752 ), .B(\Data_Mem/n6751 ), .S(N28), 
        .Z(\Data_Mem/n6753 ) );
  MUX \Data_Mem/U6760  ( .A(data_mem_out_wire[135]), .B(data_mem_out_wire[167]), .S(N29), .Z(\Data_Mem/n6752 ) );
  MUX \Data_Mem/U6759  ( .A(data_mem_out_wire[199]), .B(data_mem_out_wire[231]), .S(N29), .Z(\Data_Mem/n6751 ) );
  MUX \Data_Mem/U6758  ( .A(\Data_Mem/n6749 ), .B(\Data_Mem/n6746 ), .S(N27), 
        .Z(\Data_Mem/n6750 ) );
  MUX \Data_Mem/U6757  ( .A(\Data_Mem/n6748 ), .B(\Data_Mem/n6747 ), .S(N28), 
        .Z(\Data_Mem/n6749 ) );
  MUX \Data_Mem/U6756  ( .A(data_mem_out_wire[263]), .B(data_mem_out_wire[295]), .S(N29), .Z(\Data_Mem/n6748 ) );
  MUX \Data_Mem/U6755  ( .A(data_mem_out_wire[327]), .B(data_mem_out_wire[359]), .S(N29), .Z(\Data_Mem/n6747 ) );
  MUX \Data_Mem/U6754  ( .A(\Data_Mem/n6745 ), .B(\Data_Mem/n6744 ), .S(N28), 
        .Z(\Data_Mem/n6746 ) );
  MUX \Data_Mem/U6753  ( .A(data_mem_out_wire[391]), .B(data_mem_out_wire[423]), .S(N29), .Z(\Data_Mem/n6745 ) );
  MUX \Data_Mem/U6752  ( .A(data_mem_out_wire[455]), .B(data_mem_out_wire[487]), .S(N29), .Z(\Data_Mem/n6744 ) );
  MUX \Data_Mem/U6751  ( .A(\Data_Mem/n6742 ), .B(\Data_Mem/n6735 ), .S(N26), 
        .Z(\Data_Mem/n6743 ) );
  MUX \Data_Mem/U6750  ( .A(\Data_Mem/n6741 ), .B(\Data_Mem/n6738 ), .S(N27), 
        .Z(\Data_Mem/n6742 ) );
  MUX \Data_Mem/U6749  ( .A(\Data_Mem/n6740 ), .B(\Data_Mem/n6739 ), .S(N28), 
        .Z(\Data_Mem/n6741 ) );
  MUX \Data_Mem/U6748  ( .A(data_mem_out_wire[519]), .B(data_mem_out_wire[551]), .S(N29), .Z(\Data_Mem/n6740 ) );
  MUX \Data_Mem/U6747  ( .A(data_mem_out_wire[583]), .B(data_mem_out_wire[615]), .S(N29), .Z(\Data_Mem/n6739 ) );
  MUX \Data_Mem/U6746  ( .A(\Data_Mem/n6737 ), .B(\Data_Mem/n6736 ), .S(N28), 
        .Z(\Data_Mem/n6738 ) );
  MUX \Data_Mem/U6745  ( .A(data_mem_out_wire[647]), .B(data_mem_out_wire[679]), .S(N29), .Z(\Data_Mem/n6737 ) );
  MUX \Data_Mem/U6744  ( .A(data_mem_out_wire[711]), .B(data_mem_out_wire[743]), .S(N29), .Z(\Data_Mem/n6736 ) );
  MUX \Data_Mem/U6743  ( .A(\Data_Mem/n6734 ), .B(\Data_Mem/n6731 ), .S(N27), 
        .Z(\Data_Mem/n6735 ) );
  MUX \Data_Mem/U6742  ( .A(\Data_Mem/n6733 ), .B(\Data_Mem/n6732 ), .S(N28), 
        .Z(\Data_Mem/n6734 ) );
  MUX \Data_Mem/U6741  ( .A(data_mem_out_wire[775]), .B(data_mem_out_wire[807]), .S(N29), .Z(\Data_Mem/n6733 ) );
  MUX \Data_Mem/U6740  ( .A(data_mem_out_wire[839]), .B(data_mem_out_wire[871]), .S(N29), .Z(\Data_Mem/n6732 ) );
  MUX \Data_Mem/U6739  ( .A(\Data_Mem/n6730 ), .B(\Data_Mem/n6729 ), .S(N28), 
        .Z(\Data_Mem/n6731 ) );
  MUX \Data_Mem/U6738  ( .A(data_mem_out_wire[903]), .B(data_mem_out_wire[935]), .S(N29), .Z(\Data_Mem/n6730 ) );
  MUX \Data_Mem/U6737  ( .A(data_mem_out_wire[967]), .B(data_mem_out_wire[999]), .S(N29), .Z(\Data_Mem/n6729 ) );
  MUX \Data_Mem/U6736  ( .A(\Data_Mem/n6727 ), .B(\Data_Mem/n6712 ), .S(N25), 
        .Z(\Data_Mem/n6728 ) );
  MUX \Data_Mem/U6735  ( .A(\Data_Mem/n6726 ), .B(\Data_Mem/n6719 ), .S(N26), 
        .Z(\Data_Mem/n6727 ) );
  MUX \Data_Mem/U6734  ( .A(\Data_Mem/n6725 ), .B(\Data_Mem/n6722 ), .S(N27), 
        .Z(\Data_Mem/n6726 ) );
  MUX \Data_Mem/U6733  ( .A(\Data_Mem/n6724 ), .B(\Data_Mem/n6723 ), .S(N28), 
        .Z(\Data_Mem/n6725 ) );
  MUX \Data_Mem/U6732  ( .A(data_mem_out_wire[1031]), .B(
        data_mem_out_wire[1063]), .S(N29), .Z(\Data_Mem/n6724 ) );
  MUX \Data_Mem/U6731  ( .A(data_mem_out_wire[1095]), .B(
        data_mem_out_wire[1127]), .S(N29), .Z(\Data_Mem/n6723 ) );
  MUX \Data_Mem/U6730  ( .A(\Data_Mem/n6721 ), .B(\Data_Mem/n6720 ), .S(N28), 
        .Z(\Data_Mem/n6722 ) );
  MUX \Data_Mem/U6729  ( .A(data_mem_out_wire[1159]), .B(
        data_mem_out_wire[1191]), .S(N29), .Z(\Data_Mem/n6721 ) );
  MUX \Data_Mem/U6728  ( .A(data_mem_out_wire[1223]), .B(
        data_mem_out_wire[1255]), .S(N29), .Z(\Data_Mem/n6720 ) );
  MUX \Data_Mem/U6727  ( .A(\Data_Mem/n6718 ), .B(\Data_Mem/n6715 ), .S(N27), 
        .Z(\Data_Mem/n6719 ) );
  MUX \Data_Mem/U6726  ( .A(\Data_Mem/n6717 ), .B(\Data_Mem/n6716 ), .S(N28), 
        .Z(\Data_Mem/n6718 ) );
  MUX \Data_Mem/U6725  ( .A(data_mem_out_wire[1287]), .B(
        data_mem_out_wire[1319]), .S(N29), .Z(\Data_Mem/n6717 ) );
  MUX \Data_Mem/U6724  ( .A(data_mem_out_wire[1351]), .B(
        data_mem_out_wire[1383]), .S(N29), .Z(\Data_Mem/n6716 ) );
  MUX \Data_Mem/U6723  ( .A(\Data_Mem/n6714 ), .B(\Data_Mem/n6713 ), .S(N28), 
        .Z(\Data_Mem/n6715 ) );
  MUX \Data_Mem/U6722  ( .A(data_mem_out_wire[1415]), .B(
        data_mem_out_wire[1447]), .S(N29), .Z(\Data_Mem/n6714 ) );
  MUX \Data_Mem/U6721  ( .A(data_mem_out_wire[1479]), .B(
        data_mem_out_wire[1511]), .S(N29), .Z(\Data_Mem/n6713 ) );
  MUX \Data_Mem/U6720  ( .A(\Data_Mem/n6711 ), .B(\Data_Mem/n6704 ), .S(N26), 
        .Z(\Data_Mem/n6712 ) );
  MUX \Data_Mem/U6719  ( .A(\Data_Mem/n6710 ), .B(\Data_Mem/n6707 ), .S(N27), 
        .Z(\Data_Mem/n6711 ) );
  MUX \Data_Mem/U6718  ( .A(\Data_Mem/n6709 ), .B(\Data_Mem/n6708 ), .S(N28), 
        .Z(\Data_Mem/n6710 ) );
  MUX \Data_Mem/U6717  ( .A(data_mem_out_wire[1543]), .B(
        data_mem_out_wire[1575]), .S(N29), .Z(\Data_Mem/n6709 ) );
  MUX \Data_Mem/U6716  ( .A(data_mem_out_wire[1607]), .B(
        data_mem_out_wire[1639]), .S(N29), .Z(\Data_Mem/n6708 ) );
  MUX \Data_Mem/U6715  ( .A(\Data_Mem/n6706 ), .B(\Data_Mem/n6705 ), .S(N28), 
        .Z(\Data_Mem/n6707 ) );
  MUX \Data_Mem/U6714  ( .A(data_mem_out_wire[1671]), .B(
        data_mem_out_wire[1703]), .S(N29), .Z(\Data_Mem/n6706 ) );
  MUX \Data_Mem/U6713  ( .A(data_mem_out_wire[1735]), .B(
        data_mem_out_wire[1767]), .S(N29), .Z(\Data_Mem/n6705 ) );
  MUX \Data_Mem/U6712  ( .A(\Data_Mem/n6703 ), .B(\Data_Mem/n6700 ), .S(N27), 
        .Z(\Data_Mem/n6704 ) );
  MUX \Data_Mem/U6711  ( .A(\Data_Mem/n6702 ), .B(\Data_Mem/n6701 ), .S(N28), 
        .Z(\Data_Mem/n6703 ) );
  MUX \Data_Mem/U6710  ( .A(data_mem_out_wire[1799]), .B(
        data_mem_out_wire[1831]), .S(N29), .Z(\Data_Mem/n6702 ) );
  MUX \Data_Mem/U6709  ( .A(data_mem_out_wire[1863]), .B(
        data_mem_out_wire[1895]), .S(N29), .Z(\Data_Mem/n6701 ) );
  MUX \Data_Mem/U6708  ( .A(\Data_Mem/n6699 ), .B(\Data_Mem/n6698 ), .S(N28), 
        .Z(\Data_Mem/n6700 ) );
  MUX \Data_Mem/U6707  ( .A(data_mem_out_wire[1927]), .B(
        data_mem_out_wire[1959]), .S(N29), .Z(\Data_Mem/n6699 ) );
  MUX \Data_Mem/U6706  ( .A(data_mem_out_wire[1991]), .B(
        data_mem_out_wire[2023]), .S(N29), .Z(\Data_Mem/n6698 ) );
  MUX \Data_Mem/U6705  ( .A(\Data_Mem/n6697 ), .B(\Data_Mem/n6666 ), .S(N24), 
        .Z(c_memory[6]) );
  MUX \Data_Mem/U6704  ( .A(\Data_Mem/n6696 ), .B(\Data_Mem/n6681 ), .S(N25), 
        .Z(\Data_Mem/n6697 ) );
  MUX \Data_Mem/U6703  ( .A(\Data_Mem/n6695 ), .B(\Data_Mem/n6688 ), .S(N26), 
        .Z(\Data_Mem/n6696 ) );
  MUX \Data_Mem/U6702  ( .A(\Data_Mem/n6694 ), .B(\Data_Mem/n6691 ), .S(N27), 
        .Z(\Data_Mem/n6695 ) );
  MUX \Data_Mem/U6701  ( .A(\Data_Mem/n6693 ), .B(\Data_Mem/n6692 ), .S(N28), 
        .Z(\Data_Mem/n6694 ) );
  MUX \Data_Mem/U6700  ( .A(data_mem_out_wire[6]), .B(data_mem_out_wire[38]), 
        .S(N29), .Z(\Data_Mem/n6693 ) );
  MUX \Data_Mem/U6699  ( .A(data_mem_out_wire[70]), .B(data_mem_out_wire[102]), 
        .S(N29), .Z(\Data_Mem/n6692 ) );
  MUX \Data_Mem/U6698  ( .A(\Data_Mem/n6690 ), .B(\Data_Mem/n6689 ), .S(N28), 
        .Z(\Data_Mem/n6691 ) );
  MUX \Data_Mem/U6697  ( .A(data_mem_out_wire[134]), .B(data_mem_out_wire[166]), .S(N29), .Z(\Data_Mem/n6690 ) );
  MUX \Data_Mem/U6696  ( .A(data_mem_out_wire[198]), .B(data_mem_out_wire[230]), .S(N29), .Z(\Data_Mem/n6689 ) );
  MUX \Data_Mem/U6695  ( .A(\Data_Mem/n6687 ), .B(\Data_Mem/n6684 ), .S(N27), 
        .Z(\Data_Mem/n6688 ) );
  MUX \Data_Mem/U6694  ( .A(\Data_Mem/n6686 ), .B(\Data_Mem/n6685 ), .S(N28), 
        .Z(\Data_Mem/n6687 ) );
  MUX \Data_Mem/U6693  ( .A(data_mem_out_wire[262]), .B(data_mem_out_wire[294]), .S(N29), .Z(\Data_Mem/n6686 ) );
  MUX \Data_Mem/U6692  ( .A(data_mem_out_wire[326]), .B(data_mem_out_wire[358]), .S(N29), .Z(\Data_Mem/n6685 ) );
  MUX \Data_Mem/U6691  ( .A(\Data_Mem/n6683 ), .B(\Data_Mem/n6682 ), .S(N28), 
        .Z(\Data_Mem/n6684 ) );
  MUX \Data_Mem/U6690  ( .A(data_mem_out_wire[390]), .B(data_mem_out_wire[422]), .S(N29), .Z(\Data_Mem/n6683 ) );
  MUX \Data_Mem/U6689  ( .A(data_mem_out_wire[454]), .B(data_mem_out_wire[486]), .S(N29), .Z(\Data_Mem/n6682 ) );
  MUX \Data_Mem/U6688  ( .A(\Data_Mem/n6680 ), .B(\Data_Mem/n6673 ), .S(N26), 
        .Z(\Data_Mem/n6681 ) );
  MUX \Data_Mem/U6687  ( .A(\Data_Mem/n6679 ), .B(\Data_Mem/n6676 ), .S(N27), 
        .Z(\Data_Mem/n6680 ) );
  MUX \Data_Mem/U6686  ( .A(\Data_Mem/n6678 ), .B(\Data_Mem/n6677 ), .S(N28), 
        .Z(\Data_Mem/n6679 ) );
  MUX \Data_Mem/U6685  ( .A(data_mem_out_wire[518]), .B(data_mem_out_wire[550]), .S(N29), .Z(\Data_Mem/n6678 ) );
  MUX \Data_Mem/U6684  ( .A(data_mem_out_wire[582]), .B(data_mem_out_wire[614]), .S(N29), .Z(\Data_Mem/n6677 ) );
  MUX \Data_Mem/U6683  ( .A(\Data_Mem/n6675 ), .B(\Data_Mem/n6674 ), .S(N28), 
        .Z(\Data_Mem/n6676 ) );
  MUX \Data_Mem/U6682  ( .A(data_mem_out_wire[646]), .B(data_mem_out_wire[678]), .S(N29), .Z(\Data_Mem/n6675 ) );
  MUX \Data_Mem/U6681  ( .A(data_mem_out_wire[710]), .B(data_mem_out_wire[742]), .S(N29), .Z(\Data_Mem/n6674 ) );
  MUX \Data_Mem/U6680  ( .A(\Data_Mem/n6672 ), .B(\Data_Mem/n6669 ), .S(N27), 
        .Z(\Data_Mem/n6673 ) );
  MUX \Data_Mem/U6679  ( .A(\Data_Mem/n6671 ), .B(\Data_Mem/n6670 ), .S(N28), 
        .Z(\Data_Mem/n6672 ) );
  MUX \Data_Mem/U6678  ( .A(data_mem_out_wire[774]), .B(data_mem_out_wire[806]), .S(N29), .Z(\Data_Mem/n6671 ) );
  MUX \Data_Mem/U6677  ( .A(data_mem_out_wire[838]), .B(data_mem_out_wire[870]), .S(N29), .Z(\Data_Mem/n6670 ) );
  MUX \Data_Mem/U6676  ( .A(\Data_Mem/n6668 ), .B(\Data_Mem/n6667 ), .S(N28), 
        .Z(\Data_Mem/n6669 ) );
  MUX \Data_Mem/U6675  ( .A(data_mem_out_wire[902]), .B(data_mem_out_wire[934]), .S(N29), .Z(\Data_Mem/n6668 ) );
  MUX \Data_Mem/U6674  ( .A(data_mem_out_wire[966]), .B(data_mem_out_wire[998]), .S(N29), .Z(\Data_Mem/n6667 ) );
  MUX \Data_Mem/U6673  ( .A(\Data_Mem/n6665 ), .B(\Data_Mem/n6650 ), .S(N25), 
        .Z(\Data_Mem/n6666 ) );
  MUX \Data_Mem/U6672  ( .A(\Data_Mem/n6664 ), .B(\Data_Mem/n6657 ), .S(N26), 
        .Z(\Data_Mem/n6665 ) );
  MUX \Data_Mem/U6671  ( .A(\Data_Mem/n6663 ), .B(\Data_Mem/n6660 ), .S(N27), 
        .Z(\Data_Mem/n6664 ) );
  MUX \Data_Mem/U6670  ( .A(\Data_Mem/n6662 ), .B(\Data_Mem/n6661 ), .S(N28), 
        .Z(\Data_Mem/n6663 ) );
  MUX \Data_Mem/U6669  ( .A(data_mem_out_wire[1030]), .B(
        data_mem_out_wire[1062]), .S(N29), .Z(\Data_Mem/n6662 ) );
  MUX \Data_Mem/U6668  ( .A(data_mem_out_wire[1094]), .B(
        data_mem_out_wire[1126]), .S(N29), .Z(\Data_Mem/n6661 ) );
  MUX \Data_Mem/U6667  ( .A(\Data_Mem/n6659 ), .B(\Data_Mem/n6658 ), .S(N28), 
        .Z(\Data_Mem/n6660 ) );
  MUX \Data_Mem/U6666  ( .A(data_mem_out_wire[1158]), .B(
        data_mem_out_wire[1190]), .S(N29), .Z(\Data_Mem/n6659 ) );
  MUX \Data_Mem/U6665  ( .A(data_mem_out_wire[1222]), .B(
        data_mem_out_wire[1254]), .S(N29), .Z(\Data_Mem/n6658 ) );
  MUX \Data_Mem/U6664  ( .A(\Data_Mem/n6656 ), .B(\Data_Mem/n6653 ), .S(N27), 
        .Z(\Data_Mem/n6657 ) );
  MUX \Data_Mem/U6663  ( .A(\Data_Mem/n6655 ), .B(\Data_Mem/n6654 ), .S(N28), 
        .Z(\Data_Mem/n6656 ) );
  MUX \Data_Mem/U6662  ( .A(data_mem_out_wire[1286]), .B(
        data_mem_out_wire[1318]), .S(N29), .Z(\Data_Mem/n6655 ) );
  MUX \Data_Mem/U6661  ( .A(data_mem_out_wire[1350]), .B(
        data_mem_out_wire[1382]), .S(N29), .Z(\Data_Mem/n6654 ) );
  MUX \Data_Mem/U6660  ( .A(\Data_Mem/n6652 ), .B(\Data_Mem/n6651 ), .S(N28), 
        .Z(\Data_Mem/n6653 ) );
  MUX \Data_Mem/U6659  ( .A(data_mem_out_wire[1414]), .B(
        data_mem_out_wire[1446]), .S(N29), .Z(\Data_Mem/n6652 ) );
  MUX \Data_Mem/U6658  ( .A(data_mem_out_wire[1478]), .B(
        data_mem_out_wire[1510]), .S(N29), .Z(\Data_Mem/n6651 ) );
  MUX \Data_Mem/U6657  ( .A(\Data_Mem/n6649 ), .B(\Data_Mem/n6642 ), .S(N26), 
        .Z(\Data_Mem/n6650 ) );
  MUX \Data_Mem/U6656  ( .A(\Data_Mem/n6648 ), .B(\Data_Mem/n6645 ), .S(N27), 
        .Z(\Data_Mem/n6649 ) );
  MUX \Data_Mem/U6655  ( .A(\Data_Mem/n6647 ), .B(\Data_Mem/n6646 ), .S(N28), 
        .Z(\Data_Mem/n6648 ) );
  MUX \Data_Mem/U6654  ( .A(data_mem_out_wire[1542]), .B(
        data_mem_out_wire[1574]), .S(N29), .Z(\Data_Mem/n6647 ) );
  MUX \Data_Mem/U6653  ( .A(data_mem_out_wire[1606]), .B(
        data_mem_out_wire[1638]), .S(N29), .Z(\Data_Mem/n6646 ) );
  MUX \Data_Mem/U6652  ( .A(\Data_Mem/n6644 ), .B(\Data_Mem/n6643 ), .S(N28), 
        .Z(\Data_Mem/n6645 ) );
  MUX \Data_Mem/U6651  ( .A(data_mem_out_wire[1670]), .B(
        data_mem_out_wire[1702]), .S(N29), .Z(\Data_Mem/n6644 ) );
  MUX \Data_Mem/U6650  ( .A(data_mem_out_wire[1734]), .B(
        data_mem_out_wire[1766]), .S(N29), .Z(\Data_Mem/n6643 ) );
  MUX \Data_Mem/U6649  ( .A(\Data_Mem/n6641 ), .B(\Data_Mem/n6638 ), .S(N27), 
        .Z(\Data_Mem/n6642 ) );
  MUX \Data_Mem/U6648  ( .A(\Data_Mem/n6640 ), .B(\Data_Mem/n6639 ), .S(N28), 
        .Z(\Data_Mem/n6641 ) );
  MUX \Data_Mem/U6647  ( .A(data_mem_out_wire[1798]), .B(
        data_mem_out_wire[1830]), .S(N29), .Z(\Data_Mem/n6640 ) );
  MUX \Data_Mem/U6646  ( .A(data_mem_out_wire[1862]), .B(
        data_mem_out_wire[1894]), .S(N29), .Z(\Data_Mem/n6639 ) );
  MUX \Data_Mem/U6645  ( .A(\Data_Mem/n6637 ), .B(\Data_Mem/n6636 ), .S(N28), 
        .Z(\Data_Mem/n6638 ) );
  MUX \Data_Mem/U6644  ( .A(data_mem_out_wire[1926]), .B(
        data_mem_out_wire[1958]), .S(N29), .Z(\Data_Mem/n6637 ) );
  MUX \Data_Mem/U6643  ( .A(data_mem_out_wire[1990]), .B(
        data_mem_out_wire[2022]), .S(N29), .Z(\Data_Mem/n6636 ) );
  MUX \Data_Mem/U6642  ( .A(\Data_Mem/n6635 ), .B(\Data_Mem/n6604 ), .S(N24), 
        .Z(c_memory[5]) );
  MUX \Data_Mem/U6641  ( .A(\Data_Mem/n6634 ), .B(\Data_Mem/n6619 ), .S(N25), 
        .Z(\Data_Mem/n6635 ) );
  MUX \Data_Mem/U6640  ( .A(\Data_Mem/n6633 ), .B(\Data_Mem/n6626 ), .S(N26), 
        .Z(\Data_Mem/n6634 ) );
  MUX \Data_Mem/U6639  ( .A(\Data_Mem/n6632 ), .B(\Data_Mem/n6629 ), .S(N27), 
        .Z(\Data_Mem/n6633 ) );
  MUX \Data_Mem/U6638  ( .A(\Data_Mem/n6631 ), .B(\Data_Mem/n6630 ), .S(N28), 
        .Z(\Data_Mem/n6632 ) );
  MUX \Data_Mem/U6637  ( .A(data_mem_out_wire[5]), .B(data_mem_out_wire[37]), 
        .S(N29), .Z(\Data_Mem/n6631 ) );
  MUX \Data_Mem/U6636  ( .A(data_mem_out_wire[69]), .B(data_mem_out_wire[101]), 
        .S(N29), .Z(\Data_Mem/n6630 ) );
  MUX \Data_Mem/U6635  ( .A(\Data_Mem/n6628 ), .B(\Data_Mem/n6627 ), .S(N28), 
        .Z(\Data_Mem/n6629 ) );
  MUX \Data_Mem/U6634  ( .A(data_mem_out_wire[133]), .B(data_mem_out_wire[165]), .S(N29), .Z(\Data_Mem/n6628 ) );
  MUX \Data_Mem/U6633  ( .A(data_mem_out_wire[197]), .B(data_mem_out_wire[229]), .S(N29), .Z(\Data_Mem/n6627 ) );
  MUX \Data_Mem/U6632  ( .A(\Data_Mem/n6625 ), .B(\Data_Mem/n6622 ), .S(N27), 
        .Z(\Data_Mem/n6626 ) );
  MUX \Data_Mem/U6631  ( .A(\Data_Mem/n6624 ), .B(\Data_Mem/n6623 ), .S(N28), 
        .Z(\Data_Mem/n6625 ) );
  MUX \Data_Mem/U6630  ( .A(data_mem_out_wire[261]), .B(data_mem_out_wire[293]), .S(N29), .Z(\Data_Mem/n6624 ) );
  MUX \Data_Mem/U6629  ( .A(data_mem_out_wire[325]), .B(data_mem_out_wire[357]), .S(N29), .Z(\Data_Mem/n6623 ) );
  MUX \Data_Mem/U6628  ( .A(\Data_Mem/n6621 ), .B(\Data_Mem/n6620 ), .S(N28), 
        .Z(\Data_Mem/n6622 ) );
  MUX \Data_Mem/U6627  ( .A(data_mem_out_wire[389]), .B(data_mem_out_wire[421]), .S(N29), .Z(\Data_Mem/n6621 ) );
  MUX \Data_Mem/U6626  ( .A(data_mem_out_wire[453]), .B(data_mem_out_wire[485]), .S(N29), .Z(\Data_Mem/n6620 ) );
  MUX \Data_Mem/U6625  ( .A(\Data_Mem/n6618 ), .B(\Data_Mem/n6611 ), .S(N26), 
        .Z(\Data_Mem/n6619 ) );
  MUX \Data_Mem/U6624  ( .A(\Data_Mem/n6617 ), .B(\Data_Mem/n6614 ), .S(N27), 
        .Z(\Data_Mem/n6618 ) );
  MUX \Data_Mem/U6623  ( .A(\Data_Mem/n6616 ), .B(\Data_Mem/n6615 ), .S(N28), 
        .Z(\Data_Mem/n6617 ) );
  MUX \Data_Mem/U6622  ( .A(data_mem_out_wire[517]), .B(data_mem_out_wire[549]), .S(N29), .Z(\Data_Mem/n6616 ) );
  MUX \Data_Mem/U6621  ( .A(data_mem_out_wire[581]), .B(data_mem_out_wire[613]), .S(N29), .Z(\Data_Mem/n6615 ) );
  MUX \Data_Mem/U6620  ( .A(\Data_Mem/n6613 ), .B(\Data_Mem/n6612 ), .S(N28), 
        .Z(\Data_Mem/n6614 ) );
  MUX \Data_Mem/U6619  ( .A(data_mem_out_wire[645]), .B(data_mem_out_wire[677]), .S(N29), .Z(\Data_Mem/n6613 ) );
  MUX \Data_Mem/U6618  ( .A(data_mem_out_wire[709]), .B(data_mem_out_wire[741]), .S(N29), .Z(\Data_Mem/n6612 ) );
  MUX \Data_Mem/U6617  ( .A(\Data_Mem/n6610 ), .B(\Data_Mem/n6607 ), .S(N27), 
        .Z(\Data_Mem/n6611 ) );
  MUX \Data_Mem/U6616  ( .A(\Data_Mem/n6609 ), .B(\Data_Mem/n6608 ), .S(N28), 
        .Z(\Data_Mem/n6610 ) );
  MUX \Data_Mem/U6615  ( .A(data_mem_out_wire[773]), .B(data_mem_out_wire[805]), .S(N29), .Z(\Data_Mem/n6609 ) );
  MUX \Data_Mem/U6614  ( .A(data_mem_out_wire[837]), .B(data_mem_out_wire[869]), .S(N29), .Z(\Data_Mem/n6608 ) );
  MUX \Data_Mem/U6613  ( .A(\Data_Mem/n6606 ), .B(\Data_Mem/n6605 ), .S(N28), 
        .Z(\Data_Mem/n6607 ) );
  MUX \Data_Mem/U6612  ( .A(data_mem_out_wire[901]), .B(data_mem_out_wire[933]), .S(N29), .Z(\Data_Mem/n6606 ) );
  MUX \Data_Mem/U6611  ( .A(data_mem_out_wire[965]), .B(data_mem_out_wire[997]), .S(N29), .Z(\Data_Mem/n6605 ) );
  MUX \Data_Mem/U6610  ( .A(\Data_Mem/n6603 ), .B(\Data_Mem/n6588 ), .S(N25), 
        .Z(\Data_Mem/n6604 ) );
  MUX \Data_Mem/U6609  ( .A(\Data_Mem/n6602 ), .B(\Data_Mem/n6595 ), .S(N26), 
        .Z(\Data_Mem/n6603 ) );
  MUX \Data_Mem/U6608  ( .A(\Data_Mem/n6601 ), .B(\Data_Mem/n6598 ), .S(N27), 
        .Z(\Data_Mem/n6602 ) );
  MUX \Data_Mem/U6607  ( .A(\Data_Mem/n6600 ), .B(\Data_Mem/n6599 ), .S(N28), 
        .Z(\Data_Mem/n6601 ) );
  MUX \Data_Mem/U6606  ( .A(data_mem_out_wire[1029]), .B(
        data_mem_out_wire[1061]), .S(N29), .Z(\Data_Mem/n6600 ) );
  MUX \Data_Mem/U6605  ( .A(data_mem_out_wire[1093]), .B(
        data_mem_out_wire[1125]), .S(N29), .Z(\Data_Mem/n6599 ) );
  MUX \Data_Mem/U6604  ( .A(\Data_Mem/n6597 ), .B(\Data_Mem/n6596 ), .S(N28), 
        .Z(\Data_Mem/n6598 ) );
  MUX \Data_Mem/U6603  ( .A(data_mem_out_wire[1157]), .B(
        data_mem_out_wire[1189]), .S(N29), .Z(\Data_Mem/n6597 ) );
  MUX \Data_Mem/U6602  ( .A(data_mem_out_wire[1221]), .B(
        data_mem_out_wire[1253]), .S(N29), .Z(\Data_Mem/n6596 ) );
  MUX \Data_Mem/U6601  ( .A(\Data_Mem/n6594 ), .B(\Data_Mem/n6591 ), .S(N27), 
        .Z(\Data_Mem/n6595 ) );
  MUX \Data_Mem/U6600  ( .A(\Data_Mem/n6593 ), .B(\Data_Mem/n6592 ), .S(N28), 
        .Z(\Data_Mem/n6594 ) );
  MUX \Data_Mem/U6599  ( .A(data_mem_out_wire[1285]), .B(
        data_mem_out_wire[1317]), .S(N29), .Z(\Data_Mem/n6593 ) );
  MUX \Data_Mem/U6598  ( .A(data_mem_out_wire[1349]), .B(
        data_mem_out_wire[1381]), .S(N29), .Z(\Data_Mem/n6592 ) );
  MUX \Data_Mem/U6597  ( .A(\Data_Mem/n6590 ), .B(\Data_Mem/n6589 ), .S(N28), 
        .Z(\Data_Mem/n6591 ) );
  MUX \Data_Mem/U6596  ( .A(data_mem_out_wire[1413]), .B(
        data_mem_out_wire[1445]), .S(N29), .Z(\Data_Mem/n6590 ) );
  MUX \Data_Mem/U6595  ( .A(data_mem_out_wire[1477]), .B(
        data_mem_out_wire[1509]), .S(N29), .Z(\Data_Mem/n6589 ) );
  MUX \Data_Mem/U6594  ( .A(\Data_Mem/n6587 ), .B(\Data_Mem/n6580 ), .S(N26), 
        .Z(\Data_Mem/n6588 ) );
  MUX \Data_Mem/U6593  ( .A(\Data_Mem/n6586 ), .B(\Data_Mem/n6583 ), .S(N27), 
        .Z(\Data_Mem/n6587 ) );
  MUX \Data_Mem/U6592  ( .A(\Data_Mem/n6585 ), .B(\Data_Mem/n6584 ), .S(N28), 
        .Z(\Data_Mem/n6586 ) );
  MUX \Data_Mem/U6591  ( .A(data_mem_out_wire[1541]), .B(
        data_mem_out_wire[1573]), .S(N29), .Z(\Data_Mem/n6585 ) );
  MUX \Data_Mem/U6590  ( .A(data_mem_out_wire[1605]), .B(
        data_mem_out_wire[1637]), .S(N29), .Z(\Data_Mem/n6584 ) );
  MUX \Data_Mem/U6589  ( .A(\Data_Mem/n6582 ), .B(\Data_Mem/n6581 ), .S(N28), 
        .Z(\Data_Mem/n6583 ) );
  MUX \Data_Mem/U6588  ( .A(data_mem_out_wire[1669]), .B(
        data_mem_out_wire[1701]), .S(N29), .Z(\Data_Mem/n6582 ) );
  MUX \Data_Mem/U6587  ( .A(data_mem_out_wire[1733]), .B(
        data_mem_out_wire[1765]), .S(N29), .Z(\Data_Mem/n6581 ) );
  MUX \Data_Mem/U6586  ( .A(\Data_Mem/n6579 ), .B(\Data_Mem/n6576 ), .S(N27), 
        .Z(\Data_Mem/n6580 ) );
  MUX \Data_Mem/U6585  ( .A(\Data_Mem/n6578 ), .B(\Data_Mem/n6577 ), .S(N28), 
        .Z(\Data_Mem/n6579 ) );
  MUX \Data_Mem/U6584  ( .A(data_mem_out_wire[1797]), .B(
        data_mem_out_wire[1829]), .S(N29), .Z(\Data_Mem/n6578 ) );
  MUX \Data_Mem/U6583  ( .A(data_mem_out_wire[1861]), .B(
        data_mem_out_wire[1893]), .S(N29), .Z(\Data_Mem/n6577 ) );
  MUX \Data_Mem/U6582  ( .A(\Data_Mem/n6575 ), .B(\Data_Mem/n6574 ), .S(N28), 
        .Z(\Data_Mem/n6576 ) );
  MUX \Data_Mem/U6581  ( .A(data_mem_out_wire[1925]), .B(
        data_mem_out_wire[1957]), .S(N29), .Z(\Data_Mem/n6575 ) );
  MUX \Data_Mem/U6580  ( .A(data_mem_out_wire[1989]), .B(
        data_mem_out_wire[2021]), .S(N29), .Z(\Data_Mem/n6574 ) );
  MUX \Data_Mem/U6579  ( .A(\Data_Mem/n6573 ), .B(\Data_Mem/n6542 ), .S(N24), 
        .Z(c_memory[4]) );
  MUX \Data_Mem/U6578  ( .A(\Data_Mem/n6572 ), .B(\Data_Mem/n6557 ), .S(N25), 
        .Z(\Data_Mem/n6573 ) );
  MUX \Data_Mem/U6577  ( .A(\Data_Mem/n6571 ), .B(\Data_Mem/n6564 ), .S(N26), 
        .Z(\Data_Mem/n6572 ) );
  MUX \Data_Mem/U6576  ( .A(\Data_Mem/n6570 ), .B(\Data_Mem/n6567 ), .S(N27), 
        .Z(\Data_Mem/n6571 ) );
  MUX \Data_Mem/U6575  ( .A(\Data_Mem/n6569 ), .B(\Data_Mem/n6568 ), .S(N28), 
        .Z(\Data_Mem/n6570 ) );
  MUX \Data_Mem/U6574  ( .A(data_mem_out_wire[4]), .B(data_mem_out_wire[36]), 
        .S(N29), .Z(\Data_Mem/n6569 ) );
  MUX \Data_Mem/U6573  ( .A(data_mem_out_wire[68]), .B(data_mem_out_wire[100]), 
        .S(N29), .Z(\Data_Mem/n6568 ) );
  MUX \Data_Mem/U6572  ( .A(\Data_Mem/n6566 ), .B(\Data_Mem/n6565 ), .S(N28), 
        .Z(\Data_Mem/n6567 ) );
  MUX \Data_Mem/U6571  ( .A(data_mem_out_wire[132]), .B(data_mem_out_wire[164]), .S(N29), .Z(\Data_Mem/n6566 ) );
  MUX \Data_Mem/U6570  ( .A(data_mem_out_wire[196]), .B(data_mem_out_wire[228]), .S(N29), .Z(\Data_Mem/n6565 ) );
  MUX \Data_Mem/U6569  ( .A(\Data_Mem/n6563 ), .B(\Data_Mem/n6560 ), .S(N27), 
        .Z(\Data_Mem/n6564 ) );
  MUX \Data_Mem/U6568  ( .A(\Data_Mem/n6562 ), .B(\Data_Mem/n6561 ), .S(N28), 
        .Z(\Data_Mem/n6563 ) );
  MUX \Data_Mem/U6567  ( .A(data_mem_out_wire[260]), .B(data_mem_out_wire[292]), .S(N29), .Z(\Data_Mem/n6562 ) );
  MUX \Data_Mem/U6566  ( .A(data_mem_out_wire[324]), .B(data_mem_out_wire[356]), .S(N29), .Z(\Data_Mem/n6561 ) );
  MUX \Data_Mem/U6565  ( .A(\Data_Mem/n6559 ), .B(\Data_Mem/n6558 ), .S(N28), 
        .Z(\Data_Mem/n6560 ) );
  MUX \Data_Mem/U6564  ( .A(data_mem_out_wire[388]), .B(data_mem_out_wire[420]), .S(N29), .Z(\Data_Mem/n6559 ) );
  MUX \Data_Mem/U6563  ( .A(data_mem_out_wire[452]), .B(data_mem_out_wire[484]), .S(N29), .Z(\Data_Mem/n6558 ) );
  MUX \Data_Mem/U6562  ( .A(\Data_Mem/n6556 ), .B(\Data_Mem/n6549 ), .S(N26), 
        .Z(\Data_Mem/n6557 ) );
  MUX \Data_Mem/U6561  ( .A(\Data_Mem/n6555 ), .B(\Data_Mem/n6552 ), .S(N27), 
        .Z(\Data_Mem/n6556 ) );
  MUX \Data_Mem/U6560  ( .A(\Data_Mem/n6554 ), .B(\Data_Mem/n6553 ), .S(N28), 
        .Z(\Data_Mem/n6555 ) );
  MUX \Data_Mem/U6559  ( .A(data_mem_out_wire[516]), .B(data_mem_out_wire[548]), .S(N29), .Z(\Data_Mem/n6554 ) );
  MUX \Data_Mem/U6558  ( .A(data_mem_out_wire[580]), .B(data_mem_out_wire[612]), .S(N29), .Z(\Data_Mem/n6553 ) );
  MUX \Data_Mem/U6557  ( .A(\Data_Mem/n6551 ), .B(\Data_Mem/n6550 ), .S(N28), 
        .Z(\Data_Mem/n6552 ) );
  MUX \Data_Mem/U6556  ( .A(data_mem_out_wire[644]), .B(data_mem_out_wire[676]), .S(N29), .Z(\Data_Mem/n6551 ) );
  MUX \Data_Mem/U6555  ( .A(data_mem_out_wire[708]), .B(data_mem_out_wire[740]), .S(N29), .Z(\Data_Mem/n6550 ) );
  MUX \Data_Mem/U6554  ( .A(\Data_Mem/n6548 ), .B(\Data_Mem/n6545 ), .S(N27), 
        .Z(\Data_Mem/n6549 ) );
  MUX \Data_Mem/U6553  ( .A(\Data_Mem/n6547 ), .B(\Data_Mem/n6546 ), .S(N28), 
        .Z(\Data_Mem/n6548 ) );
  MUX \Data_Mem/U6552  ( .A(data_mem_out_wire[772]), .B(data_mem_out_wire[804]), .S(N29), .Z(\Data_Mem/n6547 ) );
  MUX \Data_Mem/U6551  ( .A(data_mem_out_wire[836]), .B(data_mem_out_wire[868]), .S(N29), .Z(\Data_Mem/n6546 ) );
  MUX \Data_Mem/U6550  ( .A(\Data_Mem/n6544 ), .B(\Data_Mem/n6543 ), .S(N28), 
        .Z(\Data_Mem/n6545 ) );
  MUX \Data_Mem/U6549  ( .A(data_mem_out_wire[900]), .B(data_mem_out_wire[932]), .S(N29), .Z(\Data_Mem/n6544 ) );
  MUX \Data_Mem/U6548  ( .A(data_mem_out_wire[964]), .B(data_mem_out_wire[996]), .S(N29), .Z(\Data_Mem/n6543 ) );
  MUX \Data_Mem/U6547  ( .A(\Data_Mem/n6541 ), .B(\Data_Mem/n6526 ), .S(N25), 
        .Z(\Data_Mem/n6542 ) );
  MUX \Data_Mem/U6546  ( .A(\Data_Mem/n6540 ), .B(\Data_Mem/n6533 ), .S(N26), 
        .Z(\Data_Mem/n6541 ) );
  MUX \Data_Mem/U6545  ( .A(\Data_Mem/n6539 ), .B(\Data_Mem/n6536 ), .S(N27), 
        .Z(\Data_Mem/n6540 ) );
  MUX \Data_Mem/U6544  ( .A(\Data_Mem/n6538 ), .B(\Data_Mem/n6537 ), .S(N28), 
        .Z(\Data_Mem/n6539 ) );
  MUX \Data_Mem/U6543  ( .A(data_mem_out_wire[1028]), .B(
        data_mem_out_wire[1060]), .S(N29), .Z(\Data_Mem/n6538 ) );
  MUX \Data_Mem/U6542  ( .A(data_mem_out_wire[1092]), .B(
        data_mem_out_wire[1124]), .S(N29), .Z(\Data_Mem/n6537 ) );
  MUX \Data_Mem/U6541  ( .A(\Data_Mem/n6535 ), .B(\Data_Mem/n6534 ), .S(N28), 
        .Z(\Data_Mem/n6536 ) );
  MUX \Data_Mem/U6540  ( .A(data_mem_out_wire[1156]), .B(
        data_mem_out_wire[1188]), .S(N29), .Z(\Data_Mem/n6535 ) );
  MUX \Data_Mem/U6539  ( .A(data_mem_out_wire[1220]), .B(
        data_mem_out_wire[1252]), .S(N29), .Z(\Data_Mem/n6534 ) );
  MUX \Data_Mem/U6538  ( .A(\Data_Mem/n6532 ), .B(\Data_Mem/n6529 ), .S(N27), 
        .Z(\Data_Mem/n6533 ) );
  MUX \Data_Mem/U6537  ( .A(\Data_Mem/n6531 ), .B(\Data_Mem/n6530 ), .S(N28), 
        .Z(\Data_Mem/n6532 ) );
  MUX \Data_Mem/U6536  ( .A(data_mem_out_wire[1284]), .B(
        data_mem_out_wire[1316]), .S(N29), .Z(\Data_Mem/n6531 ) );
  MUX \Data_Mem/U6535  ( .A(data_mem_out_wire[1348]), .B(
        data_mem_out_wire[1380]), .S(N29), .Z(\Data_Mem/n6530 ) );
  MUX \Data_Mem/U6534  ( .A(\Data_Mem/n6528 ), .B(\Data_Mem/n6527 ), .S(N28), 
        .Z(\Data_Mem/n6529 ) );
  MUX \Data_Mem/U6533  ( .A(data_mem_out_wire[1412]), .B(
        data_mem_out_wire[1444]), .S(N29), .Z(\Data_Mem/n6528 ) );
  MUX \Data_Mem/U6532  ( .A(data_mem_out_wire[1476]), .B(
        data_mem_out_wire[1508]), .S(N29), .Z(\Data_Mem/n6527 ) );
  MUX \Data_Mem/U6531  ( .A(\Data_Mem/n6525 ), .B(\Data_Mem/n6518 ), .S(N26), 
        .Z(\Data_Mem/n6526 ) );
  MUX \Data_Mem/U6530  ( .A(\Data_Mem/n6524 ), .B(\Data_Mem/n6521 ), .S(N27), 
        .Z(\Data_Mem/n6525 ) );
  MUX \Data_Mem/U6529  ( .A(\Data_Mem/n6523 ), .B(\Data_Mem/n6522 ), .S(N28), 
        .Z(\Data_Mem/n6524 ) );
  MUX \Data_Mem/U6528  ( .A(data_mem_out_wire[1540]), .B(
        data_mem_out_wire[1572]), .S(N29), .Z(\Data_Mem/n6523 ) );
  MUX \Data_Mem/U6527  ( .A(data_mem_out_wire[1604]), .B(
        data_mem_out_wire[1636]), .S(N29), .Z(\Data_Mem/n6522 ) );
  MUX \Data_Mem/U6526  ( .A(\Data_Mem/n6520 ), .B(\Data_Mem/n6519 ), .S(N28), 
        .Z(\Data_Mem/n6521 ) );
  MUX \Data_Mem/U6525  ( .A(data_mem_out_wire[1668]), .B(
        data_mem_out_wire[1700]), .S(N29), .Z(\Data_Mem/n6520 ) );
  MUX \Data_Mem/U6524  ( .A(data_mem_out_wire[1732]), .B(
        data_mem_out_wire[1764]), .S(N29), .Z(\Data_Mem/n6519 ) );
  MUX \Data_Mem/U6523  ( .A(\Data_Mem/n6517 ), .B(\Data_Mem/n6514 ), .S(N27), 
        .Z(\Data_Mem/n6518 ) );
  MUX \Data_Mem/U6522  ( .A(\Data_Mem/n6516 ), .B(\Data_Mem/n6515 ), .S(N28), 
        .Z(\Data_Mem/n6517 ) );
  MUX \Data_Mem/U6521  ( .A(data_mem_out_wire[1796]), .B(
        data_mem_out_wire[1828]), .S(N29), .Z(\Data_Mem/n6516 ) );
  MUX \Data_Mem/U6520  ( .A(data_mem_out_wire[1860]), .B(
        data_mem_out_wire[1892]), .S(N29), .Z(\Data_Mem/n6515 ) );
  MUX \Data_Mem/U6519  ( .A(\Data_Mem/n6513 ), .B(\Data_Mem/n6512 ), .S(N28), 
        .Z(\Data_Mem/n6514 ) );
  MUX \Data_Mem/U6518  ( .A(data_mem_out_wire[1924]), .B(
        data_mem_out_wire[1956]), .S(N29), .Z(\Data_Mem/n6513 ) );
  MUX \Data_Mem/U6517  ( .A(data_mem_out_wire[1988]), .B(
        data_mem_out_wire[2020]), .S(N29), .Z(\Data_Mem/n6512 ) );
  MUX \Data_Mem/U6516  ( .A(\Data_Mem/n6511 ), .B(\Data_Mem/n6480 ), .S(N24), 
        .Z(c_memory[3]) );
  MUX \Data_Mem/U6515  ( .A(\Data_Mem/n6510 ), .B(\Data_Mem/n6495 ), .S(N25), 
        .Z(\Data_Mem/n6511 ) );
  MUX \Data_Mem/U6514  ( .A(\Data_Mem/n6509 ), .B(\Data_Mem/n6502 ), .S(N26), 
        .Z(\Data_Mem/n6510 ) );
  MUX \Data_Mem/U6513  ( .A(\Data_Mem/n6508 ), .B(\Data_Mem/n6505 ), .S(N27), 
        .Z(\Data_Mem/n6509 ) );
  MUX \Data_Mem/U6512  ( .A(\Data_Mem/n6507 ), .B(\Data_Mem/n6506 ), .S(N28), 
        .Z(\Data_Mem/n6508 ) );
  MUX \Data_Mem/U6511  ( .A(data_mem_out_wire[3]), .B(data_mem_out_wire[35]), 
        .S(N29), .Z(\Data_Mem/n6507 ) );
  MUX \Data_Mem/U6510  ( .A(data_mem_out_wire[67]), .B(data_mem_out_wire[99]), 
        .S(N29), .Z(\Data_Mem/n6506 ) );
  MUX \Data_Mem/U6509  ( .A(\Data_Mem/n6504 ), .B(\Data_Mem/n6503 ), .S(N28), 
        .Z(\Data_Mem/n6505 ) );
  MUX \Data_Mem/U6508  ( .A(data_mem_out_wire[131]), .B(data_mem_out_wire[163]), .S(N29), .Z(\Data_Mem/n6504 ) );
  MUX \Data_Mem/U6507  ( .A(data_mem_out_wire[195]), .B(data_mem_out_wire[227]), .S(N29), .Z(\Data_Mem/n6503 ) );
  MUX \Data_Mem/U6506  ( .A(\Data_Mem/n6501 ), .B(\Data_Mem/n6498 ), .S(N27), 
        .Z(\Data_Mem/n6502 ) );
  MUX \Data_Mem/U6505  ( .A(\Data_Mem/n6500 ), .B(\Data_Mem/n6499 ), .S(N28), 
        .Z(\Data_Mem/n6501 ) );
  MUX \Data_Mem/U6504  ( .A(data_mem_out_wire[259]), .B(data_mem_out_wire[291]), .S(N29), .Z(\Data_Mem/n6500 ) );
  MUX \Data_Mem/U6503  ( .A(data_mem_out_wire[323]), .B(data_mem_out_wire[355]), .S(N29), .Z(\Data_Mem/n6499 ) );
  MUX \Data_Mem/U6502  ( .A(\Data_Mem/n6497 ), .B(\Data_Mem/n6496 ), .S(N28), 
        .Z(\Data_Mem/n6498 ) );
  MUX \Data_Mem/U6501  ( .A(data_mem_out_wire[387]), .B(data_mem_out_wire[419]), .S(N29), .Z(\Data_Mem/n6497 ) );
  MUX \Data_Mem/U6500  ( .A(data_mem_out_wire[451]), .B(data_mem_out_wire[483]), .S(N29), .Z(\Data_Mem/n6496 ) );
  MUX \Data_Mem/U6499  ( .A(\Data_Mem/n6494 ), .B(\Data_Mem/n6487 ), .S(N26), 
        .Z(\Data_Mem/n6495 ) );
  MUX \Data_Mem/U6498  ( .A(\Data_Mem/n6493 ), .B(\Data_Mem/n6490 ), .S(N27), 
        .Z(\Data_Mem/n6494 ) );
  MUX \Data_Mem/U6497  ( .A(\Data_Mem/n6492 ), .B(\Data_Mem/n6491 ), .S(N28), 
        .Z(\Data_Mem/n6493 ) );
  MUX \Data_Mem/U6496  ( .A(data_mem_out_wire[515]), .B(data_mem_out_wire[547]), .S(N29), .Z(\Data_Mem/n6492 ) );
  MUX \Data_Mem/U6495  ( .A(data_mem_out_wire[579]), .B(data_mem_out_wire[611]), .S(N29), .Z(\Data_Mem/n6491 ) );
  MUX \Data_Mem/U6494  ( .A(\Data_Mem/n6489 ), .B(\Data_Mem/n6488 ), .S(N28), 
        .Z(\Data_Mem/n6490 ) );
  MUX \Data_Mem/U6493  ( .A(data_mem_out_wire[643]), .B(data_mem_out_wire[675]), .S(N29), .Z(\Data_Mem/n6489 ) );
  MUX \Data_Mem/U6492  ( .A(data_mem_out_wire[707]), .B(data_mem_out_wire[739]), .S(N29), .Z(\Data_Mem/n6488 ) );
  MUX \Data_Mem/U6491  ( .A(\Data_Mem/n6486 ), .B(\Data_Mem/n6483 ), .S(N27), 
        .Z(\Data_Mem/n6487 ) );
  MUX \Data_Mem/U6490  ( .A(\Data_Mem/n6485 ), .B(\Data_Mem/n6484 ), .S(N28), 
        .Z(\Data_Mem/n6486 ) );
  MUX \Data_Mem/U6489  ( .A(data_mem_out_wire[771]), .B(data_mem_out_wire[803]), .S(N29), .Z(\Data_Mem/n6485 ) );
  MUX \Data_Mem/U6488  ( .A(data_mem_out_wire[835]), .B(data_mem_out_wire[867]), .S(N29), .Z(\Data_Mem/n6484 ) );
  MUX \Data_Mem/U6487  ( .A(\Data_Mem/n6482 ), .B(\Data_Mem/n6481 ), .S(N28), 
        .Z(\Data_Mem/n6483 ) );
  MUX \Data_Mem/U6486  ( .A(data_mem_out_wire[899]), .B(data_mem_out_wire[931]), .S(N29), .Z(\Data_Mem/n6482 ) );
  MUX \Data_Mem/U6485  ( .A(data_mem_out_wire[963]), .B(data_mem_out_wire[995]), .S(N29), .Z(\Data_Mem/n6481 ) );
  MUX \Data_Mem/U6484  ( .A(\Data_Mem/n6479 ), .B(\Data_Mem/n6464 ), .S(N25), 
        .Z(\Data_Mem/n6480 ) );
  MUX \Data_Mem/U6483  ( .A(\Data_Mem/n6478 ), .B(\Data_Mem/n6471 ), .S(N26), 
        .Z(\Data_Mem/n6479 ) );
  MUX \Data_Mem/U6482  ( .A(\Data_Mem/n6477 ), .B(\Data_Mem/n6474 ), .S(N27), 
        .Z(\Data_Mem/n6478 ) );
  MUX \Data_Mem/U6481  ( .A(\Data_Mem/n6476 ), .B(\Data_Mem/n6475 ), .S(N28), 
        .Z(\Data_Mem/n6477 ) );
  MUX \Data_Mem/U6480  ( .A(data_mem_out_wire[1027]), .B(
        data_mem_out_wire[1059]), .S(N29), .Z(\Data_Mem/n6476 ) );
  MUX \Data_Mem/U6479  ( .A(data_mem_out_wire[1091]), .B(
        data_mem_out_wire[1123]), .S(N29), .Z(\Data_Mem/n6475 ) );
  MUX \Data_Mem/U6478  ( .A(\Data_Mem/n6473 ), .B(\Data_Mem/n6472 ), .S(N28), 
        .Z(\Data_Mem/n6474 ) );
  MUX \Data_Mem/U6477  ( .A(data_mem_out_wire[1155]), .B(
        data_mem_out_wire[1187]), .S(N29), .Z(\Data_Mem/n6473 ) );
  MUX \Data_Mem/U6476  ( .A(data_mem_out_wire[1219]), .B(
        data_mem_out_wire[1251]), .S(N29), .Z(\Data_Mem/n6472 ) );
  MUX \Data_Mem/U6475  ( .A(\Data_Mem/n6470 ), .B(\Data_Mem/n6467 ), .S(N27), 
        .Z(\Data_Mem/n6471 ) );
  MUX \Data_Mem/U6474  ( .A(\Data_Mem/n6469 ), .B(\Data_Mem/n6468 ), .S(N28), 
        .Z(\Data_Mem/n6470 ) );
  MUX \Data_Mem/U6473  ( .A(data_mem_out_wire[1283]), .B(
        data_mem_out_wire[1315]), .S(N29), .Z(\Data_Mem/n6469 ) );
  MUX \Data_Mem/U6472  ( .A(data_mem_out_wire[1347]), .B(
        data_mem_out_wire[1379]), .S(N29), .Z(\Data_Mem/n6468 ) );
  MUX \Data_Mem/U6471  ( .A(\Data_Mem/n6466 ), .B(\Data_Mem/n6465 ), .S(N28), 
        .Z(\Data_Mem/n6467 ) );
  MUX \Data_Mem/U6470  ( .A(data_mem_out_wire[1411]), .B(
        data_mem_out_wire[1443]), .S(N29), .Z(\Data_Mem/n6466 ) );
  MUX \Data_Mem/U6469  ( .A(data_mem_out_wire[1475]), .B(
        data_mem_out_wire[1507]), .S(N29), .Z(\Data_Mem/n6465 ) );
  MUX \Data_Mem/U6468  ( .A(\Data_Mem/n6463 ), .B(\Data_Mem/n6456 ), .S(N26), 
        .Z(\Data_Mem/n6464 ) );
  MUX \Data_Mem/U6467  ( .A(\Data_Mem/n6462 ), .B(\Data_Mem/n6459 ), .S(N27), 
        .Z(\Data_Mem/n6463 ) );
  MUX \Data_Mem/U6466  ( .A(\Data_Mem/n6461 ), .B(\Data_Mem/n6460 ), .S(N28), 
        .Z(\Data_Mem/n6462 ) );
  MUX \Data_Mem/U6465  ( .A(data_mem_out_wire[1539]), .B(
        data_mem_out_wire[1571]), .S(N29), .Z(\Data_Mem/n6461 ) );
  MUX \Data_Mem/U6464  ( .A(data_mem_out_wire[1603]), .B(
        data_mem_out_wire[1635]), .S(N29), .Z(\Data_Mem/n6460 ) );
  MUX \Data_Mem/U6463  ( .A(\Data_Mem/n6458 ), .B(\Data_Mem/n6457 ), .S(N28), 
        .Z(\Data_Mem/n6459 ) );
  MUX \Data_Mem/U6462  ( .A(data_mem_out_wire[1667]), .B(
        data_mem_out_wire[1699]), .S(N29), .Z(\Data_Mem/n6458 ) );
  MUX \Data_Mem/U6461  ( .A(data_mem_out_wire[1731]), .B(
        data_mem_out_wire[1763]), .S(N29), .Z(\Data_Mem/n6457 ) );
  MUX \Data_Mem/U6460  ( .A(\Data_Mem/n6455 ), .B(\Data_Mem/n6452 ), .S(N27), 
        .Z(\Data_Mem/n6456 ) );
  MUX \Data_Mem/U6459  ( .A(\Data_Mem/n6454 ), .B(\Data_Mem/n6453 ), .S(N28), 
        .Z(\Data_Mem/n6455 ) );
  MUX \Data_Mem/U6458  ( .A(data_mem_out_wire[1795]), .B(
        data_mem_out_wire[1827]), .S(N29), .Z(\Data_Mem/n6454 ) );
  MUX \Data_Mem/U6457  ( .A(data_mem_out_wire[1859]), .B(
        data_mem_out_wire[1891]), .S(N29), .Z(\Data_Mem/n6453 ) );
  MUX \Data_Mem/U6456  ( .A(\Data_Mem/n6451 ), .B(\Data_Mem/n6450 ), .S(N28), 
        .Z(\Data_Mem/n6452 ) );
  MUX \Data_Mem/U6455  ( .A(data_mem_out_wire[1923]), .B(
        data_mem_out_wire[1955]), .S(N29), .Z(\Data_Mem/n6451 ) );
  MUX \Data_Mem/U6454  ( .A(data_mem_out_wire[1987]), .B(
        data_mem_out_wire[2019]), .S(N29), .Z(\Data_Mem/n6450 ) );
  MUX \Data_Mem/U6453  ( .A(\Data_Mem/n6449 ), .B(\Data_Mem/n6418 ), .S(N24), 
        .Z(c_memory[2]) );
  MUX \Data_Mem/U6452  ( .A(\Data_Mem/n6448 ), .B(\Data_Mem/n6433 ), .S(N25), 
        .Z(\Data_Mem/n6449 ) );
  MUX \Data_Mem/U6451  ( .A(\Data_Mem/n6447 ), .B(\Data_Mem/n6440 ), .S(N26), 
        .Z(\Data_Mem/n6448 ) );
  MUX \Data_Mem/U6450  ( .A(\Data_Mem/n6446 ), .B(\Data_Mem/n6443 ), .S(N27), 
        .Z(\Data_Mem/n6447 ) );
  MUX \Data_Mem/U6449  ( .A(\Data_Mem/n6445 ), .B(\Data_Mem/n6444 ), .S(N28), 
        .Z(\Data_Mem/n6446 ) );
  MUX \Data_Mem/U6448  ( .A(data_mem_out_wire[2]), .B(data_mem_out_wire[34]), 
        .S(N29), .Z(\Data_Mem/n6445 ) );
  MUX \Data_Mem/U6447  ( .A(data_mem_out_wire[66]), .B(data_mem_out_wire[98]), 
        .S(N29), .Z(\Data_Mem/n6444 ) );
  MUX \Data_Mem/U6446  ( .A(\Data_Mem/n6442 ), .B(\Data_Mem/n6441 ), .S(N28), 
        .Z(\Data_Mem/n6443 ) );
  MUX \Data_Mem/U6445  ( .A(data_mem_out_wire[130]), .B(data_mem_out_wire[162]), .S(N29), .Z(\Data_Mem/n6442 ) );
  MUX \Data_Mem/U6444  ( .A(data_mem_out_wire[194]), .B(data_mem_out_wire[226]), .S(N29), .Z(\Data_Mem/n6441 ) );
  MUX \Data_Mem/U6443  ( .A(\Data_Mem/n6439 ), .B(\Data_Mem/n6436 ), .S(N27), 
        .Z(\Data_Mem/n6440 ) );
  MUX \Data_Mem/U6442  ( .A(\Data_Mem/n6438 ), .B(\Data_Mem/n6437 ), .S(N28), 
        .Z(\Data_Mem/n6439 ) );
  MUX \Data_Mem/U6441  ( .A(data_mem_out_wire[258]), .B(data_mem_out_wire[290]), .S(N29), .Z(\Data_Mem/n6438 ) );
  MUX \Data_Mem/U6440  ( .A(data_mem_out_wire[322]), .B(data_mem_out_wire[354]), .S(N29), .Z(\Data_Mem/n6437 ) );
  MUX \Data_Mem/U6439  ( .A(\Data_Mem/n6435 ), .B(\Data_Mem/n6434 ), .S(N28), 
        .Z(\Data_Mem/n6436 ) );
  MUX \Data_Mem/U6438  ( .A(data_mem_out_wire[386]), .B(data_mem_out_wire[418]), .S(N29), .Z(\Data_Mem/n6435 ) );
  MUX \Data_Mem/U6437  ( .A(data_mem_out_wire[450]), .B(data_mem_out_wire[482]), .S(N29), .Z(\Data_Mem/n6434 ) );
  MUX \Data_Mem/U6436  ( .A(\Data_Mem/n6432 ), .B(\Data_Mem/n6425 ), .S(N26), 
        .Z(\Data_Mem/n6433 ) );
  MUX \Data_Mem/U6435  ( .A(\Data_Mem/n6431 ), .B(\Data_Mem/n6428 ), .S(N27), 
        .Z(\Data_Mem/n6432 ) );
  MUX \Data_Mem/U6434  ( .A(\Data_Mem/n6430 ), .B(\Data_Mem/n6429 ), .S(N28), 
        .Z(\Data_Mem/n6431 ) );
  MUX \Data_Mem/U6433  ( .A(data_mem_out_wire[514]), .B(data_mem_out_wire[546]), .S(N29), .Z(\Data_Mem/n6430 ) );
  MUX \Data_Mem/U6432  ( .A(data_mem_out_wire[578]), .B(data_mem_out_wire[610]), .S(N29), .Z(\Data_Mem/n6429 ) );
  MUX \Data_Mem/U6431  ( .A(\Data_Mem/n6427 ), .B(\Data_Mem/n6426 ), .S(N28), 
        .Z(\Data_Mem/n6428 ) );
  MUX \Data_Mem/U6430  ( .A(data_mem_out_wire[642]), .B(data_mem_out_wire[674]), .S(N29), .Z(\Data_Mem/n6427 ) );
  MUX \Data_Mem/U6429  ( .A(data_mem_out_wire[706]), .B(data_mem_out_wire[738]), .S(N29), .Z(\Data_Mem/n6426 ) );
  MUX \Data_Mem/U6428  ( .A(\Data_Mem/n6424 ), .B(\Data_Mem/n6421 ), .S(N27), 
        .Z(\Data_Mem/n6425 ) );
  MUX \Data_Mem/U6427  ( .A(\Data_Mem/n6423 ), .B(\Data_Mem/n6422 ), .S(N28), 
        .Z(\Data_Mem/n6424 ) );
  MUX \Data_Mem/U6426  ( .A(data_mem_out_wire[770]), .B(data_mem_out_wire[802]), .S(N29), .Z(\Data_Mem/n6423 ) );
  MUX \Data_Mem/U6425  ( .A(data_mem_out_wire[834]), .B(data_mem_out_wire[866]), .S(N29), .Z(\Data_Mem/n6422 ) );
  MUX \Data_Mem/U6424  ( .A(\Data_Mem/n6420 ), .B(\Data_Mem/n6419 ), .S(N28), 
        .Z(\Data_Mem/n6421 ) );
  MUX \Data_Mem/U6423  ( .A(data_mem_out_wire[898]), .B(data_mem_out_wire[930]), .S(N29), .Z(\Data_Mem/n6420 ) );
  MUX \Data_Mem/U6422  ( .A(data_mem_out_wire[962]), .B(data_mem_out_wire[994]), .S(N29), .Z(\Data_Mem/n6419 ) );
  MUX \Data_Mem/U6421  ( .A(\Data_Mem/n6417 ), .B(\Data_Mem/n6402 ), .S(N25), 
        .Z(\Data_Mem/n6418 ) );
  MUX \Data_Mem/U6420  ( .A(\Data_Mem/n6416 ), .B(\Data_Mem/n6409 ), .S(N26), 
        .Z(\Data_Mem/n6417 ) );
  MUX \Data_Mem/U6419  ( .A(\Data_Mem/n6415 ), .B(\Data_Mem/n6412 ), .S(N27), 
        .Z(\Data_Mem/n6416 ) );
  MUX \Data_Mem/U6418  ( .A(\Data_Mem/n6414 ), .B(\Data_Mem/n6413 ), .S(N28), 
        .Z(\Data_Mem/n6415 ) );
  MUX \Data_Mem/U6417  ( .A(data_mem_out_wire[1026]), .B(
        data_mem_out_wire[1058]), .S(N29), .Z(\Data_Mem/n6414 ) );
  MUX \Data_Mem/U6416  ( .A(data_mem_out_wire[1090]), .B(
        data_mem_out_wire[1122]), .S(N29), .Z(\Data_Mem/n6413 ) );
  MUX \Data_Mem/U6415  ( .A(\Data_Mem/n6411 ), .B(\Data_Mem/n6410 ), .S(N28), 
        .Z(\Data_Mem/n6412 ) );
  MUX \Data_Mem/U6414  ( .A(data_mem_out_wire[1154]), .B(
        data_mem_out_wire[1186]), .S(N29), .Z(\Data_Mem/n6411 ) );
  MUX \Data_Mem/U6413  ( .A(data_mem_out_wire[1218]), .B(
        data_mem_out_wire[1250]), .S(N29), .Z(\Data_Mem/n6410 ) );
  MUX \Data_Mem/U6412  ( .A(\Data_Mem/n6408 ), .B(\Data_Mem/n6405 ), .S(N27), 
        .Z(\Data_Mem/n6409 ) );
  MUX \Data_Mem/U6411  ( .A(\Data_Mem/n6407 ), .B(\Data_Mem/n6406 ), .S(N28), 
        .Z(\Data_Mem/n6408 ) );
  MUX \Data_Mem/U6410  ( .A(data_mem_out_wire[1282]), .B(
        data_mem_out_wire[1314]), .S(N29), .Z(\Data_Mem/n6407 ) );
  MUX \Data_Mem/U6409  ( .A(data_mem_out_wire[1346]), .B(
        data_mem_out_wire[1378]), .S(N29), .Z(\Data_Mem/n6406 ) );
  MUX \Data_Mem/U6408  ( .A(\Data_Mem/n6404 ), .B(\Data_Mem/n6403 ), .S(N28), 
        .Z(\Data_Mem/n6405 ) );
  MUX \Data_Mem/U6407  ( .A(data_mem_out_wire[1410]), .B(
        data_mem_out_wire[1442]), .S(N29), .Z(\Data_Mem/n6404 ) );
  MUX \Data_Mem/U6406  ( .A(data_mem_out_wire[1474]), .B(
        data_mem_out_wire[1506]), .S(N29), .Z(\Data_Mem/n6403 ) );
  MUX \Data_Mem/U6405  ( .A(\Data_Mem/n6401 ), .B(\Data_Mem/n6394 ), .S(N26), 
        .Z(\Data_Mem/n6402 ) );
  MUX \Data_Mem/U6404  ( .A(\Data_Mem/n6400 ), .B(\Data_Mem/n6397 ), .S(N27), 
        .Z(\Data_Mem/n6401 ) );
  MUX \Data_Mem/U6403  ( .A(\Data_Mem/n6399 ), .B(\Data_Mem/n6398 ), .S(N28), 
        .Z(\Data_Mem/n6400 ) );
  MUX \Data_Mem/U6402  ( .A(data_mem_out_wire[1538]), .B(
        data_mem_out_wire[1570]), .S(N29), .Z(\Data_Mem/n6399 ) );
  MUX \Data_Mem/U6401  ( .A(data_mem_out_wire[1602]), .B(
        data_mem_out_wire[1634]), .S(N29), .Z(\Data_Mem/n6398 ) );
  MUX \Data_Mem/U6400  ( .A(\Data_Mem/n6396 ), .B(\Data_Mem/n6395 ), .S(N28), 
        .Z(\Data_Mem/n6397 ) );
  MUX \Data_Mem/U6399  ( .A(data_mem_out_wire[1666]), .B(
        data_mem_out_wire[1698]), .S(N29), .Z(\Data_Mem/n6396 ) );
  MUX \Data_Mem/U6398  ( .A(data_mem_out_wire[1730]), .B(
        data_mem_out_wire[1762]), .S(N29), .Z(\Data_Mem/n6395 ) );
  MUX \Data_Mem/U6397  ( .A(\Data_Mem/n6393 ), .B(\Data_Mem/n6390 ), .S(N27), 
        .Z(\Data_Mem/n6394 ) );
  MUX \Data_Mem/U6396  ( .A(\Data_Mem/n6392 ), .B(\Data_Mem/n6391 ), .S(N28), 
        .Z(\Data_Mem/n6393 ) );
  MUX \Data_Mem/U6395  ( .A(data_mem_out_wire[1794]), .B(
        data_mem_out_wire[1826]), .S(N29), .Z(\Data_Mem/n6392 ) );
  MUX \Data_Mem/U6394  ( .A(data_mem_out_wire[1858]), .B(
        data_mem_out_wire[1890]), .S(N29), .Z(\Data_Mem/n6391 ) );
  MUX \Data_Mem/U6393  ( .A(\Data_Mem/n6389 ), .B(\Data_Mem/n6388 ), .S(N28), 
        .Z(\Data_Mem/n6390 ) );
  MUX \Data_Mem/U6392  ( .A(data_mem_out_wire[1922]), .B(
        data_mem_out_wire[1954]), .S(N29), .Z(\Data_Mem/n6389 ) );
  MUX \Data_Mem/U6391  ( .A(data_mem_out_wire[1986]), .B(
        data_mem_out_wire[2018]), .S(N29), .Z(\Data_Mem/n6388 ) );
  MUX \Data_Mem/U6390  ( .A(\Data_Mem/n6387 ), .B(\Data_Mem/n6356 ), .S(N24), 
        .Z(c_memory[1]) );
  MUX \Data_Mem/U6389  ( .A(\Data_Mem/n6386 ), .B(\Data_Mem/n6371 ), .S(N25), 
        .Z(\Data_Mem/n6387 ) );
  MUX \Data_Mem/U6388  ( .A(\Data_Mem/n6385 ), .B(\Data_Mem/n6378 ), .S(N26), 
        .Z(\Data_Mem/n6386 ) );
  MUX \Data_Mem/U6387  ( .A(\Data_Mem/n6384 ), .B(\Data_Mem/n6381 ), .S(N27), 
        .Z(\Data_Mem/n6385 ) );
  MUX \Data_Mem/U6386  ( .A(\Data_Mem/n6383 ), .B(\Data_Mem/n6382 ), .S(N28), 
        .Z(\Data_Mem/n6384 ) );
  MUX \Data_Mem/U6385  ( .A(data_mem_out_wire[1]), .B(data_mem_out_wire[33]), 
        .S(N29), .Z(\Data_Mem/n6383 ) );
  MUX \Data_Mem/U6384  ( .A(data_mem_out_wire[65]), .B(data_mem_out_wire[97]), 
        .S(N29), .Z(\Data_Mem/n6382 ) );
  MUX \Data_Mem/U6383  ( .A(\Data_Mem/n6380 ), .B(\Data_Mem/n6379 ), .S(N28), 
        .Z(\Data_Mem/n6381 ) );
  MUX \Data_Mem/U6382  ( .A(data_mem_out_wire[129]), .B(data_mem_out_wire[161]), .S(N29), .Z(\Data_Mem/n6380 ) );
  MUX \Data_Mem/U6381  ( .A(data_mem_out_wire[193]), .B(data_mem_out_wire[225]), .S(N29), .Z(\Data_Mem/n6379 ) );
  MUX \Data_Mem/U6380  ( .A(\Data_Mem/n6377 ), .B(\Data_Mem/n6374 ), .S(N27), 
        .Z(\Data_Mem/n6378 ) );
  MUX \Data_Mem/U6379  ( .A(\Data_Mem/n6376 ), .B(\Data_Mem/n6375 ), .S(N28), 
        .Z(\Data_Mem/n6377 ) );
  MUX \Data_Mem/U6378  ( .A(data_mem_out_wire[257]), .B(data_mem_out_wire[289]), .S(N29), .Z(\Data_Mem/n6376 ) );
  MUX \Data_Mem/U6377  ( .A(data_mem_out_wire[321]), .B(data_mem_out_wire[353]), .S(N29), .Z(\Data_Mem/n6375 ) );
  MUX \Data_Mem/U6376  ( .A(\Data_Mem/n6373 ), .B(\Data_Mem/n6372 ), .S(N28), 
        .Z(\Data_Mem/n6374 ) );
  MUX \Data_Mem/U6375  ( .A(data_mem_out_wire[385]), .B(data_mem_out_wire[417]), .S(N29), .Z(\Data_Mem/n6373 ) );
  MUX \Data_Mem/U6374  ( .A(data_mem_out_wire[449]), .B(data_mem_out_wire[481]), .S(N29), .Z(\Data_Mem/n6372 ) );
  MUX \Data_Mem/U6373  ( .A(\Data_Mem/n6370 ), .B(\Data_Mem/n6363 ), .S(N26), 
        .Z(\Data_Mem/n6371 ) );
  MUX \Data_Mem/U6372  ( .A(\Data_Mem/n6369 ), .B(\Data_Mem/n6366 ), .S(N27), 
        .Z(\Data_Mem/n6370 ) );
  MUX \Data_Mem/U6371  ( .A(\Data_Mem/n6368 ), .B(\Data_Mem/n6367 ), .S(N28), 
        .Z(\Data_Mem/n6369 ) );
  MUX \Data_Mem/U6370  ( .A(data_mem_out_wire[513]), .B(data_mem_out_wire[545]), .S(N29), .Z(\Data_Mem/n6368 ) );
  MUX \Data_Mem/U6369  ( .A(data_mem_out_wire[577]), .B(data_mem_out_wire[609]), .S(N29), .Z(\Data_Mem/n6367 ) );
  MUX \Data_Mem/U6368  ( .A(\Data_Mem/n6365 ), .B(\Data_Mem/n6364 ), .S(N28), 
        .Z(\Data_Mem/n6366 ) );
  MUX \Data_Mem/U6367  ( .A(data_mem_out_wire[641]), .B(data_mem_out_wire[673]), .S(N29), .Z(\Data_Mem/n6365 ) );
  MUX \Data_Mem/U6366  ( .A(data_mem_out_wire[705]), .B(data_mem_out_wire[737]), .S(N29), .Z(\Data_Mem/n6364 ) );
  MUX \Data_Mem/U6365  ( .A(\Data_Mem/n6362 ), .B(\Data_Mem/n6359 ), .S(N27), 
        .Z(\Data_Mem/n6363 ) );
  MUX \Data_Mem/U6364  ( .A(\Data_Mem/n6361 ), .B(\Data_Mem/n6360 ), .S(N28), 
        .Z(\Data_Mem/n6362 ) );
  MUX \Data_Mem/U6363  ( .A(data_mem_out_wire[769]), .B(data_mem_out_wire[801]), .S(N29), .Z(\Data_Mem/n6361 ) );
  MUX \Data_Mem/U6362  ( .A(data_mem_out_wire[833]), .B(data_mem_out_wire[865]), .S(N29), .Z(\Data_Mem/n6360 ) );
  MUX \Data_Mem/U6361  ( .A(\Data_Mem/n6358 ), .B(\Data_Mem/n6357 ), .S(N28), 
        .Z(\Data_Mem/n6359 ) );
  MUX \Data_Mem/U6360  ( .A(data_mem_out_wire[897]), .B(data_mem_out_wire[929]), .S(N29), .Z(\Data_Mem/n6358 ) );
  MUX \Data_Mem/U6359  ( .A(data_mem_out_wire[961]), .B(data_mem_out_wire[993]), .S(N29), .Z(\Data_Mem/n6357 ) );
  MUX \Data_Mem/U6358  ( .A(\Data_Mem/n6355 ), .B(\Data_Mem/n6340 ), .S(N25), 
        .Z(\Data_Mem/n6356 ) );
  MUX \Data_Mem/U6357  ( .A(\Data_Mem/n6354 ), .B(\Data_Mem/n6347 ), .S(N26), 
        .Z(\Data_Mem/n6355 ) );
  MUX \Data_Mem/U6356  ( .A(\Data_Mem/n6353 ), .B(\Data_Mem/n6350 ), .S(N27), 
        .Z(\Data_Mem/n6354 ) );
  MUX \Data_Mem/U6355  ( .A(\Data_Mem/n6352 ), .B(\Data_Mem/n6351 ), .S(N28), 
        .Z(\Data_Mem/n6353 ) );
  MUX \Data_Mem/U6354  ( .A(data_mem_out_wire[1025]), .B(
        data_mem_out_wire[1057]), .S(N29), .Z(\Data_Mem/n6352 ) );
  MUX \Data_Mem/U6353  ( .A(data_mem_out_wire[1089]), .B(
        data_mem_out_wire[1121]), .S(N29), .Z(\Data_Mem/n6351 ) );
  MUX \Data_Mem/U6352  ( .A(\Data_Mem/n6349 ), .B(\Data_Mem/n6348 ), .S(N28), 
        .Z(\Data_Mem/n6350 ) );
  MUX \Data_Mem/U6351  ( .A(data_mem_out_wire[1153]), .B(
        data_mem_out_wire[1185]), .S(N29), .Z(\Data_Mem/n6349 ) );
  MUX \Data_Mem/U6350  ( .A(data_mem_out_wire[1217]), .B(
        data_mem_out_wire[1249]), .S(N29), .Z(\Data_Mem/n6348 ) );
  MUX \Data_Mem/U6349  ( .A(\Data_Mem/n6346 ), .B(\Data_Mem/n6343 ), .S(N27), 
        .Z(\Data_Mem/n6347 ) );
  MUX \Data_Mem/U6348  ( .A(\Data_Mem/n6345 ), .B(\Data_Mem/n6344 ), .S(N28), 
        .Z(\Data_Mem/n6346 ) );
  MUX \Data_Mem/U6347  ( .A(data_mem_out_wire[1281]), .B(
        data_mem_out_wire[1313]), .S(N29), .Z(\Data_Mem/n6345 ) );
  MUX \Data_Mem/U6346  ( .A(data_mem_out_wire[1345]), .B(
        data_mem_out_wire[1377]), .S(N29), .Z(\Data_Mem/n6344 ) );
  MUX \Data_Mem/U6345  ( .A(\Data_Mem/n6342 ), .B(\Data_Mem/n6341 ), .S(N28), 
        .Z(\Data_Mem/n6343 ) );
  MUX \Data_Mem/U6344  ( .A(data_mem_out_wire[1409]), .B(
        data_mem_out_wire[1441]), .S(N29), .Z(\Data_Mem/n6342 ) );
  MUX \Data_Mem/U6343  ( .A(data_mem_out_wire[1473]), .B(
        data_mem_out_wire[1505]), .S(N29), .Z(\Data_Mem/n6341 ) );
  MUX \Data_Mem/U6342  ( .A(\Data_Mem/n6339 ), .B(\Data_Mem/n6332 ), .S(N26), 
        .Z(\Data_Mem/n6340 ) );
  MUX \Data_Mem/U6341  ( .A(\Data_Mem/n6338 ), .B(\Data_Mem/n6335 ), .S(N27), 
        .Z(\Data_Mem/n6339 ) );
  MUX \Data_Mem/U6340  ( .A(\Data_Mem/n6337 ), .B(\Data_Mem/n6336 ), .S(N28), 
        .Z(\Data_Mem/n6338 ) );
  MUX \Data_Mem/U6339  ( .A(data_mem_out_wire[1537]), .B(
        data_mem_out_wire[1569]), .S(N29), .Z(\Data_Mem/n6337 ) );
  MUX \Data_Mem/U6338  ( .A(data_mem_out_wire[1601]), .B(
        data_mem_out_wire[1633]), .S(N29), .Z(\Data_Mem/n6336 ) );
  MUX \Data_Mem/U6337  ( .A(\Data_Mem/n6334 ), .B(\Data_Mem/n6333 ), .S(N28), 
        .Z(\Data_Mem/n6335 ) );
  MUX \Data_Mem/U6336  ( .A(data_mem_out_wire[1665]), .B(
        data_mem_out_wire[1697]), .S(N29), .Z(\Data_Mem/n6334 ) );
  MUX \Data_Mem/U6335  ( .A(data_mem_out_wire[1729]), .B(
        data_mem_out_wire[1761]), .S(N29), .Z(\Data_Mem/n6333 ) );
  MUX \Data_Mem/U6334  ( .A(\Data_Mem/n6331 ), .B(\Data_Mem/n6328 ), .S(N27), 
        .Z(\Data_Mem/n6332 ) );
  MUX \Data_Mem/U6333  ( .A(\Data_Mem/n6330 ), .B(\Data_Mem/n6329 ), .S(N28), 
        .Z(\Data_Mem/n6331 ) );
  MUX \Data_Mem/U6332  ( .A(data_mem_out_wire[1793]), .B(
        data_mem_out_wire[1825]), .S(N29), .Z(\Data_Mem/n6330 ) );
  MUX \Data_Mem/U6331  ( .A(data_mem_out_wire[1857]), .B(
        data_mem_out_wire[1889]), .S(N29), .Z(\Data_Mem/n6329 ) );
  MUX \Data_Mem/U6330  ( .A(\Data_Mem/n6327 ), .B(\Data_Mem/n6326 ), .S(N28), 
        .Z(\Data_Mem/n6328 ) );
  MUX \Data_Mem/U6329  ( .A(data_mem_out_wire[1921]), .B(
        data_mem_out_wire[1953]), .S(N29), .Z(\Data_Mem/n6327 ) );
  MUX \Data_Mem/U6328  ( .A(data_mem_out_wire[1985]), .B(
        data_mem_out_wire[2017]), .S(N29), .Z(\Data_Mem/n6326 ) );
  MUX \Data_Mem/U6327  ( .A(\Data_Mem/n6325 ), .B(\Data_Mem/n6294 ), .S(N24), 
        .Z(c_memory[0]) );
  MUX \Data_Mem/U6326  ( .A(\Data_Mem/n6324 ), .B(\Data_Mem/n6309 ), .S(N25), 
        .Z(\Data_Mem/n6325 ) );
  MUX \Data_Mem/U6325  ( .A(\Data_Mem/n6323 ), .B(\Data_Mem/n6316 ), .S(N26), 
        .Z(\Data_Mem/n6324 ) );
  MUX \Data_Mem/U6324  ( .A(\Data_Mem/n6322 ), .B(\Data_Mem/n6319 ), .S(N27), 
        .Z(\Data_Mem/n6323 ) );
  MUX \Data_Mem/U6323  ( .A(\Data_Mem/n6321 ), .B(\Data_Mem/n6320 ), .S(N28), 
        .Z(\Data_Mem/n6322 ) );
  MUX \Data_Mem/U6322  ( .A(data_mem_out_wire[0]), .B(data_mem_out_wire[32]), 
        .S(N29), .Z(\Data_Mem/n6321 ) );
  MUX \Data_Mem/U6321  ( .A(data_mem_out_wire[64]), .B(data_mem_out_wire[96]), 
        .S(N29), .Z(\Data_Mem/n6320 ) );
  MUX \Data_Mem/U6320  ( .A(\Data_Mem/n6318 ), .B(\Data_Mem/n6317 ), .S(N28), 
        .Z(\Data_Mem/n6319 ) );
  MUX \Data_Mem/U6319  ( .A(data_mem_out_wire[128]), .B(data_mem_out_wire[160]), .S(N29), .Z(\Data_Mem/n6318 ) );
  MUX \Data_Mem/U6318  ( .A(data_mem_out_wire[192]), .B(data_mem_out_wire[224]), .S(N29), .Z(\Data_Mem/n6317 ) );
  MUX \Data_Mem/U6317  ( .A(\Data_Mem/n6315 ), .B(\Data_Mem/n6312 ), .S(N27), 
        .Z(\Data_Mem/n6316 ) );
  MUX \Data_Mem/U6316  ( .A(\Data_Mem/n6314 ), .B(\Data_Mem/n6313 ), .S(N28), 
        .Z(\Data_Mem/n6315 ) );
  MUX \Data_Mem/U6315  ( .A(data_mem_out_wire[256]), .B(data_mem_out_wire[288]), .S(N29), .Z(\Data_Mem/n6314 ) );
  MUX \Data_Mem/U6314  ( .A(data_mem_out_wire[320]), .B(data_mem_out_wire[352]), .S(N29), .Z(\Data_Mem/n6313 ) );
  MUX \Data_Mem/U6313  ( .A(\Data_Mem/n6311 ), .B(\Data_Mem/n6310 ), .S(N28), 
        .Z(\Data_Mem/n6312 ) );
  MUX \Data_Mem/U6312  ( .A(data_mem_out_wire[384]), .B(data_mem_out_wire[416]), .S(N29), .Z(\Data_Mem/n6311 ) );
  MUX \Data_Mem/U6311  ( .A(data_mem_out_wire[448]), .B(data_mem_out_wire[480]), .S(N29), .Z(\Data_Mem/n6310 ) );
  MUX \Data_Mem/U6310  ( .A(\Data_Mem/n6308 ), .B(\Data_Mem/n6301 ), .S(N26), 
        .Z(\Data_Mem/n6309 ) );
  MUX \Data_Mem/U6309  ( .A(\Data_Mem/n6307 ), .B(\Data_Mem/n6304 ), .S(N27), 
        .Z(\Data_Mem/n6308 ) );
  MUX \Data_Mem/U6308  ( .A(\Data_Mem/n6306 ), .B(\Data_Mem/n6305 ), .S(N28), 
        .Z(\Data_Mem/n6307 ) );
  MUX \Data_Mem/U6307  ( .A(data_mem_out_wire[512]), .B(data_mem_out_wire[544]), .S(N29), .Z(\Data_Mem/n6306 ) );
  MUX \Data_Mem/U6306  ( .A(data_mem_out_wire[576]), .B(data_mem_out_wire[608]), .S(N29), .Z(\Data_Mem/n6305 ) );
  MUX \Data_Mem/U6305  ( .A(\Data_Mem/n6303 ), .B(\Data_Mem/n6302 ), .S(N28), 
        .Z(\Data_Mem/n6304 ) );
  MUX \Data_Mem/U6304  ( .A(data_mem_out_wire[640]), .B(data_mem_out_wire[672]), .S(N29), .Z(\Data_Mem/n6303 ) );
  MUX \Data_Mem/U6303  ( .A(data_mem_out_wire[704]), .B(data_mem_out_wire[736]), .S(N29), .Z(\Data_Mem/n6302 ) );
  MUX \Data_Mem/U6302  ( .A(\Data_Mem/n6300 ), .B(\Data_Mem/n6297 ), .S(N27), 
        .Z(\Data_Mem/n6301 ) );
  MUX \Data_Mem/U6301  ( .A(\Data_Mem/n6299 ), .B(\Data_Mem/n6298 ), .S(N28), 
        .Z(\Data_Mem/n6300 ) );
  MUX \Data_Mem/U6300  ( .A(data_mem_out_wire[768]), .B(data_mem_out_wire[800]), .S(N29), .Z(\Data_Mem/n6299 ) );
  MUX \Data_Mem/U6299  ( .A(data_mem_out_wire[832]), .B(data_mem_out_wire[864]), .S(N29), .Z(\Data_Mem/n6298 ) );
  MUX \Data_Mem/U6298  ( .A(\Data_Mem/n6296 ), .B(\Data_Mem/n6295 ), .S(N28), 
        .Z(\Data_Mem/n6297 ) );
  MUX \Data_Mem/U6297  ( .A(data_mem_out_wire[896]), .B(data_mem_out_wire[928]), .S(N29), .Z(\Data_Mem/n6296 ) );
  MUX \Data_Mem/U6296  ( .A(data_mem_out_wire[960]), .B(data_mem_out_wire[992]), .S(N29), .Z(\Data_Mem/n6295 ) );
  MUX \Data_Mem/U6295  ( .A(\Data_Mem/n6293 ), .B(\Data_Mem/n6278 ), .S(N25), 
        .Z(\Data_Mem/n6294 ) );
  MUX \Data_Mem/U6294  ( .A(\Data_Mem/n6292 ), .B(\Data_Mem/n6285 ), .S(N26), 
        .Z(\Data_Mem/n6293 ) );
  MUX \Data_Mem/U6293  ( .A(\Data_Mem/n6291 ), .B(\Data_Mem/n6288 ), .S(N27), 
        .Z(\Data_Mem/n6292 ) );
  MUX \Data_Mem/U6292  ( .A(\Data_Mem/n6290 ), .B(\Data_Mem/n6289 ), .S(N28), 
        .Z(\Data_Mem/n6291 ) );
  MUX \Data_Mem/U6291  ( .A(data_mem_out_wire[1024]), .B(
        data_mem_out_wire[1056]), .S(N29), .Z(\Data_Mem/n6290 ) );
  MUX \Data_Mem/U6290  ( .A(data_mem_out_wire[1088]), .B(
        data_mem_out_wire[1120]), .S(N29), .Z(\Data_Mem/n6289 ) );
  MUX \Data_Mem/U6289  ( .A(\Data_Mem/n6287 ), .B(\Data_Mem/n6286 ), .S(N28), 
        .Z(\Data_Mem/n6288 ) );
  MUX \Data_Mem/U6288  ( .A(data_mem_out_wire[1152]), .B(
        data_mem_out_wire[1184]), .S(N29), .Z(\Data_Mem/n6287 ) );
  MUX \Data_Mem/U6287  ( .A(data_mem_out_wire[1216]), .B(
        data_mem_out_wire[1248]), .S(N29), .Z(\Data_Mem/n6286 ) );
  MUX \Data_Mem/U6286  ( .A(\Data_Mem/n6284 ), .B(\Data_Mem/n6281 ), .S(N27), 
        .Z(\Data_Mem/n6285 ) );
  MUX \Data_Mem/U6285  ( .A(\Data_Mem/n6283 ), .B(\Data_Mem/n6282 ), .S(N28), 
        .Z(\Data_Mem/n6284 ) );
  MUX \Data_Mem/U6284  ( .A(data_mem_out_wire[1280]), .B(
        data_mem_out_wire[1312]), .S(N29), .Z(\Data_Mem/n6283 ) );
  MUX \Data_Mem/U6283  ( .A(data_mem_out_wire[1344]), .B(
        data_mem_out_wire[1376]), .S(N29), .Z(\Data_Mem/n6282 ) );
  MUX \Data_Mem/U6282  ( .A(\Data_Mem/n6280 ), .B(\Data_Mem/n6279 ), .S(N28), 
        .Z(\Data_Mem/n6281 ) );
  MUX \Data_Mem/U6281  ( .A(data_mem_out_wire[1408]), .B(
        data_mem_out_wire[1440]), .S(N29), .Z(\Data_Mem/n6280 ) );
  MUX \Data_Mem/U6280  ( .A(data_mem_out_wire[1472]), .B(
        data_mem_out_wire[1504]), .S(N29), .Z(\Data_Mem/n6279 ) );
  MUX \Data_Mem/U6279  ( .A(\Data_Mem/n6277 ), .B(\Data_Mem/n6270 ), .S(N26), 
        .Z(\Data_Mem/n6278 ) );
  MUX \Data_Mem/U6278  ( .A(\Data_Mem/n6276 ), .B(\Data_Mem/n6273 ), .S(N27), 
        .Z(\Data_Mem/n6277 ) );
  MUX \Data_Mem/U6277  ( .A(\Data_Mem/n6275 ), .B(\Data_Mem/n6274 ), .S(N28), 
        .Z(\Data_Mem/n6276 ) );
  MUX \Data_Mem/U6276  ( .A(data_mem_out_wire[1536]), .B(
        data_mem_out_wire[1568]), .S(N29), .Z(\Data_Mem/n6275 ) );
  MUX \Data_Mem/U6275  ( .A(data_mem_out_wire[1600]), .B(
        data_mem_out_wire[1632]), .S(N29), .Z(\Data_Mem/n6274 ) );
  MUX \Data_Mem/U6274  ( .A(\Data_Mem/n6272 ), .B(\Data_Mem/n6271 ), .S(N28), 
        .Z(\Data_Mem/n6273 ) );
  MUX \Data_Mem/U6273  ( .A(data_mem_out_wire[1664]), .B(
        data_mem_out_wire[1696]), .S(N29), .Z(\Data_Mem/n6272 ) );
  MUX \Data_Mem/U6272  ( .A(data_mem_out_wire[1728]), .B(
        data_mem_out_wire[1760]), .S(N29), .Z(\Data_Mem/n6271 ) );
  MUX \Data_Mem/U6271  ( .A(\Data_Mem/n6269 ), .B(\Data_Mem/n6266 ), .S(N27), 
        .Z(\Data_Mem/n6270 ) );
  MUX \Data_Mem/U6270  ( .A(\Data_Mem/n6268 ), .B(\Data_Mem/n6267 ), .S(N28), 
        .Z(\Data_Mem/n6269 ) );
  MUX \Data_Mem/U6269  ( .A(data_mem_out_wire[1792]), .B(
        data_mem_out_wire[1824]), .S(N29), .Z(\Data_Mem/n6268 ) );
  MUX \Data_Mem/U6268  ( .A(data_mem_out_wire[1856]), .B(
        data_mem_out_wire[1888]), .S(N29), .Z(\Data_Mem/n6267 ) );
  MUX \Data_Mem/U6267  ( .A(\Data_Mem/n6265 ), .B(\Data_Mem/n6264 ), .S(N28), 
        .Z(\Data_Mem/n6266 ) );
  MUX \Data_Mem/U6266  ( .A(data_mem_out_wire[1920]), .B(
        data_mem_out_wire[1952]), .S(N29), .Z(\Data_Mem/n6265 ) );
  MUX \Data_Mem/U6265  ( .A(data_mem_out_wire[1984]), .B(
        data_mem_out_wire[2016]), .S(N29), .Z(\Data_Mem/n6264 ) );
  DFF \Data_Mem/memory_reg[63][0]  ( .D(\Data_Mem/n4216 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2016]), .Q(data_mem_out_wire[2016]) );
  DFF \Data_Mem/memory_reg[63][1]  ( .D(\Data_Mem/n4217 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2017]), .Q(data_mem_out_wire[2017]) );
  DFF \Data_Mem/memory_reg[63][2]  ( .D(\Data_Mem/n4218 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2018]), .Q(data_mem_out_wire[2018]) );
  DFF \Data_Mem/memory_reg[63][3]  ( .D(\Data_Mem/n4219 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2019]), .Q(data_mem_out_wire[2019]) );
  DFF \Data_Mem/memory_reg[63][4]  ( .D(\Data_Mem/n4220 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2020]), .Q(data_mem_out_wire[2020]) );
  DFF \Data_Mem/memory_reg[63][5]  ( .D(\Data_Mem/n4221 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2021]), .Q(data_mem_out_wire[2021]) );
  DFF \Data_Mem/memory_reg[63][6]  ( .D(\Data_Mem/n4222 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2022]), .Q(data_mem_out_wire[2022]) );
  DFF \Data_Mem/memory_reg[63][7]  ( .D(\Data_Mem/n4223 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2023]), .Q(data_mem_out_wire[2023]) );
  DFF \Data_Mem/memory_reg[63][8]  ( .D(\Data_Mem/n4224 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2024]), .Q(data_mem_out_wire[2024]) );
  DFF \Data_Mem/memory_reg[63][9]  ( .D(\Data_Mem/n4225 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[2025]), .Q(data_mem_out_wire[2025]) );
  DFF \Data_Mem/memory_reg[63][10]  ( .D(\Data_Mem/n4226 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2026]), .Q(data_mem_out_wire[2026]) );
  DFF \Data_Mem/memory_reg[63][11]  ( .D(\Data_Mem/n4227 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2027]), .Q(data_mem_out_wire[2027]) );
  DFF \Data_Mem/memory_reg[63][12]  ( .D(\Data_Mem/n4228 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2028]), .Q(data_mem_out_wire[2028]) );
  DFF \Data_Mem/memory_reg[63][13]  ( .D(\Data_Mem/n4229 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2029]), .Q(data_mem_out_wire[2029]) );
  DFF \Data_Mem/memory_reg[63][14]  ( .D(\Data_Mem/n4230 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2030]), .Q(data_mem_out_wire[2030]) );
  DFF \Data_Mem/memory_reg[63][15]  ( .D(\Data_Mem/n4231 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2031]), .Q(data_mem_out_wire[2031]) );
  DFF \Data_Mem/memory_reg[63][16]  ( .D(\Data_Mem/n4232 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2032]), .Q(data_mem_out_wire[2032]) );
  DFF \Data_Mem/memory_reg[63][17]  ( .D(\Data_Mem/n4233 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2033]), .Q(data_mem_out_wire[2033]) );
  DFF \Data_Mem/memory_reg[63][18]  ( .D(\Data_Mem/n4234 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2034]), .Q(data_mem_out_wire[2034]) );
  DFF \Data_Mem/memory_reg[63][19]  ( .D(\Data_Mem/n4235 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2035]), .Q(data_mem_out_wire[2035]) );
  DFF \Data_Mem/memory_reg[63][20]  ( .D(\Data_Mem/n4236 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2036]), .Q(data_mem_out_wire[2036]) );
  DFF \Data_Mem/memory_reg[63][21]  ( .D(\Data_Mem/n4237 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2037]), .Q(data_mem_out_wire[2037]) );
  DFF \Data_Mem/memory_reg[63][22]  ( .D(\Data_Mem/n4238 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2038]), .Q(data_mem_out_wire[2038]) );
  DFF \Data_Mem/memory_reg[63][23]  ( .D(\Data_Mem/n4239 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2039]), .Q(data_mem_out_wire[2039]) );
  DFF \Data_Mem/memory_reg[63][24]  ( .D(\Data_Mem/n4240 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2040]), .Q(data_mem_out_wire[2040]) );
  DFF \Data_Mem/memory_reg[63][25]  ( .D(\Data_Mem/n4241 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2041]), .Q(data_mem_out_wire[2041]) );
  DFF \Data_Mem/memory_reg[63][26]  ( .D(\Data_Mem/n4242 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2042]), .Q(data_mem_out_wire[2042]) );
  DFF \Data_Mem/memory_reg[63][27]  ( .D(\Data_Mem/n4243 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2043]), .Q(data_mem_out_wire[2043]) );
  DFF \Data_Mem/memory_reg[63][28]  ( .D(\Data_Mem/n4244 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2044]), .Q(data_mem_out_wire[2044]) );
  DFF \Data_Mem/memory_reg[63][29]  ( .D(\Data_Mem/n4245 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2045]), .Q(data_mem_out_wire[2045]) );
  DFF \Data_Mem/memory_reg[63][30]  ( .D(\Data_Mem/n4246 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2046]), .Q(data_mem_out_wire[2046]) );
  DFF \Data_Mem/memory_reg[63][31]  ( .D(\Data_Mem/n4247 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2047]), .Q(data_mem_out_wire[2047]) );
  DFF \Data_Mem/memory_reg[62][0]  ( .D(\Data_Mem/n4248 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1984]), .Q(data_mem_out_wire[1984]) );
  DFF \Data_Mem/memory_reg[62][1]  ( .D(\Data_Mem/n4249 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1985]), .Q(data_mem_out_wire[1985]) );
  DFF \Data_Mem/memory_reg[62][2]  ( .D(\Data_Mem/n4250 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1986]), .Q(data_mem_out_wire[1986]) );
  DFF \Data_Mem/memory_reg[62][3]  ( .D(\Data_Mem/n4251 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1987]), .Q(data_mem_out_wire[1987]) );
  DFF \Data_Mem/memory_reg[62][4]  ( .D(\Data_Mem/n4252 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1988]), .Q(data_mem_out_wire[1988]) );
  DFF \Data_Mem/memory_reg[62][5]  ( .D(\Data_Mem/n4253 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1989]), .Q(data_mem_out_wire[1989]) );
  DFF \Data_Mem/memory_reg[62][6]  ( .D(\Data_Mem/n4254 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1990]), .Q(data_mem_out_wire[1990]) );
  DFF \Data_Mem/memory_reg[62][7]  ( .D(\Data_Mem/n4255 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1991]), .Q(data_mem_out_wire[1991]) );
  DFF \Data_Mem/memory_reg[62][8]  ( .D(\Data_Mem/n4256 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1992]), .Q(data_mem_out_wire[1992]) );
  DFF \Data_Mem/memory_reg[62][9]  ( .D(\Data_Mem/n4257 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1993]), .Q(data_mem_out_wire[1993]) );
  DFF \Data_Mem/memory_reg[62][10]  ( .D(\Data_Mem/n4258 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1994]), .Q(data_mem_out_wire[1994]) );
  DFF \Data_Mem/memory_reg[62][11]  ( .D(\Data_Mem/n4259 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1995]), .Q(data_mem_out_wire[1995]) );
  DFF \Data_Mem/memory_reg[62][12]  ( .D(\Data_Mem/n4260 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1996]), .Q(data_mem_out_wire[1996]) );
  DFF \Data_Mem/memory_reg[62][13]  ( .D(\Data_Mem/n4261 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1997]), .Q(data_mem_out_wire[1997]) );
  DFF \Data_Mem/memory_reg[62][14]  ( .D(\Data_Mem/n4262 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1998]), .Q(data_mem_out_wire[1998]) );
  DFF \Data_Mem/memory_reg[62][15]  ( .D(\Data_Mem/n4263 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1999]), .Q(data_mem_out_wire[1999]) );
  DFF \Data_Mem/memory_reg[62][16]  ( .D(\Data_Mem/n4264 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2000]), .Q(data_mem_out_wire[2000]) );
  DFF \Data_Mem/memory_reg[62][17]  ( .D(\Data_Mem/n4265 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2001]), .Q(data_mem_out_wire[2001]) );
  DFF \Data_Mem/memory_reg[62][18]  ( .D(\Data_Mem/n4266 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2002]), .Q(data_mem_out_wire[2002]) );
  DFF \Data_Mem/memory_reg[62][19]  ( .D(\Data_Mem/n4267 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2003]), .Q(data_mem_out_wire[2003]) );
  DFF \Data_Mem/memory_reg[62][20]  ( .D(\Data_Mem/n4268 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2004]), .Q(data_mem_out_wire[2004]) );
  DFF \Data_Mem/memory_reg[62][21]  ( .D(\Data_Mem/n4269 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2005]), .Q(data_mem_out_wire[2005]) );
  DFF \Data_Mem/memory_reg[62][22]  ( .D(\Data_Mem/n4270 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2006]), .Q(data_mem_out_wire[2006]) );
  DFF \Data_Mem/memory_reg[62][23]  ( .D(\Data_Mem/n4271 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2007]), .Q(data_mem_out_wire[2007]) );
  DFF \Data_Mem/memory_reg[62][24]  ( .D(\Data_Mem/n4272 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2008]), .Q(data_mem_out_wire[2008]) );
  DFF \Data_Mem/memory_reg[62][25]  ( .D(\Data_Mem/n4273 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2009]), .Q(data_mem_out_wire[2009]) );
  DFF \Data_Mem/memory_reg[62][26]  ( .D(\Data_Mem/n4274 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2010]), .Q(data_mem_out_wire[2010]) );
  DFF \Data_Mem/memory_reg[62][27]  ( .D(\Data_Mem/n4275 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2011]), .Q(data_mem_out_wire[2011]) );
  DFF \Data_Mem/memory_reg[62][28]  ( .D(\Data_Mem/n4276 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2012]), .Q(data_mem_out_wire[2012]) );
  DFF \Data_Mem/memory_reg[62][29]  ( .D(\Data_Mem/n4277 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2013]), .Q(data_mem_out_wire[2013]) );
  DFF \Data_Mem/memory_reg[62][30]  ( .D(\Data_Mem/n4278 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2014]), .Q(data_mem_out_wire[2014]) );
  DFF \Data_Mem/memory_reg[62][31]  ( .D(\Data_Mem/n4279 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[2015]), .Q(data_mem_out_wire[2015]) );
  DFF \Data_Mem/memory_reg[61][0]  ( .D(\Data_Mem/n4280 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1952]), .Q(data_mem_out_wire[1952]) );
  DFF \Data_Mem/memory_reg[61][1]  ( .D(\Data_Mem/n4281 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1953]), .Q(data_mem_out_wire[1953]) );
  DFF \Data_Mem/memory_reg[61][2]  ( .D(\Data_Mem/n4282 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1954]), .Q(data_mem_out_wire[1954]) );
  DFF \Data_Mem/memory_reg[61][3]  ( .D(\Data_Mem/n4283 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1955]), .Q(data_mem_out_wire[1955]) );
  DFF \Data_Mem/memory_reg[61][4]  ( .D(\Data_Mem/n4284 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1956]), .Q(data_mem_out_wire[1956]) );
  DFF \Data_Mem/memory_reg[61][5]  ( .D(\Data_Mem/n4285 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1957]), .Q(data_mem_out_wire[1957]) );
  DFF \Data_Mem/memory_reg[61][6]  ( .D(\Data_Mem/n4286 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1958]), .Q(data_mem_out_wire[1958]) );
  DFF \Data_Mem/memory_reg[61][7]  ( .D(\Data_Mem/n4287 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1959]), .Q(data_mem_out_wire[1959]) );
  DFF \Data_Mem/memory_reg[61][8]  ( .D(\Data_Mem/n4288 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1960]), .Q(data_mem_out_wire[1960]) );
  DFF \Data_Mem/memory_reg[61][9]  ( .D(\Data_Mem/n4289 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1961]), .Q(data_mem_out_wire[1961]) );
  DFF \Data_Mem/memory_reg[61][10]  ( .D(\Data_Mem/n4290 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1962]), .Q(data_mem_out_wire[1962]) );
  DFF \Data_Mem/memory_reg[61][11]  ( .D(\Data_Mem/n4291 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1963]), .Q(data_mem_out_wire[1963]) );
  DFF \Data_Mem/memory_reg[61][12]  ( .D(\Data_Mem/n4292 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1964]), .Q(data_mem_out_wire[1964]) );
  DFF \Data_Mem/memory_reg[61][13]  ( .D(\Data_Mem/n4293 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1965]), .Q(data_mem_out_wire[1965]) );
  DFF \Data_Mem/memory_reg[61][14]  ( .D(\Data_Mem/n4294 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1966]), .Q(data_mem_out_wire[1966]) );
  DFF \Data_Mem/memory_reg[61][15]  ( .D(\Data_Mem/n4295 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1967]), .Q(data_mem_out_wire[1967]) );
  DFF \Data_Mem/memory_reg[61][16]  ( .D(\Data_Mem/n4296 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1968]), .Q(data_mem_out_wire[1968]) );
  DFF \Data_Mem/memory_reg[61][17]  ( .D(\Data_Mem/n4297 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1969]), .Q(data_mem_out_wire[1969]) );
  DFF \Data_Mem/memory_reg[61][18]  ( .D(\Data_Mem/n4298 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1970]), .Q(data_mem_out_wire[1970]) );
  DFF \Data_Mem/memory_reg[61][19]  ( .D(\Data_Mem/n4299 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1971]), .Q(data_mem_out_wire[1971]) );
  DFF \Data_Mem/memory_reg[61][20]  ( .D(\Data_Mem/n4300 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1972]), .Q(data_mem_out_wire[1972]) );
  DFF \Data_Mem/memory_reg[61][21]  ( .D(\Data_Mem/n4301 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1973]), .Q(data_mem_out_wire[1973]) );
  DFF \Data_Mem/memory_reg[61][22]  ( .D(\Data_Mem/n4302 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1974]), .Q(data_mem_out_wire[1974]) );
  DFF \Data_Mem/memory_reg[61][23]  ( .D(\Data_Mem/n4303 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1975]), .Q(data_mem_out_wire[1975]) );
  DFF \Data_Mem/memory_reg[61][24]  ( .D(\Data_Mem/n4304 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1976]), .Q(data_mem_out_wire[1976]) );
  DFF \Data_Mem/memory_reg[61][25]  ( .D(\Data_Mem/n4305 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1977]), .Q(data_mem_out_wire[1977]) );
  DFF \Data_Mem/memory_reg[61][26]  ( .D(\Data_Mem/n4306 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1978]), .Q(data_mem_out_wire[1978]) );
  DFF \Data_Mem/memory_reg[61][27]  ( .D(\Data_Mem/n4307 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1979]), .Q(data_mem_out_wire[1979]) );
  DFF \Data_Mem/memory_reg[61][28]  ( .D(\Data_Mem/n4308 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1980]), .Q(data_mem_out_wire[1980]) );
  DFF \Data_Mem/memory_reg[61][29]  ( .D(\Data_Mem/n4309 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1981]), .Q(data_mem_out_wire[1981]) );
  DFF \Data_Mem/memory_reg[61][30]  ( .D(\Data_Mem/n4310 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1982]), .Q(data_mem_out_wire[1982]) );
  DFF \Data_Mem/memory_reg[61][31]  ( .D(\Data_Mem/n4311 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1983]), .Q(data_mem_out_wire[1983]) );
  DFF \Data_Mem/memory_reg[60][0]  ( .D(\Data_Mem/n4312 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1920]), .Q(data_mem_out_wire[1920]) );
  DFF \Data_Mem/memory_reg[60][1]  ( .D(\Data_Mem/n4313 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1921]), .Q(data_mem_out_wire[1921]) );
  DFF \Data_Mem/memory_reg[60][2]  ( .D(\Data_Mem/n4314 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1922]), .Q(data_mem_out_wire[1922]) );
  DFF \Data_Mem/memory_reg[60][3]  ( .D(\Data_Mem/n4315 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1923]), .Q(data_mem_out_wire[1923]) );
  DFF \Data_Mem/memory_reg[60][4]  ( .D(\Data_Mem/n4316 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1924]), .Q(data_mem_out_wire[1924]) );
  DFF \Data_Mem/memory_reg[60][5]  ( .D(\Data_Mem/n4317 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1925]), .Q(data_mem_out_wire[1925]) );
  DFF \Data_Mem/memory_reg[60][6]  ( .D(\Data_Mem/n4318 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1926]), .Q(data_mem_out_wire[1926]) );
  DFF \Data_Mem/memory_reg[60][7]  ( .D(\Data_Mem/n4319 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1927]), .Q(data_mem_out_wire[1927]) );
  DFF \Data_Mem/memory_reg[60][8]  ( .D(\Data_Mem/n4320 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1928]), .Q(data_mem_out_wire[1928]) );
  DFF \Data_Mem/memory_reg[60][9]  ( .D(\Data_Mem/n4321 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1929]), .Q(data_mem_out_wire[1929]) );
  DFF \Data_Mem/memory_reg[60][10]  ( .D(\Data_Mem/n4322 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1930]), .Q(data_mem_out_wire[1930]) );
  DFF \Data_Mem/memory_reg[60][11]  ( .D(\Data_Mem/n4323 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1931]), .Q(data_mem_out_wire[1931]) );
  DFF \Data_Mem/memory_reg[60][12]  ( .D(\Data_Mem/n4324 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1932]), .Q(data_mem_out_wire[1932]) );
  DFF \Data_Mem/memory_reg[60][13]  ( .D(\Data_Mem/n4325 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1933]), .Q(data_mem_out_wire[1933]) );
  DFF \Data_Mem/memory_reg[60][14]  ( .D(\Data_Mem/n4326 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1934]), .Q(data_mem_out_wire[1934]) );
  DFF \Data_Mem/memory_reg[60][15]  ( .D(\Data_Mem/n4327 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1935]), .Q(data_mem_out_wire[1935]) );
  DFF \Data_Mem/memory_reg[60][16]  ( .D(\Data_Mem/n4328 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1936]), .Q(data_mem_out_wire[1936]) );
  DFF \Data_Mem/memory_reg[60][17]  ( .D(\Data_Mem/n4329 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1937]), .Q(data_mem_out_wire[1937]) );
  DFF \Data_Mem/memory_reg[60][18]  ( .D(\Data_Mem/n4330 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1938]), .Q(data_mem_out_wire[1938]) );
  DFF \Data_Mem/memory_reg[60][19]  ( .D(\Data_Mem/n4331 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1939]), .Q(data_mem_out_wire[1939]) );
  DFF \Data_Mem/memory_reg[60][20]  ( .D(\Data_Mem/n4332 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1940]), .Q(data_mem_out_wire[1940]) );
  DFF \Data_Mem/memory_reg[60][21]  ( .D(\Data_Mem/n4333 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1941]), .Q(data_mem_out_wire[1941]) );
  DFF \Data_Mem/memory_reg[60][22]  ( .D(\Data_Mem/n4334 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1942]), .Q(data_mem_out_wire[1942]) );
  DFF \Data_Mem/memory_reg[60][23]  ( .D(\Data_Mem/n4335 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1943]), .Q(data_mem_out_wire[1943]) );
  DFF \Data_Mem/memory_reg[60][24]  ( .D(\Data_Mem/n4336 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1944]), .Q(data_mem_out_wire[1944]) );
  DFF \Data_Mem/memory_reg[60][25]  ( .D(\Data_Mem/n4337 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1945]), .Q(data_mem_out_wire[1945]) );
  DFF \Data_Mem/memory_reg[60][26]  ( .D(\Data_Mem/n4338 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1946]), .Q(data_mem_out_wire[1946]) );
  DFF \Data_Mem/memory_reg[60][27]  ( .D(\Data_Mem/n4339 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1947]), .Q(data_mem_out_wire[1947]) );
  DFF \Data_Mem/memory_reg[60][28]  ( .D(\Data_Mem/n4340 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1948]), .Q(data_mem_out_wire[1948]) );
  DFF \Data_Mem/memory_reg[60][29]  ( .D(\Data_Mem/n4341 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1949]), .Q(data_mem_out_wire[1949]) );
  DFF \Data_Mem/memory_reg[60][30]  ( .D(\Data_Mem/n4342 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1950]), .Q(data_mem_out_wire[1950]) );
  DFF \Data_Mem/memory_reg[60][31]  ( .D(\Data_Mem/n4343 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1951]), .Q(data_mem_out_wire[1951]) );
  DFF \Data_Mem/memory_reg[59][0]  ( .D(\Data_Mem/n4344 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1888]), .Q(data_mem_out_wire[1888]) );
  DFF \Data_Mem/memory_reg[59][1]  ( .D(\Data_Mem/n4345 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1889]), .Q(data_mem_out_wire[1889]) );
  DFF \Data_Mem/memory_reg[59][2]  ( .D(\Data_Mem/n4346 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1890]), .Q(data_mem_out_wire[1890]) );
  DFF \Data_Mem/memory_reg[59][3]  ( .D(\Data_Mem/n4347 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1891]), .Q(data_mem_out_wire[1891]) );
  DFF \Data_Mem/memory_reg[59][4]  ( .D(\Data_Mem/n4348 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1892]), .Q(data_mem_out_wire[1892]) );
  DFF \Data_Mem/memory_reg[59][5]  ( .D(\Data_Mem/n4349 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1893]), .Q(data_mem_out_wire[1893]) );
  DFF \Data_Mem/memory_reg[59][6]  ( .D(\Data_Mem/n4350 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1894]), .Q(data_mem_out_wire[1894]) );
  DFF \Data_Mem/memory_reg[59][7]  ( .D(\Data_Mem/n4351 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1895]), .Q(data_mem_out_wire[1895]) );
  DFF \Data_Mem/memory_reg[59][8]  ( .D(\Data_Mem/n4352 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1896]), .Q(data_mem_out_wire[1896]) );
  DFF \Data_Mem/memory_reg[59][9]  ( .D(\Data_Mem/n4353 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1897]), .Q(data_mem_out_wire[1897]) );
  DFF \Data_Mem/memory_reg[59][10]  ( .D(\Data_Mem/n4354 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1898]), .Q(data_mem_out_wire[1898]) );
  DFF \Data_Mem/memory_reg[59][11]  ( .D(\Data_Mem/n4355 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1899]), .Q(data_mem_out_wire[1899]) );
  DFF \Data_Mem/memory_reg[59][12]  ( .D(\Data_Mem/n4356 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1900]), .Q(data_mem_out_wire[1900]) );
  DFF \Data_Mem/memory_reg[59][13]  ( .D(\Data_Mem/n4357 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1901]), .Q(data_mem_out_wire[1901]) );
  DFF \Data_Mem/memory_reg[59][14]  ( .D(\Data_Mem/n4358 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1902]), .Q(data_mem_out_wire[1902]) );
  DFF \Data_Mem/memory_reg[59][15]  ( .D(\Data_Mem/n4359 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1903]), .Q(data_mem_out_wire[1903]) );
  DFF \Data_Mem/memory_reg[59][16]  ( .D(\Data_Mem/n4360 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1904]), .Q(data_mem_out_wire[1904]) );
  DFF \Data_Mem/memory_reg[59][17]  ( .D(\Data_Mem/n4361 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1905]), .Q(data_mem_out_wire[1905]) );
  DFF \Data_Mem/memory_reg[59][18]  ( .D(\Data_Mem/n4362 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1906]), .Q(data_mem_out_wire[1906]) );
  DFF \Data_Mem/memory_reg[59][19]  ( .D(\Data_Mem/n4363 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1907]), .Q(data_mem_out_wire[1907]) );
  DFF \Data_Mem/memory_reg[59][20]  ( .D(\Data_Mem/n4364 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1908]), .Q(data_mem_out_wire[1908]) );
  DFF \Data_Mem/memory_reg[59][21]  ( .D(\Data_Mem/n4365 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1909]), .Q(data_mem_out_wire[1909]) );
  DFF \Data_Mem/memory_reg[59][22]  ( .D(\Data_Mem/n4366 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1910]), .Q(data_mem_out_wire[1910]) );
  DFF \Data_Mem/memory_reg[59][23]  ( .D(\Data_Mem/n4367 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1911]), .Q(data_mem_out_wire[1911]) );
  DFF \Data_Mem/memory_reg[59][24]  ( .D(\Data_Mem/n4368 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1912]), .Q(data_mem_out_wire[1912]) );
  DFF \Data_Mem/memory_reg[59][25]  ( .D(\Data_Mem/n4369 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1913]), .Q(data_mem_out_wire[1913]) );
  DFF \Data_Mem/memory_reg[59][26]  ( .D(\Data_Mem/n4370 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1914]), .Q(data_mem_out_wire[1914]) );
  DFF \Data_Mem/memory_reg[59][27]  ( .D(\Data_Mem/n4371 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1915]), .Q(data_mem_out_wire[1915]) );
  DFF \Data_Mem/memory_reg[59][28]  ( .D(\Data_Mem/n4372 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1916]), .Q(data_mem_out_wire[1916]) );
  DFF \Data_Mem/memory_reg[59][29]  ( .D(\Data_Mem/n4373 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1917]), .Q(data_mem_out_wire[1917]) );
  DFF \Data_Mem/memory_reg[59][30]  ( .D(\Data_Mem/n4374 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1918]), .Q(data_mem_out_wire[1918]) );
  DFF \Data_Mem/memory_reg[59][31]  ( .D(\Data_Mem/n4375 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1919]), .Q(data_mem_out_wire[1919]) );
  DFF \Data_Mem/memory_reg[58][0]  ( .D(\Data_Mem/n4376 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1856]), .Q(data_mem_out_wire[1856]) );
  DFF \Data_Mem/memory_reg[58][1]  ( .D(\Data_Mem/n4377 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1857]), .Q(data_mem_out_wire[1857]) );
  DFF \Data_Mem/memory_reg[58][2]  ( .D(\Data_Mem/n4378 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1858]), .Q(data_mem_out_wire[1858]) );
  DFF \Data_Mem/memory_reg[58][3]  ( .D(\Data_Mem/n4379 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1859]), .Q(data_mem_out_wire[1859]) );
  DFF \Data_Mem/memory_reg[58][4]  ( .D(\Data_Mem/n4380 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1860]), .Q(data_mem_out_wire[1860]) );
  DFF \Data_Mem/memory_reg[58][5]  ( .D(\Data_Mem/n4381 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1861]), .Q(data_mem_out_wire[1861]) );
  DFF \Data_Mem/memory_reg[58][6]  ( .D(\Data_Mem/n4382 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1862]), .Q(data_mem_out_wire[1862]) );
  DFF \Data_Mem/memory_reg[58][7]  ( .D(\Data_Mem/n4383 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1863]), .Q(data_mem_out_wire[1863]) );
  DFF \Data_Mem/memory_reg[58][8]  ( .D(\Data_Mem/n4384 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1864]), .Q(data_mem_out_wire[1864]) );
  DFF \Data_Mem/memory_reg[58][9]  ( .D(\Data_Mem/n4385 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1865]), .Q(data_mem_out_wire[1865]) );
  DFF \Data_Mem/memory_reg[58][10]  ( .D(\Data_Mem/n4386 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1866]), .Q(data_mem_out_wire[1866]) );
  DFF \Data_Mem/memory_reg[58][11]  ( .D(\Data_Mem/n4387 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1867]), .Q(data_mem_out_wire[1867]) );
  DFF \Data_Mem/memory_reg[58][12]  ( .D(\Data_Mem/n4388 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1868]), .Q(data_mem_out_wire[1868]) );
  DFF \Data_Mem/memory_reg[58][13]  ( .D(\Data_Mem/n4389 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1869]), .Q(data_mem_out_wire[1869]) );
  DFF \Data_Mem/memory_reg[58][14]  ( .D(\Data_Mem/n4390 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1870]), .Q(data_mem_out_wire[1870]) );
  DFF \Data_Mem/memory_reg[58][15]  ( .D(\Data_Mem/n4391 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1871]), .Q(data_mem_out_wire[1871]) );
  DFF \Data_Mem/memory_reg[58][16]  ( .D(\Data_Mem/n4392 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1872]), .Q(data_mem_out_wire[1872]) );
  DFF \Data_Mem/memory_reg[58][17]  ( .D(\Data_Mem/n4393 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1873]), .Q(data_mem_out_wire[1873]) );
  DFF \Data_Mem/memory_reg[58][18]  ( .D(\Data_Mem/n4394 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1874]), .Q(data_mem_out_wire[1874]) );
  DFF \Data_Mem/memory_reg[58][19]  ( .D(\Data_Mem/n4395 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1875]), .Q(data_mem_out_wire[1875]) );
  DFF \Data_Mem/memory_reg[58][20]  ( .D(\Data_Mem/n4396 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1876]), .Q(data_mem_out_wire[1876]) );
  DFF \Data_Mem/memory_reg[58][21]  ( .D(\Data_Mem/n4397 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1877]), .Q(data_mem_out_wire[1877]) );
  DFF \Data_Mem/memory_reg[58][22]  ( .D(\Data_Mem/n4398 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1878]), .Q(data_mem_out_wire[1878]) );
  DFF \Data_Mem/memory_reg[58][23]  ( .D(\Data_Mem/n4399 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1879]), .Q(data_mem_out_wire[1879]) );
  DFF \Data_Mem/memory_reg[58][24]  ( .D(\Data_Mem/n4400 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1880]), .Q(data_mem_out_wire[1880]) );
  DFF \Data_Mem/memory_reg[58][25]  ( .D(\Data_Mem/n4401 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1881]), .Q(data_mem_out_wire[1881]) );
  DFF \Data_Mem/memory_reg[58][26]  ( .D(\Data_Mem/n4402 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1882]), .Q(data_mem_out_wire[1882]) );
  DFF \Data_Mem/memory_reg[58][27]  ( .D(\Data_Mem/n4403 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1883]), .Q(data_mem_out_wire[1883]) );
  DFF \Data_Mem/memory_reg[58][28]  ( .D(\Data_Mem/n4404 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1884]), .Q(data_mem_out_wire[1884]) );
  DFF \Data_Mem/memory_reg[58][29]  ( .D(\Data_Mem/n4405 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1885]), .Q(data_mem_out_wire[1885]) );
  DFF \Data_Mem/memory_reg[58][30]  ( .D(\Data_Mem/n4406 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1886]), .Q(data_mem_out_wire[1886]) );
  DFF \Data_Mem/memory_reg[58][31]  ( .D(\Data_Mem/n4407 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1887]), .Q(data_mem_out_wire[1887]) );
  DFF \Data_Mem/memory_reg[57][0]  ( .D(\Data_Mem/n4408 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1824]), .Q(data_mem_out_wire[1824]) );
  DFF \Data_Mem/memory_reg[57][1]  ( .D(\Data_Mem/n4409 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1825]), .Q(data_mem_out_wire[1825]) );
  DFF \Data_Mem/memory_reg[57][2]  ( .D(\Data_Mem/n4410 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1826]), .Q(data_mem_out_wire[1826]) );
  DFF \Data_Mem/memory_reg[57][3]  ( .D(\Data_Mem/n4411 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1827]), .Q(data_mem_out_wire[1827]) );
  DFF \Data_Mem/memory_reg[57][4]  ( .D(\Data_Mem/n4412 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1828]), .Q(data_mem_out_wire[1828]) );
  DFF \Data_Mem/memory_reg[57][5]  ( .D(\Data_Mem/n4413 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1829]), .Q(data_mem_out_wire[1829]) );
  DFF \Data_Mem/memory_reg[57][6]  ( .D(\Data_Mem/n4414 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1830]), .Q(data_mem_out_wire[1830]) );
  DFF \Data_Mem/memory_reg[57][7]  ( .D(\Data_Mem/n4415 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1831]), .Q(data_mem_out_wire[1831]) );
  DFF \Data_Mem/memory_reg[57][8]  ( .D(\Data_Mem/n4416 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1832]), .Q(data_mem_out_wire[1832]) );
  DFF \Data_Mem/memory_reg[57][9]  ( .D(\Data_Mem/n4417 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1833]), .Q(data_mem_out_wire[1833]) );
  DFF \Data_Mem/memory_reg[57][10]  ( .D(\Data_Mem/n4418 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1834]), .Q(data_mem_out_wire[1834]) );
  DFF \Data_Mem/memory_reg[57][11]  ( .D(\Data_Mem/n4419 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1835]), .Q(data_mem_out_wire[1835]) );
  DFF \Data_Mem/memory_reg[57][12]  ( .D(\Data_Mem/n4420 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1836]), .Q(data_mem_out_wire[1836]) );
  DFF \Data_Mem/memory_reg[57][13]  ( .D(\Data_Mem/n4421 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1837]), .Q(data_mem_out_wire[1837]) );
  DFF \Data_Mem/memory_reg[57][14]  ( .D(\Data_Mem/n4422 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1838]), .Q(data_mem_out_wire[1838]) );
  DFF \Data_Mem/memory_reg[57][15]  ( .D(\Data_Mem/n4423 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1839]), .Q(data_mem_out_wire[1839]) );
  DFF \Data_Mem/memory_reg[57][16]  ( .D(\Data_Mem/n4424 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1840]), .Q(data_mem_out_wire[1840]) );
  DFF \Data_Mem/memory_reg[57][17]  ( .D(\Data_Mem/n4425 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1841]), .Q(data_mem_out_wire[1841]) );
  DFF \Data_Mem/memory_reg[57][18]  ( .D(\Data_Mem/n4426 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1842]), .Q(data_mem_out_wire[1842]) );
  DFF \Data_Mem/memory_reg[57][19]  ( .D(\Data_Mem/n4427 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1843]), .Q(data_mem_out_wire[1843]) );
  DFF \Data_Mem/memory_reg[57][20]  ( .D(\Data_Mem/n4428 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1844]), .Q(data_mem_out_wire[1844]) );
  DFF \Data_Mem/memory_reg[57][21]  ( .D(\Data_Mem/n4429 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1845]), .Q(data_mem_out_wire[1845]) );
  DFF \Data_Mem/memory_reg[57][22]  ( .D(\Data_Mem/n4430 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1846]), .Q(data_mem_out_wire[1846]) );
  DFF \Data_Mem/memory_reg[57][23]  ( .D(\Data_Mem/n4431 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1847]), .Q(data_mem_out_wire[1847]) );
  DFF \Data_Mem/memory_reg[57][24]  ( .D(\Data_Mem/n4432 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1848]), .Q(data_mem_out_wire[1848]) );
  DFF \Data_Mem/memory_reg[57][25]  ( .D(\Data_Mem/n4433 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1849]), .Q(data_mem_out_wire[1849]) );
  DFF \Data_Mem/memory_reg[57][26]  ( .D(\Data_Mem/n4434 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1850]), .Q(data_mem_out_wire[1850]) );
  DFF \Data_Mem/memory_reg[57][27]  ( .D(\Data_Mem/n4435 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1851]), .Q(data_mem_out_wire[1851]) );
  DFF \Data_Mem/memory_reg[57][28]  ( .D(\Data_Mem/n4436 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1852]), .Q(data_mem_out_wire[1852]) );
  DFF \Data_Mem/memory_reg[57][29]  ( .D(\Data_Mem/n4437 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1853]), .Q(data_mem_out_wire[1853]) );
  DFF \Data_Mem/memory_reg[57][30]  ( .D(\Data_Mem/n4438 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1854]), .Q(data_mem_out_wire[1854]) );
  DFF \Data_Mem/memory_reg[57][31]  ( .D(\Data_Mem/n4439 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1855]), .Q(data_mem_out_wire[1855]) );
  DFF \Data_Mem/memory_reg[56][0]  ( .D(\Data_Mem/n4440 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1792]), .Q(data_mem_out_wire[1792]) );
  DFF \Data_Mem/memory_reg[56][1]  ( .D(\Data_Mem/n4441 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1793]), .Q(data_mem_out_wire[1793]) );
  DFF \Data_Mem/memory_reg[56][2]  ( .D(\Data_Mem/n4442 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1794]), .Q(data_mem_out_wire[1794]) );
  DFF \Data_Mem/memory_reg[56][3]  ( .D(\Data_Mem/n4443 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1795]), .Q(data_mem_out_wire[1795]) );
  DFF \Data_Mem/memory_reg[56][4]  ( .D(\Data_Mem/n4444 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1796]), .Q(data_mem_out_wire[1796]) );
  DFF \Data_Mem/memory_reg[56][5]  ( .D(\Data_Mem/n4445 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1797]), .Q(data_mem_out_wire[1797]) );
  DFF \Data_Mem/memory_reg[56][6]  ( .D(\Data_Mem/n4446 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1798]), .Q(data_mem_out_wire[1798]) );
  DFF \Data_Mem/memory_reg[56][7]  ( .D(\Data_Mem/n4447 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1799]), .Q(data_mem_out_wire[1799]) );
  DFF \Data_Mem/memory_reg[56][8]  ( .D(\Data_Mem/n4448 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1800]), .Q(data_mem_out_wire[1800]) );
  DFF \Data_Mem/memory_reg[56][9]  ( .D(\Data_Mem/n4449 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1801]), .Q(data_mem_out_wire[1801]) );
  DFF \Data_Mem/memory_reg[56][10]  ( .D(\Data_Mem/n4450 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1802]), .Q(data_mem_out_wire[1802]) );
  DFF \Data_Mem/memory_reg[56][11]  ( .D(\Data_Mem/n4451 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1803]), .Q(data_mem_out_wire[1803]) );
  DFF \Data_Mem/memory_reg[56][12]  ( .D(\Data_Mem/n4452 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1804]), .Q(data_mem_out_wire[1804]) );
  DFF \Data_Mem/memory_reg[56][13]  ( .D(\Data_Mem/n4453 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1805]), .Q(data_mem_out_wire[1805]) );
  DFF \Data_Mem/memory_reg[56][14]  ( .D(\Data_Mem/n4454 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1806]), .Q(data_mem_out_wire[1806]) );
  DFF \Data_Mem/memory_reg[56][15]  ( .D(\Data_Mem/n4455 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1807]), .Q(data_mem_out_wire[1807]) );
  DFF \Data_Mem/memory_reg[56][16]  ( .D(\Data_Mem/n4456 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1808]), .Q(data_mem_out_wire[1808]) );
  DFF \Data_Mem/memory_reg[56][17]  ( .D(\Data_Mem/n4457 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1809]), .Q(data_mem_out_wire[1809]) );
  DFF \Data_Mem/memory_reg[56][18]  ( .D(\Data_Mem/n4458 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1810]), .Q(data_mem_out_wire[1810]) );
  DFF \Data_Mem/memory_reg[56][19]  ( .D(\Data_Mem/n4459 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1811]), .Q(data_mem_out_wire[1811]) );
  DFF \Data_Mem/memory_reg[56][20]  ( .D(\Data_Mem/n4460 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1812]), .Q(data_mem_out_wire[1812]) );
  DFF \Data_Mem/memory_reg[56][21]  ( .D(\Data_Mem/n4461 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1813]), .Q(data_mem_out_wire[1813]) );
  DFF \Data_Mem/memory_reg[56][22]  ( .D(\Data_Mem/n4462 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1814]), .Q(data_mem_out_wire[1814]) );
  DFF \Data_Mem/memory_reg[56][23]  ( .D(\Data_Mem/n4463 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1815]), .Q(data_mem_out_wire[1815]) );
  DFF \Data_Mem/memory_reg[56][24]  ( .D(\Data_Mem/n4464 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1816]), .Q(data_mem_out_wire[1816]) );
  DFF \Data_Mem/memory_reg[56][25]  ( .D(\Data_Mem/n4465 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1817]), .Q(data_mem_out_wire[1817]) );
  DFF \Data_Mem/memory_reg[56][26]  ( .D(\Data_Mem/n4466 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1818]), .Q(data_mem_out_wire[1818]) );
  DFF \Data_Mem/memory_reg[56][27]  ( .D(\Data_Mem/n4467 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1819]), .Q(data_mem_out_wire[1819]) );
  DFF \Data_Mem/memory_reg[56][28]  ( .D(\Data_Mem/n4468 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1820]), .Q(data_mem_out_wire[1820]) );
  DFF \Data_Mem/memory_reg[56][29]  ( .D(\Data_Mem/n4469 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1821]), .Q(data_mem_out_wire[1821]) );
  DFF \Data_Mem/memory_reg[56][30]  ( .D(\Data_Mem/n4470 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1822]), .Q(data_mem_out_wire[1822]) );
  DFF \Data_Mem/memory_reg[56][31]  ( .D(\Data_Mem/n4471 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1823]), .Q(data_mem_out_wire[1823]) );
  DFF \Data_Mem/memory_reg[55][0]  ( .D(\Data_Mem/n4472 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1760]), .Q(data_mem_out_wire[1760]) );
  DFF \Data_Mem/memory_reg[55][1]  ( .D(\Data_Mem/n4473 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1761]), .Q(data_mem_out_wire[1761]) );
  DFF \Data_Mem/memory_reg[55][2]  ( .D(\Data_Mem/n4474 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1762]), .Q(data_mem_out_wire[1762]) );
  DFF \Data_Mem/memory_reg[55][3]  ( .D(\Data_Mem/n4475 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1763]), .Q(data_mem_out_wire[1763]) );
  DFF \Data_Mem/memory_reg[55][4]  ( .D(\Data_Mem/n4476 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1764]), .Q(data_mem_out_wire[1764]) );
  DFF \Data_Mem/memory_reg[55][5]  ( .D(\Data_Mem/n4477 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1765]), .Q(data_mem_out_wire[1765]) );
  DFF \Data_Mem/memory_reg[55][6]  ( .D(\Data_Mem/n4478 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1766]), .Q(data_mem_out_wire[1766]) );
  DFF \Data_Mem/memory_reg[55][7]  ( .D(\Data_Mem/n4479 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1767]), .Q(data_mem_out_wire[1767]) );
  DFF \Data_Mem/memory_reg[55][8]  ( .D(\Data_Mem/n4480 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1768]), .Q(data_mem_out_wire[1768]) );
  DFF \Data_Mem/memory_reg[55][9]  ( .D(\Data_Mem/n4481 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1769]), .Q(data_mem_out_wire[1769]) );
  DFF \Data_Mem/memory_reg[55][10]  ( .D(\Data_Mem/n4482 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1770]), .Q(data_mem_out_wire[1770]) );
  DFF \Data_Mem/memory_reg[55][11]  ( .D(\Data_Mem/n4483 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1771]), .Q(data_mem_out_wire[1771]) );
  DFF \Data_Mem/memory_reg[55][12]  ( .D(\Data_Mem/n4484 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1772]), .Q(data_mem_out_wire[1772]) );
  DFF \Data_Mem/memory_reg[55][13]  ( .D(\Data_Mem/n4485 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1773]), .Q(data_mem_out_wire[1773]) );
  DFF \Data_Mem/memory_reg[55][14]  ( .D(\Data_Mem/n4486 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1774]), .Q(data_mem_out_wire[1774]) );
  DFF \Data_Mem/memory_reg[55][15]  ( .D(\Data_Mem/n4487 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1775]), .Q(data_mem_out_wire[1775]) );
  DFF \Data_Mem/memory_reg[55][16]  ( .D(\Data_Mem/n4488 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1776]), .Q(data_mem_out_wire[1776]) );
  DFF \Data_Mem/memory_reg[55][17]  ( .D(\Data_Mem/n4489 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1777]), .Q(data_mem_out_wire[1777]) );
  DFF \Data_Mem/memory_reg[55][18]  ( .D(\Data_Mem/n4490 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1778]), .Q(data_mem_out_wire[1778]) );
  DFF \Data_Mem/memory_reg[55][19]  ( .D(\Data_Mem/n4491 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1779]), .Q(data_mem_out_wire[1779]) );
  DFF \Data_Mem/memory_reg[55][20]  ( .D(\Data_Mem/n4492 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1780]), .Q(data_mem_out_wire[1780]) );
  DFF \Data_Mem/memory_reg[55][21]  ( .D(\Data_Mem/n4493 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1781]), .Q(data_mem_out_wire[1781]) );
  DFF \Data_Mem/memory_reg[55][22]  ( .D(\Data_Mem/n4494 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1782]), .Q(data_mem_out_wire[1782]) );
  DFF \Data_Mem/memory_reg[55][23]  ( .D(\Data_Mem/n4495 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1783]), .Q(data_mem_out_wire[1783]) );
  DFF \Data_Mem/memory_reg[55][24]  ( .D(\Data_Mem/n4496 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1784]), .Q(data_mem_out_wire[1784]) );
  DFF \Data_Mem/memory_reg[55][25]  ( .D(\Data_Mem/n4497 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1785]), .Q(data_mem_out_wire[1785]) );
  DFF \Data_Mem/memory_reg[55][26]  ( .D(\Data_Mem/n4498 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1786]), .Q(data_mem_out_wire[1786]) );
  DFF \Data_Mem/memory_reg[55][27]  ( .D(\Data_Mem/n4499 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1787]), .Q(data_mem_out_wire[1787]) );
  DFF \Data_Mem/memory_reg[55][28]  ( .D(\Data_Mem/n4500 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1788]), .Q(data_mem_out_wire[1788]) );
  DFF \Data_Mem/memory_reg[55][29]  ( .D(\Data_Mem/n4501 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1789]), .Q(data_mem_out_wire[1789]) );
  DFF \Data_Mem/memory_reg[55][30]  ( .D(\Data_Mem/n4502 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1790]), .Q(data_mem_out_wire[1790]) );
  DFF \Data_Mem/memory_reg[55][31]  ( .D(\Data_Mem/n4503 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1791]), .Q(data_mem_out_wire[1791]) );
  DFF \Data_Mem/memory_reg[54][0]  ( .D(\Data_Mem/n4504 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1728]), .Q(data_mem_out_wire[1728]) );
  DFF \Data_Mem/memory_reg[54][1]  ( .D(\Data_Mem/n4505 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1729]), .Q(data_mem_out_wire[1729]) );
  DFF \Data_Mem/memory_reg[54][2]  ( .D(\Data_Mem/n4506 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1730]), .Q(data_mem_out_wire[1730]) );
  DFF \Data_Mem/memory_reg[54][3]  ( .D(\Data_Mem/n4507 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1731]), .Q(data_mem_out_wire[1731]) );
  DFF \Data_Mem/memory_reg[54][4]  ( .D(\Data_Mem/n4508 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1732]), .Q(data_mem_out_wire[1732]) );
  DFF \Data_Mem/memory_reg[54][5]  ( .D(\Data_Mem/n4509 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1733]), .Q(data_mem_out_wire[1733]) );
  DFF \Data_Mem/memory_reg[54][6]  ( .D(\Data_Mem/n4510 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1734]), .Q(data_mem_out_wire[1734]) );
  DFF \Data_Mem/memory_reg[54][7]  ( .D(\Data_Mem/n4511 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1735]), .Q(data_mem_out_wire[1735]) );
  DFF \Data_Mem/memory_reg[54][8]  ( .D(\Data_Mem/n4512 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1736]), .Q(data_mem_out_wire[1736]) );
  DFF \Data_Mem/memory_reg[54][9]  ( .D(\Data_Mem/n4513 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1737]), .Q(data_mem_out_wire[1737]) );
  DFF \Data_Mem/memory_reg[54][10]  ( .D(\Data_Mem/n4514 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1738]), .Q(data_mem_out_wire[1738]) );
  DFF \Data_Mem/memory_reg[54][11]  ( .D(\Data_Mem/n4515 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1739]), .Q(data_mem_out_wire[1739]) );
  DFF \Data_Mem/memory_reg[54][12]  ( .D(\Data_Mem/n4516 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1740]), .Q(data_mem_out_wire[1740]) );
  DFF \Data_Mem/memory_reg[54][13]  ( .D(\Data_Mem/n4517 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1741]), .Q(data_mem_out_wire[1741]) );
  DFF \Data_Mem/memory_reg[54][14]  ( .D(\Data_Mem/n4518 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1742]), .Q(data_mem_out_wire[1742]) );
  DFF \Data_Mem/memory_reg[54][15]  ( .D(\Data_Mem/n4519 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1743]), .Q(data_mem_out_wire[1743]) );
  DFF \Data_Mem/memory_reg[54][16]  ( .D(\Data_Mem/n4520 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1744]), .Q(data_mem_out_wire[1744]) );
  DFF \Data_Mem/memory_reg[54][17]  ( .D(\Data_Mem/n4521 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1745]), .Q(data_mem_out_wire[1745]) );
  DFF \Data_Mem/memory_reg[54][18]  ( .D(\Data_Mem/n4522 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1746]), .Q(data_mem_out_wire[1746]) );
  DFF \Data_Mem/memory_reg[54][19]  ( .D(\Data_Mem/n4523 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1747]), .Q(data_mem_out_wire[1747]) );
  DFF \Data_Mem/memory_reg[54][20]  ( .D(\Data_Mem/n4524 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1748]), .Q(data_mem_out_wire[1748]) );
  DFF \Data_Mem/memory_reg[54][21]  ( .D(\Data_Mem/n4525 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1749]), .Q(data_mem_out_wire[1749]) );
  DFF \Data_Mem/memory_reg[54][22]  ( .D(\Data_Mem/n4526 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1750]), .Q(data_mem_out_wire[1750]) );
  DFF \Data_Mem/memory_reg[54][23]  ( .D(\Data_Mem/n4527 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1751]), .Q(data_mem_out_wire[1751]) );
  DFF \Data_Mem/memory_reg[54][24]  ( .D(\Data_Mem/n4528 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1752]), .Q(data_mem_out_wire[1752]) );
  DFF \Data_Mem/memory_reg[54][25]  ( .D(\Data_Mem/n4529 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1753]), .Q(data_mem_out_wire[1753]) );
  DFF \Data_Mem/memory_reg[54][26]  ( .D(\Data_Mem/n4530 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1754]), .Q(data_mem_out_wire[1754]) );
  DFF \Data_Mem/memory_reg[54][27]  ( .D(\Data_Mem/n4531 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1755]), .Q(data_mem_out_wire[1755]) );
  DFF \Data_Mem/memory_reg[54][28]  ( .D(\Data_Mem/n4532 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1756]), .Q(data_mem_out_wire[1756]) );
  DFF \Data_Mem/memory_reg[54][29]  ( .D(\Data_Mem/n4533 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1757]), .Q(data_mem_out_wire[1757]) );
  DFF \Data_Mem/memory_reg[54][30]  ( .D(\Data_Mem/n4534 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1758]), .Q(data_mem_out_wire[1758]) );
  DFF \Data_Mem/memory_reg[54][31]  ( .D(\Data_Mem/n4535 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1759]), .Q(data_mem_out_wire[1759]) );
  DFF \Data_Mem/memory_reg[53][0]  ( .D(\Data_Mem/n4536 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1696]), .Q(data_mem_out_wire[1696]) );
  DFF \Data_Mem/memory_reg[53][1]  ( .D(\Data_Mem/n4537 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1697]), .Q(data_mem_out_wire[1697]) );
  DFF \Data_Mem/memory_reg[53][2]  ( .D(\Data_Mem/n4538 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1698]), .Q(data_mem_out_wire[1698]) );
  DFF \Data_Mem/memory_reg[53][3]  ( .D(\Data_Mem/n4539 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1699]), .Q(data_mem_out_wire[1699]) );
  DFF \Data_Mem/memory_reg[53][4]  ( .D(\Data_Mem/n4540 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1700]), .Q(data_mem_out_wire[1700]) );
  DFF \Data_Mem/memory_reg[53][5]  ( .D(\Data_Mem/n4541 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1701]), .Q(data_mem_out_wire[1701]) );
  DFF \Data_Mem/memory_reg[53][6]  ( .D(\Data_Mem/n4542 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1702]), .Q(data_mem_out_wire[1702]) );
  DFF \Data_Mem/memory_reg[53][7]  ( .D(\Data_Mem/n4543 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1703]), .Q(data_mem_out_wire[1703]) );
  DFF \Data_Mem/memory_reg[53][8]  ( .D(\Data_Mem/n4544 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1704]), .Q(data_mem_out_wire[1704]) );
  DFF \Data_Mem/memory_reg[53][9]  ( .D(\Data_Mem/n4545 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1705]), .Q(data_mem_out_wire[1705]) );
  DFF \Data_Mem/memory_reg[53][10]  ( .D(\Data_Mem/n4546 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1706]), .Q(data_mem_out_wire[1706]) );
  DFF \Data_Mem/memory_reg[53][11]  ( .D(\Data_Mem/n4547 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1707]), .Q(data_mem_out_wire[1707]) );
  DFF \Data_Mem/memory_reg[53][12]  ( .D(\Data_Mem/n4548 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1708]), .Q(data_mem_out_wire[1708]) );
  DFF \Data_Mem/memory_reg[53][13]  ( .D(\Data_Mem/n4549 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1709]), .Q(data_mem_out_wire[1709]) );
  DFF \Data_Mem/memory_reg[53][14]  ( .D(\Data_Mem/n4550 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1710]), .Q(data_mem_out_wire[1710]) );
  DFF \Data_Mem/memory_reg[53][15]  ( .D(\Data_Mem/n4551 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1711]), .Q(data_mem_out_wire[1711]) );
  DFF \Data_Mem/memory_reg[53][16]  ( .D(\Data_Mem/n4552 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1712]), .Q(data_mem_out_wire[1712]) );
  DFF \Data_Mem/memory_reg[53][17]  ( .D(\Data_Mem/n4553 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1713]), .Q(data_mem_out_wire[1713]) );
  DFF \Data_Mem/memory_reg[53][18]  ( .D(\Data_Mem/n4554 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1714]), .Q(data_mem_out_wire[1714]) );
  DFF \Data_Mem/memory_reg[53][19]  ( .D(\Data_Mem/n4555 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1715]), .Q(data_mem_out_wire[1715]) );
  DFF \Data_Mem/memory_reg[53][20]  ( .D(\Data_Mem/n4556 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1716]), .Q(data_mem_out_wire[1716]) );
  DFF \Data_Mem/memory_reg[53][21]  ( .D(\Data_Mem/n4557 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1717]), .Q(data_mem_out_wire[1717]) );
  DFF \Data_Mem/memory_reg[53][22]  ( .D(\Data_Mem/n4558 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1718]), .Q(data_mem_out_wire[1718]) );
  DFF \Data_Mem/memory_reg[53][23]  ( .D(\Data_Mem/n4559 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1719]), .Q(data_mem_out_wire[1719]) );
  DFF \Data_Mem/memory_reg[53][24]  ( .D(\Data_Mem/n4560 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1720]), .Q(data_mem_out_wire[1720]) );
  DFF \Data_Mem/memory_reg[53][25]  ( .D(\Data_Mem/n4561 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1721]), .Q(data_mem_out_wire[1721]) );
  DFF \Data_Mem/memory_reg[53][26]  ( .D(\Data_Mem/n4562 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1722]), .Q(data_mem_out_wire[1722]) );
  DFF \Data_Mem/memory_reg[53][27]  ( .D(\Data_Mem/n4563 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1723]), .Q(data_mem_out_wire[1723]) );
  DFF \Data_Mem/memory_reg[53][28]  ( .D(\Data_Mem/n4564 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1724]), .Q(data_mem_out_wire[1724]) );
  DFF \Data_Mem/memory_reg[53][29]  ( .D(\Data_Mem/n4565 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1725]), .Q(data_mem_out_wire[1725]) );
  DFF \Data_Mem/memory_reg[53][30]  ( .D(\Data_Mem/n4566 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1726]), .Q(data_mem_out_wire[1726]) );
  DFF \Data_Mem/memory_reg[53][31]  ( .D(\Data_Mem/n4567 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1727]), .Q(data_mem_out_wire[1727]) );
  DFF \Data_Mem/memory_reg[52][0]  ( .D(\Data_Mem/n4568 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1664]), .Q(data_mem_out_wire[1664]) );
  DFF \Data_Mem/memory_reg[52][1]  ( .D(\Data_Mem/n4569 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1665]), .Q(data_mem_out_wire[1665]) );
  DFF \Data_Mem/memory_reg[52][2]  ( .D(\Data_Mem/n4570 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1666]), .Q(data_mem_out_wire[1666]) );
  DFF \Data_Mem/memory_reg[52][3]  ( .D(\Data_Mem/n4571 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1667]), .Q(data_mem_out_wire[1667]) );
  DFF \Data_Mem/memory_reg[52][4]  ( .D(\Data_Mem/n4572 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1668]), .Q(data_mem_out_wire[1668]) );
  DFF \Data_Mem/memory_reg[52][5]  ( .D(\Data_Mem/n4573 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1669]), .Q(data_mem_out_wire[1669]) );
  DFF \Data_Mem/memory_reg[52][6]  ( .D(\Data_Mem/n4574 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1670]), .Q(data_mem_out_wire[1670]) );
  DFF \Data_Mem/memory_reg[52][7]  ( .D(\Data_Mem/n4575 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1671]), .Q(data_mem_out_wire[1671]) );
  DFF \Data_Mem/memory_reg[52][8]  ( .D(\Data_Mem/n4576 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1672]), .Q(data_mem_out_wire[1672]) );
  DFF \Data_Mem/memory_reg[52][9]  ( .D(\Data_Mem/n4577 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1673]), .Q(data_mem_out_wire[1673]) );
  DFF \Data_Mem/memory_reg[52][10]  ( .D(\Data_Mem/n4578 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1674]), .Q(data_mem_out_wire[1674]) );
  DFF \Data_Mem/memory_reg[52][11]  ( .D(\Data_Mem/n4579 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1675]), .Q(data_mem_out_wire[1675]) );
  DFF \Data_Mem/memory_reg[52][12]  ( .D(\Data_Mem/n4580 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1676]), .Q(data_mem_out_wire[1676]) );
  DFF \Data_Mem/memory_reg[52][13]  ( .D(\Data_Mem/n4581 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1677]), .Q(data_mem_out_wire[1677]) );
  DFF \Data_Mem/memory_reg[52][14]  ( .D(\Data_Mem/n4582 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1678]), .Q(data_mem_out_wire[1678]) );
  DFF \Data_Mem/memory_reg[52][15]  ( .D(\Data_Mem/n4583 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1679]), .Q(data_mem_out_wire[1679]) );
  DFF \Data_Mem/memory_reg[52][16]  ( .D(\Data_Mem/n4584 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1680]), .Q(data_mem_out_wire[1680]) );
  DFF \Data_Mem/memory_reg[52][17]  ( .D(\Data_Mem/n4585 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1681]), .Q(data_mem_out_wire[1681]) );
  DFF \Data_Mem/memory_reg[52][18]  ( .D(\Data_Mem/n4586 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1682]), .Q(data_mem_out_wire[1682]) );
  DFF \Data_Mem/memory_reg[52][19]  ( .D(\Data_Mem/n4587 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1683]), .Q(data_mem_out_wire[1683]) );
  DFF \Data_Mem/memory_reg[52][20]  ( .D(\Data_Mem/n4588 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1684]), .Q(data_mem_out_wire[1684]) );
  DFF \Data_Mem/memory_reg[52][21]  ( .D(\Data_Mem/n4589 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1685]), .Q(data_mem_out_wire[1685]) );
  DFF \Data_Mem/memory_reg[52][22]  ( .D(\Data_Mem/n4590 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1686]), .Q(data_mem_out_wire[1686]) );
  DFF \Data_Mem/memory_reg[52][23]  ( .D(\Data_Mem/n4591 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1687]), .Q(data_mem_out_wire[1687]) );
  DFF \Data_Mem/memory_reg[52][24]  ( .D(\Data_Mem/n4592 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1688]), .Q(data_mem_out_wire[1688]) );
  DFF \Data_Mem/memory_reg[52][25]  ( .D(\Data_Mem/n4593 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1689]), .Q(data_mem_out_wire[1689]) );
  DFF \Data_Mem/memory_reg[52][26]  ( .D(\Data_Mem/n4594 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1690]), .Q(data_mem_out_wire[1690]) );
  DFF \Data_Mem/memory_reg[52][27]  ( .D(\Data_Mem/n4595 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1691]), .Q(data_mem_out_wire[1691]) );
  DFF \Data_Mem/memory_reg[52][28]  ( .D(\Data_Mem/n4596 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1692]), .Q(data_mem_out_wire[1692]) );
  DFF \Data_Mem/memory_reg[52][29]  ( .D(\Data_Mem/n4597 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1693]), .Q(data_mem_out_wire[1693]) );
  DFF \Data_Mem/memory_reg[52][30]  ( .D(\Data_Mem/n4598 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1694]), .Q(data_mem_out_wire[1694]) );
  DFF \Data_Mem/memory_reg[52][31]  ( .D(\Data_Mem/n4599 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1695]), .Q(data_mem_out_wire[1695]) );
  DFF \Data_Mem/memory_reg[51][0]  ( .D(\Data_Mem/n4600 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1632]), .Q(data_mem_out_wire[1632]) );
  DFF \Data_Mem/memory_reg[51][1]  ( .D(\Data_Mem/n4601 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1633]), .Q(data_mem_out_wire[1633]) );
  DFF \Data_Mem/memory_reg[51][2]  ( .D(\Data_Mem/n4602 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1634]), .Q(data_mem_out_wire[1634]) );
  DFF \Data_Mem/memory_reg[51][3]  ( .D(\Data_Mem/n4603 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1635]), .Q(data_mem_out_wire[1635]) );
  DFF \Data_Mem/memory_reg[51][4]  ( .D(\Data_Mem/n4604 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1636]), .Q(data_mem_out_wire[1636]) );
  DFF \Data_Mem/memory_reg[51][5]  ( .D(\Data_Mem/n4605 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1637]), .Q(data_mem_out_wire[1637]) );
  DFF \Data_Mem/memory_reg[51][6]  ( .D(\Data_Mem/n4606 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1638]), .Q(data_mem_out_wire[1638]) );
  DFF \Data_Mem/memory_reg[51][7]  ( .D(\Data_Mem/n4607 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1639]), .Q(data_mem_out_wire[1639]) );
  DFF \Data_Mem/memory_reg[51][8]  ( .D(\Data_Mem/n4608 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1640]), .Q(data_mem_out_wire[1640]) );
  DFF \Data_Mem/memory_reg[51][9]  ( .D(\Data_Mem/n4609 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1641]), .Q(data_mem_out_wire[1641]) );
  DFF \Data_Mem/memory_reg[51][10]  ( .D(\Data_Mem/n4610 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1642]), .Q(data_mem_out_wire[1642]) );
  DFF \Data_Mem/memory_reg[51][11]  ( .D(\Data_Mem/n4611 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1643]), .Q(data_mem_out_wire[1643]) );
  DFF \Data_Mem/memory_reg[51][12]  ( .D(\Data_Mem/n4612 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1644]), .Q(data_mem_out_wire[1644]) );
  DFF \Data_Mem/memory_reg[51][13]  ( .D(\Data_Mem/n4613 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1645]), .Q(data_mem_out_wire[1645]) );
  DFF \Data_Mem/memory_reg[51][14]  ( .D(\Data_Mem/n4614 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1646]), .Q(data_mem_out_wire[1646]) );
  DFF \Data_Mem/memory_reg[51][15]  ( .D(\Data_Mem/n4615 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1647]), .Q(data_mem_out_wire[1647]) );
  DFF \Data_Mem/memory_reg[51][16]  ( .D(\Data_Mem/n4616 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1648]), .Q(data_mem_out_wire[1648]) );
  DFF \Data_Mem/memory_reg[51][17]  ( .D(\Data_Mem/n4617 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1649]), .Q(data_mem_out_wire[1649]) );
  DFF \Data_Mem/memory_reg[51][18]  ( .D(\Data_Mem/n4618 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1650]), .Q(data_mem_out_wire[1650]) );
  DFF \Data_Mem/memory_reg[51][19]  ( .D(\Data_Mem/n4619 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1651]), .Q(data_mem_out_wire[1651]) );
  DFF \Data_Mem/memory_reg[51][20]  ( .D(\Data_Mem/n4620 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1652]), .Q(data_mem_out_wire[1652]) );
  DFF \Data_Mem/memory_reg[51][21]  ( .D(\Data_Mem/n4621 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1653]), .Q(data_mem_out_wire[1653]) );
  DFF \Data_Mem/memory_reg[51][22]  ( .D(\Data_Mem/n4622 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1654]), .Q(data_mem_out_wire[1654]) );
  DFF \Data_Mem/memory_reg[51][23]  ( .D(\Data_Mem/n4623 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1655]), .Q(data_mem_out_wire[1655]) );
  DFF \Data_Mem/memory_reg[51][24]  ( .D(\Data_Mem/n4624 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1656]), .Q(data_mem_out_wire[1656]) );
  DFF \Data_Mem/memory_reg[51][25]  ( .D(\Data_Mem/n4625 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1657]), .Q(data_mem_out_wire[1657]) );
  DFF \Data_Mem/memory_reg[51][26]  ( .D(\Data_Mem/n4626 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1658]), .Q(data_mem_out_wire[1658]) );
  DFF \Data_Mem/memory_reg[51][27]  ( .D(\Data_Mem/n4627 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1659]), .Q(data_mem_out_wire[1659]) );
  DFF \Data_Mem/memory_reg[51][28]  ( .D(\Data_Mem/n4628 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1660]), .Q(data_mem_out_wire[1660]) );
  DFF \Data_Mem/memory_reg[51][29]  ( .D(\Data_Mem/n4629 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1661]), .Q(data_mem_out_wire[1661]) );
  DFF \Data_Mem/memory_reg[51][30]  ( .D(\Data_Mem/n4630 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1662]), .Q(data_mem_out_wire[1662]) );
  DFF \Data_Mem/memory_reg[51][31]  ( .D(\Data_Mem/n4631 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1663]), .Q(data_mem_out_wire[1663]) );
  DFF \Data_Mem/memory_reg[50][0]  ( .D(\Data_Mem/n4632 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1600]), .Q(data_mem_out_wire[1600]) );
  DFF \Data_Mem/memory_reg[50][1]  ( .D(\Data_Mem/n4633 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1601]), .Q(data_mem_out_wire[1601]) );
  DFF \Data_Mem/memory_reg[50][2]  ( .D(\Data_Mem/n4634 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1602]), .Q(data_mem_out_wire[1602]) );
  DFF \Data_Mem/memory_reg[50][3]  ( .D(\Data_Mem/n4635 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1603]), .Q(data_mem_out_wire[1603]) );
  DFF \Data_Mem/memory_reg[50][4]  ( .D(\Data_Mem/n4636 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1604]), .Q(data_mem_out_wire[1604]) );
  DFF \Data_Mem/memory_reg[50][5]  ( .D(\Data_Mem/n4637 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1605]), .Q(data_mem_out_wire[1605]) );
  DFF \Data_Mem/memory_reg[50][6]  ( .D(\Data_Mem/n4638 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1606]), .Q(data_mem_out_wire[1606]) );
  DFF \Data_Mem/memory_reg[50][7]  ( .D(\Data_Mem/n4639 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1607]), .Q(data_mem_out_wire[1607]) );
  DFF \Data_Mem/memory_reg[50][8]  ( .D(\Data_Mem/n4640 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1608]), .Q(data_mem_out_wire[1608]) );
  DFF \Data_Mem/memory_reg[50][9]  ( .D(\Data_Mem/n4641 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1609]), .Q(data_mem_out_wire[1609]) );
  DFF \Data_Mem/memory_reg[50][10]  ( .D(\Data_Mem/n4642 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1610]), .Q(data_mem_out_wire[1610]) );
  DFF \Data_Mem/memory_reg[50][11]  ( .D(\Data_Mem/n4643 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1611]), .Q(data_mem_out_wire[1611]) );
  DFF \Data_Mem/memory_reg[50][12]  ( .D(\Data_Mem/n4644 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1612]), .Q(data_mem_out_wire[1612]) );
  DFF \Data_Mem/memory_reg[50][13]  ( .D(\Data_Mem/n4645 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1613]), .Q(data_mem_out_wire[1613]) );
  DFF \Data_Mem/memory_reg[50][14]  ( .D(\Data_Mem/n4646 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1614]), .Q(data_mem_out_wire[1614]) );
  DFF \Data_Mem/memory_reg[50][15]  ( .D(\Data_Mem/n4647 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1615]), .Q(data_mem_out_wire[1615]) );
  DFF \Data_Mem/memory_reg[50][16]  ( .D(\Data_Mem/n4648 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1616]), .Q(data_mem_out_wire[1616]) );
  DFF \Data_Mem/memory_reg[50][17]  ( .D(\Data_Mem/n4649 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1617]), .Q(data_mem_out_wire[1617]) );
  DFF \Data_Mem/memory_reg[50][18]  ( .D(\Data_Mem/n4650 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1618]), .Q(data_mem_out_wire[1618]) );
  DFF \Data_Mem/memory_reg[50][19]  ( .D(\Data_Mem/n4651 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1619]), .Q(data_mem_out_wire[1619]) );
  DFF \Data_Mem/memory_reg[50][20]  ( .D(\Data_Mem/n4652 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1620]), .Q(data_mem_out_wire[1620]) );
  DFF \Data_Mem/memory_reg[50][21]  ( .D(\Data_Mem/n4653 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1621]), .Q(data_mem_out_wire[1621]) );
  DFF \Data_Mem/memory_reg[50][22]  ( .D(\Data_Mem/n4654 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1622]), .Q(data_mem_out_wire[1622]) );
  DFF \Data_Mem/memory_reg[50][23]  ( .D(\Data_Mem/n4655 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1623]), .Q(data_mem_out_wire[1623]) );
  DFF \Data_Mem/memory_reg[50][24]  ( .D(\Data_Mem/n4656 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1624]), .Q(data_mem_out_wire[1624]) );
  DFF \Data_Mem/memory_reg[50][25]  ( .D(\Data_Mem/n4657 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1625]), .Q(data_mem_out_wire[1625]) );
  DFF \Data_Mem/memory_reg[50][26]  ( .D(\Data_Mem/n4658 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1626]), .Q(data_mem_out_wire[1626]) );
  DFF \Data_Mem/memory_reg[50][27]  ( .D(\Data_Mem/n4659 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1627]), .Q(data_mem_out_wire[1627]) );
  DFF \Data_Mem/memory_reg[50][28]  ( .D(\Data_Mem/n4660 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1628]), .Q(data_mem_out_wire[1628]) );
  DFF \Data_Mem/memory_reg[50][29]  ( .D(\Data_Mem/n4661 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1629]), .Q(data_mem_out_wire[1629]) );
  DFF \Data_Mem/memory_reg[50][30]  ( .D(\Data_Mem/n4662 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1630]), .Q(data_mem_out_wire[1630]) );
  DFF \Data_Mem/memory_reg[50][31]  ( .D(\Data_Mem/n4663 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1631]), .Q(data_mem_out_wire[1631]) );
  DFF \Data_Mem/memory_reg[49][0]  ( .D(\Data_Mem/n4664 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1568]), .Q(data_mem_out_wire[1568]) );
  DFF \Data_Mem/memory_reg[49][1]  ( .D(\Data_Mem/n4665 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1569]), .Q(data_mem_out_wire[1569]) );
  DFF \Data_Mem/memory_reg[49][2]  ( .D(\Data_Mem/n4666 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1570]), .Q(data_mem_out_wire[1570]) );
  DFF \Data_Mem/memory_reg[49][3]  ( .D(\Data_Mem/n4667 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1571]), .Q(data_mem_out_wire[1571]) );
  DFF \Data_Mem/memory_reg[49][4]  ( .D(\Data_Mem/n4668 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1572]), .Q(data_mem_out_wire[1572]) );
  DFF \Data_Mem/memory_reg[49][5]  ( .D(\Data_Mem/n4669 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1573]), .Q(data_mem_out_wire[1573]) );
  DFF \Data_Mem/memory_reg[49][6]  ( .D(\Data_Mem/n4670 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1574]), .Q(data_mem_out_wire[1574]) );
  DFF \Data_Mem/memory_reg[49][7]  ( .D(\Data_Mem/n4671 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1575]), .Q(data_mem_out_wire[1575]) );
  DFF \Data_Mem/memory_reg[49][8]  ( .D(\Data_Mem/n4672 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1576]), .Q(data_mem_out_wire[1576]) );
  DFF \Data_Mem/memory_reg[49][9]  ( .D(\Data_Mem/n4673 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1577]), .Q(data_mem_out_wire[1577]) );
  DFF \Data_Mem/memory_reg[49][10]  ( .D(\Data_Mem/n4674 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1578]), .Q(data_mem_out_wire[1578]) );
  DFF \Data_Mem/memory_reg[49][11]  ( .D(\Data_Mem/n4675 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1579]), .Q(data_mem_out_wire[1579]) );
  DFF \Data_Mem/memory_reg[49][12]  ( .D(\Data_Mem/n4676 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1580]), .Q(data_mem_out_wire[1580]) );
  DFF \Data_Mem/memory_reg[49][13]  ( .D(\Data_Mem/n4677 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1581]), .Q(data_mem_out_wire[1581]) );
  DFF \Data_Mem/memory_reg[49][14]  ( .D(\Data_Mem/n4678 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1582]), .Q(data_mem_out_wire[1582]) );
  DFF \Data_Mem/memory_reg[49][15]  ( .D(\Data_Mem/n4679 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1583]), .Q(data_mem_out_wire[1583]) );
  DFF \Data_Mem/memory_reg[49][16]  ( .D(\Data_Mem/n4680 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1584]), .Q(data_mem_out_wire[1584]) );
  DFF \Data_Mem/memory_reg[49][17]  ( .D(\Data_Mem/n4681 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1585]), .Q(data_mem_out_wire[1585]) );
  DFF \Data_Mem/memory_reg[49][18]  ( .D(\Data_Mem/n4682 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1586]), .Q(data_mem_out_wire[1586]) );
  DFF \Data_Mem/memory_reg[49][19]  ( .D(\Data_Mem/n4683 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1587]), .Q(data_mem_out_wire[1587]) );
  DFF \Data_Mem/memory_reg[49][20]  ( .D(\Data_Mem/n4684 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1588]), .Q(data_mem_out_wire[1588]) );
  DFF \Data_Mem/memory_reg[49][21]  ( .D(\Data_Mem/n4685 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1589]), .Q(data_mem_out_wire[1589]) );
  DFF \Data_Mem/memory_reg[49][22]  ( .D(\Data_Mem/n4686 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1590]), .Q(data_mem_out_wire[1590]) );
  DFF \Data_Mem/memory_reg[49][23]  ( .D(\Data_Mem/n4687 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1591]), .Q(data_mem_out_wire[1591]) );
  DFF \Data_Mem/memory_reg[49][24]  ( .D(\Data_Mem/n4688 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1592]), .Q(data_mem_out_wire[1592]) );
  DFF \Data_Mem/memory_reg[49][25]  ( .D(\Data_Mem/n4689 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1593]), .Q(data_mem_out_wire[1593]) );
  DFF \Data_Mem/memory_reg[49][26]  ( .D(\Data_Mem/n4690 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1594]), .Q(data_mem_out_wire[1594]) );
  DFF \Data_Mem/memory_reg[49][27]  ( .D(\Data_Mem/n4691 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1595]), .Q(data_mem_out_wire[1595]) );
  DFF \Data_Mem/memory_reg[49][28]  ( .D(\Data_Mem/n4692 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1596]), .Q(data_mem_out_wire[1596]) );
  DFF \Data_Mem/memory_reg[49][29]  ( .D(\Data_Mem/n4693 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1597]), .Q(data_mem_out_wire[1597]) );
  DFF \Data_Mem/memory_reg[49][30]  ( .D(\Data_Mem/n4694 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1598]), .Q(data_mem_out_wire[1598]) );
  DFF \Data_Mem/memory_reg[49][31]  ( .D(\Data_Mem/n4695 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1599]), .Q(data_mem_out_wire[1599]) );
  DFF \Data_Mem/memory_reg[48][0]  ( .D(\Data_Mem/n4696 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1536]), .Q(data_mem_out_wire[1536]) );
  DFF \Data_Mem/memory_reg[48][1]  ( .D(\Data_Mem/n4697 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1537]), .Q(data_mem_out_wire[1537]) );
  DFF \Data_Mem/memory_reg[48][2]  ( .D(\Data_Mem/n4698 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1538]), .Q(data_mem_out_wire[1538]) );
  DFF \Data_Mem/memory_reg[48][3]  ( .D(\Data_Mem/n4699 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1539]), .Q(data_mem_out_wire[1539]) );
  DFF \Data_Mem/memory_reg[48][4]  ( .D(\Data_Mem/n4700 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1540]), .Q(data_mem_out_wire[1540]) );
  DFF \Data_Mem/memory_reg[48][5]  ( .D(\Data_Mem/n4701 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1541]), .Q(data_mem_out_wire[1541]) );
  DFF \Data_Mem/memory_reg[48][6]  ( .D(\Data_Mem/n4702 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1542]), .Q(data_mem_out_wire[1542]) );
  DFF \Data_Mem/memory_reg[48][7]  ( .D(\Data_Mem/n4703 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1543]), .Q(data_mem_out_wire[1543]) );
  DFF \Data_Mem/memory_reg[48][8]  ( .D(\Data_Mem/n4704 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1544]), .Q(data_mem_out_wire[1544]) );
  DFF \Data_Mem/memory_reg[48][9]  ( .D(\Data_Mem/n4705 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1545]), .Q(data_mem_out_wire[1545]) );
  DFF \Data_Mem/memory_reg[48][10]  ( .D(\Data_Mem/n4706 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1546]), .Q(data_mem_out_wire[1546]) );
  DFF \Data_Mem/memory_reg[48][11]  ( .D(\Data_Mem/n4707 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1547]), .Q(data_mem_out_wire[1547]) );
  DFF \Data_Mem/memory_reg[48][12]  ( .D(\Data_Mem/n4708 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1548]), .Q(data_mem_out_wire[1548]) );
  DFF \Data_Mem/memory_reg[48][13]  ( .D(\Data_Mem/n4709 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1549]), .Q(data_mem_out_wire[1549]) );
  DFF \Data_Mem/memory_reg[48][14]  ( .D(\Data_Mem/n4710 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1550]), .Q(data_mem_out_wire[1550]) );
  DFF \Data_Mem/memory_reg[48][15]  ( .D(\Data_Mem/n4711 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1551]), .Q(data_mem_out_wire[1551]) );
  DFF \Data_Mem/memory_reg[48][16]  ( .D(\Data_Mem/n4712 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1552]), .Q(data_mem_out_wire[1552]) );
  DFF \Data_Mem/memory_reg[48][17]  ( .D(\Data_Mem/n4713 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1553]), .Q(data_mem_out_wire[1553]) );
  DFF \Data_Mem/memory_reg[48][18]  ( .D(\Data_Mem/n4714 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1554]), .Q(data_mem_out_wire[1554]) );
  DFF \Data_Mem/memory_reg[48][19]  ( .D(\Data_Mem/n4715 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1555]), .Q(data_mem_out_wire[1555]) );
  DFF \Data_Mem/memory_reg[48][20]  ( .D(\Data_Mem/n4716 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1556]), .Q(data_mem_out_wire[1556]) );
  DFF \Data_Mem/memory_reg[48][21]  ( .D(\Data_Mem/n4717 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1557]), .Q(data_mem_out_wire[1557]) );
  DFF \Data_Mem/memory_reg[48][22]  ( .D(\Data_Mem/n4718 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1558]), .Q(data_mem_out_wire[1558]) );
  DFF \Data_Mem/memory_reg[48][23]  ( .D(\Data_Mem/n4719 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1559]), .Q(data_mem_out_wire[1559]) );
  DFF \Data_Mem/memory_reg[48][24]  ( .D(\Data_Mem/n4720 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1560]), .Q(data_mem_out_wire[1560]) );
  DFF \Data_Mem/memory_reg[48][25]  ( .D(\Data_Mem/n4721 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1561]), .Q(data_mem_out_wire[1561]) );
  DFF \Data_Mem/memory_reg[48][26]  ( .D(\Data_Mem/n4722 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1562]), .Q(data_mem_out_wire[1562]) );
  DFF \Data_Mem/memory_reg[48][27]  ( .D(\Data_Mem/n4723 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1563]), .Q(data_mem_out_wire[1563]) );
  DFF \Data_Mem/memory_reg[48][28]  ( .D(\Data_Mem/n4724 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1564]), .Q(data_mem_out_wire[1564]) );
  DFF \Data_Mem/memory_reg[48][29]  ( .D(\Data_Mem/n4725 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1565]), .Q(data_mem_out_wire[1565]) );
  DFF \Data_Mem/memory_reg[48][30]  ( .D(\Data_Mem/n4726 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1566]), .Q(data_mem_out_wire[1566]) );
  DFF \Data_Mem/memory_reg[48][31]  ( .D(\Data_Mem/n4727 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1567]), .Q(data_mem_out_wire[1567]) );
  DFF \Data_Mem/memory_reg[47][0]  ( .D(\Data_Mem/n4728 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1504]), .Q(data_mem_out_wire[1504]) );
  DFF \Data_Mem/memory_reg[47][1]  ( .D(\Data_Mem/n4729 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1505]), .Q(data_mem_out_wire[1505]) );
  DFF \Data_Mem/memory_reg[47][2]  ( .D(\Data_Mem/n4730 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1506]), .Q(data_mem_out_wire[1506]) );
  DFF \Data_Mem/memory_reg[47][3]  ( .D(\Data_Mem/n4731 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1507]), .Q(data_mem_out_wire[1507]) );
  DFF \Data_Mem/memory_reg[47][4]  ( .D(\Data_Mem/n4732 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1508]), .Q(data_mem_out_wire[1508]) );
  DFF \Data_Mem/memory_reg[47][5]  ( .D(\Data_Mem/n4733 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1509]), .Q(data_mem_out_wire[1509]) );
  DFF \Data_Mem/memory_reg[47][6]  ( .D(\Data_Mem/n4734 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1510]), .Q(data_mem_out_wire[1510]) );
  DFF \Data_Mem/memory_reg[47][7]  ( .D(\Data_Mem/n4735 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1511]), .Q(data_mem_out_wire[1511]) );
  DFF \Data_Mem/memory_reg[47][8]  ( .D(\Data_Mem/n4736 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1512]), .Q(data_mem_out_wire[1512]) );
  DFF \Data_Mem/memory_reg[47][9]  ( .D(\Data_Mem/n4737 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1513]), .Q(data_mem_out_wire[1513]) );
  DFF \Data_Mem/memory_reg[47][10]  ( .D(\Data_Mem/n4738 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1514]), .Q(data_mem_out_wire[1514]) );
  DFF \Data_Mem/memory_reg[47][11]  ( .D(\Data_Mem/n4739 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1515]), .Q(data_mem_out_wire[1515]) );
  DFF \Data_Mem/memory_reg[47][12]  ( .D(\Data_Mem/n4740 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1516]), .Q(data_mem_out_wire[1516]) );
  DFF \Data_Mem/memory_reg[47][13]  ( .D(\Data_Mem/n4741 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1517]), .Q(data_mem_out_wire[1517]) );
  DFF \Data_Mem/memory_reg[47][14]  ( .D(\Data_Mem/n4742 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1518]), .Q(data_mem_out_wire[1518]) );
  DFF \Data_Mem/memory_reg[47][15]  ( .D(\Data_Mem/n4743 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1519]), .Q(data_mem_out_wire[1519]) );
  DFF \Data_Mem/memory_reg[47][16]  ( .D(\Data_Mem/n4744 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1520]), .Q(data_mem_out_wire[1520]) );
  DFF \Data_Mem/memory_reg[47][17]  ( .D(\Data_Mem/n4745 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1521]), .Q(data_mem_out_wire[1521]) );
  DFF \Data_Mem/memory_reg[47][18]  ( .D(\Data_Mem/n4746 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1522]), .Q(data_mem_out_wire[1522]) );
  DFF \Data_Mem/memory_reg[47][19]  ( .D(\Data_Mem/n4747 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1523]), .Q(data_mem_out_wire[1523]) );
  DFF \Data_Mem/memory_reg[47][20]  ( .D(\Data_Mem/n4748 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1524]), .Q(data_mem_out_wire[1524]) );
  DFF \Data_Mem/memory_reg[47][21]  ( .D(\Data_Mem/n4749 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1525]), .Q(data_mem_out_wire[1525]) );
  DFF \Data_Mem/memory_reg[47][22]  ( .D(\Data_Mem/n4750 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1526]), .Q(data_mem_out_wire[1526]) );
  DFF \Data_Mem/memory_reg[47][23]  ( .D(\Data_Mem/n4751 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1527]), .Q(data_mem_out_wire[1527]) );
  DFF \Data_Mem/memory_reg[47][24]  ( .D(\Data_Mem/n4752 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1528]), .Q(data_mem_out_wire[1528]) );
  DFF \Data_Mem/memory_reg[47][25]  ( .D(\Data_Mem/n4753 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1529]), .Q(data_mem_out_wire[1529]) );
  DFF \Data_Mem/memory_reg[47][26]  ( .D(\Data_Mem/n4754 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1530]), .Q(data_mem_out_wire[1530]) );
  DFF \Data_Mem/memory_reg[47][27]  ( .D(\Data_Mem/n4755 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1531]), .Q(data_mem_out_wire[1531]) );
  DFF \Data_Mem/memory_reg[47][28]  ( .D(\Data_Mem/n4756 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1532]), .Q(data_mem_out_wire[1532]) );
  DFF \Data_Mem/memory_reg[47][29]  ( .D(\Data_Mem/n4757 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1533]), .Q(data_mem_out_wire[1533]) );
  DFF \Data_Mem/memory_reg[47][30]  ( .D(\Data_Mem/n4758 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1534]), .Q(data_mem_out_wire[1534]) );
  DFF \Data_Mem/memory_reg[47][31]  ( .D(\Data_Mem/n4759 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1535]), .Q(data_mem_out_wire[1535]) );
  DFF \Data_Mem/memory_reg[46][0]  ( .D(\Data_Mem/n4760 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1472]), .Q(data_mem_out_wire[1472]) );
  DFF \Data_Mem/memory_reg[46][1]  ( .D(\Data_Mem/n4761 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1473]), .Q(data_mem_out_wire[1473]) );
  DFF \Data_Mem/memory_reg[46][2]  ( .D(\Data_Mem/n4762 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1474]), .Q(data_mem_out_wire[1474]) );
  DFF \Data_Mem/memory_reg[46][3]  ( .D(\Data_Mem/n4763 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1475]), .Q(data_mem_out_wire[1475]) );
  DFF \Data_Mem/memory_reg[46][4]  ( .D(\Data_Mem/n4764 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1476]), .Q(data_mem_out_wire[1476]) );
  DFF \Data_Mem/memory_reg[46][5]  ( .D(\Data_Mem/n4765 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1477]), .Q(data_mem_out_wire[1477]) );
  DFF \Data_Mem/memory_reg[46][6]  ( .D(\Data_Mem/n4766 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1478]), .Q(data_mem_out_wire[1478]) );
  DFF \Data_Mem/memory_reg[46][7]  ( .D(\Data_Mem/n4767 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1479]), .Q(data_mem_out_wire[1479]) );
  DFF \Data_Mem/memory_reg[46][8]  ( .D(\Data_Mem/n4768 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1480]), .Q(data_mem_out_wire[1480]) );
  DFF \Data_Mem/memory_reg[46][9]  ( .D(\Data_Mem/n4769 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1481]), .Q(data_mem_out_wire[1481]) );
  DFF \Data_Mem/memory_reg[46][10]  ( .D(\Data_Mem/n4770 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1482]), .Q(data_mem_out_wire[1482]) );
  DFF \Data_Mem/memory_reg[46][11]  ( .D(\Data_Mem/n4771 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1483]), .Q(data_mem_out_wire[1483]) );
  DFF \Data_Mem/memory_reg[46][12]  ( .D(\Data_Mem/n4772 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1484]), .Q(data_mem_out_wire[1484]) );
  DFF \Data_Mem/memory_reg[46][13]  ( .D(\Data_Mem/n4773 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1485]), .Q(data_mem_out_wire[1485]) );
  DFF \Data_Mem/memory_reg[46][14]  ( .D(\Data_Mem/n4774 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1486]), .Q(data_mem_out_wire[1486]) );
  DFF \Data_Mem/memory_reg[46][15]  ( .D(\Data_Mem/n4775 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1487]), .Q(data_mem_out_wire[1487]) );
  DFF \Data_Mem/memory_reg[46][16]  ( .D(\Data_Mem/n4776 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1488]), .Q(data_mem_out_wire[1488]) );
  DFF \Data_Mem/memory_reg[46][17]  ( .D(\Data_Mem/n4777 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1489]), .Q(data_mem_out_wire[1489]) );
  DFF \Data_Mem/memory_reg[46][18]  ( .D(\Data_Mem/n4778 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1490]), .Q(data_mem_out_wire[1490]) );
  DFF \Data_Mem/memory_reg[46][19]  ( .D(\Data_Mem/n4779 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1491]), .Q(data_mem_out_wire[1491]) );
  DFF \Data_Mem/memory_reg[46][20]  ( .D(\Data_Mem/n4780 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1492]), .Q(data_mem_out_wire[1492]) );
  DFF \Data_Mem/memory_reg[46][21]  ( .D(\Data_Mem/n4781 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1493]), .Q(data_mem_out_wire[1493]) );
  DFF \Data_Mem/memory_reg[46][22]  ( .D(\Data_Mem/n4782 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1494]), .Q(data_mem_out_wire[1494]) );
  DFF \Data_Mem/memory_reg[46][23]  ( .D(\Data_Mem/n4783 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1495]), .Q(data_mem_out_wire[1495]) );
  DFF \Data_Mem/memory_reg[46][24]  ( .D(\Data_Mem/n4784 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1496]), .Q(data_mem_out_wire[1496]) );
  DFF \Data_Mem/memory_reg[46][25]  ( .D(\Data_Mem/n4785 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1497]), .Q(data_mem_out_wire[1497]) );
  DFF \Data_Mem/memory_reg[46][26]  ( .D(\Data_Mem/n4786 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1498]), .Q(data_mem_out_wire[1498]) );
  DFF \Data_Mem/memory_reg[46][27]  ( .D(\Data_Mem/n4787 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1499]), .Q(data_mem_out_wire[1499]) );
  DFF \Data_Mem/memory_reg[46][28]  ( .D(\Data_Mem/n4788 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1500]), .Q(data_mem_out_wire[1500]) );
  DFF \Data_Mem/memory_reg[46][29]  ( .D(\Data_Mem/n4789 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1501]), .Q(data_mem_out_wire[1501]) );
  DFF \Data_Mem/memory_reg[46][30]  ( .D(\Data_Mem/n4790 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1502]), .Q(data_mem_out_wire[1502]) );
  DFF \Data_Mem/memory_reg[46][31]  ( .D(\Data_Mem/n4791 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1503]), .Q(data_mem_out_wire[1503]) );
  DFF \Data_Mem/memory_reg[45][0]  ( .D(\Data_Mem/n4792 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1440]), .Q(data_mem_out_wire[1440]) );
  DFF \Data_Mem/memory_reg[45][1]  ( .D(\Data_Mem/n4793 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1441]), .Q(data_mem_out_wire[1441]) );
  DFF \Data_Mem/memory_reg[45][2]  ( .D(\Data_Mem/n4794 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1442]), .Q(data_mem_out_wire[1442]) );
  DFF \Data_Mem/memory_reg[45][3]  ( .D(\Data_Mem/n4795 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1443]), .Q(data_mem_out_wire[1443]) );
  DFF \Data_Mem/memory_reg[45][4]  ( .D(\Data_Mem/n4796 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1444]), .Q(data_mem_out_wire[1444]) );
  DFF \Data_Mem/memory_reg[45][5]  ( .D(\Data_Mem/n4797 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1445]), .Q(data_mem_out_wire[1445]) );
  DFF \Data_Mem/memory_reg[45][6]  ( .D(\Data_Mem/n4798 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1446]), .Q(data_mem_out_wire[1446]) );
  DFF \Data_Mem/memory_reg[45][7]  ( .D(\Data_Mem/n4799 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1447]), .Q(data_mem_out_wire[1447]) );
  DFF \Data_Mem/memory_reg[45][8]  ( .D(\Data_Mem/n4800 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1448]), .Q(data_mem_out_wire[1448]) );
  DFF \Data_Mem/memory_reg[45][9]  ( .D(\Data_Mem/n4801 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1449]), .Q(data_mem_out_wire[1449]) );
  DFF \Data_Mem/memory_reg[45][10]  ( .D(\Data_Mem/n4802 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1450]), .Q(data_mem_out_wire[1450]) );
  DFF \Data_Mem/memory_reg[45][11]  ( .D(\Data_Mem/n4803 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1451]), .Q(data_mem_out_wire[1451]) );
  DFF \Data_Mem/memory_reg[45][12]  ( .D(\Data_Mem/n4804 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1452]), .Q(data_mem_out_wire[1452]) );
  DFF \Data_Mem/memory_reg[45][13]  ( .D(\Data_Mem/n4805 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1453]), .Q(data_mem_out_wire[1453]) );
  DFF \Data_Mem/memory_reg[45][14]  ( .D(\Data_Mem/n4806 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1454]), .Q(data_mem_out_wire[1454]) );
  DFF \Data_Mem/memory_reg[45][15]  ( .D(\Data_Mem/n4807 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1455]), .Q(data_mem_out_wire[1455]) );
  DFF \Data_Mem/memory_reg[45][16]  ( .D(\Data_Mem/n4808 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1456]), .Q(data_mem_out_wire[1456]) );
  DFF \Data_Mem/memory_reg[45][17]  ( .D(\Data_Mem/n4809 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1457]), .Q(data_mem_out_wire[1457]) );
  DFF \Data_Mem/memory_reg[45][18]  ( .D(\Data_Mem/n4810 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1458]), .Q(data_mem_out_wire[1458]) );
  DFF \Data_Mem/memory_reg[45][19]  ( .D(\Data_Mem/n4811 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1459]), .Q(data_mem_out_wire[1459]) );
  DFF \Data_Mem/memory_reg[45][20]  ( .D(\Data_Mem/n4812 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1460]), .Q(data_mem_out_wire[1460]) );
  DFF \Data_Mem/memory_reg[45][21]  ( .D(\Data_Mem/n4813 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1461]), .Q(data_mem_out_wire[1461]) );
  DFF \Data_Mem/memory_reg[45][22]  ( .D(\Data_Mem/n4814 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1462]), .Q(data_mem_out_wire[1462]) );
  DFF \Data_Mem/memory_reg[45][23]  ( .D(\Data_Mem/n4815 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1463]), .Q(data_mem_out_wire[1463]) );
  DFF \Data_Mem/memory_reg[45][24]  ( .D(\Data_Mem/n4816 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1464]), .Q(data_mem_out_wire[1464]) );
  DFF \Data_Mem/memory_reg[45][25]  ( .D(\Data_Mem/n4817 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1465]), .Q(data_mem_out_wire[1465]) );
  DFF \Data_Mem/memory_reg[45][26]  ( .D(\Data_Mem/n4818 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1466]), .Q(data_mem_out_wire[1466]) );
  DFF \Data_Mem/memory_reg[45][27]  ( .D(\Data_Mem/n4819 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1467]), .Q(data_mem_out_wire[1467]) );
  DFF \Data_Mem/memory_reg[45][28]  ( .D(\Data_Mem/n4820 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1468]), .Q(data_mem_out_wire[1468]) );
  DFF \Data_Mem/memory_reg[45][29]  ( .D(\Data_Mem/n4821 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1469]), .Q(data_mem_out_wire[1469]) );
  DFF \Data_Mem/memory_reg[45][30]  ( .D(\Data_Mem/n4822 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1470]), .Q(data_mem_out_wire[1470]) );
  DFF \Data_Mem/memory_reg[45][31]  ( .D(\Data_Mem/n4823 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1471]), .Q(data_mem_out_wire[1471]) );
  DFF \Data_Mem/memory_reg[44][0]  ( .D(\Data_Mem/n4824 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1408]), .Q(data_mem_out_wire[1408]) );
  DFF \Data_Mem/memory_reg[44][1]  ( .D(\Data_Mem/n4825 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1409]), .Q(data_mem_out_wire[1409]) );
  DFF \Data_Mem/memory_reg[44][2]  ( .D(\Data_Mem/n4826 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1410]), .Q(data_mem_out_wire[1410]) );
  DFF \Data_Mem/memory_reg[44][3]  ( .D(\Data_Mem/n4827 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1411]), .Q(data_mem_out_wire[1411]) );
  DFF \Data_Mem/memory_reg[44][4]  ( .D(\Data_Mem/n4828 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1412]), .Q(data_mem_out_wire[1412]) );
  DFF \Data_Mem/memory_reg[44][5]  ( .D(\Data_Mem/n4829 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1413]), .Q(data_mem_out_wire[1413]) );
  DFF \Data_Mem/memory_reg[44][6]  ( .D(\Data_Mem/n4830 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1414]), .Q(data_mem_out_wire[1414]) );
  DFF \Data_Mem/memory_reg[44][7]  ( .D(\Data_Mem/n4831 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1415]), .Q(data_mem_out_wire[1415]) );
  DFF \Data_Mem/memory_reg[44][8]  ( .D(\Data_Mem/n4832 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1416]), .Q(data_mem_out_wire[1416]) );
  DFF \Data_Mem/memory_reg[44][9]  ( .D(\Data_Mem/n4833 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1417]), .Q(data_mem_out_wire[1417]) );
  DFF \Data_Mem/memory_reg[44][10]  ( .D(\Data_Mem/n4834 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1418]), .Q(data_mem_out_wire[1418]) );
  DFF \Data_Mem/memory_reg[44][11]  ( .D(\Data_Mem/n4835 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1419]), .Q(data_mem_out_wire[1419]) );
  DFF \Data_Mem/memory_reg[44][12]  ( .D(\Data_Mem/n4836 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1420]), .Q(data_mem_out_wire[1420]) );
  DFF \Data_Mem/memory_reg[44][13]  ( .D(\Data_Mem/n4837 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1421]), .Q(data_mem_out_wire[1421]) );
  DFF \Data_Mem/memory_reg[44][14]  ( .D(\Data_Mem/n4838 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1422]), .Q(data_mem_out_wire[1422]) );
  DFF \Data_Mem/memory_reg[44][15]  ( .D(\Data_Mem/n4839 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1423]), .Q(data_mem_out_wire[1423]) );
  DFF \Data_Mem/memory_reg[44][16]  ( .D(\Data_Mem/n4840 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1424]), .Q(data_mem_out_wire[1424]) );
  DFF \Data_Mem/memory_reg[44][17]  ( .D(\Data_Mem/n4841 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1425]), .Q(data_mem_out_wire[1425]) );
  DFF \Data_Mem/memory_reg[44][18]  ( .D(\Data_Mem/n4842 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1426]), .Q(data_mem_out_wire[1426]) );
  DFF \Data_Mem/memory_reg[44][19]  ( .D(\Data_Mem/n4843 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1427]), .Q(data_mem_out_wire[1427]) );
  DFF \Data_Mem/memory_reg[44][20]  ( .D(\Data_Mem/n4844 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1428]), .Q(data_mem_out_wire[1428]) );
  DFF \Data_Mem/memory_reg[44][21]  ( .D(\Data_Mem/n4845 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1429]), .Q(data_mem_out_wire[1429]) );
  DFF \Data_Mem/memory_reg[44][22]  ( .D(\Data_Mem/n4846 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1430]), .Q(data_mem_out_wire[1430]) );
  DFF \Data_Mem/memory_reg[44][23]  ( .D(\Data_Mem/n4847 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1431]), .Q(data_mem_out_wire[1431]) );
  DFF \Data_Mem/memory_reg[44][24]  ( .D(\Data_Mem/n4848 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1432]), .Q(data_mem_out_wire[1432]) );
  DFF \Data_Mem/memory_reg[44][25]  ( .D(\Data_Mem/n4849 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1433]), .Q(data_mem_out_wire[1433]) );
  DFF \Data_Mem/memory_reg[44][26]  ( .D(\Data_Mem/n4850 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1434]), .Q(data_mem_out_wire[1434]) );
  DFF \Data_Mem/memory_reg[44][27]  ( .D(\Data_Mem/n4851 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1435]), .Q(data_mem_out_wire[1435]) );
  DFF \Data_Mem/memory_reg[44][28]  ( .D(\Data_Mem/n4852 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1436]), .Q(data_mem_out_wire[1436]) );
  DFF \Data_Mem/memory_reg[44][29]  ( .D(\Data_Mem/n4853 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1437]), .Q(data_mem_out_wire[1437]) );
  DFF \Data_Mem/memory_reg[44][30]  ( .D(\Data_Mem/n4854 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1438]), .Q(data_mem_out_wire[1438]) );
  DFF \Data_Mem/memory_reg[44][31]  ( .D(\Data_Mem/n4855 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1439]), .Q(data_mem_out_wire[1439]) );
  DFF \Data_Mem/memory_reg[43][0]  ( .D(\Data_Mem/n4856 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1376]), .Q(data_mem_out_wire[1376]) );
  DFF \Data_Mem/memory_reg[43][1]  ( .D(\Data_Mem/n4857 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1377]), .Q(data_mem_out_wire[1377]) );
  DFF \Data_Mem/memory_reg[43][2]  ( .D(\Data_Mem/n4858 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1378]), .Q(data_mem_out_wire[1378]) );
  DFF \Data_Mem/memory_reg[43][3]  ( .D(\Data_Mem/n4859 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1379]), .Q(data_mem_out_wire[1379]) );
  DFF \Data_Mem/memory_reg[43][4]  ( .D(\Data_Mem/n4860 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1380]), .Q(data_mem_out_wire[1380]) );
  DFF \Data_Mem/memory_reg[43][5]  ( .D(\Data_Mem/n4861 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1381]), .Q(data_mem_out_wire[1381]) );
  DFF \Data_Mem/memory_reg[43][6]  ( .D(\Data_Mem/n4862 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1382]), .Q(data_mem_out_wire[1382]) );
  DFF \Data_Mem/memory_reg[43][7]  ( .D(\Data_Mem/n4863 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1383]), .Q(data_mem_out_wire[1383]) );
  DFF \Data_Mem/memory_reg[43][8]  ( .D(\Data_Mem/n4864 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1384]), .Q(data_mem_out_wire[1384]) );
  DFF \Data_Mem/memory_reg[43][9]  ( .D(\Data_Mem/n4865 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1385]), .Q(data_mem_out_wire[1385]) );
  DFF \Data_Mem/memory_reg[43][10]  ( .D(\Data_Mem/n4866 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1386]), .Q(data_mem_out_wire[1386]) );
  DFF \Data_Mem/memory_reg[43][11]  ( .D(\Data_Mem/n4867 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1387]), .Q(data_mem_out_wire[1387]) );
  DFF \Data_Mem/memory_reg[43][12]  ( .D(\Data_Mem/n4868 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1388]), .Q(data_mem_out_wire[1388]) );
  DFF \Data_Mem/memory_reg[43][13]  ( .D(\Data_Mem/n4869 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1389]), .Q(data_mem_out_wire[1389]) );
  DFF \Data_Mem/memory_reg[43][14]  ( .D(\Data_Mem/n4870 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1390]), .Q(data_mem_out_wire[1390]) );
  DFF \Data_Mem/memory_reg[43][15]  ( .D(\Data_Mem/n4871 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1391]), .Q(data_mem_out_wire[1391]) );
  DFF \Data_Mem/memory_reg[43][16]  ( .D(\Data_Mem/n4872 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1392]), .Q(data_mem_out_wire[1392]) );
  DFF \Data_Mem/memory_reg[43][17]  ( .D(\Data_Mem/n4873 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1393]), .Q(data_mem_out_wire[1393]) );
  DFF \Data_Mem/memory_reg[43][18]  ( .D(\Data_Mem/n4874 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1394]), .Q(data_mem_out_wire[1394]) );
  DFF \Data_Mem/memory_reg[43][19]  ( .D(\Data_Mem/n4875 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1395]), .Q(data_mem_out_wire[1395]) );
  DFF \Data_Mem/memory_reg[43][20]  ( .D(\Data_Mem/n4876 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1396]), .Q(data_mem_out_wire[1396]) );
  DFF \Data_Mem/memory_reg[43][21]  ( .D(\Data_Mem/n4877 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1397]), .Q(data_mem_out_wire[1397]) );
  DFF \Data_Mem/memory_reg[43][22]  ( .D(\Data_Mem/n4878 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1398]), .Q(data_mem_out_wire[1398]) );
  DFF \Data_Mem/memory_reg[43][23]  ( .D(\Data_Mem/n4879 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1399]), .Q(data_mem_out_wire[1399]) );
  DFF \Data_Mem/memory_reg[43][24]  ( .D(\Data_Mem/n4880 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1400]), .Q(data_mem_out_wire[1400]) );
  DFF \Data_Mem/memory_reg[43][25]  ( .D(\Data_Mem/n4881 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1401]), .Q(data_mem_out_wire[1401]) );
  DFF \Data_Mem/memory_reg[43][26]  ( .D(\Data_Mem/n4882 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1402]), .Q(data_mem_out_wire[1402]) );
  DFF \Data_Mem/memory_reg[43][27]  ( .D(\Data_Mem/n4883 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1403]), .Q(data_mem_out_wire[1403]) );
  DFF \Data_Mem/memory_reg[43][28]  ( .D(\Data_Mem/n4884 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1404]), .Q(data_mem_out_wire[1404]) );
  DFF \Data_Mem/memory_reg[43][29]  ( .D(\Data_Mem/n4885 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1405]), .Q(data_mem_out_wire[1405]) );
  DFF \Data_Mem/memory_reg[43][30]  ( .D(\Data_Mem/n4886 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1406]), .Q(data_mem_out_wire[1406]) );
  DFF \Data_Mem/memory_reg[43][31]  ( .D(\Data_Mem/n4887 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1407]), .Q(data_mem_out_wire[1407]) );
  DFF \Data_Mem/memory_reg[42][0]  ( .D(\Data_Mem/n4888 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1344]), .Q(data_mem_out_wire[1344]) );
  DFF \Data_Mem/memory_reg[42][1]  ( .D(\Data_Mem/n4889 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1345]), .Q(data_mem_out_wire[1345]) );
  DFF \Data_Mem/memory_reg[42][2]  ( .D(\Data_Mem/n4890 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1346]), .Q(data_mem_out_wire[1346]) );
  DFF \Data_Mem/memory_reg[42][3]  ( .D(\Data_Mem/n4891 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1347]), .Q(data_mem_out_wire[1347]) );
  DFF \Data_Mem/memory_reg[42][4]  ( .D(\Data_Mem/n4892 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1348]), .Q(data_mem_out_wire[1348]) );
  DFF \Data_Mem/memory_reg[42][5]  ( .D(\Data_Mem/n4893 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1349]), .Q(data_mem_out_wire[1349]) );
  DFF \Data_Mem/memory_reg[42][6]  ( .D(\Data_Mem/n4894 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1350]), .Q(data_mem_out_wire[1350]) );
  DFF \Data_Mem/memory_reg[42][7]  ( .D(\Data_Mem/n4895 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1351]), .Q(data_mem_out_wire[1351]) );
  DFF \Data_Mem/memory_reg[42][8]  ( .D(\Data_Mem/n4896 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1352]), .Q(data_mem_out_wire[1352]) );
  DFF \Data_Mem/memory_reg[42][9]  ( .D(\Data_Mem/n4897 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1353]), .Q(data_mem_out_wire[1353]) );
  DFF \Data_Mem/memory_reg[42][10]  ( .D(\Data_Mem/n4898 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1354]), .Q(data_mem_out_wire[1354]) );
  DFF \Data_Mem/memory_reg[42][11]  ( .D(\Data_Mem/n4899 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1355]), .Q(data_mem_out_wire[1355]) );
  DFF \Data_Mem/memory_reg[42][12]  ( .D(\Data_Mem/n4900 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1356]), .Q(data_mem_out_wire[1356]) );
  DFF \Data_Mem/memory_reg[42][13]  ( .D(\Data_Mem/n4901 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1357]), .Q(data_mem_out_wire[1357]) );
  DFF \Data_Mem/memory_reg[42][14]  ( .D(\Data_Mem/n4902 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1358]), .Q(data_mem_out_wire[1358]) );
  DFF \Data_Mem/memory_reg[42][15]  ( .D(\Data_Mem/n4903 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1359]), .Q(data_mem_out_wire[1359]) );
  DFF \Data_Mem/memory_reg[42][16]  ( .D(\Data_Mem/n4904 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1360]), .Q(data_mem_out_wire[1360]) );
  DFF \Data_Mem/memory_reg[42][17]  ( .D(\Data_Mem/n4905 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1361]), .Q(data_mem_out_wire[1361]) );
  DFF \Data_Mem/memory_reg[42][18]  ( .D(\Data_Mem/n4906 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1362]), .Q(data_mem_out_wire[1362]) );
  DFF \Data_Mem/memory_reg[42][19]  ( .D(\Data_Mem/n4907 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1363]), .Q(data_mem_out_wire[1363]) );
  DFF \Data_Mem/memory_reg[42][20]  ( .D(\Data_Mem/n4908 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1364]), .Q(data_mem_out_wire[1364]) );
  DFF \Data_Mem/memory_reg[42][21]  ( .D(\Data_Mem/n4909 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1365]), .Q(data_mem_out_wire[1365]) );
  DFF \Data_Mem/memory_reg[42][22]  ( .D(\Data_Mem/n4910 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1366]), .Q(data_mem_out_wire[1366]) );
  DFF \Data_Mem/memory_reg[42][23]  ( .D(\Data_Mem/n4911 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1367]), .Q(data_mem_out_wire[1367]) );
  DFF \Data_Mem/memory_reg[42][24]  ( .D(\Data_Mem/n4912 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1368]), .Q(data_mem_out_wire[1368]) );
  DFF \Data_Mem/memory_reg[42][25]  ( .D(\Data_Mem/n4913 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1369]), .Q(data_mem_out_wire[1369]) );
  DFF \Data_Mem/memory_reg[42][26]  ( .D(\Data_Mem/n4914 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1370]), .Q(data_mem_out_wire[1370]) );
  DFF \Data_Mem/memory_reg[42][27]  ( .D(\Data_Mem/n4915 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1371]), .Q(data_mem_out_wire[1371]) );
  DFF \Data_Mem/memory_reg[42][28]  ( .D(\Data_Mem/n4916 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1372]), .Q(data_mem_out_wire[1372]) );
  DFF \Data_Mem/memory_reg[42][29]  ( .D(\Data_Mem/n4917 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1373]), .Q(data_mem_out_wire[1373]) );
  DFF \Data_Mem/memory_reg[42][30]  ( .D(\Data_Mem/n4918 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1374]), .Q(data_mem_out_wire[1374]) );
  DFF \Data_Mem/memory_reg[42][31]  ( .D(\Data_Mem/n4919 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1375]), .Q(data_mem_out_wire[1375]) );
  DFF \Data_Mem/memory_reg[41][0]  ( .D(\Data_Mem/n4920 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1312]), .Q(data_mem_out_wire[1312]) );
  DFF \Data_Mem/memory_reg[41][1]  ( .D(\Data_Mem/n4921 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1313]), .Q(data_mem_out_wire[1313]) );
  DFF \Data_Mem/memory_reg[41][2]  ( .D(\Data_Mem/n4922 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1314]), .Q(data_mem_out_wire[1314]) );
  DFF \Data_Mem/memory_reg[41][3]  ( .D(\Data_Mem/n4923 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1315]), .Q(data_mem_out_wire[1315]) );
  DFF \Data_Mem/memory_reg[41][4]  ( .D(\Data_Mem/n4924 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1316]), .Q(data_mem_out_wire[1316]) );
  DFF \Data_Mem/memory_reg[41][5]  ( .D(\Data_Mem/n4925 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1317]), .Q(data_mem_out_wire[1317]) );
  DFF \Data_Mem/memory_reg[41][6]  ( .D(\Data_Mem/n4926 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1318]), .Q(data_mem_out_wire[1318]) );
  DFF \Data_Mem/memory_reg[41][7]  ( .D(\Data_Mem/n4927 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1319]), .Q(data_mem_out_wire[1319]) );
  DFF \Data_Mem/memory_reg[41][8]  ( .D(\Data_Mem/n4928 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1320]), .Q(data_mem_out_wire[1320]) );
  DFF \Data_Mem/memory_reg[41][9]  ( .D(\Data_Mem/n4929 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1321]), .Q(data_mem_out_wire[1321]) );
  DFF \Data_Mem/memory_reg[41][10]  ( .D(\Data_Mem/n4930 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1322]), .Q(data_mem_out_wire[1322]) );
  DFF \Data_Mem/memory_reg[41][11]  ( .D(\Data_Mem/n4931 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1323]), .Q(data_mem_out_wire[1323]) );
  DFF \Data_Mem/memory_reg[41][12]  ( .D(\Data_Mem/n4932 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1324]), .Q(data_mem_out_wire[1324]) );
  DFF \Data_Mem/memory_reg[41][13]  ( .D(\Data_Mem/n4933 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1325]), .Q(data_mem_out_wire[1325]) );
  DFF \Data_Mem/memory_reg[41][14]  ( .D(\Data_Mem/n4934 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1326]), .Q(data_mem_out_wire[1326]) );
  DFF \Data_Mem/memory_reg[41][15]  ( .D(\Data_Mem/n4935 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1327]), .Q(data_mem_out_wire[1327]) );
  DFF \Data_Mem/memory_reg[41][16]  ( .D(\Data_Mem/n4936 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1328]), .Q(data_mem_out_wire[1328]) );
  DFF \Data_Mem/memory_reg[41][17]  ( .D(\Data_Mem/n4937 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1329]), .Q(data_mem_out_wire[1329]) );
  DFF \Data_Mem/memory_reg[41][18]  ( .D(\Data_Mem/n4938 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1330]), .Q(data_mem_out_wire[1330]) );
  DFF \Data_Mem/memory_reg[41][19]  ( .D(\Data_Mem/n4939 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1331]), .Q(data_mem_out_wire[1331]) );
  DFF \Data_Mem/memory_reg[41][20]  ( .D(\Data_Mem/n4940 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1332]), .Q(data_mem_out_wire[1332]) );
  DFF \Data_Mem/memory_reg[41][21]  ( .D(\Data_Mem/n4941 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1333]), .Q(data_mem_out_wire[1333]) );
  DFF \Data_Mem/memory_reg[41][22]  ( .D(\Data_Mem/n4942 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1334]), .Q(data_mem_out_wire[1334]) );
  DFF \Data_Mem/memory_reg[41][23]  ( .D(\Data_Mem/n4943 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1335]), .Q(data_mem_out_wire[1335]) );
  DFF \Data_Mem/memory_reg[41][24]  ( .D(\Data_Mem/n4944 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1336]), .Q(data_mem_out_wire[1336]) );
  DFF \Data_Mem/memory_reg[41][25]  ( .D(\Data_Mem/n4945 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1337]), .Q(data_mem_out_wire[1337]) );
  DFF \Data_Mem/memory_reg[41][26]  ( .D(\Data_Mem/n4946 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1338]), .Q(data_mem_out_wire[1338]) );
  DFF \Data_Mem/memory_reg[41][27]  ( .D(\Data_Mem/n4947 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1339]), .Q(data_mem_out_wire[1339]) );
  DFF \Data_Mem/memory_reg[41][28]  ( .D(\Data_Mem/n4948 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1340]), .Q(data_mem_out_wire[1340]) );
  DFF \Data_Mem/memory_reg[41][29]  ( .D(\Data_Mem/n4949 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1341]), .Q(data_mem_out_wire[1341]) );
  DFF \Data_Mem/memory_reg[41][30]  ( .D(\Data_Mem/n4950 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1342]), .Q(data_mem_out_wire[1342]) );
  DFF \Data_Mem/memory_reg[41][31]  ( .D(\Data_Mem/n4951 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1343]), .Q(data_mem_out_wire[1343]) );
  DFF \Data_Mem/memory_reg[40][0]  ( .D(\Data_Mem/n4952 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1280]), .Q(data_mem_out_wire[1280]) );
  DFF \Data_Mem/memory_reg[40][1]  ( .D(\Data_Mem/n4953 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1281]), .Q(data_mem_out_wire[1281]) );
  DFF \Data_Mem/memory_reg[40][2]  ( .D(\Data_Mem/n4954 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1282]), .Q(data_mem_out_wire[1282]) );
  DFF \Data_Mem/memory_reg[40][3]  ( .D(\Data_Mem/n4955 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1283]), .Q(data_mem_out_wire[1283]) );
  DFF \Data_Mem/memory_reg[40][4]  ( .D(\Data_Mem/n4956 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1284]), .Q(data_mem_out_wire[1284]) );
  DFF \Data_Mem/memory_reg[40][5]  ( .D(\Data_Mem/n4957 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1285]), .Q(data_mem_out_wire[1285]) );
  DFF \Data_Mem/memory_reg[40][6]  ( .D(\Data_Mem/n4958 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1286]), .Q(data_mem_out_wire[1286]) );
  DFF \Data_Mem/memory_reg[40][7]  ( .D(\Data_Mem/n4959 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1287]), .Q(data_mem_out_wire[1287]) );
  DFF \Data_Mem/memory_reg[40][8]  ( .D(\Data_Mem/n4960 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1288]), .Q(data_mem_out_wire[1288]) );
  DFF \Data_Mem/memory_reg[40][9]  ( .D(\Data_Mem/n4961 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1289]), .Q(data_mem_out_wire[1289]) );
  DFF \Data_Mem/memory_reg[40][10]  ( .D(\Data_Mem/n4962 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1290]), .Q(data_mem_out_wire[1290]) );
  DFF \Data_Mem/memory_reg[40][11]  ( .D(\Data_Mem/n4963 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1291]), .Q(data_mem_out_wire[1291]) );
  DFF \Data_Mem/memory_reg[40][12]  ( .D(\Data_Mem/n4964 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1292]), .Q(data_mem_out_wire[1292]) );
  DFF \Data_Mem/memory_reg[40][13]  ( .D(\Data_Mem/n4965 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1293]), .Q(data_mem_out_wire[1293]) );
  DFF \Data_Mem/memory_reg[40][14]  ( .D(\Data_Mem/n4966 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1294]), .Q(data_mem_out_wire[1294]) );
  DFF \Data_Mem/memory_reg[40][15]  ( .D(\Data_Mem/n4967 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1295]), .Q(data_mem_out_wire[1295]) );
  DFF \Data_Mem/memory_reg[40][16]  ( .D(\Data_Mem/n4968 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1296]), .Q(data_mem_out_wire[1296]) );
  DFF \Data_Mem/memory_reg[40][17]  ( .D(\Data_Mem/n4969 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1297]), .Q(data_mem_out_wire[1297]) );
  DFF \Data_Mem/memory_reg[40][18]  ( .D(\Data_Mem/n4970 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1298]), .Q(data_mem_out_wire[1298]) );
  DFF \Data_Mem/memory_reg[40][19]  ( .D(\Data_Mem/n4971 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1299]), .Q(data_mem_out_wire[1299]) );
  DFF \Data_Mem/memory_reg[40][20]  ( .D(\Data_Mem/n4972 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1300]), .Q(data_mem_out_wire[1300]) );
  DFF \Data_Mem/memory_reg[40][21]  ( .D(\Data_Mem/n4973 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1301]), .Q(data_mem_out_wire[1301]) );
  DFF \Data_Mem/memory_reg[40][22]  ( .D(\Data_Mem/n4974 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1302]), .Q(data_mem_out_wire[1302]) );
  DFF \Data_Mem/memory_reg[40][23]  ( .D(\Data_Mem/n4975 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1303]), .Q(data_mem_out_wire[1303]) );
  DFF \Data_Mem/memory_reg[40][24]  ( .D(\Data_Mem/n4976 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1304]), .Q(data_mem_out_wire[1304]) );
  DFF \Data_Mem/memory_reg[40][25]  ( .D(\Data_Mem/n4977 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1305]), .Q(data_mem_out_wire[1305]) );
  DFF \Data_Mem/memory_reg[40][26]  ( .D(\Data_Mem/n4978 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1306]), .Q(data_mem_out_wire[1306]) );
  DFF \Data_Mem/memory_reg[40][27]  ( .D(\Data_Mem/n4979 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1307]), .Q(data_mem_out_wire[1307]) );
  DFF \Data_Mem/memory_reg[40][28]  ( .D(\Data_Mem/n4980 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1308]), .Q(data_mem_out_wire[1308]) );
  DFF \Data_Mem/memory_reg[40][29]  ( .D(\Data_Mem/n4981 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1309]), .Q(data_mem_out_wire[1309]) );
  DFF \Data_Mem/memory_reg[40][30]  ( .D(\Data_Mem/n4982 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1310]), .Q(data_mem_out_wire[1310]) );
  DFF \Data_Mem/memory_reg[40][31]  ( .D(\Data_Mem/n4983 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1311]), .Q(data_mem_out_wire[1311]) );
  DFF \Data_Mem/memory_reg[39][0]  ( .D(\Data_Mem/n4984 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1248]), .Q(data_mem_out_wire[1248]) );
  DFF \Data_Mem/memory_reg[39][1]  ( .D(\Data_Mem/n4985 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1249]), .Q(data_mem_out_wire[1249]) );
  DFF \Data_Mem/memory_reg[39][2]  ( .D(\Data_Mem/n4986 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1250]), .Q(data_mem_out_wire[1250]) );
  DFF \Data_Mem/memory_reg[39][3]  ( .D(\Data_Mem/n4987 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1251]), .Q(data_mem_out_wire[1251]) );
  DFF \Data_Mem/memory_reg[39][4]  ( .D(\Data_Mem/n4988 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1252]), .Q(data_mem_out_wire[1252]) );
  DFF \Data_Mem/memory_reg[39][5]  ( .D(\Data_Mem/n4989 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1253]), .Q(data_mem_out_wire[1253]) );
  DFF \Data_Mem/memory_reg[39][6]  ( .D(\Data_Mem/n4990 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1254]), .Q(data_mem_out_wire[1254]) );
  DFF \Data_Mem/memory_reg[39][7]  ( .D(\Data_Mem/n4991 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1255]), .Q(data_mem_out_wire[1255]) );
  DFF \Data_Mem/memory_reg[39][8]  ( .D(\Data_Mem/n4992 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1256]), .Q(data_mem_out_wire[1256]) );
  DFF \Data_Mem/memory_reg[39][9]  ( .D(\Data_Mem/n4993 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1257]), .Q(data_mem_out_wire[1257]) );
  DFF \Data_Mem/memory_reg[39][10]  ( .D(\Data_Mem/n4994 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1258]), .Q(data_mem_out_wire[1258]) );
  DFF \Data_Mem/memory_reg[39][11]  ( .D(\Data_Mem/n4995 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1259]), .Q(data_mem_out_wire[1259]) );
  DFF \Data_Mem/memory_reg[39][12]  ( .D(\Data_Mem/n4996 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1260]), .Q(data_mem_out_wire[1260]) );
  DFF \Data_Mem/memory_reg[39][13]  ( .D(\Data_Mem/n4997 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1261]), .Q(data_mem_out_wire[1261]) );
  DFF \Data_Mem/memory_reg[39][14]  ( .D(\Data_Mem/n4998 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1262]), .Q(data_mem_out_wire[1262]) );
  DFF \Data_Mem/memory_reg[39][15]  ( .D(\Data_Mem/n4999 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1263]), .Q(data_mem_out_wire[1263]) );
  DFF \Data_Mem/memory_reg[39][16]  ( .D(\Data_Mem/n5000 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1264]), .Q(data_mem_out_wire[1264]) );
  DFF \Data_Mem/memory_reg[39][17]  ( .D(\Data_Mem/n5001 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1265]), .Q(data_mem_out_wire[1265]) );
  DFF \Data_Mem/memory_reg[39][18]  ( .D(\Data_Mem/n5002 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1266]), .Q(data_mem_out_wire[1266]) );
  DFF \Data_Mem/memory_reg[39][19]  ( .D(\Data_Mem/n5003 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1267]), .Q(data_mem_out_wire[1267]) );
  DFF \Data_Mem/memory_reg[39][20]  ( .D(\Data_Mem/n5004 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1268]), .Q(data_mem_out_wire[1268]) );
  DFF \Data_Mem/memory_reg[39][21]  ( .D(\Data_Mem/n5005 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1269]), .Q(data_mem_out_wire[1269]) );
  DFF \Data_Mem/memory_reg[39][22]  ( .D(\Data_Mem/n5006 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1270]), .Q(data_mem_out_wire[1270]) );
  DFF \Data_Mem/memory_reg[39][23]  ( .D(\Data_Mem/n5007 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1271]), .Q(data_mem_out_wire[1271]) );
  DFF \Data_Mem/memory_reg[39][24]  ( .D(\Data_Mem/n5008 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1272]), .Q(data_mem_out_wire[1272]) );
  DFF \Data_Mem/memory_reg[39][25]  ( .D(\Data_Mem/n5009 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1273]), .Q(data_mem_out_wire[1273]) );
  DFF \Data_Mem/memory_reg[39][26]  ( .D(\Data_Mem/n5010 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1274]), .Q(data_mem_out_wire[1274]) );
  DFF \Data_Mem/memory_reg[39][27]  ( .D(\Data_Mem/n5011 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1275]), .Q(data_mem_out_wire[1275]) );
  DFF \Data_Mem/memory_reg[39][28]  ( .D(\Data_Mem/n5012 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1276]), .Q(data_mem_out_wire[1276]) );
  DFF \Data_Mem/memory_reg[39][29]  ( .D(\Data_Mem/n5013 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1277]), .Q(data_mem_out_wire[1277]) );
  DFF \Data_Mem/memory_reg[39][30]  ( .D(\Data_Mem/n5014 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1278]), .Q(data_mem_out_wire[1278]) );
  DFF \Data_Mem/memory_reg[39][31]  ( .D(\Data_Mem/n5015 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1279]), .Q(data_mem_out_wire[1279]) );
  DFF \Data_Mem/memory_reg[38][0]  ( .D(\Data_Mem/n5016 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1216]), .Q(data_mem_out_wire[1216]) );
  DFF \Data_Mem/memory_reg[38][1]  ( .D(\Data_Mem/n5017 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1217]), .Q(data_mem_out_wire[1217]) );
  DFF \Data_Mem/memory_reg[38][2]  ( .D(\Data_Mem/n5018 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1218]), .Q(data_mem_out_wire[1218]) );
  DFF \Data_Mem/memory_reg[38][3]  ( .D(\Data_Mem/n5019 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1219]), .Q(data_mem_out_wire[1219]) );
  DFF \Data_Mem/memory_reg[38][4]  ( .D(\Data_Mem/n5020 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1220]), .Q(data_mem_out_wire[1220]) );
  DFF \Data_Mem/memory_reg[38][5]  ( .D(\Data_Mem/n5021 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1221]), .Q(data_mem_out_wire[1221]) );
  DFF \Data_Mem/memory_reg[38][6]  ( .D(\Data_Mem/n5022 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1222]), .Q(data_mem_out_wire[1222]) );
  DFF \Data_Mem/memory_reg[38][7]  ( .D(\Data_Mem/n5023 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1223]), .Q(data_mem_out_wire[1223]) );
  DFF \Data_Mem/memory_reg[38][8]  ( .D(\Data_Mem/n5024 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1224]), .Q(data_mem_out_wire[1224]) );
  DFF \Data_Mem/memory_reg[38][9]  ( .D(\Data_Mem/n5025 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1225]), .Q(data_mem_out_wire[1225]) );
  DFF \Data_Mem/memory_reg[38][10]  ( .D(\Data_Mem/n5026 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1226]), .Q(data_mem_out_wire[1226]) );
  DFF \Data_Mem/memory_reg[38][11]  ( .D(\Data_Mem/n5027 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1227]), .Q(data_mem_out_wire[1227]) );
  DFF \Data_Mem/memory_reg[38][12]  ( .D(\Data_Mem/n5028 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1228]), .Q(data_mem_out_wire[1228]) );
  DFF \Data_Mem/memory_reg[38][13]  ( .D(\Data_Mem/n5029 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1229]), .Q(data_mem_out_wire[1229]) );
  DFF \Data_Mem/memory_reg[38][14]  ( .D(\Data_Mem/n5030 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1230]), .Q(data_mem_out_wire[1230]) );
  DFF \Data_Mem/memory_reg[38][15]  ( .D(\Data_Mem/n5031 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1231]), .Q(data_mem_out_wire[1231]) );
  DFF \Data_Mem/memory_reg[38][16]  ( .D(\Data_Mem/n5032 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1232]), .Q(data_mem_out_wire[1232]) );
  DFF \Data_Mem/memory_reg[38][17]  ( .D(\Data_Mem/n5033 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1233]), .Q(data_mem_out_wire[1233]) );
  DFF \Data_Mem/memory_reg[38][18]  ( .D(\Data_Mem/n5034 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1234]), .Q(data_mem_out_wire[1234]) );
  DFF \Data_Mem/memory_reg[38][19]  ( .D(\Data_Mem/n5035 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1235]), .Q(data_mem_out_wire[1235]) );
  DFF \Data_Mem/memory_reg[38][20]  ( .D(\Data_Mem/n5036 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1236]), .Q(data_mem_out_wire[1236]) );
  DFF \Data_Mem/memory_reg[38][21]  ( .D(\Data_Mem/n5037 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1237]), .Q(data_mem_out_wire[1237]) );
  DFF \Data_Mem/memory_reg[38][22]  ( .D(\Data_Mem/n5038 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1238]), .Q(data_mem_out_wire[1238]) );
  DFF \Data_Mem/memory_reg[38][23]  ( .D(\Data_Mem/n5039 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1239]), .Q(data_mem_out_wire[1239]) );
  DFF \Data_Mem/memory_reg[38][24]  ( .D(\Data_Mem/n5040 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1240]), .Q(data_mem_out_wire[1240]) );
  DFF \Data_Mem/memory_reg[38][25]  ( .D(\Data_Mem/n5041 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1241]), .Q(data_mem_out_wire[1241]) );
  DFF \Data_Mem/memory_reg[38][26]  ( .D(\Data_Mem/n5042 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1242]), .Q(data_mem_out_wire[1242]) );
  DFF \Data_Mem/memory_reg[38][27]  ( .D(\Data_Mem/n5043 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1243]), .Q(data_mem_out_wire[1243]) );
  DFF \Data_Mem/memory_reg[38][28]  ( .D(\Data_Mem/n5044 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1244]), .Q(data_mem_out_wire[1244]) );
  DFF \Data_Mem/memory_reg[38][29]  ( .D(\Data_Mem/n5045 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1245]), .Q(data_mem_out_wire[1245]) );
  DFF \Data_Mem/memory_reg[38][30]  ( .D(\Data_Mem/n5046 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1246]), .Q(data_mem_out_wire[1246]) );
  DFF \Data_Mem/memory_reg[38][31]  ( .D(\Data_Mem/n5047 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1247]), .Q(data_mem_out_wire[1247]) );
  DFF \Data_Mem/memory_reg[37][0]  ( .D(\Data_Mem/n5048 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1184]), .Q(data_mem_out_wire[1184]) );
  DFF \Data_Mem/memory_reg[37][1]  ( .D(\Data_Mem/n5049 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1185]), .Q(data_mem_out_wire[1185]) );
  DFF \Data_Mem/memory_reg[37][2]  ( .D(\Data_Mem/n5050 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1186]), .Q(data_mem_out_wire[1186]) );
  DFF \Data_Mem/memory_reg[37][3]  ( .D(\Data_Mem/n5051 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1187]), .Q(data_mem_out_wire[1187]) );
  DFF \Data_Mem/memory_reg[37][4]  ( .D(\Data_Mem/n5052 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1188]), .Q(data_mem_out_wire[1188]) );
  DFF \Data_Mem/memory_reg[37][5]  ( .D(\Data_Mem/n5053 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1189]), .Q(data_mem_out_wire[1189]) );
  DFF \Data_Mem/memory_reg[37][6]  ( .D(\Data_Mem/n5054 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1190]), .Q(data_mem_out_wire[1190]) );
  DFF \Data_Mem/memory_reg[37][7]  ( .D(\Data_Mem/n5055 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1191]), .Q(data_mem_out_wire[1191]) );
  DFF \Data_Mem/memory_reg[37][8]  ( .D(\Data_Mem/n5056 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1192]), .Q(data_mem_out_wire[1192]) );
  DFF \Data_Mem/memory_reg[37][9]  ( .D(\Data_Mem/n5057 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1193]), .Q(data_mem_out_wire[1193]) );
  DFF \Data_Mem/memory_reg[37][10]  ( .D(\Data_Mem/n5058 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1194]), .Q(data_mem_out_wire[1194]) );
  DFF \Data_Mem/memory_reg[37][11]  ( .D(\Data_Mem/n5059 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1195]), .Q(data_mem_out_wire[1195]) );
  DFF \Data_Mem/memory_reg[37][12]  ( .D(\Data_Mem/n5060 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1196]), .Q(data_mem_out_wire[1196]) );
  DFF \Data_Mem/memory_reg[37][13]  ( .D(\Data_Mem/n5061 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1197]), .Q(data_mem_out_wire[1197]) );
  DFF \Data_Mem/memory_reg[37][14]  ( .D(\Data_Mem/n5062 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1198]), .Q(data_mem_out_wire[1198]) );
  DFF \Data_Mem/memory_reg[37][15]  ( .D(\Data_Mem/n5063 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1199]), .Q(data_mem_out_wire[1199]) );
  DFF \Data_Mem/memory_reg[37][16]  ( .D(\Data_Mem/n5064 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1200]), .Q(data_mem_out_wire[1200]) );
  DFF \Data_Mem/memory_reg[37][17]  ( .D(\Data_Mem/n5065 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1201]), .Q(data_mem_out_wire[1201]) );
  DFF \Data_Mem/memory_reg[37][18]  ( .D(\Data_Mem/n5066 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1202]), .Q(data_mem_out_wire[1202]) );
  DFF \Data_Mem/memory_reg[37][19]  ( .D(\Data_Mem/n5067 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1203]), .Q(data_mem_out_wire[1203]) );
  DFF \Data_Mem/memory_reg[37][20]  ( .D(\Data_Mem/n5068 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1204]), .Q(data_mem_out_wire[1204]) );
  DFF \Data_Mem/memory_reg[37][21]  ( .D(\Data_Mem/n5069 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1205]), .Q(data_mem_out_wire[1205]) );
  DFF \Data_Mem/memory_reg[37][22]  ( .D(\Data_Mem/n5070 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1206]), .Q(data_mem_out_wire[1206]) );
  DFF \Data_Mem/memory_reg[37][23]  ( .D(\Data_Mem/n5071 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1207]), .Q(data_mem_out_wire[1207]) );
  DFF \Data_Mem/memory_reg[37][24]  ( .D(\Data_Mem/n5072 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1208]), .Q(data_mem_out_wire[1208]) );
  DFF \Data_Mem/memory_reg[37][25]  ( .D(\Data_Mem/n5073 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1209]), .Q(data_mem_out_wire[1209]) );
  DFF \Data_Mem/memory_reg[37][26]  ( .D(\Data_Mem/n5074 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1210]), .Q(data_mem_out_wire[1210]) );
  DFF \Data_Mem/memory_reg[37][27]  ( .D(\Data_Mem/n5075 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1211]), .Q(data_mem_out_wire[1211]) );
  DFF \Data_Mem/memory_reg[37][28]  ( .D(\Data_Mem/n5076 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1212]), .Q(data_mem_out_wire[1212]) );
  DFF \Data_Mem/memory_reg[37][29]  ( .D(\Data_Mem/n5077 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1213]), .Q(data_mem_out_wire[1213]) );
  DFF \Data_Mem/memory_reg[37][30]  ( .D(\Data_Mem/n5078 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1214]), .Q(data_mem_out_wire[1214]) );
  DFF \Data_Mem/memory_reg[37][31]  ( .D(\Data_Mem/n5079 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1215]), .Q(data_mem_out_wire[1215]) );
  DFF \Data_Mem/memory_reg[36][0]  ( .D(\Data_Mem/n5080 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1152]), .Q(data_mem_out_wire[1152]) );
  DFF \Data_Mem/memory_reg[36][1]  ( .D(\Data_Mem/n5081 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1153]), .Q(data_mem_out_wire[1153]) );
  DFF \Data_Mem/memory_reg[36][2]  ( .D(\Data_Mem/n5082 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1154]), .Q(data_mem_out_wire[1154]) );
  DFF \Data_Mem/memory_reg[36][3]  ( .D(\Data_Mem/n5083 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1155]), .Q(data_mem_out_wire[1155]) );
  DFF \Data_Mem/memory_reg[36][4]  ( .D(\Data_Mem/n5084 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1156]), .Q(data_mem_out_wire[1156]) );
  DFF \Data_Mem/memory_reg[36][5]  ( .D(\Data_Mem/n5085 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1157]), .Q(data_mem_out_wire[1157]) );
  DFF \Data_Mem/memory_reg[36][6]  ( .D(\Data_Mem/n5086 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1158]), .Q(data_mem_out_wire[1158]) );
  DFF \Data_Mem/memory_reg[36][7]  ( .D(\Data_Mem/n5087 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1159]), .Q(data_mem_out_wire[1159]) );
  DFF \Data_Mem/memory_reg[36][8]  ( .D(\Data_Mem/n5088 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1160]), .Q(data_mem_out_wire[1160]) );
  DFF \Data_Mem/memory_reg[36][9]  ( .D(\Data_Mem/n5089 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1161]), .Q(data_mem_out_wire[1161]) );
  DFF \Data_Mem/memory_reg[36][10]  ( .D(\Data_Mem/n5090 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1162]), .Q(data_mem_out_wire[1162]) );
  DFF \Data_Mem/memory_reg[36][11]  ( .D(\Data_Mem/n5091 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1163]), .Q(data_mem_out_wire[1163]) );
  DFF \Data_Mem/memory_reg[36][12]  ( .D(\Data_Mem/n5092 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1164]), .Q(data_mem_out_wire[1164]) );
  DFF \Data_Mem/memory_reg[36][13]  ( .D(\Data_Mem/n5093 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1165]), .Q(data_mem_out_wire[1165]) );
  DFF \Data_Mem/memory_reg[36][14]  ( .D(\Data_Mem/n5094 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1166]), .Q(data_mem_out_wire[1166]) );
  DFF \Data_Mem/memory_reg[36][15]  ( .D(\Data_Mem/n5095 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1167]), .Q(data_mem_out_wire[1167]) );
  DFF \Data_Mem/memory_reg[36][16]  ( .D(\Data_Mem/n5096 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1168]), .Q(data_mem_out_wire[1168]) );
  DFF \Data_Mem/memory_reg[36][17]  ( .D(\Data_Mem/n5097 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1169]), .Q(data_mem_out_wire[1169]) );
  DFF \Data_Mem/memory_reg[36][18]  ( .D(\Data_Mem/n5098 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1170]), .Q(data_mem_out_wire[1170]) );
  DFF \Data_Mem/memory_reg[36][19]  ( .D(\Data_Mem/n5099 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1171]), .Q(data_mem_out_wire[1171]) );
  DFF \Data_Mem/memory_reg[36][20]  ( .D(\Data_Mem/n5100 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1172]), .Q(data_mem_out_wire[1172]) );
  DFF \Data_Mem/memory_reg[36][21]  ( .D(\Data_Mem/n5101 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1173]), .Q(data_mem_out_wire[1173]) );
  DFF \Data_Mem/memory_reg[36][22]  ( .D(\Data_Mem/n5102 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1174]), .Q(data_mem_out_wire[1174]) );
  DFF \Data_Mem/memory_reg[36][23]  ( .D(\Data_Mem/n5103 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1175]), .Q(data_mem_out_wire[1175]) );
  DFF \Data_Mem/memory_reg[36][24]  ( .D(\Data_Mem/n5104 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1176]), .Q(data_mem_out_wire[1176]) );
  DFF \Data_Mem/memory_reg[36][25]  ( .D(\Data_Mem/n5105 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1177]), .Q(data_mem_out_wire[1177]) );
  DFF \Data_Mem/memory_reg[36][26]  ( .D(\Data_Mem/n5106 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1178]), .Q(data_mem_out_wire[1178]) );
  DFF \Data_Mem/memory_reg[36][27]  ( .D(\Data_Mem/n5107 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1179]), .Q(data_mem_out_wire[1179]) );
  DFF \Data_Mem/memory_reg[36][28]  ( .D(\Data_Mem/n5108 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1180]), .Q(data_mem_out_wire[1180]) );
  DFF \Data_Mem/memory_reg[36][29]  ( .D(\Data_Mem/n5109 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1181]), .Q(data_mem_out_wire[1181]) );
  DFF \Data_Mem/memory_reg[36][30]  ( .D(\Data_Mem/n5110 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1182]), .Q(data_mem_out_wire[1182]) );
  DFF \Data_Mem/memory_reg[36][31]  ( .D(\Data_Mem/n5111 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1183]), .Q(data_mem_out_wire[1183]) );
  DFF \Data_Mem/memory_reg[35][0]  ( .D(\Data_Mem/n5112 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1120]), .Q(data_mem_out_wire[1120]) );
  DFF \Data_Mem/memory_reg[35][1]  ( .D(\Data_Mem/n5113 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1121]), .Q(data_mem_out_wire[1121]) );
  DFF \Data_Mem/memory_reg[35][2]  ( .D(\Data_Mem/n5114 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1122]), .Q(data_mem_out_wire[1122]) );
  DFF \Data_Mem/memory_reg[35][3]  ( .D(\Data_Mem/n5115 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1123]), .Q(data_mem_out_wire[1123]) );
  DFF \Data_Mem/memory_reg[35][4]  ( .D(\Data_Mem/n5116 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1124]), .Q(data_mem_out_wire[1124]) );
  DFF \Data_Mem/memory_reg[35][5]  ( .D(\Data_Mem/n5117 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1125]), .Q(data_mem_out_wire[1125]) );
  DFF \Data_Mem/memory_reg[35][6]  ( .D(\Data_Mem/n5118 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1126]), .Q(data_mem_out_wire[1126]) );
  DFF \Data_Mem/memory_reg[35][7]  ( .D(\Data_Mem/n5119 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1127]), .Q(data_mem_out_wire[1127]) );
  DFF \Data_Mem/memory_reg[35][8]  ( .D(\Data_Mem/n5120 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1128]), .Q(data_mem_out_wire[1128]) );
  DFF \Data_Mem/memory_reg[35][9]  ( .D(\Data_Mem/n5121 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1129]), .Q(data_mem_out_wire[1129]) );
  DFF \Data_Mem/memory_reg[35][10]  ( .D(\Data_Mem/n5122 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1130]), .Q(data_mem_out_wire[1130]) );
  DFF \Data_Mem/memory_reg[35][11]  ( .D(\Data_Mem/n5123 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1131]), .Q(data_mem_out_wire[1131]) );
  DFF \Data_Mem/memory_reg[35][12]  ( .D(\Data_Mem/n5124 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1132]), .Q(data_mem_out_wire[1132]) );
  DFF \Data_Mem/memory_reg[35][13]  ( .D(\Data_Mem/n5125 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1133]), .Q(data_mem_out_wire[1133]) );
  DFF \Data_Mem/memory_reg[35][14]  ( .D(\Data_Mem/n5126 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1134]), .Q(data_mem_out_wire[1134]) );
  DFF \Data_Mem/memory_reg[35][15]  ( .D(\Data_Mem/n5127 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1135]), .Q(data_mem_out_wire[1135]) );
  DFF \Data_Mem/memory_reg[35][16]  ( .D(\Data_Mem/n5128 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1136]), .Q(data_mem_out_wire[1136]) );
  DFF \Data_Mem/memory_reg[35][17]  ( .D(\Data_Mem/n5129 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1137]), .Q(data_mem_out_wire[1137]) );
  DFF \Data_Mem/memory_reg[35][18]  ( .D(\Data_Mem/n5130 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1138]), .Q(data_mem_out_wire[1138]) );
  DFF \Data_Mem/memory_reg[35][19]  ( .D(\Data_Mem/n5131 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1139]), .Q(data_mem_out_wire[1139]) );
  DFF \Data_Mem/memory_reg[35][20]  ( .D(\Data_Mem/n5132 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1140]), .Q(data_mem_out_wire[1140]) );
  DFF \Data_Mem/memory_reg[35][21]  ( .D(\Data_Mem/n5133 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1141]), .Q(data_mem_out_wire[1141]) );
  DFF \Data_Mem/memory_reg[35][22]  ( .D(\Data_Mem/n5134 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1142]), .Q(data_mem_out_wire[1142]) );
  DFF \Data_Mem/memory_reg[35][23]  ( .D(\Data_Mem/n5135 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1143]), .Q(data_mem_out_wire[1143]) );
  DFF \Data_Mem/memory_reg[35][24]  ( .D(\Data_Mem/n5136 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1144]), .Q(data_mem_out_wire[1144]) );
  DFF \Data_Mem/memory_reg[35][25]  ( .D(\Data_Mem/n5137 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1145]), .Q(data_mem_out_wire[1145]) );
  DFF \Data_Mem/memory_reg[35][26]  ( .D(\Data_Mem/n5138 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1146]), .Q(data_mem_out_wire[1146]) );
  DFF \Data_Mem/memory_reg[35][27]  ( .D(\Data_Mem/n5139 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1147]), .Q(data_mem_out_wire[1147]) );
  DFF \Data_Mem/memory_reg[35][28]  ( .D(\Data_Mem/n5140 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1148]), .Q(data_mem_out_wire[1148]) );
  DFF \Data_Mem/memory_reg[35][29]  ( .D(\Data_Mem/n5141 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1149]), .Q(data_mem_out_wire[1149]) );
  DFF \Data_Mem/memory_reg[35][30]  ( .D(\Data_Mem/n5142 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1150]), .Q(data_mem_out_wire[1150]) );
  DFF \Data_Mem/memory_reg[35][31]  ( .D(\Data_Mem/n5143 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1151]), .Q(data_mem_out_wire[1151]) );
  DFF \Data_Mem/memory_reg[34][0]  ( .D(\Data_Mem/n5144 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1088]), .Q(data_mem_out_wire[1088]) );
  DFF \Data_Mem/memory_reg[34][1]  ( .D(\Data_Mem/n5145 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1089]), .Q(data_mem_out_wire[1089]) );
  DFF \Data_Mem/memory_reg[34][2]  ( .D(\Data_Mem/n5146 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1090]), .Q(data_mem_out_wire[1090]) );
  DFF \Data_Mem/memory_reg[34][3]  ( .D(\Data_Mem/n5147 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1091]), .Q(data_mem_out_wire[1091]) );
  DFF \Data_Mem/memory_reg[34][4]  ( .D(\Data_Mem/n5148 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1092]), .Q(data_mem_out_wire[1092]) );
  DFF \Data_Mem/memory_reg[34][5]  ( .D(\Data_Mem/n5149 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1093]), .Q(data_mem_out_wire[1093]) );
  DFF \Data_Mem/memory_reg[34][6]  ( .D(\Data_Mem/n5150 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1094]), .Q(data_mem_out_wire[1094]) );
  DFF \Data_Mem/memory_reg[34][7]  ( .D(\Data_Mem/n5151 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1095]), .Q(data_mem_out_wire[1095]) );
  DFF \Data_Mem/memory_reg[34][8]  ( .D(\Data_Mem/n5152 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1096]), .Q(data_mem_out_wire[1096]) );
  DFF \Data_Mem/memory_reg[34][9]  ( .D(\Data_Mem/n5153 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1097]), .Q(data_mem_out_wire[1097]) );
  DFF \Data_Mem/memory_reg[34][10]  ( .D(\Data_Mem/n5154 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1098]), .Q(data_mem_out_wire[1098]) );
  DFF \Data_Mem/memory_reg[34][11]  ( .D(\Data_Mem/n5155 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1099]), .Q(data_mem_out_wire[1099]) );
  DFF \Data_Mem/memory_reg[34][12]  ( .D(\Data_Mem/n5156 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1100]), .Q(data_mem_out_wire[1100]) );
  DFF \Data_Mem/memory_reg[34][13]  ( .D(\Data_Mem/n5157 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1101]), .Q(data_mem_out_wire[1101]) );
  DFF \Data_Mem/memory_reg[34][14]  ( .D(\Data_Mem/n5158 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1102]), .Q(data_mem_out_wire[1102]) );
  DFF \Data_Mem/memory_reg[34][15]  ( .D(\Data_Mem/n5159 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1103]), .Q(data_mem_out_wire[1103]) );
  DFF \Data_Mem/memory_reg[34][16]  ( .D(\Data_Mem/n5160 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1104]), .Q(data_mem_out_wire[1104]) );
  DFF \Data_Mem/memory_reg[34][17]  ( .D(\Data_Mem/n5161 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1105]), .Q(data_mem_out_wire[1105]) );
  DFF \Data_Mem/memory_reg[34][18]  ( .D(\Data_Mem/n5162 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1106]), .Q(data_mem_out_wire[1106]) );
  DFF \Data_Mem/memory_reg[34][19]  ( .D(\Data_Mem/n5163 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1107]), .Q(data_mem_out_wire[1107]) );
  DFF \Data_Mem/memory_reg[34][20]  ( .D(\Data_Mem/n5164 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1108]), .Q(data_mem_out_wire[1108]) );
  DFF \Data_Mem/memory_reg[34][21]  ( .D(\Data_Mem/n5165 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1109]), .Q(data_mem_out_wire[1109]) );
  DFF \Data_Mem/memory_reg[34][22]  ( .D(\Data_Mem/n5166 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1110]), .Q(data_mem_out_wire[1110]) );
  DFF \Data_Mem/memory_reg[34][23]  ( .D(\Data_Mem/n5167 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1111]), .Q(data_mem_out_wire[1111]) );
  DFF \Data_Mem/memory_reg[34][24]  ( .D(\Data_Mem/n5168 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1112]), .Q(data_mem_out_wire[1112]) );
  DFF \Data_Mem/memory_reg[34][25]  ( .D(\Data_Mem/n5169 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1113]), .Q(data_mem_out_wire[1113]) );
  DFF \Data_Mem/memory_reg[34][26]  ( .D(\Data_Mem/n5170 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1114]), .Q(data_mem_out_wire[1114]) );
  DFF \Data_Mem/memory_reg[34][27]  ( .D(\Data_Mem/n5171 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1115]), .Q(data_mem_out_wire[1115]) );
  DFF \Data_Mem/memory_reg[34][28]  ( .D(\Data_Mem/n5172 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1116]), .Q(data_mem_out_wire[1116]) );
  DFF \Data_Mem/memory_reg[34][29]  ( .D(\Data_Mem/n5173 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1117]), .Q(data_mem_out_wire[1117]) );
  DFF \Data_Mem/memory_reg[34][30]  ( .D(\Data_Mem/n5174 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1118]), .Q(data_mem_out_wire[1118]) );
  DFF \Data_Mem/memory_reg[34][31]  ( .D(\Data_Mem/n5175 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1119]), .Q(data_mem_out_wire[1119]) );
  DFF \Data_Mem/memory_reg[33][0]  ( .D(\Data_Mem/n5176 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1056]), .Q(data_mem_out_wire[1056]) );
  DFF \Data_Mem/memory_reg[33][1]  ( .D(\Data_Mem/n5177 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1057]), .Q(data_mem_out_wire[1057]) );
  DFF \Data_Mem/memory_reg[33][2]  ( .D(\Data_Mem/n5178 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1058]), .Q(data_mem_out_wire[1058]) );
  DFF \Data_Mem/memory_reg[33][3]  ( .D(\Data_Mem/n5179 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1059]), .Q(data_mem_out_wire[1059]) );
  DFF \Data_Mem/memory_reg[33][4]  ( .D(\Data_Mem/n5180 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1060]), .Q(data_mem_out_wire[1060]) );
  DFF \Data_Mem/memory_reg[33][5]  ( .D(\Data_Mem/n5181 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1061]), .Q(data_mem_out_wire[1061]) );
  DFF \Data_Mem/memory_reg[33][6]  ( .D(\Data_Mem/n5182 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1062]), .Q(data_mem_out_wire[1062]) );
  DFF \Data_Mem/memory_reg[33][7]  ( .D(\Data_Mem/n5183 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1063]), .Q(data_mem_out_wire[1063]) );
  DFF \Data_Mem/memory_reg[33][8]  ( .D(\Data_Mem/n5184 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1064]), .Q(data_mem_out_wire[1064]) );
  DFF \Data_Mem/memory_reg[33][9]  ( .D(\Data_Mem/n5185 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1065]), .Q(data_mem_out_wire[1065]) );
  DFF \Data_Mem/memory_reg[33][10]  ( .D(\Data_Mem/n5186 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1066]), .Q(data_mem_out_wire[1066]) );
  DFF \Data_Mem/memory_reg[33][11]  ( .D(\Data_Mem/n5187 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1067]), .Q(data_mem_out_wire[1067]) );
  DFF \Data_Mem/memory_reg[33][12]  ( .D(\Data_Mem/n5188 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1068]), .Q(data_mem_out_wire[1068]) );
  DFF \Data_Mem/memory_reg[33][13]  ( .D(\Data_Mem/n5189 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1069]), .Q(data_mem_out_wire[1069]) );
  DFF \Data_Mem/memory_reg[33][14]  ( .D(\Data_Mem/n5190 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1070]), .Q(data_mem_out_wire[1070]) );
  DFF \Data_Mem/memory_reg[33][15]  ( .D(\Data_Mem/n5191 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1071]), .Q(data_mem_out_wire[1071]) );
  DFF \Data_Mem/memory_reg[33][16]  ( .D(\Data_Mem/n5192 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1072]), .Q(data_mem_out_wire[1072]) );
  DFF \Data_Mem/memory_reg[33][17]  ( .D(\Data_Mem/n5193 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1073]), .Q(data_mem_out_wire[1073]) );
  DFF \Data_Mem/memory_reg[33][18]  ( .D(\Data_Mem/n5194 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1074]), .Q(data_mem_out_wire[1074]) );
  DFF \Data_Mem/memory_reg[33][19]  ( .D(\Data_Mem/n5195 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1075]), .Q(data_mem_out_wire[1075]) );
  DFF \Data_Mem/memory_reg[33][20]  ( .D(\Data_Mem/n5196 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1076]), .Q(data_mem_out_wire[1076]) );
  DFF \Data_Mem/memory_reg[33][21]  ( .D(\Data_Mem/n5197 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1077]), .Q(data_mem_out_wire[1077]) );
  DFF \Data_Mem/memory_reg[33][22]  ( .D(\Data_Mem/n5198 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1078]), .Q(data_mem_out_wire[1078]) );
  DFF \Data_Mem/memory_reg[33][23]  ( .D(\Data_Mem/n5199 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1079]), .Q(data_mem_out_wire[1079]) );
  DFF \Data_Mem/memory_reg[33][24]  ( .D(\Data_Mem/n5200 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1080]), .Q(data_mem_out_wire[1080]) );
  DFF \Data_Mem/memory_reg[33][25]  ( .D(\Data_Mem/n5201 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1081]), .Q(data_mem_out_wire[1081]) );
  DFF \Data_Mem/memory_reg[33][26]  ( .D(\Data_Mem/n5202 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1082]), .Q(data_mem_out_wire[1082]) );
  DFF \Data_Mem/memory_reg[33][27]  ( .D(\Data_Mem/n5203 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1083]), .Q(data_mem_out_wire[1083]) );
  DFF \Data_Mem/memory_reg[33][28]  ( .D(\Data_Mem/n5204 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1084]), .Q(data_mem_out_wire[1084]) );
  DFF \Data_Mem/memory_reg[33][29]  ( .D(\Data_Mem/n5205 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1085]), .Q(data_mem_out_wire[1085]) );
  DFF \Data_Mem/memory_reg[33][30]  ( .D(\Data_Mem/n5206 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1086]), .Q(data_mem_out_wire[1086]) );
  DFF \Data_Mem/memory_reg[33][31]  ( .D(\Data_Mem/n5207 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1087]), .Q(data_mem_out_wire[1087]) );
  DFF \Data_Mem/memory_reg[32][0]  ( .D(\Data_Mem/n5208 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1024]), .Q(data_mem_out_wire[1024]) );
  DFF \Data_Mem/memory_reg[32][1]  ( .D(\Data_Mem/n5209 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1025]), .Q(data_mem_out_wire[1025]) );
  DFF \Data_Mem/memory_reg[32][2]  ( .D(\Data_Mem/n5210 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1026]), .Q(data_mem_out_wire[1026]) );
  DFF \Data_Mem/memory_reg[32][3]  ( .D(\Data_Mem/n5211 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1027]), .Q(data_mem_out_wire[1027]) );
  DFF \Data_Mem/memory_reg[32][4]  ( .D(\Data_Mem/n5212 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1028]), .Q(data_mem_out_wire[1028]) );
  DFF \Data_Mem/memory_reg[32][5]  ( .D(\Data_Mem/n5213 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1029]), .Q(data_mem_out_wire[1029]) );
  DFF \Data_Mem/memory_reg[32][6]  ( .D(\Data_Mem/n5214 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1030]), .Q(data_mem_out_wire[1030]) );
  DFF \Data_Mem/memory_reg[32][7]  ( .D(\Data_Mem/n5215 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1031]), .Q(data_mem_out_wire[1031]) );
  DFF \Data_Mem/memory_reg[32][8]  ( .D(\Data_Mem/n5216 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1032]), .Q(data_mem_out_wire[1032]) );
  DFF \Data_Mem/memory_reg[32][9]  ( .D(\Data_Mem/n5217 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1033]), .Q(data_mem_out_wire[1033]) );
  DFF \Data_Mem/memory_reg[32][10]  ( .D(\Data_Mem/n5218 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1034]), .Q(data_mem_out_wire[1034]) );
  DFF \Data_Mem/memory_reg[32][11]  ( .D(\Data_Mem/n5219 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1035]), .Q(data_mem_out_wire[1035]) );
  DFF \Data_Mem/memory_reg[32][12]  ( .D(\Data_Mem/n5220 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1036]), .Q(data_mem_out_wire[1036]) );
  DFF \Data_Mem/memory_reg[32][13]  ( .D(\Data_Mem/n5221 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1037]), .Q(data_mem_out_wire[1037]) );
  DFF \Data_Mem/memory_reg[32][14]  ( .D(\Data_Mem/n5222 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1038]), .Q(data_mem_out_wire[1038]) );
  DFF \Data_Mem/memory_reg[32][15]  ( .D(\Data_Mem/n5223 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1039]), .Q(data_mem_out_wire[1039]) );
  DFF \Data_Mem/memory_reg[32][16]  ( .D(\Data_Mem/n5224 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1040]), .Q(data_mem_out_wire[1040]) );
  DFF \Data_Mem/memory_reg[32][17]  ( .D(\Data_Mem/n5225 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1041]), .Q(data_mem_out_wire[1041]) );
  DFF \Data_Mem/memory_reg[32][18]  ( .D(\Data_Mem/n5226 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1042]), .Q(data_mem_out_wire[1042]) );
  DFF \Data_Mem/memory_reg[32][19]  ( .D(\Data_Mem/n5227 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1043]), .Q(data_mem_out_wire[1043]) );
  DFF \Data_Mem/memory_reg[32][20]  ( .D(\Data_Mem/n5228 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1044]), .Q(data_mem_out_wire[1044]) );
  DFF \Data_Mem/memory_reg[32][21]  ( .D(\Data_Mem/n5229 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1045]), .Q(data_mem_out_wire[1045]) );
  DFF \Data_Mem/memory_reg[32][22]  ( .D(\Data_Mem/n5230 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1046]), .Q(data_mem_out_wire[1046]) );
  DFF \Data_Mem/memory_reg[32][23]  ( .D(\Data_Mem/n5231 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1047]), .Q(data_mem_out_wire[1047]) );
  DFF \Data_Mem/memory_reg[32][24]  ( .D(\Data_Mem/n5232 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1048]), .Q(data_mem_out_wire[1048]) );
  DFF \Data_Mem/memory_reg[32][25]  ( .D(\Data_Mem/n5233 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1049]), .Q(data_mem_out_wire[1049]) );
  DFF \Data_Mem/memory_reg[32][26]  ( .D(\Data_Mem/n5234 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1050]), .Q(data_mem_out_wire[1050]) );
  DFF \Data_Mem/memory_reg[32][27]  ( .D(\Data_Mem/n5235 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1051]), .Q(data_mem_out_wire[1051]) );
  DFF \Data_Mem/memory_reg[32][28]  ( .D(\Data_Mem/n5236 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1052]), .Q(data_mem_out_wire[1052]) );
  DFF \Data_Mem/memory_reg[32][29]  ( .D(\Data_Mem/n5237 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1053]), .Q(data_mem_out_wire[1053]) );
  DFF \Data_Mem/memory_reg[32][30]  ( .D(\Data_Mem/n5238 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1054]), .Q(data_mem_out_wire[1054]) );
  DFF \Data_Mem/memory_reg[32][31]  ( .D(\Data_Mem/n5239 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1055]), .Q(data_mem_out_wire[1055]) );
  DFF \Data_Mem/memory_reg[31][0]  ( .D(\Data_Mem/n5240 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[992]), .Q(data_mem_out_wire[992]) );
  DFF \Data_Mem/memory_reg[31][1]  ( .D(\Data_Mem/n5241 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[993]), .Q(data_mem_out_wire[993]) );
  DFF \Data_Mem/memory_reg[31][2]  ( .D(\Data_Mem/n5242 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[994]), .Q(data_mem_out_wire[994]) );
  DFF \Data_Mem/memory_reg[31][3]  ( .D(\Data_Mem/n5243 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[995]), .Q(data_mem_out_wire[995]) );
  DFF \Data_Mem/memory_reg[31][4]  ( .D(\Data_Mem/n5244 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[996]), .Q(data_mem_out_wire[996]) );
  DFF \Data_Mem/memory_reg[31][5]  ( .D(\Data_Mem/n5245 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[997]), .Q(data_mem_out_wire[997]) );
  DFF \Data_Mem/memory_reg[31][6]  ( .D(\Data_Mem/n5246 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[998]), .Q(data_mem_out_wire[998]) );
  DFF \Data_Mem/memory_reg[31][7]  ( .D(\Data_Mem/n5247 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[999]), .Q(data_mem_out_wire[999]) );
  DFF \Data_Mem/memory_reg[31][8]  ( .D(\Data_Mem/n5248 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1000]), .Q(data_mem_out_wire[1000]) );
  DFF \Data_Mem/memory_reg[31][9]  ( .D(\Data_Mem/n5249 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[1001]), .Q(data_mem_out_wire[1001]) );
  DFF \Data_Mem/memory_reg[31][10]  ( .D(\Data_Mem/n5250 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1002]), .Q(data_mem_out_wire[1002]) );
  DFF \Data_Mem/memory_reg[31][11]  ( .D(\Data_Mem/n5251 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1003]), .Q(data_mem_out_wire[1003]) );
  DFF \Data_Mem/memory_reg[31][12]  ( .D(\Data_Mem/n5252 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1004]), .Q(data_mem_out_wire[1004]) );
  DFF \Data_Mem/memory_reg[31][13]  ( .D(\Data_Mem/n5253 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1005]), .Q(data_mem_out_wire[1005]) );
  DFF \Data_Mem/memory_reg[31][14]  ( .D(\Data_Mem/n5254 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1006]), .Q(data_mem_out_wire[1006]) );
  DFF \Data_Mem/memory_reg[31][15]  ( .D(\Data_Mem/n5255 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1007]), .Q(data_mem_out_wire[1007]) );
  DFF \Data_Mem/memory_reg[31][16]  ( .D(\Data_Mem/n5256 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1008]), .Q(data_mem_out_wire[1008]) );
  DFF \Data_Mem/memory_reg[31][17]  ( .D(\Data_Mem/n5257 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1009]), .Q(data_mem_out_wire[1009]) );
  DFF \Data_Mem/memory_reg[31][18]  ( .D(\Data_Mem/n5258 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1010]), .Q(data_mem_out_wire[1010]) );
  DFF \Data_Mem/memory_reg[31][19]  ( .D(\Data_Mem/n5259 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1011]), .Q(data_mem_out_wire[1011]) );
  DFF \Data_Mem/memory_reg[31][20]  ( .D(\Data_Mem/n5260 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1012]), .Q(data_mem_out_wire[1012]) );
  DFF \Data_Mem/memory_reg[31][21]  ( .D(\Data_Mem/n5261 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1013]), .Q(data_mem_out_wire[1013]) );
  DFF \Data_Mem/memory_reg[31][22]  ( .D(\Data_Mem/n5262 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1014]), .Q(data_mem_out_wire[1014]) );
  DFF \Data_Mem/memory_reg[31][23]  ( .D(\Data_Mem/n5263 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1015]), .Q(data_mem_out_wire[1015]) );
  DFF \Data_Mem/memory_reg[31][24]  ( .D(\Data_Mem/n5264 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1016]), .Q(data_mem_out_wire[1016]) );
  DFF \Data_Mem/memory_reg[31][25]  ( .D(\Data_Mem/n5265 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1017]), .Q(data_mem_out_wire[1017]) );
  DFF \Data_Mem/memory_reg[31][26]  ( .D(\Data_Mem/n5266 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1018]), .Q(data_mem_out_wire[1018]) );
  DFF \Data_Mem/memory_reg[31][27]  ( .D(\Data_Mem/n5267 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1019]), .Q(data_mem_out_wire[1019]) );
  DFF \Data_Mem/memory_reg[31][28]  ( .D(\Data_Mem/n5268 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1020]), .Q(data_mem_out_wire[1020]) );
  DFF \Data_Mem/memory_reg[31][29]  ( .D(\Data_Mem/n5269 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1021]), .Q(data_mem_out_wire[1021]) );
  DFF \Data_Mem/memory_reg[31][30]  ( .D(\Data_Mem/n5270 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1022]), .Q(data_mem_out_wire[1022]) );
  DFF \Data_Mem/memory_reg[31][31]  ( .D(\Data_Mem/n5271 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[1023]), .Q(data_mem_out_wire[1023]) );
  DFF \Data_Mem/memory_reg[30][0]  ( .D(\Data_Mem/n5272 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[960]), .Q(data_mem_out_wire[960]) );
  DFF \Data_Mem/memory_reg[30][1]  ( .D(\Data_Mem/n5273 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[961]), .Q(data_mem_out_wire[961]) );
  DFF \Data_Mem/memory_reg[30][2]  ( .D(\Data_Mem/n5274 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[962]), .Q(data_mem_out_wire[962]) );
  DFF \Data_Mem/memory_reg[30][3]  ( .D(\Data_Mem/n5275 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[963]), .Q(data_mem_out_wire[963]) );
  DFF \Data_Mem/memory_reg[30][4]  ( .D(\Data_Mem/n5276 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[964]), .Q(data_mem_out_wire[964]) );
  DFF \Data_Mem/memory_reg[30][5]  ( .D(\Data_Mem/n5277 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[965]), .Q(data_mem_out_wire[965]) );
  DFF \Data_Mem/memory_reg[30][6]  ( .D(\Data_Mem/n5278 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[966]), .Q(data_mem_out_wire[966]) );
  DFF \Data_Mem/memory_reg[30][7]  ( .D(\Data_Mem/n5279 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[967]), .Q(data_mem_out_wire[967]) );
  DFF \Data_Mem/memory_reg[30][8]  ( .D(\Data_Mem/n5280 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[968]), .Q(data_mem_out_wire[968]) );
  DFF \Data_Mem/memory_reg[30][9]  ( .D(\Data_Mem/n5281 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[969]), .Q(data_mem_out_wire[969]) );
  DFF \Data_Mem/memory_reg[30][10]  ( .D(\Data_Mem/n5282 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[970]), .Q(data_mem_out_wire[970]) );
  DFF \Data_Mem/memory_reg[30][11]  ( .D(\Data_Mem/n5283 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[971]), .Q(data_mem_out_wire[971]) );
  DFF \Data_Mem/memory_reg[30][12]  ( .D(\Data_Mem/n5284 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[972]), .Q(data_mem_out_wire[972]) );
  DFF \Data_Mem/memory_reg[30][13]  ( .D(\Data_Mem/n5285 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[973]), .Q(data_mem_out_wire[973]) );
  DFF \Data_Mem/memory_reg[30][14]  ( .D(\Data_Mem/n5286 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[974]), .Q(data_mem_out_wire[974]) );
  DFF \Data_Mem/memory_reg[30][15]  ( .D(\Data_Mem/n5287 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[975]), .Q(data_mem_out_wire[975]) );
  DFF \Data_Mem/memory_reg[30][16]  ( .D(\Data_Mem/n5288 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[976]), .Q(data_mem_out_wire[976]) );
  DFF \Data_Mem/memory_reg[30][17]  ( .D(\Data_Mem/n5289 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[977]), .Q(data_mem_out_wire[977]) );
  DFF \Data_Mem/memory_reg[30][18]  ( .D(\Data_Mem/n5290 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[978]), .Q(data_mem_out_wire[978]) );
  DFF \Data_Mem/memory_reg[30][19]  ( .D(\Data_Mem/n5291 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[979]), .Q(data_mem_out_wire[979]) );
  DFF \Data_Mem/memory_reg[30][20]  ( .D(\Data_Mem/n5292 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[980]), .Q(data_mem_out_wire[980]) );
  DFF \Data_Mem/memory_reg[30][21]  ( .D(\Data_Mem/n5293 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[981]), .Q(data_mem_out_wire[981]) );
  DFF \Data_Mem/memory_reg[30][22]  ( .D(\Data_Mem/n5294 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[982]), .Q(data_mem_out_wire[982]) );
  DFF \Data_Mem/memory_reg[30][23]  ( .D(\Data_Mem/n5295 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[983]), .Q(data_mem_out_wire[983]) );
  DFF \Data_Mem/memory_reg[30][24]  ( .D(\Data_Mem/n5296 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[984]), .Q(data_mem_out_wire[984]) );
  DFF \Data_Mem/memory_reg[30][25]  ( .D(\Data_Mem/n5297 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[985]), .Q(data_mem_out_wire[985]) );
  DFF \Data_Mem/memory_reg[30][26]  ( .D(\Data_Mem/n5298 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[986]), .Q(data_mem_out_wire[986]) );
  DFF \Data_Mem/memory_reg[30][27]  ( .D(\Data_Mem/n5299 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[987]), .Q(data_mem_out_wire[987]) );
  DFF \Data_Mem/memory_reg[30][28]  ( .D(\Data_Mem/n5300 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[988]), .Q(data_mem_out_wire[988]) );
  DFF \Data_Mem/memory_reg[30][29]  ( .D(\Data_Mem/n5301 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[989]), .Q(data_mem_out_wire[989]) );
  DFF \Data_Mem/memory_reg[30][30]  ( .D(\Data_Mem/n5302 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[990]), .Q(data_mem_out_wire[990]) );
  DFF \Data_Mem/memory_reg[30][31]  ( .D(\Data_Mem/n5303 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[991]), .Q(data_mem_out_wire[991]) );
  DFF \Data_Mem/memory_reg[29][0]  ( .D(\Data_Mem/n5304 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[928]), .Q(data_mem_out_wire[928]) );
  DFF \Data_Mem/memory_reg[29][1]  ( .D(\Data_Mem/n5305 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[929]), .Q(data_mem_out_wire[929]) );
  DFF \Data_Mem/memory_reg[29][2]  ( .D(\Data_Mem/n5306 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[930]), .Q(data_mem_out_wire[930]) );
  DFF \Data_Mem/memory_reg[29][3]  ( .D(\Data_Mem/n5307 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[931]), .Q(data_mem_out_wire[931]) );
  DFF \Data_Mem/memory_reg[29][4]  ( .D(\Data_Mem/n5308 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[932]), .Q(data_mem_out_wire[932]) );
  DFF \Data_Mem/memory_reg[29][5]  ( .D(\Data_Mem/n5309 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[933]), .Q(data_mem_out_wire[933]) );
  DFF \Data_Mem/memory_reg[29][6]  ( .D(\Data_Mem/n5310 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[934]), .Q(data_mem_out_wire[934]) );
  DFF \Data_Mem/memory_reg[29][7]  ( .D(\Data_Mem/n5311 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[935]), .Q(data_mem_out_wire[935]) );
  DFF \Data_Mem/memory_reg[29][8]  ( .D(\Data_Mem/n5312 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[936]), .Q(data_mem_out_wire[936]) );
  DFF \Data_Mem/memory_reg[29][9]  ( .D(\Data_Mem/n5313 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[937]), .Q(data_mem_out_wire[937]) );
  DFF \Data_Mem/memory_reg[29][10]  ( .D(\Data_Mem/n5314 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[938]), .Q(data_mem_out_wire[938]) );
  DFF \Data_Mem/memory_reg[29][11]  ( .D(\Data_Mem/n5315 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[939]), .Q(data_mem_out_wire[939]) );
  DFF \Data_Mem/memory_reg[29][12]  ( .D(\Data_Mem/n5316 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[940]), .Q(data_mem_out_wire[940]) );
  DFF \Data_Mem/memory_reg[29][13]  ( .D(\Data_Mem/n5317 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[941]), .Q(data_mem_out_wire[941]) );
  DFF \Data_Mem/memory_reg[29][14]  ( .D(\Data_Mem/n5318 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[942]), .Q(data_mem_out_wire[942]) );
  DFF \Data_Mem/memory_reg[29][15]  ( .D(\Data_Mem/n5319 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[943]), .Q(data_mem_out_wire[943]) );
  DFF \Data_Mem/memory_reg[29][16]  ( .D(\Data_Mem/n5320 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[944]), .Q(data_mem_out_wire[944]) );
  DFF \Data_Mem/memory_reg[29][17]  ( .D(\Data_Mem/n5321 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[945]), .Q(data_mem_out_wire[945]) );
  DFF \Data_Mem/memory_reg[29][18]  ( .D(\Data_Mem/n5322 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[946]), .Q(data_mem_out_wire[946]) );
  DFF \Data_Mem/memory_reg[29][19]  ( .D(\Data_Mem/n5323 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[947]), .Q(data_mem_out_wire[947]) );
  DFF \Data_Mem/memory_reg[29][20]  ( .D(\Data_Mem/n5324 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[948]), .Q(data_mem_out_wire[948]) );
  DFF \Data_Mem/memory_reg[29][21]  ( .D(\Data_Mem/n5325 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[949]), .Q(data_mem_out_wire[949]) );
  DFF \Data_Mem/memory_reg[29][22]  ( .D(\Data_Mem/n5326 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[950]), .Q(data_mem_out_wire[950]) );
  DFF \Data_Mem/memory_reg[29][23]  ( .D(\Data_Mem/n5327 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[951]), .Q(data_mem_out_wire[951]) );
  DFF \Data_Mem/memory_reg[29][24]  ( .D(\Data_Mem/n5328 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[952]), .Q(data_mem_out_wire[952]) );
  DFF \Data_Mem/memory_reg[29][25]  ( .D(\Data_Mem/n5329 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[953]), .Q(data_mem_out_wire[953]) );
  DFF \Data_Mem/memory_reg[29][26]  ( .D(\Data_Mem/n5330 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[954]), .Q(data_mem_out_wire[954]) );
  DFF \Data_Mem/memory_reg[29][27]  ( .D(\Data_Mem/n5331 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[955]), .Q(data_mem_out_wire[955]) );
  DFF \Data_Mem/memory_reg[29][28]  ( .D(\Data_Mem/n5332 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[956]), .Q(data_mem_out_wire[956]) );
  DFF \Data_Mem/memory_reg[29][29]  ( .D(\Data_Mem/n5333 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[957]), .Q(data_mem_out_wire[957]) );
  DFF \Data_Mem/memory_reg[29][30]  ( .D(\Data_Mem/n5334 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[958]), .Q(data_mem_out_wire[958]) );
  DFF \Data_Mem/memory_reg[29][31]  ( .D(\Data_Mem/n5335 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[959]), .Q(data_mem_out_wire[959]) );
  DFF \Data_Mem/memory_reg[28][0]  ( .D(\Data_Mem/n5336 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[896]), .Q(data_mem_out_wire[896]) );
  DFF \Data_Mem/memory_reg[28][1]  ( .D(\Data_Mem/n5337 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[897]), .Q(data_mem_out_wire[897]) );
  DFF \Data_Mem/memory_reg[28][2]  ( .D(\Data_Mem/n5338 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[898]), .Q(data_mem_out_wire[898]) );
  DFF \Data_Mem/memory_reg[28][3]  ( .D(\Data_Mem/n5339 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[899]), .Q(data_mem_out_wire[899]) );
  DFF \Data_Mem/memory_reg[28][4]  ( .D(\Data_Mem/n5340 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[900]), .Q(data_mem_out_wire[900]) );
  DFF \Data_Mem/memory_reg[28][5]  ( .D(\Data_Mem/n5341 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[901]), .Q(data_mem_out_wire[901]) );
  DFF \Data_Mem/memory_reg[28][6]  ( .D(\Data_Mem/n5342 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[902]), .Q(data_mem_out_wire[902]) );
  DFF \Data_Mem/memory_reg[28][7]  ( .D(\Data_Mem/n5343 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[903]), .Q(data_mem_out_wire[903]) );
  DFF \Data_Mem/memory_reg[28][8]  ( .D(\Data_Mem/n5344 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[904]), .Q(data_mem_out_wire[904]) );
  DFF \Data_Mem/memory_reg[28][9]  ( .D(\Data_Mem/n5345 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[905]), .Q(data_mem_out_wire[905]) );
  DFF \Data_Mem/memory_reg[28][10]  ( .D(\Data_Mem/n5346 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[906]), .Q(data_mem_out_wire[906]) );
  DFF \Data_Mem/memory_reg[28][11]  ( .D(\Data_Mem/n5347 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[907]), .Q(data_mem_out_wire[907]) );
  DFF \Data_Mem/memory_reg[28][12]  ( .D(\Data_Mem/n5348 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[908]), .Q(data_mem_out_wire[908]) );
  DFF \Data_Mem/memory_reg[28][13]  ( .D(\Data_Mem/n5349 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[909]), .Q(data_mem_out_wire[909]) );
  DFF \Data_Mem/memory_reg[28][14]  ( .D(\Data_Mem/n5350 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[910]), .Q(data_mem_out_wire[910]) );
  DFF \Data_Mem/memory_reg[28][15]  ( .D(\Data_Mem/n5351 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[911]), .Q(data_mem_out_wire[911]) );
  DFF \Data_Mem/memory_reg[28][16]  ( .D(\Data_Mem/n5352 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[912]), .Q(data_mem_out_wire[912]) );
  DFF \Data_Mem/memory_reg[28][17]  ( .D(\Data_Mem/n5353 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[913]), .Q(data_mem_out_wire[913]) );
  DFF \Data_Mem/memory_reg[28][18]  ( .D(\Data_Mem/n5354 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[914]), .Q(data_mem_out_wire[914]) );
  DFF \Data_Mem/memory_reg[28][19]  ( .D(\Data_Mem/n5355 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[915]), .Q(data_mem_out_wire[915]) );
  DFF \Data_Mem/memory_reg[28][20]  ( .D(\Data_Mem/n5356 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[916]), .Q(data_mem_out_wire[916]) );
  DFF \Data_Mem/memory_reg[28][21]  ( .D(\Data_Mem/n5357 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[917]), .Q(data_mem_out_wire[917]) );
  DFF \Data_Mem/memory_reg[28][22]  ( .D(\Data_Mem/n5358 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[918]), .Q(data_mem_out_wire[918]) );
  DFF \Data_Mem/memory_reg[28][23]  ( .D(\Data_Mem/n5359 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[919]), .Q(data_mem_out_wire[919]) );
  DFF \Data_Mem/memory_reg[28][24]  ( .D(\Data_Mem/n5360 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[920]), .Q(data_mem_out_wire[920]) );
  DFF \Data_Mem/memory_reg[28][25]  ( .D(\Data_Mem/n5361 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[921]), .Q(data_mem_out_wire[921]) );
  DFF \Data_Mem/memory_reg[28][26]  ( .D(\Data_Mem/n5362 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[922]), .Q(data_mem_out_wire[922]) );
  DFF \Data_Mem/memory_reg[28][27]  ( .D(\Data_Mem/n5363 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[923]), .Q(data_mem_out_wire[923]) );
  DFF \Data_Mem/memory_reg[28][28]  ( .D(\Data_Mem/n5364 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[924]), .Q(data_mem_out_wire[924]) );
  DFF \Data_Mem/memory_reg[28][29]  ( .D(\Data_Mem/n5365 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[925]), .Q(data_mem_out_wire[925]) );
  DFF \Data_Mem/memory_reg[28][30]  ( .D(\Data_Mem/n5366 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[926]), .Q(data_mem_out_wire[926]) );
  DFF \Data_Mem/memory_reg[28][31]  ( .D(\Data_Mem/n5367 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[927]), .Q(data_mem_out_wire[927]) );
  DFF \Data_Mem/memory_reg[27][0]  ( .D(\Data_Mem/n5368 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[864]), .Q(data_mem_out_wire[864]) );
  DFF \Data_Mem/memory_reg[27][1]  ( .D(\Data_Mem/n5369 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[865]), .Q(data_mem_out_wire[865]) );
  DFF \Data_Mem/memory_reg[27][2]  ( .D(\Data_Mem/n5370 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[866]), .Q(data_mem_out_wire[866]) );
  DFF \Data_Mem/memory_reg[27][3]  ( .D(\Data_Mem/n5371 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[867]), .Q(data_mem_out_wire[867]) );
  DFF \Data_Mem/memory_reg[27][4]  ( .D(\Data_Mem/n5372 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[868]), .Q(data_mem_out_wire[868]) );
  DFF \Data_Mem/memory_reg[27][5]  ( .D(\Data_Mem/n5373 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[869]), .Q(data_mem_out_wire[869]) );
  DFF \Data_Mem/memory_reg[27][6]  ( .D(\Data_Mem/n5374 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[870]), .Q(data_mem_out_wire[870]) );
  DFF \Data_Mem/memory_reg[27][7]  ( .D(\Data_Mem/n5375 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[871]), .Q(data_mem_out_wire[871]) );
  DFF \Data_Mem/memory_reg[27][8]  ( .D(\Data_Mem/n5376 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[872]), .Q(data_mem_out_wire[872]) );
  DFF \Data_Mem/memory_reg[27][9]  ( .D(\Data_Mem/n5377 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[873]), .Q(data_mem_out_wire[873]) );
  DFF \Data_Mem/memory_reg[27][10]  ( .D(\Data_Mem/n5378 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[874]), .Q(data_mem_out_wire[874]) );
  DFF \Data_Mem/memory_reg[27][11]  ( .D(\Data_Mem/n5379 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[875]), .Q(data_mem_out_wire[875]) );
  DFF \Data_Mem/memory_reg[27][12]  ( .D(\Data_Mem/n5380 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[876]), .Q(data_mem_out_wire[876]) );
  DFF \Data_Mem/memory_reg[27][13]  ( .D(\Data_Mem/n5381 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[877]), .Q(data_mem_out_wire[877]) );
  DFF \Data_Mem/memory_reg[27][14]  ( .D(\Data_Mem/n5382 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[878]), .Q(data_mem_out_wire[878]) );
  DFF \Data_Mem/memory_reg[27][15]  ( .D(\Data_Mem/n5383 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[879]), .Q(data_mem_out_wire[879]) );
  DFF \Data_Mem/memory_reg[27][16]  ( .D(\Data_Mem/n5384 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[880]), .Q(data_mem_out_wire[880]) );
  DFF \Data_Mem/memory_reg[27][17]  ( .D(\Data_Mem/n5385 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[881]), .Q(data_mem_out_wire[881]) );
  DFF \Data_Mem/memory_reg[27][18]  ( .D(\Data_Mem/n5386 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[882]), .Q(data_mem_out_wire[882]) );
  DFF \Data_Mem/memory_reg[27][19]  ( .D(\Data_Mem/n5387 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[883]), .Q(data_mem_out_wire[883]) );
  DFF \Data_Mem/memory_reg[27][20]  ( .D(\Data_Mem/n5388 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[884]), .Q(data_mem_out_wire[884]) );
  DFF \Data_Mem/memory_reg[27][21]  ( .D(\Data_Mem/n5389 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[885]), .Q(data_mem_out_wire[885]) );
  DFF \Data_Mem/memory_reg[27][22]  ( .D(\Data_Mem/n5390 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[886]), .Q(data_mem_out_wire[886]) );
  DFF \Data_Mem/memory_reg[27][23]  ( .D(\Data_Mem/n5391 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[887]), .Q(data_mem_out_wire[887]) );
  DFF \Data_Mem/memory_reg[27][24]  ( .D(\Data_Mem/n5392 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[888]), .Q(data_mem_out_wire[888]) );
  DFF \Data_Mem/memory_reg[27][25]  ( .D(\Data_Mem/n5393 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[889]), .Q(data_mem_out_wire[889]) );
  DFF \Data_Mem/memory_reg[27][26]  ( .D(\Data_Mem/n5394 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[890]), .Q(data_mem_out_wire[890]) );
  DFF \Data_Mem/memory_reg[27][27]  ( .D(\Data_Mem/n5395 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[891]), .Q(data_mem_out_wire[891]) );
  DFF \Data_Mem/memory_reg[27][28]  ( .D(\Data_Mem/n5396 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[892]), .Q(data_mem_out_wire[892]) );
  DFF \Data_Mem/memory_reg[27][29]  ( .D(\Data_Mem/n5397 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[893]), .Q(data_mem_out_wire[893]) );
  DFF \Data_Mem/memory_reg[27][30]  ( .D(\Data_Mem/n5398 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[894]), .Q(data_mem_out_wire[894]) );
  DFF \Data_Mem/memory_reg[27][31]  ( .D(\Data_Mem/n5399 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[895]), .Q(data_mem_out_wire[895]) );
  DFF \Data_Mem/memory_reg[26][0]  ( .D(\Data_Mem/n5400 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[832]), .Q(data_mem_out_wire[832]) );
  DFF \Data_Mem/memory_reg[26][1]  ( .D(\Data_Mem/n5401 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[833]), .Q(data_mem_out_wire[833]) );
  DFF \Data_Mem/memory_reg[26][2]  ( .D(\Data_Mem/n5402 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[834]), .Q(data_mem_out_wire[834]) );
  DFF \Data_Mem/memory_reg[26][3]  ( .D(\Data_Mem/n5403 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[835]), .Q(data_mem_out_wire[835]) );
  DFF \Data_Mem/memory_reg[26][4]  ( .D(\Data_Mem/n5404 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[836]), .Q(data_mem_out_wire[836]) );
  DFF \Data_Mem/memory_reg[26][5]  ( .D(\Data_Mem/n5405 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[837]), .Q(data_mem_out_wire[837]) );
  DFF \Data_Mem/memory_reg[26][6]  ( .D(\Data_Mem/n5406 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[838]), .Q(data_mem_out_wire[838]) );
  DFF \Data_Mem/memory_reg[26][7]  ( .D(\Data_Mem/n5407 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[839]), .Q(data_mem_out_wire[839]) );
  DFF \Data_Mem/memory_reg[26][8]  ( .D(\Data_Mem/n5408 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[840]), .Q(data_mem_out_wire[840]) );
  DFF \Data_Mem/memory_reg[26][9]  ( .D(\Data_Mem/n5409 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[841]), .Q(data_mem_out_wire[841]) );
  DFF \Data_Mem/memory_reg[26][10]  ( .D(\Data_Mem/n5410 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[842]), .Q(data_mem_out_wire[842]) );
  DFF \Data_Mem/memory_reg[26][11]  ( .D(\Data_Mem/n5411 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[843]), .Q(data_mem_out_wire[843]) );
  DFF \Data_Mem/memory_reg[26][12]  ( .D(\Data_Mem/n5412 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[844]), .Q(data_mem_out_wire[844]) );
  DFF \Data_Mem/memory_reg[26][13]  ( .D(\Data_Mem/n5413 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[845]), .Q(data_mem_out_wire[845]) );
  DFF \Data_Mem/memory_reg[26][14]  ( .D(\Data_Mem/n5414 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[846]), .Q(data_mem_out_wire[846]) );
  DFF \Data_Mem/memory_reg[26][15]  ( .D(\Data_Mem/n5415 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[847]), .Q(data_mem_out_wire[847]) );
  DFF \Data_Mem/memory_reg[26][16]  ( .D(\Data_Mem/n5416 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[848]), .Q(data_mem_out_wire[848]) );
  DFF \Data_Mem/memory_reg[26][17]  ( .D(\Data_Mem/n5417 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[849]), .Q(data_mem_out_wire[849]) );
  DFF \Data_Mem/memory_reg[26][18]  ( .D(\Data_Mem/n5418 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[850]), .Q(data_mem_out_wire[850]) );
  DFF \Data_Mem/memory_reg[26][19]  ( .D(\Data_Mem/n5419 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[851]), .Q(data_mem_out_wire[851]) );
  DFF \Data_Mem/memory_reg[26][20]  ( .D(\Data_Mem/n5420 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[852]), .Q(data_mem_out_wire[852]) );
  DFF \Data_Mem/memory_reg[26][21]  ( .D(\Data_Mem/n5421 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[853]), .Q(data_mem_out_wire[853]) );
  DFF \Data_Mem/memory_reg[26][22]  ( .D(\Data_Mem/n5422 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[854]), .Q(data_mem_out_wire[854]) );
  DFF \Data_Mem/memory_reg[26][23]  ( .D(\Data_Mem/n5423 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[855]), .Q(data_mem_out_wire[855]) );
  DFF \Data_Mem/memory_reg[26][24]  ( .D(\Data_Mem/n5424 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[856]), .Q(data_mem_out_wire[856]) );
  DFF \Data_Mem/memory_reg[26][25]  ( .D(\Data_Mem/n5425 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[857]), .Q(data_mem_out_wire[857]) );
  DFF \Data_Mem/memory_reg[26][26]  ( .D(\Data_Mem/n5426 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[858]), .Q(data_mem_out_wire[858]) );
  DFF \Data_Mem/memory_reg[26][27]  ( .D(\Data_Mem/n5427 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[859]), .Q(data_mem_out_wire[859]) );
  DFF \Data_Mem/memory_reg[26][28]  ( .D(\Data_Mem/n5428 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[860]), .Q(data_mem_out_wire[860]) );
  DFF \Data_Mem/memory_reg[26][29]  ( .D(\Data_Mem/n5429 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[861]), .Q(data_mem_out_wire[861]) );
  DFF \Data_Mem/memory_reg[26][30]  ( .D(\Data_Mem/n5430 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[862]), .Q(data_mem_out_wire[862]) );
  DFF \Data_Mem/memory_reg[26][31]  ( .D(\Data_Mem/n5431 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[863]), .Q(data_mem_out_wire[863]) );
  DFF \Data_Mem/memory_reg[25][0]  ( .D(\Data_Mem/n5432 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[800]), .Q(data_mem_out_wire[800]) );
  DFF \Data_Mem/memory_reg[25][1]  ( .D(\Data_Mem/n5433 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[801]), .Q(data_mem_out_wire[801]) );
  DFF \Data_Mem/memory_reg[25][2]  ( .D(\Data_Mem/n5434 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[802]), .Q(data_mem_out_wire[802]) );
  DFF \Data_Mem/memory_reg[25][3]  ( .D(\Data_Mem/n5435 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[803]), .Q(data_mem_out_wire[803]) );
  DFF \Data_Mem/memory_reg[25][4]  ( .D(\Data_Mem/n5436 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[804]), .Q(data_mem_out_wire[804]) );
  DFF \Data_Mem/memory_reg[25][5]  ( .D(\Data_Mem/n5437 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[805]), .Q(data_mem_out_wire[805]) );
  DFF \Data_Mem/memory_reg[25][6]  ( .D(\Data_Mem/n5438 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[806]), .Q(data_mem_out_wire[806]) );
  DFF \Data_Mem/memory_reg[25][7]  ( .D(\Data_Mem/n5439 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[807]), .Q(data_mem_out_wire[807]) );
  DFF \Data_Mem/memory_reg[25][8]  ( .D(\Data_Mem/n5440 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[808]), .Q(data_mem_out_wire[808]) );
  DFF \Data_Mem/memory_reg[25][9]  ( .D(\Data_Mem/n5441 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[809]), .Q(data_mem_out_wire[809]) );
  DFF \Data_Mem/memory_reg[25][10]  ( .D(\Data_Mem/n5442 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[810]), .Q(data_mem_out_wire[810]) );
  DFF \Data_Mem/memory_reg[25][11]  ( .D(\Data_Mem/n5443 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[811]), .Q(data_mem_out_wire[811]) );
  DFF \Data_Mem/memory_reg[25][12]  ( .D(\Data_Mem/n5444 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[812]), .Q(data_mem_out_wire[812]) );
  DFF \Data_Mem/memory_reg[25][13]  ( .D(\Data_Mem/n5445 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[813]), .Q(data_mem_out_wire[813]) );
  DFF \Data_Mem/memory_reg[25][14]  ( .D(\Data_Mem/n5446 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[814]), .Q(data_mem_out_wire[814]) );
  DFF \Data_Mem/memory_reg[25][15]  ( .D(\Data_Mem/n5447 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[815]), .Q(data_mem_out_wire[815]) );
  DFF \Data_Mem/memory_reg[25][16]  ( .D(\Data_Mem/n5448 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[816]), .Q(data_mem_out_wire[816]) );
  DFF \Data_Mem/memory_reg[25][17]  ( .D(\Data_Mem/n5449 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[817]), .Q(data_mem_out_wire[817]) );
  DFF \Data_Mem/memory_reg[25][18]  ( .D(\Data_Mem/n5450 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[818]), .Q(data_mem_out_wire[818]) );
  DFF \Data_Mem/memory_reg[25][19]  ( .D(\Data_Mem/n5451 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[819]), .Q(data_mem_out_wire[819]) );
  DFF \Data_Mem/memory_reg[25][20]  ( .D(\Data_Mem/n5452 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[820]), .Q(data_mem_out_wire[820]) );
  DFF \Data_Mem/memory_reg[25][21]  ( .D(\Data_Mem/n5453 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[821]), .Q(data_mem_out_wire[821]) );
  DFF \Data_Mem/memory_reg[25][22]  ( .D(\Data_Mem/n5454 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[822]), .Q(data_mem_out_wire[822]) );
  DFF \Data_Mem/memory_reg[25][23]  ( .D(\Data_Mem/n5455 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[823]), .Q(data_mem_out_wire[823]) );
  DFF \Data_Mem/memory_reg[25][24]  ( .D(\Data_Mem/n5456 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[824]), .Q(data_mem_out_wire[824]) );
  DFF \Data_Mem/memory_reg[25][25]  ( .D(\Data_Mem/n5457 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[825]), .Q(data_mem_out_wire[825]) );
  DFF \Data_Mem/memory_reg[25][26]  ( .D(\Data_Mem/n5458 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[826]), .Q(data_mem_out_wire[826]) );
  DFF \Data_Mem/memory_reg[25][27]  ( .D(\Data_Mem/n5459 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[827]), .Q(data_mem_out_wire[827]) );
  DFF \Data_Mem/memory_reg[25][28]  ( .D(\Data_Mem/n5460 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[828]), .Q(data_mem_out_wire[828]) );
  DFF \Data_Mem/memory_reg[25][29]  ( .D(\Data_Mem/n5461 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[829]), .Q(data_mem_out_wire[829]) );
  DFF \Data_Mem/memory_reg[25][30]  ( .D(\Data_Mem/n5462 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[830]), .Q(data_mem_out_wire[830]) );
  DFF \Data_Mem/memory_reg[25][31]  ( .D(\Data_Mem/n5463 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[831]), .Q(data_mem_out_wire[831]) );
  DFF \Data_Mem/memory_reg[24][0]  ( .D(\Data_Mem/n5464 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[768]), .Q(data_mem_out_wire[768]) );
  DFF \Data_Mem/memory_reg[24][1]  ( .D(\Data_Mem/n5465 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[769]), .Q(data_mem_out_wire[769]) );
  DFF \Data_Mem/memory_reg[24][2]  ( .D(\Data_Mem/n5466 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[770]), .Q(data_mem_out_wire[770]) );
  DFF \Data_Mem/memory_reg[24][3]  ( .D(\Data_Mem/n5467 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[771]), .Q(data_mem_out_wire[771]) );
  DFF \Data_Mem/memory_reg[24][4]  ( .D(\Data_Mem/n5468 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[772]), .Q(data_mem_out_wire[772]) );
  DFF \Data_Mem/memory_reg[24][5]  ( .D(\Data_Mem/n5469 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[773]), .Q(data_mem_out_wire[773]) );
  DFF \Data_Mem/memory_reg[24][6]  ( .D(\Data_Mem/n5470 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[774]), .Q(data_mem_out_wire[774]) );
  DFF \Data_Mem/memory_reg[24][7]  ( .D(\Data_Mem/n5471 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[775]), .Q(data_mem_out_wire[775]) );
  DFF \Data_Mem/memory_reg[24][8]  ( .D(\Data_Mem/n5472 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[776]), .Q(data_mem_out_wire[776]) );
  DFF \Data_Mem/memory_reg[24][9]  ( .D(\Data_Mem/n5473 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[777]), .Q(data_mem_out_wire[777]) );
  DFF \Data_Mem/memory_reg[24][10]  ( .D(\Data_Mem/n5474 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[778]), .Q(data_mem_out_wire[778]) );
  DFF \Data_Mem/memory_reg[24][11]  ( .D(\Data_Mem/n5475 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[779]), .Q(data_mem_out_wire[779]) );
  DFF \Data_Mem/memory_reg[24][12]  ( .D(\Data_Mem/n5476 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[780]), .Q(data_mem_out_wire[780]) );
  DFF \Data_Mem/memory_reg[24][13]  ( .D(\Data_Mem/n5477 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[781]), .Q(data_mem_out_wire[781]) );
  DFF \Data_Mem/memory_reg[24][14]  ( .D(\Data_Mem/n5478 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[782]), .Q(data_mem_out_wire[782]) );
  DFF \Data_Mem/memory_reg[24][15]  ( .D(\Data_Mem/n5479 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[783]), .Q(data_mem_out_wire[783]) );
  DFF \Data_Mem/memory_reg[24][16]  ( .D(\Data_Mem/n5480 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[784]), .Q(data_mem_out_wire[784]) );
  DFF \Data_Mem/memory_reg[24][17]  ( .D(\Data_Mem/n5481 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[785]), .Q(data_mem_out_wire[785]) );
  DFF \Data_Mem/memory_reg[24][18]  ( .D(\Data_Mem/n5482 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[786]), .Q(data_mem_out_wire[786]) );
  DFF \Data_Mem/memory_reg[24][19]  ( .D(\Data_Mem/n5483 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[787]), .Q(data_mem_out_wire[787]) );
  DFF \Data_Mem/memory_reg[24][20]  ( .D(\Data_Mem/n5484 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[788]), .Q(data_mem_out_wire[788]) );
  DFF \Data_Mem/memory_reg[24][21]  ( .D(\Data_Mem/n5485 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[789]), .Q(data_mem_out_wire[789]) );
  DFF \Data_Mem/memory_reg[24][22]  ( .D(\Data_Mem/n5486 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[790]), .Q(data_mem_out_wire[790]) );
  DFF \Data_Mem/memory_reg[24][23]  ( .D(\Data_Mem/n5487 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[791]), .Q(data_mem_out_wire[791]) );
  DFF \Data_Mem/memory_reg[24][24]  ( .D(\Data_Mem/n5488 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[792]), .Q(data_mem_out_wire[792]) );
  DFF \Data_Mem/memory_reg[24][25]  ( .D(\Data_Mem/n5489 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[793]), .Q(data_mem_out_wire[793]) );
  DFF \Data_Mem/memory_reg[24][26]  ( .D(\Data_Mem/n5490 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[794]), .Q(data_mem_out_wire[794]) );
  DFF \Data_Mem/memory_reg[24][27]  ( .D(\Data_Mem/n5491 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[795]), .Q(data_mem_out_wire[795]) );
  DFF \Data_Mem/memory_reg[24][28]  ( .D(\Data_Mem/n5492 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[796]), .Q(data_mem_out_wire[796]) );
  DFF \Data_Mem/memory_reg[24][29]  ( .D(\Data_Mem/n5493 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[797]), .Q(data_mem_out_wire[797]) );
  DFF \Data_Mem/memory_reg[24][30]  ( .D(\Data_Mem/n5494 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[798]), .Q(data_mem_out_wire[798]) );
  DFF \Data_Mem/memory_reg[24][31]  ( .D(\Data_Mem/n5495 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[799]), .Q(data_mem_out_wire[799]) );
  DFF \Data_Mem/memory_reg[23][0]  ( .D(\Data_Mem/n5496 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[736]), .Q(data_mem_out_wire[736]) );
  DFF \Data_Mem/memory_reg[23][1]  ( .D(\Data_Mem/n5497 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[737]), .Q(data_mem_out_wire[737]) );
  DFF \Data_Mem/memory_reg[23][2]  ( .D(\Data_Mem/n5498 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[738]), .Q(data_mem_out_wire[738]) );
  DFF \Data_Mem/memory_reg[23][3]  ( .D(\Data_Mem/n5499 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[739]), .Q(data_mem_out_wire[739]) );
  DFF \Data_Mem/memory_reg[23][4]  ( .D(\Data_Mem/n5500 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[740]), .Q(data_mem_out_wire[740]) );
  DFF \Data_Mem/memory_reg[23][5]  ( .D(\Data_Mem/n5501 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[741]), .Q(data_mem_out_wire[741]) );
  DFF \Data_Mem/memory_reg[23][6]  ( .D(\Data_Mem/n5502 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[742]), .Q(data_mem_out_wire[742]) );
  DFF \Data_Mem/memory_reg[23][7]  ( .D(\Data_Mem/n5503 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[743]), .Q(data_mem_out_wire[743]) );
  DFF \Data_Mem/memory_reg[23][8]  ( .D(\Data_Mem/n5504 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[744]), .Q(data_mem_out_wire[744]) );
  DFF \Data_Mem/memory_reg[23][9]  ( .D(\Data_Mem/n5505 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[745]), .Q(data_mem_out_wire[745]) );
  DFF \Data_Mem/memory_reg[23][10]  ( .D(\Data_Mem/n5506 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[746]), .Q(data_mem_out_wire[746]) );
  DFF \Data_Mem/memory_reg[23][11]  ( .D(\Data_Mem/n5507 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[747]), .Q(data_mem_out_wire[747]) );
  DFF \Data_Mem/memory_reg[23][12]  ( .D(\Data_Mem/n5508 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[748]), .Q(data_mem_out_wire[748]) );
  DFF \Data_Mem/memory_reg[23][13]  ( .D(\Data_Mem/n5509 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[749]), .Q(data_mem_out_wire[749]) );
  DFF \Data_Mem/memory_reg[23][14]  ( .D(\Data_Mem/n5510 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[750]), .Q(data_mem_out_wire[750]) );
  DFF \Data_Mem/memory_reg[23][15]  ( .D(\Data_Mem/n5511 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[751]), .Q(data_mem_out_wire[751]) );
  DFF \Data_Mem/memory_reg[23][16]  ( .D(\Data_Mem/n5512 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[752]), .Q(data_mem_out_wire[752]) );
  DFF \Data_Mem/memory_reg[23][17]  ( .D(\Data_Mem/n5513 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[753]), .Q(data_mem_out_wire[753]) );
  DFF \Data_Mem/memory_reg[23][18]  ( .D(\Data_Mem/n5514 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[754]), .Q(data_mem_out_wire[754]) );
  DFF \Data_Mem/memory_reg[23][19]  ( .D(\Data_Mem/n5515 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[755]), .Q(data_mem_out_wire[755]) );
  DFF \Data_Mem/memory_reg[23][20]  ( .D(\Data_Mem/n5516 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[756]), .Q(data_mem_out_wire[756]) );
  DFF \Data_Mem/memory_reg[23][21]  ( .D(\Data_Mem/n5517 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[757]), .Q(data_mem_out_wire[757]) );
  DFF \Data_Mem/memory_reg[23][22]  ( .D(\Data_Mem/n5518 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[758]), .Q(data_mem_out_wire[758]) );
  DFF \Data_Mem/memory_reg[23][23]  ( .D(\Data_Mem/n5519 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[759]), .Q(data_mem_out_wire[759]) );
  DFF \Data_Mem/memory_reg[23][24]  ( .D(\Data_Mem/n5520 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[760]), .Q(data_mem_out_wire[760]) );
  DFF \Data_Mem/memory_reg[23][25]  ( .D(\Data_Mem/n5521 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[761]), .Q(data_mem_out_wire[761]) );
  DFF \Data_Mem/memory_reg[23][26]  ( .D(\Data_Mem/n5522 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[762]), .Q(data_mem_out_wire[762]) );
  DFF \Data_Mem/memory_reg[23][27]  ( .D(\Data_Mem/n5523 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[763]), .Q(data_mem_out_wire[763]) );
  DFF \Data_Mem/memory_reg[23][28]  ( .D(\Data_Mem/n5524 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[764]), .Q(data_mem_out_wire[764]) );
  DFF \Data_Mem/memory_reg[23][29]  ( .D(\Data_Mem/n5525 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[765]), .Q(data_mem_out_wire[765]) );
  DFF \Data_Mem/memory_reg[23][30]  ( .D(\Data_Mem/n5526 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[766]), .Q(data_mem_out_wire[766]) );
  DFF \Data_Mem/memory_reg[23][31]  ( .D(\Data_Mem/n5527 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[767]), .Q(data_mem_out_wire[767]) );
  DFF \Data_Mem/memory_reg[22][0]  ( .D(\Data_Mem/n5528 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[704]), .Q(data_mem_out_wire[704]) );
  DFF \Data_Mem/memory_reg[22][1]  ( .D(\Data_Mem/n5529 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[705]), .Q(data_mem_out_wire[705]) );
  DFF \Data_Mem/memory_reg[22][2]  ( .D(\Data_Mem/n5530 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[706]), .Q(data_mem_out_wire[706]) );
  DFF \Data_Mem/memory_reg[22][3]  ( .D(\Data_Mem/n5531 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[707]), .Q(data_mem_out_wire[707]) );
  DFF \Data_Mem/memory_reg[22][4]  ( .D(\Data_Mem/n5532 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[708]), .Q(data_mem_out_wire[708]) );
  DFF \Data_Mem/memory_reg[22][5]  ( .D(\Data_Mem/n5533 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[709]), .Q(data_mem_out_wire[709]) );
  DFF \Data_Mem/memory_reg[22][6]  ( .D(\Data_Mem/n5534 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[710]), .Q(data_mem_out_wire[710]) );
  DFF \Data_Mem/memory_reg[22][7]  ( .D(\Data_Mem/n5535 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[711]), .Q(data_mem_out_wire[711]) );
  DFF \Data_Mem/memory_reg[22][8]  ( .D(\Data_Mem/n5536 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[712]), .Q(data_mem_out_wire[712]) );
  DFF \Data_Mem/memory_reg[22][9]  ( .D(\Data_Mem/n5537 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[713]), .Q(data_mem_out_wire[713]) );
  DFF \Data_Mem/memory_reg[22][10]  ( .D(\Data_Mem/n5538 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[714]), .Q(data_mem_out_wire[714]) );
  DFF \Data_Mem/memory_reg[22][11]  ( .D(\Data_Mem/n5539 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[715]), .Q(data_mem_out_wire[715]) );
  DFF \Data_Mem/memory_reg[22][12]  ( .D(\Data_Mem/n5540 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[716]), .Q(data_mem_out_wire[716]) );
  DFF \Data_Mem/memory_reg[22][13]  ( .D(\Data_Mem/n5541 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[717]), .Q(data_mem_out_wire[717]) );
  DFF \Data_Mem/memory_reg[22][14]  ( .D(\Data_Mem/n5542 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[718]), .Q(data_mem_out_wire[718]) );
  DFF \Data_Mem/memory_reg[22][15]  ( .D(\Data_Mem/n5543 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[719]), .Q(data_mem_out_wire[719]) );
  DFF \Data_Mem/memory_reg[22][16]  ( .D(\Data_Mem/n5544 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[720]), .Q(data_mem_out_wire[720]) );
  DFF \Data_Mem/memory_reg[22][17]  ( .D(\Data_Mem/n5545 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[721]), .Q(data_mem_out_wire[721]) );
  DFF \Data_Mem/memory_reg[22][18]  ( .D(\Data_Mem/n5546 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[722]), .Q(data_mem_out_wire[722]) );
  DFF \Data_Mem/memory_reg[22][19]  ( .D(\Data_Mem/n5547 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[723]), .Q(data_mem_out_wire[723]) );
  DFF \Data_Mem/memory_reg[22][20]  ( .D(\Data_Mem/n5548 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[724]), .Q(data_mem_out_wire[724]) );
  DFF \Data_Mem/memory_reg[22][21]  ( .D(\Data_Mem/n5549 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[725]), .Q(data_mem_out_wire[725]) );
  DFF \Data_Mem/memory_reg[22][22]  ( .D(\Data_Mem/n5550 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[726]), .Q(data_mem_out_wire[726]) );
  DFF \Data_Mem/memory_reg[22][23]  ( .D(\Data_Mem/n5551 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[727]), .Q(data_mem_out_wire[727]) );
  DFF \Data_Mem/memory_reg[22][24]  ( .D(\Data_Mem/n5552 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[728]), .Q(data_mem_out_wire[728]) );
  DFF \Data_Mem/memory_reg[22][25]  ( .D(\Data_Mem/n5553 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[729]), .Q(data_mem_out_wire[729]) );
  DFF \Data_Mem/memory_reg[22][26]  ( .D(\Data_Mem/n5554 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[730]), .Q(data_mem_out_wire[730]) );
  DFF \Data_Mem/memory_reg[22][27]  ( .D(\Data_Mem/n5555 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[731]), .Q(data_mem_out_wire[731]) );
  DFF \Data_Mem/memory_reg[22][28]  ( .D(\Data_Mem/n5556 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[732]), .Q(data_mem_out_wire[732]) );
  DFF \Data_Mem/memory_reg[22][29]  ( .D(\Data_Mem/n5557 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[733]), .Q(data_mem_out_wire[733]) );
  DFF \Data_Mem/memory_reg[22][30]  ( .D(\Data_Mem/n5558 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[734]), .Q(data_mem_out_wire[734]) );
  DFF \Data_Mem/memory_reg[22][31]  ( .D(\Data_Mem/n5559 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[735]), .Q(data_mem_out_wire[735]) );
  DFF \Data_Mem/memory_reg[21][0]  ( .D(\Data_Mem/n5560 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[672]), .Q(data_mem_out_wire[672]) );
  DFF \Data_Mem/memory_reg[21][1]  ( .D(\Data_Mem/n5561 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[673]), .Q(data_mem_out_wire[673]) );
  DFF \Data_Mem/memory_reg[21][2]  ( .D(\Data_Mem/n5562 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[674]), .Q(data_mem_out_wire[674]) );
  DFF \Data_Mem/memory_reg[21][3]  ( .D(\Data_Mem/n5563 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[675]), .Q(data_mem_out_wire[675]) );
  DFF \Data_Mem/memory_reg[21][4]  ( .D(\Data_Mem/n5564 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[676]), .Q(data_mem_out_wire[676]) );
  DFF \Data_Mem/memory_reg[21][5]  ( .D(\Data_Mem/n5565 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[677]), .Q(data_mem_out_wire[677]) );
  DFF \Data_Mem/memory_reg[21][6]  ( .D(\Data_Mem/n5566 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[678]), .Q(data_mem_out_wire[678]) );
  DFF \Data_Mem/memory_reg[21][7]  ( .D(\Data_Mem/n5567 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[679]), .Q(data_mem_out_wire[679]) );
  DFF \Data_Mem/memory_reg[21][8]  ( .D(\Data_Mem/n5568 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[680]), .Q(data_mem_out_wire[680]) );
  DFF \Data_Mem/memory_reg[21][9]  ( .D(\Data_Mem/n5569 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[681]), .Q(data_mem_out_wire[681]) );
  DFF \Data_Mem/memory_reg[21][10]  ( .D(\Data_Mem/n5570 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[682]), .Q(data_mem_out_wire[682]) );
  DFF \Data_Mem/memory_reg[21][11]  ( .D(\Data_Mem/n5571 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[683]), .Q(data_mem_out_wire[683]) );
  DFF \Data_Mem/memory_reg[21][12]  ( .D(\Data_Mem/n5572 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[684]), .Q(data_mem_out_wire[684]) );
  DFF \Data_Mem/memory_reg[21][13]  ( .D(\Data_Mem/n5573 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[685]), .Q(data_mem_out_wire[685]) );
  DFF \Data_Mem/memory_reg[21][14]  ( .D(\Data_Mem/n5574 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[686]), .Q(data_mem_out_wire[686]) );
  DFF \Data_Mem/memory_reg[21][15]  ( .D(\Data_Mem/n5575 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[687]), .Q(data_mem_out_wire[687]) );
  DFF \Data_Mem/memory_reg[21][16]  ( .D(\Data_Mem/n5576 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[688]), .Q(data_mem_out_wire[688]) );
  DFF \Data_Mem/memory_reg[21][17]  ( .D(\Data_Mem/n5577 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[689]), .Q(data_mem_out_wire[689]) );
  DFF \Data_Mem/memory_reg[21][18]  ( .D(\Data_Mem/n5578 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[690]), .Q(data_mem_out_wire[690]) );
  DFF \Data_Mem/memory_reg[21][19]  ( .D(\Data_Mem/n5579 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[691]), .Q(data_mem_out_wire[691]) );
  DFF \Data_Mem/memory_reg[21][20]  ( .D(\Data_Mem/n5580 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[692]), .Q(data_mem_out_wire[692]) );
  DFF \Data_Mem/memory_reg[21][21]  ( .D(\Data_Mem/n5581 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[693]), .Q(data_mem_out_wire[693]) );
  DFF \Data_Mem/memory_reg[21][22]  ( .D(\Data_Mem/n5582 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[694]), .Q(data_mem_out_wire[694]) );
  DFF \Data_Mem/memory_reg[21][23]  ( .D(\Data_Mem/n5583 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[695]), .Q(data_mem_out_wire[695]) );
  DFF \Data_Mem/memory_reg[21][24]  ( .D(\Data_Mem/n5584 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[696]), .Q(data_mem_out_wire[696]) );
  DFF \Data_Mem/memory_reg[21][25]  ( .D(\Data_Mem/n5585 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[697]), .Q(data_mem_out_wire[697]) );
  DFF \Data_Mem/memory_reg[21][26]  ( .D(\Data_Mem/n5586 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[698]), .Q(data_mem_out_wire[698]) );
  DFF \Data_Mem/memory_reg[21][27]  ( .D(\Data_Mem/n5587 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[699]), .Q(data_mem_out_wire[699]) );
  DFF \Data_Mem/memory_reg[21][28]  ( .D(\Data_Mem/n5588 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[700]), .Q(data_mem_out_wire[700]) );
  DFF \Data_Mem/memory_reg[21][29]  ( .D(\Data_Mem/n5589 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[701]), .Q(data_mem_out_wire[701]) );
  DFF \Data_Mem/memory_reg[21][30]  ( .D(\Data_Mem/n5590 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[702]), .Q(data_mem_out_wire[702]) );
  DFF \Data_Mem/memory_reg[21][31]  ( .D(\Data_Mem/n5591 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[703]), .Q(data_mem_out_wire[703]) );
  DFF \Data_Mem/memory_reg[20][0]  ( .D(\Data_Mem/n5592 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[640]), .Q(data_mem_out_wire[640]) );
  DFF \Data_Mem/memory_reg[20][1]  ( .D(\Data_Mem/n5593 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[641]), .Q(data_mem_out_wire[641]) );
  DFF \Data_Mem/memory_reg[20][2]  ( .D(\Data_Mem/n5594 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[642]), .Q(data_mem_out_wire[642]) );
  DFF \Data_Mem/memory_reg[20][3]  ( .D(\Data_Mem/n5595 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[643]), .Q(data_mem_out_wire[643]) );
  DFF \Data_Mem/memory_reg[20][4]  ( .D(\Data_Mem/n5596 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[644]), .Q(data_mem_out_wire[644]) );
  DFF \Data_Mem/memory_reg[20][5]  ( .D(\Data_Mem/n5597 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[645]), .Q(data_mem_out_wire[645]) );
  DFF \Data_Mem/memory_reg[20][6]  ( .D(\Data_Mem/n5598 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[646]), .Q(data_mem_out_wire[646]) );
  DFF \Data_Mem/memory_reg[20][7]  ( .D(\Data_Mem/n5599 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[647]), .Q(data_mem_out_wire[647]) );
  DFF \Data_Mem/memory_reg[20][8]  ( .D(\Data_Mem/n5600 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[648]), .Q(data_mem_out_wire[648]) );
  DFF \Data_Mem/memory_reg[20][9]  ( .D(\Data_Mem/n5601 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[649]), .Q(data_mem_out_wire[649]) );
  DFF \Data_Mem/memory_reg[20][10]  ( .D(\Data_Mem/n5602 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[650]), .Q(data_mem_out_wire[650]) );
  DFF \Data_Mem/memory_reg[20][11]  ( .D(\Data_Mem/n5603 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[651]), .Q(data_mem_out_wire[651]) );
  DFF \Data_Mem/memory_reg[20][12]  ( .D(\Data_Mem/n5604 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[652]), .Q(data_mem_out_wire[652]) );
  DFF \Data_Mem/memory_reg[20][13]  ( .D(\Data_Mem/n5605 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[653]), .Q(data_mem_out_wire[653]) );
  DFF \Data_Mem/memory_reg[20][14]  ( .D(\Data_Mem/n5606 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[654]), .Q(data_mem_out_wire[654]) );
  DFF \Data_Mem/memory_reg[20][15]  ( .D(\Data_Mem/n5607 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[655]), .Q(data_mem_out_wire[655]) );
  DFF \Data_Mem/memory_reg[20][16]  ( .D(\Data_Mem/n5608 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[656]), .Q(data_mem_out_wire[656]) );
  DFF \Data_Mem/memory_reg[20][17]  ( .D(\Data_Mem/n5609 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[657]), .Q(data_mem_out_wire[657]) );
  DFF \Data_Mem/memory_reg[20][18]  ( .D(\Data_Mem/n5610 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[658]), .Q(data_mem_out_wire[658]) );
  DFF \Data_Mem/memory_reg[20][19]  ( .D(\Data_Mem/n5611 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[659]), .Q(data_mem_out_wire[659]) );
  DFF \Data_Mem/memory_reg[20][20]  ( .D(\Data_Mem/n5612 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[660]), .Q(data_mem_out_wire[660]) );
  DFF \Data_Mem/memory_reg[20][21]  ( .D(\Data_Mem/n5613 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[661]), .Q(data_mem_out_wire[661]) );
  DFF \Data_Mem/memory_reg[20][22]  ( .D(\Data_Mem/n5614 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[662]), .Q(data_mem_out_wire[662]) );
  DFF \Data_Mem/memory_reg[20][23]  ( .D(\Data_Mem/n5615 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[663]), .Q(data_mem_out_wire[663]) );
  DFF \Data_Mem/memory_reg[20][24]  ( .D(\Data_Mem/n5616 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[664]), .Q(data_mem_out_wire[664]) );
  DFF \Data_Mem/memory_reg[20][25]  ( .D(\Data_Mem/n5617 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[665]), .Q(data_mem_out_wire[665]) );
  DFF \Data_Mem/memory_reg[20][26]  ( .D(\Data_Mem/n5618 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[666]), .Q(data_mem_out_wire[666]) );
  DFF \Data_Mem/memory_reg[20][27]  ( .D(\Data_Mem/n5619 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[667]), .Q(data_mem_out_wire[667]) );
  DFF \Data_Mem/memory_reg[20][28]  ( .D(\Data_Mem/n5620 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[668]), .Q(data_mem_out_wire[668]) );
  DFF \Data_Mem/memory_reg[20][29]  ( .D(\Data_Mem/n5621 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[669]), .Q(data_mem_out_wire[669]) );
  DFF \Data_Mem/memory_reg[20][30]  ( .D(\Data_Mem/n5622 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[670]), .Q(data_mem_out_wire[670]) );
  DFF \Data_Mem/memory_reg[20][31]  ( .D(\Data_Mem/n5623 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[671]), .Q(data_mem_out_wire[671]) );
  DFF \Data_Mem/memory_reg[19][0]  ( .D(\Data_Mem/n5624 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[608]), .Q(data_mem_out_wire[608]) );
  DFF \Data_Mem/memory_reg[19][1]  ( .D(\Data_Mem/n5625 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[609]), .Q(data_mem_out_wire[609]) );
  DFF \Data_Mem/memory_reg[19][2]  ( .D(\Data_Mem/n5626 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[610]), .Q(data_mem_out_wire[610]) );
  DFF \Data_Mem/memory_reg[19][3]  ( .D(\Data_Mem/n5627 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[611]), .Q(data_mem_out_wire[611]) );
  DFF \Data_Mem/memory_reg[19][4]  ( .D(\Data_Mem/n5628 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[612]), .Q(data_mem_out_wire[612]) );
  DFF \Data_Mem/memory_reg[19][5]  ( .D(\Data_Mem/n5629 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[613]), .Q(data_mem_out_wire[613]) );
  DFF \Data_Mem/memory_reg[19][6]  ( .D(\Data_Mem/n5630 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[614]), .Q(data_mem_out_wire[614]) );
  DFF \Data_Mem/memory_reg[19][7]  ( .D(\Data_Mem/n5631 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[615]), .Q(data_mem_out_wire[615]) );
  DFF \Data_Mem/memory_reg[19][8]  ( .D(\Data_Mem/n5632 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[616]), .Q(data_mem_out_wire[616]) );
  DFF \Data_Mem/memory_reg[19][9]  ( .D(\Data_Mem/n5633 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[617]), .Q(data_mem_out_wire[617]) );
  DFF \Data_Mem/memory_reg[19][10]  ( .D(\Data_Mem/n5634 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[618]), .Q(data_mem_out_wire[618]) );
  DFF \Data_Mem/memory_reg[19][11]  ( .D(\Data_Mem/n5635 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[619]), .Q(data_mem_out_wire[619]) );
  DFF \Data_Mem/memory_reg[19][12]  ( .D(\Data_Mem/n5636 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[620]), .Q(data_mem_out_wire[620]) );
  DFF \Data_Mem/memory_reg[19][13]  ( .D(\Data_Mem/n5637 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[621]), .Q(data_mem_out_wire[621]) );
  DFF \Data_Mem/memory_reg[19][14]  ( .D(\Data_Mem/n5638 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[622]), .Q(data_mem_out_wire[622]) );
  DFF \Data_Mem/memory_reg[19][15]  ( .D(\Data_Mem/n5639 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[623]), .Q(data_mem_out_wire[623]) );
  DFF \Data_Mem/memory_reg[19][16]  ( .D(\Data_Mem/n5640 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[624]), .Q(data_mem_out_wire[624]) );
  DFF \Data_Mem/memory_reg[19][17]  ( .D(\Data_Mem/n5641 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[625]), .Q(data_mem_out_wire[625]) );
  DFF \Data_Mem/memory_reg[19][18]  ( .D(\Data_Mem/n5642 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[626]), .Q(data_mem_out_wire[626]) );
  DFF \Data_Mem/memory_reg[19][19]  ( .D(\Data_Mem/n5643 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[627]), .Q(data_mem_out_wire[627]) );
  DFF \Data_Mem/memory_reg[19][20]  ( .D(\Data_Mem/n5644 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[628]), .Q(data_mem_out_wire[628]) );
  DFF \Data_Mem/memory_reg[19][21]  ( .D(\Data_Mem/n5645 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[629]), .Q(data_mem_out_wire[629]) );
  DFF \Data_Mem/memory_reg[19][22]  ( .D(\Data_Mem/n5646 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[630]), .Q(data_mem_out_wire[630]) );
  DFF \Data_Mem/memory_reg[19][23]  ( .D(\Data_Mem/n5647 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[631]), .Q(data_mem_out_wire[631]) );
  DFF \Data_Mem/memory_reg[19][24]  ( .D(\Data_Mem/n5648 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[632]), .Q(data_mem_out_wire[632]) );
  DFF \Data_Mem/memory_reg[19][25]  ( .D(\Data_Mem/n5649 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[633]), .Q(data_mem_out_wire[633]) );
  DFF \Data_Mem/memory_reg[19][26]  ( .D(\Data_Mem/n5650 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[634]), .Q(data_mem_out_wire[634]) );
  DFF \Data_Mem/memory_reg[19][27]  ( .D(\Data_Mem/n5651 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[635]), .Q(data_mem_out_wire[635]) );
  DFF \Data_Mem/memory_reg[19][28]  ( .D(\Data_Mem/n5652 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[636]), .Q(data_mem_out_wire[636]) );
  DFF \Data_Mem/memory_reg[19][29]  ( .D(\Data_Mem/n5653 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[637]), .Q(data_mem_out_wire[637]) );
  DFF \Data_Mem/memory_reg[19][30]  ( .D(\Data_Mem/n5654 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[638]), .Q(data_mem_out_wire[638]) );
  DFF \Data_Mem/memory_reg[19][31]  ( .D(\Data_Mem/n5655 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[639]), .Q(data_mem_out_wire[639]) );
  DFF \Data_Mem/memory_reg[18][0]  ( .D(\Data_Mem/n5656 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[576]), .Q(data_mem_out_wire[576]) );
  DFF \Data_Mem/memory_reg[18][1]  ( .D(\Data_Mem/n5657 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[577]), .Q(data_mem_out_wire[577]) );
  DFF \Data_Mem/memory_reg[18][2]  ( .D(\Data_Mem/n5658 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[578]), .Q(data_mem_out_wire[578]) );
  DFF \Data_Mem/memory_reg[18][3]  ( .D(\Data_Mem/n5659 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[579]), .Q(data_mem_out_wire[579]) );
  DFF \Data_Mem/memory_reg[18][4]  ( .D(\Data_Mem/n5660 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[580]), .Q(data_mem_out_wire[580]) );
  DFF \Data_Mem/memory_reg[18][5]  ( .D(\Data_Mem/n5661 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[581]), .Q(data_mem_out_wire[581]) );
  DFF \Data_Mem/memory_reg[18][6]  ( .D(\Data_Mem/n5662 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[582]), .Q(data_mem_out_wire[582]) );
  DFF \Data_Mem/memory_reg[18][7]  ( .D(\Data_Mem/n5663 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[583]), .Q(data_mem_out_wire[583]) );
  DFF \Data_Mem/memory_reg[18][8]  ( .D(\Data_Mem/n5664 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[584]), .Q(data_mem_out_wire[584]) );
  DFF \Data_Mem/memory_reg[18][9]  ( .D(\Data_Mem/n5665 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[585]), .Q(data_mem_out_wire[585]) );
  DFF \Data_Mem/memory_reg[18][10]  ( .D(\Data_Mem/n5666 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[586]), .Q(data_mem_out_wire[586]) );
  DFF \Data_Mem/memory_reg[18][11]  ( .D(\Data_Mem/n5667 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[587]), .Q(data_mem_out_wire[587]) );
  DFF \Data_Mem/memory_reg[18][12]  ( .D(\Data_Mem/n5668 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[588]), .Q(data_mem_out_wire[588]) );
  DFF \Data_Mem/memory_reg[18][13]  ( .D(\Data_Mem/n5669 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[589]), .Q(data_mem_out_wire[589]) );
  DFF \Data_Mem/memory_reg[18][14]  ( .D(\Data_Mem/n5670 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[590]), .Q(data_mem_out_wire[590]) );
  DFF \Data_Mem/memory_reg[18][15]  ( .D(\Data_Mem/n5671 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[591]), .Q(data_mem_out_wire[591]) );
  DFF \Data_Mem/memory_reg[18][16]  ( .D(\Data_Mem/n5672 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[592]), .Q(data_mem_out_wire[592]) );
  DFF \Data_Mem/memory_reg[18][17]  ( .D(\Data_Mem/n5673 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[593]), .Q(data_mem_out_wire[593]) );
  DFF \Data_Mem/memory_reg[18][18]  ( .D(\Data_Mem/n5674 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[594]), .Q(data_mem_out_wire[594]) );
  DFF \Data_Mem/memory_reg[18][19]  ( .D(\Data_Mem/n5675 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[595]), .Q(data_mem_out_wire[595]) );
  DFF \Data_Mem/memory_reg[18][20]  ( .D(\Data_Mem/n5676 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[596]), .Q(data_mem_out_wire[596]) );
  DFF \Data_Mem/memory_reg[18][21]  ( .D(\Data_Mem/n5677 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[597]), .Q(data_mem_out_wire[597]) );
  DFF \Data_Mem/memory_reg[18][22]  ( .D(\Data_Mem/n5678 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[598]), .Q(data_mem_out_wire[598]) );
  DFF \Data_Mem/memory_reg[18][23]  ( .D(\Data_Mem/n5679 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[599]), .Q(data_mem_out_wire[599]) );
  DFF \Data_Mem/memory_reg[18][24]  ( .D(\Data_Mem/n5680 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[600]), .Q(data_mem_out_wire[600]) );
  DFF \Data_Mem/memory_reg[18][25]  ( .D(\Data_Mem/n5681 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[601]), .Q(data_mem_out_wire[601]) );
  DFF \Data_Mem/memory_reg[18][26]  ( .D(\Data_Mem/n5682 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[602]), .Q(data_mem_out_wire[602]) );
  DFF \Data_Mem/memory_reg[18][27]  ( .D(\Data_Mem/n5683 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[603]), .Q(data_mem_out_wire[603]) );
  DFF \Data_Mem/memory_reg[18][28]  ( .D(\Data_Mem/n5684 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[604]), .Q(data_mem_out_wire[604]) );
  DFF \Data_Mem/memory_reg[18][29]  ( .D(\Data_Mem/n5685 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[605]), .Q(data_mem_out_wire[605]) );
  DFF \Data_Mem/memory_reg[18][30]  ( .D(\Data_Mem/n5686 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[606]), .Q(data_mem_out_wire[606]) );
  DFF \Data_Mem/memory_reg[18][31]  ( .D(\Data_Mem/n5687 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[607]), .Q(data_mem_out_wire[607]) );
  DFF \Data_Mem/memory_reg[17][0]  ( .D(\Data_Mem/n5688 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[544]), .Q(data_mem_out_wire[544]) );
  DFF \Data_Mem/memory_reg[17][1]  ( .D(\Data_Mem/n5689 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[545]), .Q(data_mem_out_wire[545]) );
  DFF \Data_Mem/memory_reg[17][2]  ( .D(\Data_Mem/n5690 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[546]), .Q(data_mem_out_wire[546]) );
  DFF \Data_Mem/memory_reg[17][3]  ( .D(\Data_Mem/n5691 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[547]), .Q(data_mem_out_wire[547]) );
  DFF \Data_Mem/memory_reg[17][4]  ( .D(\Data_Mem/n5692 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[548]), .Q(data_mem_out_wire[548]) );
  DFF \Data_Mem/memory_reg[17][5]  ( .D(\Data_Mem/n5693 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[549]), .Q(data_mem_out_wire[549]) );
  DFF \Data_Mem/memory_reg[17][6]  ( .D(\Data_Mem/n5694 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[550]), .Q(data_mem_out_wire[550]) );
  DFF \Data_Mem/memory_reg[17][7]  ( .D(\Data_Mem/n5695 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[551]), .Q(data_mem_out_wire[551]) );
  DFF \Data_Mem/memory_reg[17][8]  ( .D(\Data_Mem/n5696 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[552]), .Q(data_mem_out_wire[552]) );
  DFF \Data_Mem/memory_reg[17][9]  ( .D(\Data_Mem/n5697 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[553]), .Q(data_mem_out_wire[553]) );
  DFF \Data_Mem/memory_reg[17][10]  ( .D(\Data_Mem/n5698 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[554]), .Q(data_mem_out_wire[554]) );
  DFF \Data_Mem/memory_reg[17][11]  ( .D(\Data_Mem/n5699 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[555]), .Q(data_mem_out_wire[555]) );
  DFF \Data_Mem/memory_reg[17][12]  ( .D(\Data_Mem/n5700 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[556]), .Q(data_mem_out_wire[556]) );
  DFF \Data_Mem/memory_reg[17][13]  ( .D(\Data_Mem/n5701 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[557]), .Q(data_mem_out_wire[557]) );
  DFF \Data_Mem/memory_reg[17][14]  ( .D(\Data_Mem/n5702 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[558]), .Q(data_mem_out_wire[558]) );
  DFF \Data_Mem/memory_reg[17][15]  ( .D(\Data_Mem/n5703 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[559]), .Q(data_mem_out_wire[559]) );
  DFF \Data_Mem/memory_reg[17][16]  ( .D(\Data_Mem/n5704 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[560]), .Q(data_mem_out_wire[560]) );
  DFF \Data_Mem/memory_reg[17][17]  ( .D(\Data_Mem/n5705 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[561]), .Q(data_mem_out_wire[561]) );
  DFF \Data_Mem/memory_reg[17][18]  ( .D(\Data_Mem/n5706 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[562]), .Q(data_mem_out_wire[562]) );
  DFF \Data_Mem/memory_reg[17][19]  ( .D(\Data_Mem/n5707 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[563]), .Q(data_mem_out_wire[563]) );
  DFF \Data_Mem/memory_reg[17][20]  ( .D(\Data_Mem/n5708 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[564]), .Q(data_mem_out_wire[564]) );
  DFF \Data_Mem/memory_reg[17][21]  ( .D(\Data_Mem/n5709 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[565]), .Q(data_mem_out_wire[565]) );
  DFF \Data_Mem/memory_reg[17][22]  ( .D(\Data_Mem/n5710 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[566]), .Q(data_mem_out_wire[566]) );
  DFF \Data_Mem/memory_reg[17][23]  ( .D(\Data_Mem/n5711 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[567]), .Q(data_mem_out_wire[567]) );
  DFF \Data_Mem/memory_reg[17][24]  ( .D(\Data_Mem/n5712 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[568]), .Q(data_mem_out_wire[568]) );
  DFF \Data_Mem/memory_reg[17][25]  ( .D(\Data_Mem/n5713 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[569]), .Q(data_mem_out_wire[569]) );
  DFF \Data_Mem/memory_reg[17][26]  ( .D(\Data_Mem/n5714 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[570]), .Q(data_mem_out_wire[570]) );
  DFF \Data_Mem/memory_reg[17][27]  ( .D(\Data_Mem/n5715 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[571]), .Q(data_mem_out_wire[571]) );
  DFF \Data_Mem/memory_reg[17][28]  ( .D(\Data_Mem/n5716 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[572]), .Q(data_mem_out_wire[572]) );
  DFF \Data_Mem/memory_reg[17][29]  ( .D(\Data_Mem/n5717 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[573]), .Q(data_mem_out_wire[573]) );
  DFF \Data_Mem/memory_reg[17][30]  ( .D(\Data_Mem/n5718 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[574]), .Q(data_mem_out_wire[574]) );
  DFF \Data_Mem/memory_reg[17][31]  ( .D(\Data_Mem/n5719 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[575]), .Q(data_mem_out_wire[575]) );
  DFF \Data_Mem/memory_reg[16][0]  ( .D(\Data_Mem/n5720 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[512]), .Q(data_mem_out_wire[512]) );
  DFF \Data_Mem/memory_reg[16][1]  ( .D(\Data_Mem/n5721 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[513]), .Q(data_mem_out_wire[513]) );
  DFF \Data_Mem/memory_reg[16][2]  ( .D(\Data_Mem/n5722 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[514]), .Q(data_mem_out_wire[514]) );
  DFF \Data_Mem/memory_reg[16][3]  ( .D(\Data_Mem/n5723 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[515]), .Q(data_mem_out_wire[515]) );
  DFF \Data_Mem/memory_reg[16][4]  ( .D(\Data_Mem/n5724 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[516]), .Q(data_mem_out_wire[516]) );
  DFF \Data_Mem/memory_reg[16][5]  ( .D(\Data_Mem/n5725 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[517]), .Q(data_mem_out_wire[517]) );
  DFF \Data_Mem/memory_reg[16][6]  ( .D(\Data_Mem/n5726 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[518]), .Q(data_mem_out_wire[518]) );
  DFF \Data_Mem/memory_reg[16][7]  ( .D(\Data_Mem/n5727 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[519]), .Q(data_mem_out_wire[519]) );
  DFF \Data_Mem/memory_reg[16][8]  ( .D(\Data_Mem/n5728 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[520]), .Q(data_mem_out_wire[520]) );
  DFF \Data_Mem/memory_reg[16][9]  ( .D(\Data_Mem/n5729 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[521]), .Q(data_mem_out_wire[521]) );
  DFF \Data_Mem/memory_reg[16][10]  ( .D(\Data_Mem/n5730 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[522]), .Q(data_mem_out_wire[522]) );
  DFF \Data_Mem/memory_reg[16][11]  ( .D(\Data_Mem/n5731 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[523]), .Q(data_mem_out_wire[523]) );
  DFF \Data_Mem/memory_reg[16][12]  ( .D(\Data_Mem/n5732 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[524]), .Q(data_mem_out_wire[524]) );
  DFF \Data_Mem/memory_reg[16][13]  ( .D(\Data_Mem/n5733 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[525]), .Q(data_mem_out_wire[525]) );
  DFF \Data_Mem/memory_reg[16][14]  ( .D(\Data_Mem/n5734 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[526]), .Q(data_mem_out_wire[526]) );
  DFF \Data_Mem/memory_reg[16][15]  ( .D(\Data_Mem/n5735 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[527]), .Q(data_mem_out_wire[527]) );
  DFF \Data_Mem/memory_reg[16][16]  ( .D(\Data_Mem/n5736 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[528]), .Q(data_mem_out_wire[528]) );
  DFF \Data_Mem/memory_reg[16][17]  ( .D(\Data_Mem/n5737 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[529]), .Q(data_mem_out_wire[529]) );
  DFF \Data_Mem/memory_reg[16][18]  ( .D(\Data_Mem/n5738 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[530]), .Q(data_mem_out_wire[530]) );
  DFF \Data_Mem/memory_reg[16][19]  ( .D(\Data_Mem/n5739 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[531]), .Q(data_mem_out_wire[531]) );
  DFF \Data_Mem/memory_reg[16][20]  ( .D(\Data_Mem/n5740 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[532]), .Q(data_mem_out_wire[532]) );
  DFF \Data_Mem/memory_reg[16][21]  ( .D(\Data_Mem/n5741 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[533]), .Q(data_mem_out_wire[533]) );
  DFF \Data_Mem/memory_reg[16][22]  ( .D(\Data_Mem/n5742 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[534]), .Q(data_mem_out_wire[534]) );
  DFF \Data_Mem/memory_reg[16][23]  ( .D(\Data_Mem/n5743 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[535]), .Q(data_mem_out_wire[535]) );
  DFF \Data_Mem/memory_reg[16][24]  ( .D(\Data_Mem/n5744 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[536]), .Q(data_mem_out_wire[536]) );
  DFF \Data_Mem/memory_reg[16][25]  ( .D(\Data_Mem/n5745 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[537]), .Q(data_mem_out_wire[537]) );
  DFF \Data_Mem/memory_reg[16][26]  ( .D(\Data_Mem/n5746 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[538]), .Q(data_mem_out_wire[538]) );
  DFF \Data_Mem/memory_reg[16][27]  ( .D(\Data_Mem/n5747 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[539]), .Q(data_mem_out_wire[539]) );
  DFF \Data_Mem/memory_reg[16][28]  ( .D(\Data_Mem/n5748 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[540]), .Q(data_mem_out_wire[540]) );
  DFF \Data_Mem/memory_reg[16][29]  ( .D(\Data_Mem/n5749 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[541]), .Q(data_mem_out_wire[541]) );
  DFF \Data_Mem/memory_reg[16][30]  ( .D(\Data_Mem/n5750 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[542]), .Q(data_mem_out_wire[542]) );
  DFF \Data_Mem/memory_reg[16][31]  ( .D(\Data_Mem/n5751 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[543]), .Q(data_mem_out_wire[543]) );
  DFF \Data_Mem/memory_reg[15][0]  ( .D(\Data_Mem/n5752 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[480]), .Q(data_mem_out_wire[480]) );
  DFF \Data_Mem/memory_reg[15][1]  ( .D(\Data_Mem/n5753 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[481]), .Q(data_mem_out_wire[481]) );
  DFF \Data_Mem/memory_reg[15][2]  ( .D(\Data_Mem/n5754 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[482]), .Q(data_mem_out_wire[482]) );
  DFF \Data_Mem/memory_reg[15][3]  ( .D(\Data_Mem/n5755 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[483]), .Q(data_mem_out_wire[483]) );
  DFF \Data_Mem/memory_reg[15][4]  ( .D(\Data_Mem/n5756 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[484]), .Q(data_mem_out_wire[484]) );
  DFF \Data_Mem/memory_reg[15][5]  ( .D(\Data_Mem/n5757 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[485]), .Q(data_mem_out_wire[485]) );
  DFF \Data_Mem/memory_reg[15][6]  ( .D(\Data_Mem/n5758 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[486]), .Q(data_mem_out_wire[486]) );
  DFF \Data_Mem/memory_reg[15][7]  ( .D(\Data_Mem/n5759 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[487]), .Q(data_mem_out_wire[487]) );
  DFF \Data_Mem/memory_reg[15][8]  ( .D(\Data_Mem/n5760 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[488]), .Q(data_mem_out_wire[488]) );
  DFF \Data_Mem/memory_reg[15][9]  ( .D(\Data_Mem/n5761 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[489]), .Q(data_mem_out_wire[489]) );
  DFF \Data_Mem/memory_reg[15][10]  ( .D(\Data_Mem/n5762 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[490]), .Q(data_mem_out_wire[490]) );
  DFF \Data_Mem/memory_reg[15][11]  ( .D(\Data_Mem/n5763 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[491]), .Q(data_mem_out_wire[491]) );
  DFF \Data_Mem/memory_reg[15][12]  ( .D(\Data_Mem/n5764 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[492]), .Q(data_mem_out_wire[492]) );
  DFF \Data_Mem/memory_reg[15][13]  ( .D(\Data_Mem/n5765 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[493]), .Q(data_mem_out_wire[493]) );
  DFF \Data_Mem/memory_reg[15][14]  ( .D(\Data_Mem/n5766 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[494]), .Q(data_mem_out_wire[494]) );
  DFF \Data_Mem/memory_reg[15][15]  ( .D(\Data_Mem/n5767 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[495]), .Q(data_mem_out_wire[495]) );
  DFF \Data_Mem/memory_reg[15][16]  ( .D(\Data_Mem/n5768 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[496]), .Q(data_mem_out_wire[496]) );
  DFF \Data_Mem/memory_reg[15][17]  ( .D(\Data_Mem/n5769 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[497]), .Q(data_mem_out_wire[497]) );
  DFF \Data_Mem/memory_reg[15][18]  ( .D(\Data_Mem/n5770 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[498]), .Q(data_mem_out_wire[498]) );
  DFF \Data_Mem/memory_reg[15][19]  ( .D(\Data_Mem/n5771 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[499]), .Q(data_mem_out_wire[499]) );
  DFF \Data_Mem/memory_reg[15][20]  ( .D(\Data_Mem/n5772 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[500]), .Q(data_mem_out_wire[500]) );
  DFF \Data_Mem/memory_reg[15][21]  ( .D(\Data_Mem/n5773 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[501]), .Q(data_mem_out_wire[501]) );
  DFF \Data_Mem/memory_reg[15][22]  ( .D(\Data_Mem/n5774 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[502]), .Q(data_mem_out_wire[502]) );
  DFF \Data_Mem/memory_reg[15][23]  ( .D(\Data_Mem/n5775 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[503]), .Q(data_mem_out_wire[503]) );
  DFF \Data_Mem/memory_reg[15][24]  ( .D(\Data_Mem/n5776 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[504]), .Q(data_mem_out_wire[504]) );
  DFF \Data_Mem/memory_reg[15][25]  ( .D(\Data_Mem/n5777 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[505]), .Q(data_mem_out_wire[505]) );
  DFF \Data_Mem/memory_reg[15][26]  ( .D(\Data_Mem/n5778 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[506]), .Q(data_mem_out_wire[506]) );
  DFF \Data_Mem/memory_reg[15][27]  ( .D(\Data_Mem/n5779 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[507]), .Q(data_mem_out_wire[507]) );
  DFF \Data_Mem/memory_reg[15][28]  ( .D(\Data_Mem/n5780 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[508]), .Q(data_mem_out_wire[508]) );
  DFF \Data_Mem/memory_reg[15][29]  ( .D(\Data_Mem/n5781 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[509]), .Q(data_mem_out_wire[509]) );
  DFF \Data_Mem/memory_reg[15][30]  ( .D(\Data_Mem/n5782 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[510]), .Q(data_mem_out_wire[510]) );
  DFF \Data_Mem/memory_reg[15][31]  ( .D(\Data_Mem/n5783 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[511]), .Q(data_mem_out_wire[511]) );
  DFF \Data_Mem/memory_reg[14][0]  ( .D(\Data_Mem/n5784 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[448]), .Q(data_mem_out_wire[448]) );
  DFF \Data_Mem/memory_reg[14][1]  ( .D(\Data_Mem/n5785 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[449]), .Q(data_mem_out_wire[449]) );
  DFF \Data_Mem/memory_reg[14][2]  ( .D(\Data_Mem/n5786 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[450]), .Q(data_mem_out_wire[450]) );
  DFF \Data_Mem/memory_reg[14][3]  ( .D(\Data_Mem/n5787 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[451]), .Q(data_mem_out_wire[451]) );
  DFF \Data_Mem/memory_reg[14][4]  ( .D(\Data_Mem/n5788 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[452]), .Q(data_mem_out_wire[452]) );
  DFF \Data_Mem/memory_reg[14][5]  ( .D(\Data_Mem/n5789 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[453]), .Q(data_mem_out_wire[453]) );
  DFF \Data_Mem/memory_reg[14][6]  ( .D(\Data_Mem/n5790 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[454]), .Q(data_mem_out_wire[454]) );
  DFF \Data_Mem/memory_reg[14][7]  ( .D(\Data_Mem/n5791 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[455]), .Q(data_mem_out_wire[455]) );
  DFF \Data_Mem/memory_reg[14][8]  ( .D(\Data_Mem/n5792 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[456]), .Q(data_mem_out_wire[456]) );
  DFF \Data_Mem/memory_reg[14][9]  ( .D(\Data_Mem/n5793 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[457]), .Q(data_mem_out_wire[457]) );
  DFF \Data_Mem/memory_reg[14][10]  ( .D(\Data_Mem/n5794 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[458]), .Q(data_mem_out_wire[458]) );
  DFF \Data_Mem/memory_reg[14][11]  ( .D(\Data_Mem/n5795 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[459]), .Q(data_mem_out_wire[459]) );
  DFF \Data_Mem/memory_reg[14][12]  ( .D(\Data_Mem/n5796 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[460]), .Q(data_mem_out_wire[460]) );
  DFF \Data_Mem/memory_reg[14][13]  ( .D(\Data_Mem/n5797 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[461]), .Q(data_mem_out_wire[461]) );
  DFF \Data_Mem/memory_reg[14][14]  ( .D(\Data_Mem/n5798 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[462]), .Q(data_mem_out_wire[462]) );
  DFF \Data_Mem/memory_reg[14][15]  ( .D(\Data_Mem/n5799 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[463]), .Q(data_mem_out_wire[463]) );
  DFF \Data_Mem/memory_reg[14][16]  ( .D(\Data_Mem/n5800 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[464]), .Q(data_mem_out_wire[464]) );
  DFF \Data_Mem/memory_reg[14][17]  ( .D(\Data_Mem/n5801 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[465]), .Q(data_mem_out_wire[465]) );
  DFF \Data_Mem/memory_reg[14][18]  ( .D(\Data_Mem/n5802 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[466]), .Q(data_mem_out_wire[466]) );
  DFF \Data_Mem/memory_reg[14][19]  ( .D(\Data_Mem/n5803 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[467]), .Q(data_mem_out_wire[467]) );
  DFF \Data_Mem/memory_reg[14][20]  ( .D(\Data_Mem/n5804 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[468]), .Q(data_mem_out_wire[468]) );
  DFF \Data_Mem/memory_reg[14][21]  ( .D(\Data_Mem/n5805 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[469]), .Q(data_mem_out_wire[469]) );
  DFF \Data_Mem/memory_reg[14][22]  ( .D(\Data_Mem/n5806 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[470]), .Q(data_mem_out_wire[470]) );
  DFF \Data_Mem/memory_reg[14][23]  ( .D(\Data_Mem/n5807 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[471]), .Q(data_mem_out_wire[471]) );
  DFF \Data_Mem/memory_reg[14][24]  ( .D(\Data_Mem/n5808 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[472]), .Q(data_mem_out_wire[472]) );
  DFF \Data_Mem/memory_reg[14][25]  ( .D(\Data_Mem/n5809 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[473]), .Q(data_mem_out_wire[473]) );
  DFF \Data_Mem/memory_reg[14][26]  ( .D(\Data_Mem/n5810 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[474]), .Q(data_mem_out_wire[474]) );
  DFF \Data_Mem/memory_reg[14][27]  ( .D(\Data_Mem/n5811 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[475]), .Q(data_mem_out_wire[475]) );
  DFF \Data_Mem/memory_reg[14][28]  ( .D(\Data_Mem/n5812 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[476]), .Q(data_mem_out_wire[476]) );
  DFF \Data_Mem/memory_reg[14][29]  ( .D(\Data_Mem/n5813 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[477]), .Q(data_mem_out_wire[477]) );
  DFF \Data_Mem/memory_reg[14][30]  ( .D(\Data_Mem/n5814 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[478]), .Q(data_mem_out_wire[478]) );
  DFF \Data_Mem/memory_reg[14][31]  ( .D(\Data_Mem/n5815 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[479]), .Q(data_mem_out_wire[479]) );
  DFF \Data_Mem/memory_reg[13][0]  ( .D(\Data_Mem/n5816 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[416]), .Q(data_mem_out_wire[416]) );
  DFF \Data_Mem/memory_reg[13][1]  ( .D(\Data_Mem/n5817 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[417]), .Q(data_mem_out_wire[417]) );
  DFF \Data_Mem/memory_reg[13][2]  ( .D(\Data_Mem/n5818 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[418]), .Q(data_mem_out_wire[418]) );
  DFF \Data_Mem/memory_reg[13][3]  ( .D(\Data_Mem/n5819 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[419]), .Q(data_mem_out_wire[419]) );
  DFF \Data_Mem/memory_reg[13][4]  ( .D(\Data_Mem/n5820 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[420]), .Q(data_mem_out_wire[420]) );
  DFF \Data_Mem/memory_reg[13][5]  ( .D(\Data_Mem/n5821 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[421]), .Q(data_mem_out_wire[421]) );
  DFF \Data_Mem/memory_reg[13][6]  ( .D(\Data_Mem/n5822 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[422]), .Q(data_mem_out_wire[422]) );
  DFF \Data_Mem/memory_reg[13][7]  ( .D(\Data_Mem/n5823 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[423]), .Q(data_mem_out_wire[423]) );
  DFF \Data_Mem/memory_reg[13][8]  ( .D(\Data_Mem/n5824 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[424]), .Q(data_mem_out_wire[424]) );
  DFF \Data_Mem/memory_reg[13][9]  ( .D(\Data_Mem/n5825 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[425]), .Q(data_mem_out_wire[425]) );
  DFF \Data_Mem/memory_reg[13][10]  ( .D(\Data_Mem/n5826 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[426]), .Q(data_mem_out_wire[426]) );
  DFF \Data_Mem/memory_reg[13][11]  ( .D(\Data_Mem/n5827 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[427]), .Q(data_mem_out_wire[427]) );
  DFF \Data_Mem/memory_reg[13][12]  ( .D(\Data_Mem/n5828 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[428]), .Q(data_mem_out_wire[428]) );
  DFF \Data_Mem/memory_reg[13][13]  ( .D(\Data_Mem/n5829 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[429]), .Q(data_mem_out_wire[429]) );
  DFF \Data_Mem/memory_reg[13][14]  ( .D(\Data_Mem/n5830 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[430]), .Q(data_mem_out_wire[430]) );
  DFF \Data_Mem/memory_reg[13][15]  ( .D(\Data_Mem/n5831 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[431]), .Q(data_mem_out_wire[431]) );
  DFF \Data_Mem/memory_reg[13][16]  ( .D(\Data_Mem/n5832 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[432]), .Q(data_mem_out_wire[432]) );
  DFF \Data_Mem/memory_reg[13][17]  ( .D(\Data_Mem/n5833 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[433]), .Q(data_mem_out_wire[433]) );
  DFF \Data_Mem/memory_reg[13][18]  ( .D(\Data_Mem/n5834 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[434]), .Q(data_mem_out_wire[434]) );
  DFF \Data_Mem/memory_reg[13][19]  ( .D(\Data_Mem/n5835 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[435]), .Q(data_mem_out_wire[435]) );
  DFF \Data_Mem/memory_reg[13][20]  ( .D(\Data_Mem/n5836 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[436]), .Q(data_mem_out_wire[436]) );
  DFF \Data_Mem/memory_reg[13][21]  ( .D(\Data_Mem/n5837 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[437]), .Q(data_mem_out_wire[437]) );
  DFF \Data_Mem/memory_reg[13][22]  ( .D(\Data_Mem/n5838 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[438]), .Q(data_mem_out_wire[438]) );
  DFF \Data_Mem/memory_reg[13][23]  ( .D(\Data_Mem/n5839 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[439]), .Q(data_mem_out_wire[439]) );
  DFF \Data_Mem/memory_reg[13][24]  ( .D(\Data_Mem/n5840 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[440]), .Q(data_mem_out_wire[440]) );
  DFF \Data_Mem/memory_reg[13][25]  ( .D(\Data_Mem/n5841 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[441]), .Q(data_mem_out_wire[441]) );
  DFF \Data_Mem/memory_reg[13][26]  ( .D(\Data_Mem/n5842 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[442]), .Q(data_mem_out_wire[442]) );
  DFF \Data_Mem/memory_reg[13][27]  ( .D(\Data_Mem/n5843 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[443]), .Q(data_mem_out_wire[443]) );
  DFF \Data_Mem/memory_reg[13][28]  ( .D(\Data_Mem/n5844 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[444]), .Q(data_mem_out_wire[444]) );
  DFF \Data_Mem/memory_reg[13][29]  ( .D(\Data_Mem/n5845 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[445]), .Q(data_mem_out_wire[445]) );
  DFF \Data_Mem/memory_reg[13][30]  ( .D(\Data_Mem/n5846 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[446]), .Q(data_mem_out_wire[446]) );
  DFF \Data_Mem/memory_reg[13][31]  ( .D(\Data_Mem/n5847 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[447]), .Q(data_mem_out_wire[447]) );
  DFF \Data_Mem/memory_reg[12][0]  ( .D(\Data_Mem/n5848 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[384]), .Q(data_mem_out_wire[384]) );
  DFF \Data_Mem/memory_reg[12][1]  ( .D(\Data_Mem/n5849 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[385]), .Q(data_mem_out_wire[385]) );
  DFF \Data_Mem/memory_reg[12][2]  ( .D(\Data_Mem/n5850 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[386]), .Q(data_mem_out_wire[386]) );
  DFF \Data_Mem/memory_reg[12][3]  ( .D(\Data_Mem/n5851 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[387]), .Q(data_mem_out_wire[387]) );
  DFF \Data_Mem/memory_reg[12][4]  ( .D(\Data_Mem/n5852 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[388]), .Q(data_mem_out_wire[388]) );
  DFF \Data_Mem/memory_reg[12][5]  ( .D(\Data_Mem/n5853 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[389]), .Q(data_mem_out_wire[389]) );
  DFF \Data_Mem/memory_reg[12][6]  ( .D(\Data_Mem/n5854 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[390]), .Q(data_mem_out_wire[390]) );
  DFF \Data_Mem/memory_reg[12][7]  ( .D(\Data_Mem/n5855 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[391]), .Q(data_mem_out_wire[391]) );
  DFF \Data_Mem/memory_reg[12][8]  ( .D(\Data_Mem/n5856 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[392]), .Q(data_mem_out_wire[392]) );
  DFF \Data_Mem/memory_reg[12][9]  ( .D(\Data_Mem/n5857 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[393]), .Q(data_mem_out_wire[393]) );
  DFF \Data_Mem/memory_reg[12][10]  ( .D(\Data_Mem/n5858 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[394]), .Q(data_mem_out_wire[394]) );
  DFF \Data_Mem/memory_reg[12][11]  ( .D(\Data_Mem/n5859 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[395]), .Q(data_mem_out_wire[395]) );
  DFF \Data_Mem/memory_reg[12][12]  ( .D(\Data_Mem/n5860 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[396]), .Q(data_mem_out_wire[396]) );
  DFF \Data_Mem/memory_reg[12][13]  ( .D(\Data_Mem/n5861 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[397]), .Q(data_mem_out_wire[397]) );
  DFF \Data_Mem/memory_reg[12][14]  ( .D(\Data_Mem/n5862 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[398]), .Q(data_mem_out_wire[398]) );
  DFF \Data_Mem/memory_reg[12][15]  ( .D(\Data_Mem/n5863 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[399]), .Q(data_mem_out_wire[399]) );
  DFF \Data_Mem/memory_reg[12][16]  ( .D(\Data_Mem/n5864 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[400]), .Q(data_mem_out_wire[400]) );
  DFF \Data_Mem/memory_reg[12][17]  ( .D(\Data_Mem/n5865 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[401]), .Q(data_mem_out_wire[401]) );
  DFF \Data_Mem/memory_reg[12][18]  ( .D(\Data_Mem/n5866 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[402]), .Q(data_mem_out_wire[402]) );
  DFF \Data_Mem/memory_reg[12][19]  ( .D(\Data_Mem/n5867 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[403]), .Q(data_mem_out_wire[403]) );
  DFF \Data_Mem/memory_reg[12][20]  ( .D(\Data_Mem/n5868 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[404]), .Q(data_mem_out_wire[404]) );
  DFF \Data_Mem/memory_reg[12][21]  ( .D(\Data_Mem/n5869 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[405]), .Q(data_mem_out_wire[405]) );
  DFF \Data_Mem/memory_reg[12][22]  ( .D(\Data_Mem/n5870 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[406]), .Q(data_mem_out_wire[406]) );
  DFF \Data_Mem/memory_reg[12][23]  ( .D(\Data_Mem/n5871 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[407]), .Q(data_mem_out_wire[407]) );
  DFF \Data_Mem/memory_reg[12][24]  ( .D(\Data_Mem/n5872 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[408]), .Q(data_mem_out_wire[408]) );
  DFF \Data_Mem/memory_reg[12][25]  ( .D(\Data_Mem/n5873 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[409]), .Q(data_mem_out_wire[409]) );
  DFF \Data_Mem/memory_reg[12][26]  ( .D(\Data_Mem/n5874 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[410]), .Q(data_mem_out_wire[410]) );
  DFF \Data_Mem/memory_reg[12][27]  ( .D(\Data_Mem/n5875 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[411]), .Q(data_mem_out_wire[411]) );
  DFF \Data_Mem/memory_reg[12][28]  ( .D(\Data_Mem/n5876 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[412]), .Q(data_mem_out_wire[412]) );
  DFF \Data_Mem/memory_reg[12][29]  ( .D(\Data_Mem/n5877 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[413]), .Q(data_mem_out_wire[413]) );
  DFF \Data_Mem/memory_reg[12][30]  ( .D(\Data_Mem/n5878 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[414]), .Q(data_mem_out_wire[414]) );
  DFF \Data_Mem/memory_reg[12][31]  ( .D(\Data_Mem/n5879 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[415]), .Q(data_mem_out_wire[415]) );
  DFF \Data_Mem/memory_reg[11][0]  ( .D(\Data_Mem/n5880 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[352]), .Q(data_mem_out_wire[352]) );
  DFF \Data_Mem/memory_reg[11][1]  ( .D(\Data_Mem/n5881 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[353]), .Q(data_mem_out_wire[353]) );
  DFF \Data_Mem/memory_reg[11][2]  ( .D(\Data_Mem/n5882 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[354]), .Q(data_mem_out_wire[354]) );
  DFF \Data_Mem/memory_reg[11][3]  ( .D(\Data_Mem/n5883 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[355]), .Q(data_mem_out_wire[355]) );
  DFF \Data_Mem/memory_reg[11][4]  ( .D(\Data_Mem/n5884 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[356]), .Q(data_mem_out_wire[356]) );
  DFF \Data_Mem/memory_reg[11][5]  ( .D(\Data_Mem/n5885 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[357]), .Q(data_mem_out_wire[357]) );
  DFF \Data_Mem/memory_reg[11][6]  ( .D(\Data_Mem/n5886 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[358]), .Q(data_mem_out_wire[358]) );
  DFF \Data_Mem/memory_reg[11][7]  ( .D(\Data_Mem/n5887 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[359]), .Q(data_mem_out_wire[359]) );
  DFF \Data_Mem/memory_reg[11][8]  ( .D(\Data_Mem/n5888 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[360]), .Q(data_mem_out_wire[360]) );
  DFF \Data_Mem/memory_reg[11][9]  ( .D(\Data_Mem/n5889 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[361]), .Q(data_mem_out_wire[361]) );
  DFF \Data_Mem/memory_reg[11][10]  ( .D(\Data_Mem/n5890 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[362]), .Q(data_mem_out_wire[362]) );
  DFF \Data_Mem/memory_reg[11][11]  ( .D(\Data_Mem/n5891 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[363]), .Q(data_mem_out_wire[363]) );
  DFF \Data_Mem/memory_reg[11][12]  ( .D(\Data_Mem/n5892 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[364]), .Q(data_mem_out_wire[364]) );
  DFF \Data_Mem/memory_reg[11][13]  ( .D(\Data_Mem/n5893 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[365]), .Q(data_mem_out_wire[365]) );
  DFF \Data_Mem/memory_reg[11][14]  ( .D(\Data_Mem/n5894 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[366]), .Q(data_mem_out_wire[366]) );
  DFF \Data_Mem/memory_reg[11][15]  ( .D(\Data_Mem/n5895 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[367]), .Q(data_mem_out_wire[367]) );
  DFF \Data_Mem/memory_reg[11][16]  ( .D(\Data_Mem/n5896 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[368]), .Q(data_mem_out_wire[368]) );
  DFF \Data_Mem/memory_reg[11][17]  ( .D(\Data_Mem/n5897 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[369]), .Q(data_mem_out_wire[369]) );
  DFF \Data_Mem/memory_reg[11][18]  ( .D(\Data_Mem/n5898 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[370]), .Q(data_mem_out_wire[370]) );
  DFF \Data_Mem/memory_reg[11][19]  ( .D(\Data_Mem/n5899 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[371]), .Q(data_mem_out_wire[371]) );
  DFF \Data_Mem/memory_reg[11][20]  ( .D(\Data_Mem/n5900 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[372]), .Q(data_mem_out_wire[372]) );
  DFF \Data_Mem/memory_reg[11][21]  ( .D(\Data_Mem/n5901 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[373]), .Q(data_mem_out_wire[373]) );
  DFF \Data_Mem/memory_reg[11][22]  ( .D(\Data_Mem/n5902 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[374]), .Q(data_mem_out_wire[374]) );
  DFF \Data_Mem/memory_reg[11][23]  ( .D(\Data_Mem/n5903 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[375]), .Q(data_mem_out_wire[375]) );
  DFF \Data_Mem/memory_reg[11][24]  ( .D(\Data_Mem/n5904 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[376]), .Q(data_mem_out_wire[376]) );
  DFF \Data_Mem/memory_reg[11][25]  ( .D(\Data_Mem/n5905 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[377]), .Q(data_mem_out_wire[377]) );
  DFF \Data_Mem/memory_reg[11][26]  ( .D(\Data_Mem/n5906 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[378]), .Q(data_mem_out_wire[378]) );
  DFF \Data_Mem/memory_reg[11][27]  ( .D(\Data_Mem/n5907 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[379]), .Q(data_mem_out_wire[379]) );
  DFF \Data_Mem/memory_reg[11][28]  ( .D(\Data_Mem/n5908 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[380]), .Q(data_mem_out_wire[380]) );
  DFF \Data_Mem/memory_reg[11][29]  ( .D(\Data_Mem/n5909 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[381]), .Q(data_mem_out_wire[381]) );
  DFF \Data_Mem/memory_reg[11][30]  ( .D(\Data_Mem/n5910 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[382]), .Q(data_mem_out_wire[382]) );
  DFF \Data_Mem/memory_reg[11][31]  ( .D(\Data_Mem/n5911 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[383]), .Q(data_mem_out_wire[383]) );
  DFF \Data_Mem/memory_reg[10][0]  ( .D(\Data_Mem/n5912 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[320]), .Q(data_mem_out_wire[320]) );
  DFF \Data_Mem/memory_reg[10][1]  ( .D(\Data_Mem/n5913 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[321]), .Q(data_mem_out_wire[321]) );
  DFF \Data_Mem/memory_reg[10][2]  ( .D(\Data_Mem/n5914 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[322]), .Q(data_mem_out_wire[322]) );
  DFF \Data_Mem/memory_reg[10][3]  ( .D(\Data_Mem/n5915 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[323]), .Q(data_mem_out_wire[323]) );
  DFF \Data_Mem/memory_reg[10][4]  ( .D(\Data_Mem/n5916 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[324]), .Q(data_mem_out_wire[324]) );
  DFF \Data_Mem/memory_reg[10][5]  ( .D(\Data_Mem/n5917 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[325]), .Q(data_mem_out_wire[325]) );
  DFF \Data_Mem/memory_reg[10][6]  ( .D(\Data_Mem/n5918 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[326]), .Q(data_mem_out_wire[326]) );
  DFF \Data_Mem/memory_reg[10][7]  ( .D(\Data_Mem/n5919 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[327]), .Q(data_mem_out_wire[327]) );
  DFF \Data_Mem/memory_reg[10][8]  ( .D(\Data_Mem/n5920 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[328]), .Q(data_mem_out_wire[328]) );
  DFF \Data_Mem/memory_reg[10][9]  ( .D(\Data_Mem/n5921 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[329]), .Q(data_mem_out_wire[329]) );
  DFF \Data_Mem/memory_reg[10][10]  ( .D(\Data_Mem/n5922 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[330]), .Q(data_mem_out_wire[330]) );
  DFF \Data_Mem/memory_reg[10][11]  ( .D(\Data_Mem/n5923 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[331]), .Q(data_mem_out_wire[331]) );
  DFF \Data_Mem/memory_reg[10][12]  ( .D(\Data_Mem/n5924 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[332]), .Q(data_mem_out_wire[332]) );
  DFF \Data_Mem/memory_reg[10][13]  ( .D(\Data_Mem/n5925 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[333]), .Q(data_mem_out_wire[333]) );
  DFF \Data_Mem/memory_reg[10][14]  ( .D(\Data_Mem/n5926 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[334]), .Q(data_mem_out_wire[334]) );
  DFF \Data_Mem/memory_reg[10][15]  ( .D(\Data_Mem/n5927 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[335]), .Q(data_mem_out_wire[335]) );
  DFF \Data_Mem/memory_reg[10][16]  ( .D(\Data_Mem/n5928 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[336]), .Q(data_mem_out_wire[336]) );
  DFF \Data_Mem/memory_reg[10][17]  ( .D(\Data_Mem/n5929 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[337]), .Q(data_mem_out_wire[337]) );
  DFF \Data_Mem/memory_reg[10][18]  ( .D(\Data_Mem/n5930 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[338]), .Q(data_mem_out_wire[338]) );
  DFF \Data_Mem/memory_reg[10][19]  ( .D(\Data_Mem/n5931 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[339]), .Q(data_mem_out_wire[339]) );
  DFF \Data_Mem/memory_reg[10][20]  ( .D(\Data_Mem/n5932 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[340]), .Q(data_mem_out_wire[340]) );
  DFF \Data_Mem/memory_reg[10][21]  ( .D(\Data_Mem/n5933 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[341]), .Q(data_mem_out_wire[341]) );
  DFF \Data_Mem/memory_reg[10][22]  ( .D(\Data_Mem/n5934 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[342]), .Q(data_mem_out_wire[342]) );
  DFF \Data_Mem/memory_reg[10][23]  ( .D(\Data_Mem/n5935 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[343]), .Q(data_mem_out_wire[343]) );
  DFF \Data_Mem/memory_reg[10][24]  ( .D(\Data_Mem/n5936 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[344]), .Q(data_mem_out_wire[344]) );
  DFF \Data_Mem/memory_reg[10][25]  ( .D(\Data_Mem/n5937 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[345]), .Q(data_mem_out_wire[345]) );
  DFF \Data_Mem/memory_reg[10][26]  ( .D(\Data_Mem/n5938 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[346]), .Q(data_mem_out_wire[346]) );
  DFF \Data_Mem/memory_reg[10][27]  ( .D(\Data_Mem/n5939 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[347]), .Q(data_mem_out_wire[347]) );
  DFF \Data_Mem/memory_reg[10][28]  ( .D(\Data_Mem/n5940 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[348]), .Q(data_mem_out_wire[348]) );
  DFF \Data_Mem/memory_reg[10][29]  ( .D(\Data_Mem/n5941 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[349]), .Q(data_mem_out_wire[349]) );
  DFF \Data_Mem/memory_reg[10][30]  ( .D(\Data_Mem/n5942 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[350]), .Q(data_mem_out_wire[350]) );
  DFF \Data_Mem/memory_reg[10][31]  ( .D(\Data_Mem/n5943 ), .CLK(clk), .RST(
        rst), .I(data_mem_in_wire[351]), .Q(data_mem_out_wire[351]) );
  DFF \Data_Mem/memory_reg[9][0]  ( .D(\Data_Mem/n5944 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[288]), .Q(data_mem_out_wire[288]) );
  DFF \Data_Mem/memory_reg[9][1]  ( .D(\Data_Mem/n5945 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[289]), .Q(data_mem_out_wire[289]) );
  DFF \Data_Mem/memory_reg[9][2]  ( .D(\Data_Mem/n5946 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[290]), .Q(data_mem_out_wire[290]) );
  DFF \Data_Mem/memory_reg[9][3]  ( .D(\Data_Mem/n5947 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[291]), .Q(data_mem_out_wire[291]) );
  DFF \Data_Mem/memory_reg[9][4]  ( .D(\Data_Mem/n5948 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[292]), .Q(data_mem_out_wire[292]) );
  DFF \Data_Mem/memory_reg[9][5]  ( .D(\Data_Mem/n5949 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[293]), .Q(data_mem_out_wire[293]) );
  DFF \Data_Mem/memory_reg[9][6]  ( .D(\Data_Mem/n5950 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[294]), .Q(data_mem_out_wire[294]) );
  DFF \Data_Mem/memory_reg[9][7]  ( .D(\Data_Mem/n5951 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[295]), .Q(data_mem_out_wire[295]) );
  DFF \Data_Mem/memory_reg[9][8]  ( .D(\Data_Mem/n5952 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[296]), .Q(data_mem_out_wire[296]) );
  DFF \Data_Mem/memory_reg[9][9]  ( .D(\Data_Mem/n5953 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[297]), .Q(data_mem_out_wire[297]) );
  DFF \Data_Mem/memory_reg[9][10]  ( .D(\Data_Mem/n5954 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[298]), .Q(data_mem_out_wire[298]) );
  DFF \Data_Mem/memory_reg[9][11]  ( .D(\Data_Mem/n5955 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[299]), .Q(data_mem_out_wire[299]) );
  DFF \Data_Mem/memory_reg[9][12]  ( .D(\Data_Mem/n5956 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[300]), .Q(data_mem_out_wire[300]) );
  DFF \Data_Mem/memory_reg[9][13]  ( .D(\Data_Mem/n5957 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[301]), .Q(data_mem_out_wire[301]) );
  DFF \Data_Mem/memory_reg[9][14]  ( .D(\Data_Mem/n5958 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[302]), .Q(data_mem_out_wire[302]) );
  DFF \Data_Mem/memory_reg[9][15]  ( .D(\Data_Mem/n5959 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[303]), .Q(data_mem_out_wire[303]) );
  DFF \Data_Mem/memory_reg[9][16]  ( .D(\Data_Mem/n5960 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[304]), .Q(data_mem_out_wire[304]) );
  DFF \Data_Mem/memory_reg[9][17]  ( .D(\Data_Mem/n5961 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[305]), .Q(data_mem_out_wire[305]) );
  DFF \Data_Mem/memory_reg[9][18]  ( .D(\Data_Mem/n5962 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[306]), .Q(data_mem_out_wire[306]) );
  DFF \Data_Mem/memory_reg[9][19]  ( .D(\Data_Mem/n5963 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[307]), .Q(data_mem_out_wire[307]) );
  DFF \Data_Mem/memory_reg[9][20]  ( .D(\Data_Mem/n5964 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[308]), .Q(data_mem_out_wire[308]) );
  DFF \Data_Mem/memory_reg[9][21]  ( .D(\Data_Mem/n5965 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[309]), .Q(data_mem_out_wire[309]) );
  DFF \Data_Mem/memory_reg[9][22]  ( .D(\Data_Mem/n5966 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[310]), .Q(data_mem_out_wire[310]) );
  DFF \Data_Mem/memory_reg[9][23]  ( .D(\Data_Mem/n5967 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[311]), .Q(data_mem_out_wire[311]) );
  DFF \Data_Mem/memory_reg[9][24]  ( .D(\Data_Mem/n5968 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[312]), .Q(data_mem_out_wire[312]) );
  DFF \Data_Mem/memory_reg[9][25]  ( .D(\Data_Mem/n5969 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[313]), .Q(data_mem_out_wire[313]) );
  DFF \Data_Mem/memory_reg[9][26]  ( .D(\Data_Mem/n5970 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[314]), .Q(data_mem_out_wire[314]) );
  DFF \Data_Mem/memory_reg[9][27]  ( .D(\Data_Mem/n5971 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[315]), .Q(data_mem_out_wire[315]) );
  DFF \Data_Mem/memory_reg[9][28]  ( .D(\Data_Mem/n5972 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[316]), .Q(data_mem_out_wire[316]) );
  DFF \Data_Mem/memory_reg[9][29]  ( .D(\Data_Mem/n5973 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[317]), .Q(data_mem_out_wire[317]) );
  DFF \Data_Mem/memory_reg[9][30]  ( .D(\Data_Mem/n5974 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[318]), .Q(data_mem_out_wire[318]) );
  DFF \Data_Mem/memory_reg[9][31]  ( .D(\Data_Mem/n5975 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[319]), .Q(data_mem_out_wire[319]) );
  DFF \Data_Mem/memory_reg[8][0]  ( .D(\Data_Mem/n5976 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[256]), .Q(data_mem_out_wire[256]) );
  DFF \Data_Mem/memory_reg[8][1]  ( .D(\Data_Mem/n5977 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[257]), .Q(data_mem_out_wire[257]) );
  DFF \Data_Mem/memory_reg[8][2]  ( .D(\Data_Mem/n5978 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[258]), .Q(data_mem_out_wire[258]) );
  DFF \Data_Mem/memory_reg[8][3]  ( .D(\Data_Mem/n5979 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[259]), .Q(data_mem_out_wire[259]) );
  DFF \Data_Mem/memory_reg[8][4]  ( .D(\Data_Mem/n5980 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[260]), .Q(data_mem_out_wire[260]) );
  DFF \Data_Mem/memory_reg[8][5]  ( .D(\Data_Mem/n5981 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[261]), .Q(data_mem_out_wire[261]) );
  DFF \Data_Mem/memory_reg[8][6]  ( .D(\Data_Mem/n5982 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[262]), .Q(data_mem_out_wire[262]) );
  DFF \Data_Mem/memory_reg[8][7]  ( .D(\Data_Mem/n5983 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[263]), .Q(data_mem_out_wire[263]) );
  DFF \Data_Mem/memory_reg[8][8]  ( .D(\Data_Mem/n5984 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[264]), .Q(data_mem_out_wire[264]) );
  DFF \Data_Mem/memory_reg[8][9]  ( .D(\Data_Mem/n5985 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[265]), .Q(data_mem_out_wire[265]) );
  DFF \Data_Mem/memory_reg[8][10]  ( .D(\Data_Mem/n5986 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[266]), .Q(data_mem_out_wire[266]) );
  DFF \Data_Mem/memory_reg[8][11]  ( .D(\Data_Mem/n5987 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[267]), .Q(data_mem_out_wire[267]) );
  DFF \Data_Mem/memory_reg[8][12]  ( .D(\Data_Mem/n5988 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[268]), .Q(data_mem_out_wire[268]) );
  DFF \Data_Mem/memory_reg[8][13]  ( .D(\Data_Mem/n5989 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[269]), .Q(data_mem_out_wire[269]) );
  DFF \Data_Mem/memory_reg[8][14]  ( .D(\Data_Mem/n5990 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[270]), .Q(data_mem_out_wire[270]) );
  DFF \Data_Mem/memory_reg[8][15]  ( .D(\Data_Mem/n5991 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[271]), .Q(data_mem_out_wire[271]) );
  DFF \Data_Mem/memory_reg[8][16]  ( .D(\Data_Mem/n5992 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[272]), .Q(data_mem_out_wire[272]) );
  DFF \Data_Mem/memory_reg[8][17]  ( .D(\Data_Mem/n5993 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[273]), .Q(data_mem_out_wire[273]) );
  DFF \Data_Mem/memory_reg[8][18]  ( .D(\Data_Mem/n5994 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[274]), .Q(data_mem_out_wire[274]) );
  DFF \Data_Mem/memory_reg[8][19]  ( .D(\Data_Mem/n5995 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[275]), .Q(data_mem_out_wire[275]) );
  DFF \Data_Mem/memory_reg[8][20]  ( .D(\Data_Mem/n5996 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[276]), .Q(data_mem_out_wire[276]) );
  DFF \Data_Mem/memory_reg[8][21]  ( .D(\Data_Mem/n5997 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[277]), .Q(data_mem_out_wire[277]) );
  DFF \Data_Mem/memory_reg[8][22]  ( .D(\Data_Mem/n5998 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[278]), .Q(data_mem_out_wire[278]) );
  DFF \Data_Mem/memory_reg[8][23]  ( .D(\Data_Mem/n5999 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[279]), .Q(data_mem_out_wire[279]) );
  DFF \Data_Mem/memory_reg[8][24]  ( .D(\Data_Mem/n6000 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[280]), .Q(data_mem_out_wire[280]) );
  DFF \Data_Mem/memory_reg[8][25]  ( .D(\Data_Mem/n6001 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[281]), .Q(data_mem_out_wire[281]) );
  DFF \Data_Mem/memory_reg[8][26]  ( .D(\Data_Mem/n6002 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[282]), .Q(data_mem_out_wire[282]) );
  DFF \Data_Mem/memory_reg[8][27]  ( .D(\Data_Mem/n6003 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[283]), .Q(data_mem_out_wire[283]) );
  DFF \Data_Mem/memory_reg[8][28]  ( .D(\Data_Mem/n6004 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[284]), .Q(data_mem_out_wire[284]) );
  DFF \Data_Mem/memory_reg[8][29]  ( .D(\Data_Mem/n6005 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[285]), .Q(data_mem_out_wire[285]) );
  DFF \Data_Mem/memory_reg[8][30]  ( .D(\Data_Mem/n6006 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[286]), .Q(data_mem_out_wire[286]) );
  DFF \Data_Mem/memory_reg[8][31]  ( .D(\Data_Mem/n6007 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[287]), .Q(data_mem_out_wire[287]) );
  DFF \Data_Mem/memory_reg[7][0]  ( .D(\Data_Mem/n6008 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[224]), .Q(data_mem_out_wire[224]) );
  DFF \Data_Mem/memory_reg[7][1]  ( .D(\Data_Mem/n6009 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[225]), .Q(data_mem_out_wire[225]) );
  DFF \Data_Mem/memory_reg[7][2]  ( .D(\Data_Mem/n6010 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[226]), .Q(data_mem_out_wire[226]) );
  DFF \Data_Mem/memory_reg[7][3]  ( .D(\Data_Mem/n6011 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[227]), .Q(data_mem_out_wire[227]) );
  DFF \Data_Mem/memory_reg[7][4]  ( .D(\Data_Mem/n6012 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[228]), .Q(data_mem_out_wire[228]) );
  DFF \Data_Mem/memory_reg[7][5]  ( .D(\Data_Mem/n6013 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[229]), .Q(data_mem_out_wire[229]) );
  DFF \Data_Mem/memory_reg[7][6]  ( .D(\Data_Mem/n6014 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[230]), .Q(data_mem_out_wire[230]) );
  DFF \Data_Mem/memory_reg[7][7]  ( .D(\Data_Mem/n6015 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[231]), .Q(data_mem_out_wire[231]) );
  DFF \Data_Mem/memory_reg[7][8]  ( .D(\Data_Mem/n6016 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[232]), .Q(data_mem_out_wire[232]) );
  DFF \Data_Mem/memory_reg[7][9]  ( .D(\Data_Mem/n6017 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[233]), .Q(data_mem_out_wire[233]) );
  DFF \Data_Mem/memory_reg[7][10]  ( .D(\Data_Mem/n6018 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[234]), .Q(data_mem_out_wire[234]) );
  DFF \Data_Mem/memory_reg[7][11]  ( .D(\Data_Mem/n6019 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[235]), .Q(data_mem_out_wire[235]) );
  DFF \Data_Mem/memory_reg[7][12]  ( .D(\Data_Mem/n6020 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[236]), .Q(data_mem_out_wire[236]) );
  DFF \Data_Mem/memory_reg[7][13]  ( .D(\Data_Mem/n6021 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[237]), .Q(data_mem_out_wire[237]) );
  DFF \Data_Mem/memory_reg[7][14]  ( .D(\Data_Mem/n6022 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[238]), .Q(data_mem_out_wire[238]) );
  DFF \Data_Mem/memory_reg[7][15]  ( .D(\Data_Mem/n6023 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[239]), .Q(data_mem_out_wire[239]) );
  DFF \Data_Mem/memory_reg[7][16]  ( .D(\Data_Mem/n6024 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[240]), .Q(data_mem_out_wire[240]) );
  DFF \Data_Mem/memory_reg[7][17]  ( .D(\Data_Mem/n6025 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[241]), .Q(data_mem_out_wire[241]) );
  DFF \Data_Mem/memory_reg[7][18]  ( .D(\Data_Mem/n6026 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[242]), .Q(data_mem_out_wire[242]) );
  DFF \Data_Mem/memory_reg[7][19]  ( .D(\Data_Mem/n6027 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[243]), .Q(data_mem_out_wire[243]) );
  DFF \Data_Mem/memory_reg[7][20]  ( .D(\Data_Mem/n6028 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[244]), .Q(data_mem_out_wire[244]) );
  DFF \Data_Mem/memory_reg[7][21]  ( .D(\Data_Mem/n6029 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[245]), .Q(data_mem_out_wire[245]) );
  DFF \Data_Mem/memory_reg[7][22]  ( .D(\Data_Mem/n6030 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[246]), .Q(data_mem_out_wire[246]) );
  DFF \Data_Mem/memory_reg[7][23]  ( .D(\Data_Mem/n6031 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[247]), .Q(data_mem_out_wire[247]) );
  DFF \Data_Mem/memory_reg[7][24]  ( .D(\Data_Mem/n6032 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[248]), .Q(data_mem_out_wire[248]) );
  DFF \Data_Mem/memory_reg[7][25]  ( .D(\Data_Mem/n6033 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[249]), .Q(data_mem_out_wire[249]) );
  DFF \Data_Mem/memory_reg[7][26]  ( .D(\Data_Mem/n6034 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[250]), .Q(data_mem_out_wire[250]) );
  DFF \Data_Mem/memory_reg[7][27]  ( .D(\Data_Mem/n6035 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[251]), .Q(data_mem_out_wire[251]) );
  DFF \Data_Mem/memory_reg[7][28]  ( .D(\Data_Mem/n6036 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[252]), .Q(data_mem_out_wire[252]) );
  DFF \Data_Mem/memory_reg[7][29]  ( .D(\Data_Mem/n6037 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[253]), .Q(data_mem_out_wire[253]) );
  DFF \Data_Mem/memory_reg[7][30]  ( .D(\Data_Mem/n6038 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[254]), .Q(data_mem_out_wire[254]) );
  DFF \Data_Mem/memory_reg[7][31]  ( .D(\Data_Mem/n6039 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[255]), .Q(data_mem_out_wire[255]) );
  DFF \Data_Mem/memory_reg[6][0]  ( .D(\Data_Mem/n6040 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[192]), .Q(data_mem_out_wire[192]) );
  DFF \Data_Mem/memory_reg[6][1]  ( .D(\Data_Mem/n6041 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[193]), .Q(data_mem_out_wire[193]) );
  DFF \Data_Mem/memory_reg[6][2]  ( .D(\Data_Mem/n6042 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[194]), .Q(data_mem_out_wire[194]) );
  DFF \Data_Mem/memory_reg[6][3]  ( .D(\Data_Mem/n6043 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[195]), .Q(data_mem_out_wire[195]) );
  DFF \Data_Mem/memory_reg[6][4]  ( .D(\Data_Mem/n6044 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[196]), .Q(data_mem_out_wire[196]) );
  DFF \Data_Mem/memory_reg[6][5]  ( .D(\Data_Mem/n6045 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[197]), .Q(data_mem_out_wire[197]) );
  DFF \Data_Mem/memory_reg[6][6]  ( .D(\Data_Mem/n6046 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[198]), .Q(data_mem_out_wire[198]) );
  DFF \Data_Mem/memory_reg[6][7]  ( .D(\Data_Mem/n6047 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[199]), .Q(data_mem_out_wire[199]) );
  DFF \Data_Mem/memory_reg[6][8]  ( .D(\Data_Mem/n6048 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[200]), .Q(data_mem_out_wire[200]) );
  DFF \Data_Mem/memory_reg[6][9]  ( .D(\Data_Mem/n6049 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[201]), .Q(data_mem_out_wire[201]) );
  DFF \Data_Mem/memory_reg[6][10]  ( .D(\Data_Mem/n6050 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[202]), .Q(data_mem_out_wire[202]) );
  DFF \Data_Mem/memory_reg[6][11]  ( .D(\Data_Mem/n6051 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[203]), .Q(data_mem_out_wire[203]) );
  DFF \Data_Mem/memory_reg[6][12]  ( .D(\Data_Mem/n6052 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[204]), .Q(data_mem_out_wire[204]) );
  DFF \Data_Mem/memory_reg[6][13]  ( .D(\Data_Mem/n6053 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[205]), .Q(data_mem_out_wire[205]) );
  DFF \Data_Mem/memory_reg[6][14]  ( .D(\Data_Mem/n6054 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[206]), .Q(data_mem_out_wire[206]) );
  DFF \Data_Mem/memory_reg[6][15]  ( .D(\Data_Mem/n6055 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[207]), .Q(data_mem_out_wire[207]) );
  DFF \Data_Mem/memory_reg[6][16]  ( .D(\Data_Mem/n6056 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[208]), .Q(data_mem_out_wire[208]) );
  DFF \Data_Mem/memory_reg[6][17]  ( .D(\Data_Mem/n6057 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[209]), .Q(data_mem_out_wire[209]) );
  DFF \Data_Mem/memory_reg[6][18]  ( .D(\Data_Mem/n6058 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[210]), .Q(data_mem_out_wire[210]) );
  DFF \Data_Mem/memory_reg[6][19]  ( .D(\Data_Mem/n6059 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[211]), .Q(data_mem_out_wire[211]) );
  DFF \Data_Mem/memory_reg[6][20]  ( .D(\Data_Mem/n6060 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[212]), .Q(data_mem_out_wire[212]) );
  DFF \Data_Mem/memory_reg[6][21]  ( .D(\Data_Mem/n6061 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[213]), .Q(data_mem_out_wire[213]) );
  DFF \Data_Mem/memory_reg[6][22]  ( .D(\Data_Mem/n6062 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[214]), .Q(data_mem_out_wire[214]) );
  DFF \Data_Mem/memory_reg[6][23]  ( .D(\Data_Mem/n6063 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[215]), .Q(data_mem_out_wire[215]) );
  DFF \Data_Mem/memory_reg[6][24]  ( .D(\Data_Mem/n6064 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[216]), .Q(data_mem_out_wire[216]) );
  DFF \Data_Mem/memory_reg[6][25]  ( .D(\Data_Mem/n6065 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[217]), .Q(data_mem_out_wire[217]) );
  DFF \Data_Mem/memory_reg[6][26]  ( .D(\Data_Mem/n6066 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[218]), .Q(data_mem_out_wire[218]) );
  DFF \Data_Mem/memory_reg[6][27]  ( .D(\Data_Mem/n6067 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[219]), .Q(data_mem_out_wire[219]) );
  DFF \Data_Mem/memory_reg[6][28]  ( .D(\Data_Mem/n6068 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[220]), .Q(data_mem_out_wire[220]) );
  DFF \Data_Mem/memory_reg[6][29]  ( .D(\Data_Mem/n6069 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[221]), .Q(data_mem_out_wire[221]) );
  DFF \Data_Mem/memory_reg[6][30]  ( .D(\Data_Mem/n6070 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[222]), .Q(data_mem_out_wire[222]) );
  DFF \Data_Mem/memory_reg[6][31]  ( .D(\Data_Mem/n6071 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[223]), .Q(data_mem_out_wire[223]) );
  DFF \Data_Mem/memory_reg[5][0]  ( .D(\Data_Mem/n6072 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[160]), .Q(data_mem_out_wire[160]) );
  DFF \Data_Mem/memory_reg[5][1]  ( .D(\Data_Mem/n6073 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[161]), .Q(data_mem_out_wire[161]) );
  DFF \Data_Mem/memory_reg[5][2]  ( .D(\Data_Mem/n6074 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[162]), .Q(data_mem_out_wire[162]) );
  DFF \Data_Mem/memory_reg[5][3]  ( .D(\Data_Mem/n6075 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[163]), .Q(data_mem_out_wire[163]) );
  DFF \Data_Mem/memory_reg[5][4]  ( .D(\Data_Mem/n6076 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[164]), .Q(data_mem_out_wire[164]) );
  DFF \Data_Mem/memory_reg[5][5]  ( .D(\Data_Mem/n6077 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[165]), .Q(data_mem_out_wire[165]) );
  DFF \Data_Mem/memory_reg[5][6]  ( .D(\Data_Mem/n6078 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[166]), .Q(data_mem_out_wire[166]) );
  DFF \Data_Mem/memory_reg[5][7]  ( .D(\Data_Mem/n6079 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[167]), .Q(data_mem_out_wire[167]) );
  DFF \Data_Mem/memory_reg[5][8]  ( .D(\Data_Mem/n6080 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[168]), .Q(data_mem_out_wire[168]) );
  DFF \Data_Mem/memory_reg[5][9]  ( .D(\Data_Mem/n6081 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[169]), .Q(data_mem_out_wire[169]) );
  DFF \Data_Mem/memory_reg[5][10]  ( .D(\Data_Mem/n6082 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[170]), .Q(data_mem_out_wire[170]) );
  DFF \Data_Mem/memory_reg[5][11]  ( .D(\Data_Mem/n6083 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[171]), .Q(data_mem_out_wire[171]) );
  DFF \Data_Mem/memory_reg[5][12]  ( .D(\Data_Mem/n6084 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[172]), .Q(data_mem_out_wire[172]) );
  DFF \Data_Mem/memory_reg[5][13]  ( .D(\Data_Mem/n6085 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[173]), .Q(data_mem_out_wire[173]) );
  DFF \Data_Mem/memory_reg[5][14]  ( .D(\Data_Mem/n6086 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[174]), .Q(data_mem_out_wire[174]) );
  DFF \Data_Mem/memory_reg[5][15]  ( .D(\Data_Mem/n6087 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[175]), .Q(data_mem_out_wire[175]) );
  DFF \Data_Mem/memory_reg[5][16]  ( .D(\Data_Mem/n6088 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[176]), .Q(data_mem_out_wire[176]) );
  DFF \Data_Mem/memory_reg[5][17]  ( .D(\Data_Mem/n6089 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[177]), .Q(data_mem_out_wire[177]) );
  DFF \Data_Mem/memory_reg[5][18]  ( .D(\Data_Mem/n6090 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[178]), .Q(data_mem_out_wire[178]) );
  DFF \Data_Mem/memory_reg[5][19]  ( .D(\Data_Mem/n6091 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[179]), .Q(data_mem_out_wire[179]) );
  DFF \Data_Mem/memory_reg[5][20]  ( .D(\Data_Mem/n6092 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[180]), .Q(data_mem_out_wire[180]) );
  DFF \Data_Mem/memory_reg[5][21]  ( .D(\Data_Mem/n6093 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[181]), .Q(data_mem_out_wire[181]) );
  DFF \Data_Mem/memory_reg[5][22]  ( .D(\Data_Mem/n6094 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[182]), .Q(data_mem_out_wire[182]) );
  DFF \Data_Mem/memory_reg[5][23]  ( .D(\Data_Mem/n6095 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[183]), .Q(data_mem_out_wire[183]) );
  DFF \Data_Mem/memory_reg[5][24]  ( .D(\Data_Mem/n6096 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[184]), .Q(data_mem_out_wire[184]) );
  DFF \Data_Mem/memory_reg[5][25]  ( .D(\Data_Mem/n6097 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[185]), .Q(data_mem_out_wire[185]) );
  DFF \Data_Mem/memory_reg[5][26]  ( .D(\Data_Mem/n6098 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[186]), .Q(data_mem_out_wire[186]) );
  DFF \Data_Mem/memory_reg[5][27]  ( .D(\Data_Mem/n6099 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[187]), .Q(data_mem_out_wire[187]) );
  DFF \Data_Mem/memory_reg[5][28]  ( .D(\Data_Mem/n6100 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[188]), .Q(data_mem_out_wire[188]) );
  DFF \Data_Mem/memory_reg[5][29]  ( .D(\Data_Mem/n6101 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[189]), .Q(data_mem_out_wire[189]) );
  DFF \Data_Mem/memory_reg[5][30]  ( .D(\Data_Mem/n6102 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[190]), .Q(data_mem_out_wire[190]) );
  DFF \Data_Mem/memory_reg[5][31]  ( .D(\Data_Mem/n6103 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[191]), .Q(data_mem_out_wire[191]) );
  DFF \Data_Mem/memory_reg[4][0]  ( .D(\Data_Mem/n6104 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[128]), .Q(data_mem_out_wire[128]) );
  DFF \Data_Mem/memory_reg[4][1]  ( .D(\Data_Mem/n6105 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[129]), .Q(data_mem_out_wire[129]) );
  DFF \Data_Mem/memory_reg[4][2]  ( .D(\Data_Mem/n6106 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[130]), .Q(data_mem_out_wire[130]) );
  DFF \Data_Mem/memory_reg[4][3]  ( .D(\Data_Mem/n6107 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[131]), .Q(data_mem_out_wire[131]) );
  DFF \Data_Mem/memory_reg[4][4]  ( .D(\Data_Mem/n6108 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[132]), .Q(data_mem_out_wire[132]) );
  DFF \Data_Mem/memory_reg[4][5]  ( .D(\Data_Mem/n6109 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[133]), .Q(data_mem_out_wire[133]) );
  DFF \Data_Mem/memory_reg[4][6]  ( .D(\Data_Mem/n6110 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[134]), .Q(data_mem_out_wire[134]) );
  DFF \Data_Mem/memory_reg[4][7]  ( .D(\Data_Mem/n6111 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[135]), .Q(data_mem_out_wire[135]) );
  DFF \Data_Mem/memory_reg[4][8]  ( .D(\Data_Mem/n6112 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[136]), .Q(data_mem_out_wire[136]) );
  DFF \Data_Mem/memory_reg[4][9]  ( .D(\Data_Mem/n6113 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[137]), .Q(data_mem_out_wire[137]) );
  DFF \Data_Mem/memory_reg[4][10]  ( .D(\Data_Mem/n6114 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[138]), .Q(data_mem_out_wire[138]) );
  DFF \Data_Mem/memory_reg[4][11]  ( .D(\Data_Mem/n6115 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[139]), .Q(data_mem_out_wire[139]) );
  DFF \Data_Mem/memory_reg[4][12]  ( .D(\Data_Mem/n6116 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[140]), .Q(data_mem_out_wire[140]) );
  DFF \Data_Mem/memory_reg[4][13]  ( .D(\Data_Mem/n6117 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[141]), .Q(data_mem_out_wire[141]) );
  DFF \Data_Mem/memory_reg[4][14]  ( .D(\Data_Mem/n6118 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[142]), .Q(data_mem_out_wire[142]) );
  DFF \Data_Mem/memory_reg[4][15]  ( .D(\Data_Mem/n6119 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[143]), .Q(data_mem_out_wire[143]) );
  DFF \Data_Mem/memory_reg[4][16]  ( .D(\Data_Mem/n6120 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[144]), .Q(data_mem_out_wire[144]) );
  DFF \Data_Mem/memory_reg[4][17]  ( .D(\Data_Mem/n6121 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[145]), .Q(data_mem_out_wire[145]) );
  DFF \Data_Mem/memory_reg[4][18]  ( .D(\Data_Mem/n6122 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[146]), .Q(data_mem_out_wire[146]) );
  DFF \Data_Mem/memory_reg[4][19]  ( .D(\Data_Mem/n6123 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[147]), .Q(data_mem_out_wire[147]) );
  DFF \Data_Mem/memory_reg[4][20]  ( .D(\Data_Mem/n6124 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[148]), .Q(data_mem_out_wire[148]) );
  DFF \Data_Mem/memory_reg[4][21]  ( .D(\Data_Mem/n6125 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[149]), .Q(data_mem_out_wire[149]) );
  DFF \Data_Mem/memory_reg[4][22]  ( .D(\Data_Mem/n6126 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[150]), .Q(data_mem_out_wire[150]) );
  DFF \Data_Mem/memory_reg[4][23]  ( .D(\Data_Mem/n6127 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[151]), .Q(data_mem_out_wire[151]) );
  DFF \Data_Mem/memory_reg[4][24]  ( .D(\Data_Mem/n6128 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[152]), .Q(data_mem_out_wire[152]) );
  DFF \Data_Mem/memory_reg[4][25]  ( .D(\Data_Mem/n6129 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[153]), .Q(data_mem_out_wire[153]) );
  DFF \Data_Mem/memory_reg[4][26]  ( .D(\Data_Mem/n6130 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[154]), .Q(data_mem_out_wire[154]) );
  DFF \Data_Mem/memory_reg[4][27]  ( .D(\Data_Mem/n6131 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[155]), .Q(data_mem_out_wire[155]) );
  DFF \Data_Mem/memory_reg[4][28]  ( .D(\Data_Mem/n6132 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[156]), .Q(data_mem_out_wire[156]) );
  DFF \Data_Mem/memory_reg[4][29]  ( .D(\Data_Mem/n6133 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[157]), .Q(data_mem_out_wire[157]) );
  DFF \Data_Mem/memory_reg[4][30]  ( .D(\Data_Mem/n6134 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[158]), .Q(data_mem_out_wire[158]) );
  DFF \Data_Mem/memory_reg[4][31]  ( .D(\Data_Mem/n6135 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[159]), .Q(data_mem_out_wire[159]) );
  DFF \Data_Mem/memory_reg[3][0]  ( .D(\Data_Mem/n6136 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[96]), .Q(data_mem_out_wire[96]) );
  DFF \Data_Mem/memory_reg[3][1]  ( .D(\Data_Mem/n6137 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[97]), .Q(data_mem_out_wire[97]) );
  DFF \Data_Mem/memory_reg[3][2]  ( .D(\Data_Mem/n6138 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[98]), .Q(data_mem_out_wire[98]) );
  DFF \Data_Mem/memory_reg[3][3]  ( .D(\Data_Mem/n6139 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[99]), .Q(data_mem_out_wire[99]) );
  DFF \Data_Mem/memory_reg[3][4]  ( .D(\Data_Mem/n6140 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[100]), .Q(data_mem_out_wire[100]) );
  DFF \Data_Mem/memory_reg[3][5]  ( .D(\Data_Mem/n6141 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[101]), .Q(data_mem_out_wire[101]) );
  DFF \Data_Mem/memory_reg[3][6]  ( .D(\Data_Mem/n6142 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[102]), .Q(data_mem_out_wire[102]) );
  DFF \Data_Mem/memory_reg[3][7]  ( .D(\Data_Mem/n6143 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[103]), .Q(data_mem_out_wire[103]) );
  DFF \Data_Mem/memory_reg[3][8]  ( .D(\Data_Mem/n6144 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[104]), .Q(data_mem_out_wire[104]) );
  DFF \Data_Mem/memory_reg[3][9]  ( .D(\Data_Mem/n6145 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[105]), .Q(data_mem_out_wire[105]) );
  DFF \Data_Mem/memory_reg[3][10]  ( .D(\Data_Mem/n6146 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[106]), .Q(data_mem_out_wire[106]) );
  DFF \Data_Mem/memory_reg[3][11]  ( .D(\Data_Mem/n6147 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[107]), .Q(data_mem_out_wire[107]) );
  DFF \Data_Mem/memory_reg[3][12]  ( .D(\Data_Mem/n6148 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[108]), .Q(data_mem_out_wire[108]) );
  DFF \Data_Mem/memory_reg[3][13]  ( .D(\Data_Mem/n6149 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[109]), .Q(data_mem_out_wire[109]) );
  DFF \Data_Mem/memory_reg[3][14]  ( .D(\Data_Mem/n6150 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[110]), .Q(data_mem_out_wire[110]) );
  DFF \Data_Mem/memory_reg[3][15]  ( .D(\Data_Mem/n6151 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[111]), .Q(data_mem_out_wire[111]) );
  DFF \Data_Mem/memory_reg[3][16]  ( .D(\Data_Mem/n6152 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[112]), .Q(data_mem_out_wire[112]) );
  DFF \Data_Mem/memory_reg[3][17]  ( .D(\Data_Mem/n6153 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[113]), .Q(data_mem_out_wire[113]) );
  DFF \Data_Mem/memory_reg[3][18]  ( .D(\Data_Mem/n6154 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[114]), .Q(data_mem_out_wire[114]) );
  DFF \Data_Mem/memory_reg[3][19]  ( .D(\Data_Mem/n6155 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[115]), .Q(data_mem_out_wire[115]) );
  DFF \Data_Mem/memory_reg[3][20]  ( .D(\Data_Mem/n6156 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[116]), .Q(data_mem_out_wire[116]) );
  DFF \Data_Mem/memory_reg[3][21]  ( .D(\Data_Mem/n6157 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[117]), .Q(data_mem_out_wire[117]) );
  DFF \Data_Mem/memory_reg[3][22]  ( .D(\Data_Mem/n6158 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[118]), .Q(data_mem_out_wire[118]) );
  DFF \Data_Mem/memory_reg[3][23]  ( .D(\Data_Mem/n6159 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[119]), .Q(data_mem_out_wire[119]) );
  DFF \Data_Mem/memory_reg[3][24]  ( .D(\Data_Mem/n6160 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[120]), .Q(data_mem_out_wire[120]) );
  DFF \Data_Mem/memory_reg[3][25]  ( .D(\Data_Mem/n6161 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[121]), .Q(data_mem_out_wire[121]) );
  DFF \Data_Mem/memory_reg[3][26]  ( .D(\Data_Mem/n6162 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[122]), .Q(data_mem_out_wire[122]) );
  DFF \Data_Mem/memory_reg[3][27]  ( .D(\Data_Mem/n6163 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[123]), .Q(data_mem_out_wire[123]) );
  DFF \Data_Mem/memory_reg[3][28]  ( .D(\Data_Mem/n6164 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[124]), .Q(data_mem_out_wire[124]) );
  DFF \Data_Mem/memory_reg[3][29]  ( .D(\Data_Mem/n6165 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[125]), .Q(data_mem_out_wire[125]) );
  DFF \Data_Mem/memory_reg[3][30]  ( .D(\Data_Mem/n6166 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[126]), .Q(data_mem_out_wire[126]) );
  DFF \Data_Mem/memory_reg[3][31]  ( .D(\Data_Mem/n6167 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[127]), .Q(data_mem_out_wire[127]) );
  DFF \Data_Mem/memory_reg[2][0]  ( .D(\Data_Mem/n6168 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[64]), .Q(data_mem_out_wire[64]) );
  DFF \Data_Mem/memory_reg[2][1]  ( .D(\Data_Mem/n6169 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[65]), .Q(data_mem_out_wire[65]) );
  DFF \Data_Mem/memory_reg[2][2]  ( .D(\Data_Mem/n6170 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[66]), .Q(data_mem_out_wire[66]) );
  DFF \Data_Mem/memory_reg[2][3]  ( .D(\Data_Mem/n6171 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[67]), .Q(data_mem_out_wire[67]) );
  DFF \Data_Mem/memory_reg[2][4]  ( .D(\Data_Mem/n6172 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[68]), .Q(data_mem_out_wire[68]) );
  DFF \Data_Mem/memory_reg[2][5]  ( .D(\Data_Mem/n6173 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[69]), .Q(data_mem_out_wire[69]) );
  DFF \Data_Mem/memory_reg[2][6]  ( .D(\Data_Mem/n6174 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[70]), .Q(data_mem_out_wire[70]) );
  DFF \Data_Mem/memory_reg[2][7]  ( .D(\Data_Mem/n6175 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[71]), .Q(data_mem_out_wire[71]) );
  DFF \Data_Mem/memory_reg[2][8]  ( .D(\Data_Mem/n6176 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[72]), .Q(data_mem_out_wire[72]) );
  DFF \Data_Mem/memory_reg[2][9]  ( .D(\Data_Mem/n6177 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[73]), .Q(data_mem_out_wire[73]) );
  DFF \Data_Mem/memory_reg[2][10]  ( .D(\Data_Mem/n6178 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[74]), .Q(data_mem_out_wire[74]) );
  DFF \Data_Mem/memory_reg[2][11]  ( .D(\Data_Mem/n6179 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[75]), .Q(data_mem_out_wire[75]) );
  DFF \Data_Mem/memory_reg[2][12]  ( .D(\Data_Mem/n6180 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[76]), .Q(data_mem_out_wire[76]) );
  DFF \Data_Mem/memory_reg[2][13]  ( .D(\Data_Mem/n6181 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[77]), .Q(data_mem_out_wire[77]) );
  DFF \Data_Mem/memory_reg[2][14]  ( .D(\Data_Mem/n6182 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[78]), .Q(data_mem_out_wire[78]) );
  DFF \Data_Mem/memory_reg[2][15]  ( .D(\Data_Mem/n6183 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[79]), .Q(data_mem_out_wire[79]) );
  DFF \Data_Mem/memory_reg[2][16]  ( .D(\Data_Mem/n6184 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[80]), .Q(data_mem_out_wire[80]) );
  DFF \Data_Mem/memory_reg[2][17]  ( .D(\Data_Mem/n6185 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[81]), .Q(data_mem_out_wire[81]) );
  DFF \Data_Mem/memory_reg[2][18]  ( .D(\Data_Mem/n6186 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[82]), .Q(data_mem_out_wire[82]) );
  DFF \Data_Mem/memory_reg[2][19]  ( .D(\Data_Mem/n6187 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[83]), .Q(data_mem_out_wire[83]) );
  DFF \Data_Mem/memory_reg[2][20]  ( .D(\Data_Mem/n6188 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[84]), .Q(data_mem_out_wire[84]) );
  DFF \Data_Mem/memory_reg[2][21]  ( .D(\Data_Mem/n6189 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[85]), .Q(data_mem_out_wire[85]) );
  DFF \Data_Mem/memory_reg[2][22]  ( .D(\Data_Mem/n6190 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[86]), .Q(data_mem_out_wire[86]) );
  DFF \Data_Mem/memory_reg[2][23]  ( .D(\Data_Mem/n6191 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[87]), .Q(data_mem_out_wire[87]) );
  DFF \Data_Mem/memory_reg[2][24]  ( .D(\Data_Mem/n6192 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[88]), .Q(data_mem_out_wire[88]) );
  DFF \Data_Mem/memory_reg[2][25]  ( .D(\Data_Mem/n6193 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[89]), .Q(data_mem_out_wire[89]) );
  DFF \Data_Mem/memory_reg[2][26]  ( .D(\Data_Mem/n6194 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[90]), .Q(data_mem_out_wire[90]) );
  DFF \Data_Mem/memory_reg[2][27]  ( .D(\Data_Mem/n6195 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[91]), .Q(data_mem_out_wire[91]) );
  DFF \Data_Mem/memory_reg[2][28]  ( .D(\Data_Mem/n6196 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[92]), .Q(data_mem_out_wire[92]) );
  DFF \Data_Mem/memory_reg[2][29]  ( .D(\Data_Mem/n6197 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[93]), .Q(data_mem_out_wire[93]) );
  DFF \Data_Mem/memory_reg[2][30]  ( .D(\Data_Mem/n6198 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[94]), .Q(data_mem_out_wire[94]) );
  DFF \Data_Mem/memory_reg[2][31]  ( .D(\Data_Mem/n6199 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[95]), .Q(data_mem_out_wire[95]) );
  DFF \Data_Mem/memory_reg[1][0]  ( .D(\Data_Mem/n6200 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[32]), .Q(data_mem_out_wire[32]) );
  DFF \Data_Mem/memory_reg[1][1]  ( .D(\Data_Mem/n6201 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[33]), .Q(data_mem_out_wire[33]) );
  DFF \Data_Mem/memory_reg[1][2]  ( .D(\Data_Mem/n6202 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[34]), .Q(data_mem_out_wire[34]) );
  DFF \Data_Mem/memory_reg[1][3]  ( .D(\Data_Mem/n6203 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[35]), .Q(data_mem_out_wire[35]) );
  DFF \Data_Mem/memory_reg[1][4]  ( .D(\Data_Mem/n6204 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[36]), .Q(data_mem_out_wire[36]) );
  DFF \Data_Mem/memory_reg[1][5]  ( .D(\Data_Mem/n6205 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[37]), .Q(data_mem_out_wire[37]) );
  DFF \Data_Mem/memory_reg[1][6]  ( .D(\Data_Mem/n6206 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[38]), .Q(data_mem_out_wire[38]) );
  DFF \Data_Mem/memory_reg[1][7]  ( .D(\Data_Mem/n6207 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[39]), .Q(data_mem_out_wire[39]) );
  DFF \Data_Mem/memory_reg[1][8]  ( .D(\Data_Mem/n6208 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[40]), .Q(data_mem_out_wire[40]) );
  DFF \Data_Mem/memory_reg[1][9]  ( .D(\Data_Mem/n6209 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[41]), .Q(data_mem_out_wire[41]) );
  DFF \Data_Mem/memory_reg[1][10]  ( .D(\Data_Mem/n6210 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[42]), .Q(data_mem_out_wire[42]) );
  DFF \Data_Mem/memory_reg[1][11]  ( .D(\Data_Mem/n6211 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[43]), .Q(data_mem_out_wire[43]) );
  DFF \Data_Mem/memory_reg[1][12]  ( .D(\Data_Mem/n6212 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[44]), .Q(data_mem_out_wire[44]) );
  DFF \Data_Mem/memory_reg[1][13]  ( .D(\Data_Mem/n6213 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[45]), .Q(data_mem_out_wire[45]) );
  DFF \Data_Mem/memory_reg[1][14]  ( .D(\Data_Mem/n6214 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[46]), .Q(data_mem_out_wire[46]) );
  DFF \Data_Mem/memory_reg[1][15]  ( .D(\Data_Mem/n6215 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[47]), .Q(data_mem_out_wire[47]) );
  DFF \Data_Mem/memory_reg[1][16]  ( .D(\Data_Mem/n6216 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[48]), .Q(data_mem_out_wire[48]) );
  DFF \Data_Mem/memory_reg[1][17]  ( .D(\Data_Mem/n6217 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[49]), .Q(data_mem_out_wire[49]) );
  DFF \Data_Mem/memory_reg[1][18]  ( .D(\Data_Mem/n6218 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[50]), .Q(data_mem_out_wire[50]) );
  DFF \Data_Mem/memory_reg[1][19]  ( .D(\Data_Mem/n6219 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[51]), .Q(data_mem_out_wire[51]) );
  DFF \Data_Mem/memory_reg[1][20]  ( .D(\Data_Mem/n6220 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[52]), .Q(data_mem_out_wire[52]) );
  DFF \Data_Mem/memory_reg[1][21]  ( .D(\Data_Mem/n6221 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[53]), .Q(data_mem_out_wire[53]) );
  DFF \Data_Mem/memory_reg[1][22]  ( .D(\Data_Mem/n6222 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[54]), .Q(data_mem_out_wire[54]) );
  DFF \Data_Mem/memory_reg[1][23]  ( .D(\Data_Mem/n6223 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[55]), .Q(data_mem_out_wire[55]) );
  DFF \Data_Mem/memory_reg[1][24]  ( .D(\Data_Mem/n6224 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[56]), .Q(data_mem_out_wire[56]) );
  DFF \Data_Mem/memory_reg[1][25]  ( .D(\Data_Mem/n6225 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[57]), .Q(data_mem_out_wire[57]) );
  DFF \Data_Mem/memory_reg[1][26]  ( .D(\Data_Mem/n6226 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[58]), .Q(data_mem_out_wire[58]) );
  DFF \Data_Mem/memory_reg[1][27]  ( .D(\Data_Mem/n6227 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[59]), .Q(data_mem_out_wire[59]) );
  DFF \Data_Mem/memory_reg[1][28]  ( .D(\Data_Mem/n6228 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[60]), .Q(data_mem_out_wire[60]) );
  DFF \Data_Mem/memory_reg[1][29]  ( .D(\Data_Mem/n6229 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[61]), .Q(data_mem_out_wire[61]) );
  DFF \Data_Mem/memory_reg[1][30]  ( .D(\Data_Mem/n6230 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[62]), .Q(data_mem_out_wire[62]) );
  DFF \Data_Mem/memory_reg[1][31]  ( .D(\Data_Mem/n6231 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[63]), .Q(data_mem_out_wire[63]) );
  DFF \Data_Mem/memory_reg[0][0]  ( .D(\Data_Mem/n6232 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[0]), .Q(data_mem_out_wire[0]) );
  DFF \Data_Mem/memory_reg[0][1]  ( .D(\Data_Mem/n6233 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[1]), .Q(data_mem_out_wire[1]) );
  DFF \Data_Mem/memory_reg[0][2]  ( .D(\Data_Mem/n6234 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[2]), .Q(data_mem_out_wire[2]) );
  DFF \Data_Mem/memory_reg[0][3]  ( .D(\Data_Mem/n6235 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[3]), .Q(data_mem_out_wire[3]) );
  DFF \Data_Mem/memory_reg[0][4]  ( .D(\Data_Mem/n6236 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[4]), .Q(data_mem_out_wire[4]) );
  DFF \Data_Mem/memory_reg[0][5]  ( .D(\Data_Mem/n6237 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[5]), .Q(data_mem_out_wire[5]) );
  DFF \Data_Mem/memory_reg[0][6]  ( .D(\Data_Mem/n6238 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[6]), .Q(data_mem_out_wire[6]) );
  DFF \Data_Mem/memory_reg[0][7]  ( .D(\Data_Mem/n6239 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[7]), .Q(data_mem_out_wire[7]) );
  DFF \Data_Mem/memory_reg[0][8]  ( .D(\Data_Mem/n6240 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[8]), .Q(data_mem_out_wire[8]) );
  DFF \Data_Mem/memory_reg[0][9]  ( .D(\Data_Mem/n6241 ), .CLK(clk), .RST(rst), 
        .I(data_mem_in_wire[9]), .Q(data_mem_out_wire[9]) );
  DFF \Data_Mem/memory_reg[0][10]  ( .D(\Data_Mem/n6242 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[10]), .Q(data_mem_out_wire[10]) );
  DFF \Data_Mem/memory_reg[0][11]  ( .D(\Data_Mem/n6243 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[11]), .Q(data_mem_out_wire[11]) );
  DFF \Data_Mem/memory_reg[0][12]  ( .D(\Data_Mem/n6244 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[12]), .Q(data_mem_out_wire[12]) );
  DFF \Data_Mem/memory_reg[0][13]  ( .D(\Data_Mem/n6245 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[13]), .Q(data_mem_out_wire[13]) );
  DFF \Data_Mem/memory_reg[0][14]  ( .D(\Data_Mem/n6246 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[14]), .Q(data_mem_out_wire[14]) );
  DFF \Data_Mem/memory_reg[0][15]  ( .D(\Data_Mem/n6247 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[15]), .Q(data_mem_out_wire[15]) );
  DFF \Data_Mem/memory_reg[0][16]  ( .D(\Data_Mem/n6248 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[16]), .Q(data_mem_out_wire[16]) );
  DFF \Data_Mem/memory_reg[0][17]  ( .D(\Data_Mem/n6249 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[17]), .Q(data_mem_out_wire[17]) );
  DFF \Data_Mem/memory_reg[0][18]  ( .D(\Data_Mem/n6250 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[18]), .Q(data_mem_out_wire[18]) );
  DFF \Data_Mem/memory_reg[0][19]  ( .D(\Data_Mem/n6251 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[19]), .Q(data_mem_out_wire[19]) );
  DFF \Data_Mem/memory_reg[0][20]  ( .D(\Data_Mem/n6252 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[20]), .Q(data_mem_out_wire[20]) );
  DFF \Data_Mem/memory_reg[0][21]  ( .D(\Data_Mem/n6253 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[21]), .Q(data_mem_out_wire[21]) );
  DFF \Data_Mem/memory_reg[0][22]  ( .D(\Data_Mem/n6254 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[22]), .Q(data_mem_out_wire[22]) );
  DFF \Data_Mem/memory_reg[0][23]  ( .D(\Data_Mem/n6255 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[23]), .Q(data_mem_out_wire[23]) );
  DFF \Data_Mem/memory_reg[0][24]  ( .D(\Data_Mem/n6256 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[24]), .Q(data_mem_out_wire[24]) );
  DFF \Data_Mem/memory_reg[0][25]  ( .D(\Data_Mem/n6257 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[25]), .Q(data_mem_out_wire[25]) );
  DFF \Data_Mem/memory_reg[0][26]  ( .D(\Data_Mem/n6258 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[26]), .Q(data_mem_out_wire[26]) );
  DFF \Data_Mem/memory_reg[0][27]  ( .D(\Data_Mem/n6259 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[27]), .Q(data_mem_out_wire[27]) );
  DFF \Data_Mem/memory_reg[0][28]  ( .D(\Data_Mem/n6260 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[28]), .Q(data_mem_out_wire[28]) );
  DFF \Data_Mem/memory_reg[0][29]  ( .D(\Data_Mem/n6261 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[29]), .Q(data_mem_out_wire[29]) );
  DFF \Data_Mem/memory_reg[0][30]  ( .D(\Data_Mem/n6262 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[30]), .Q(data_mem_out_wire[30]) );
  DFF \Data_Mem/memory_reg[0][31]  ( .D(\Data_Mem/n6263 ), .CLK(clk), .RST(rst), .I(data_mem_in_wire[31]), .Q(data_mem_out_wire[31]) );
  MUX \Reg_Bank/U6038  ( .A(\Reg_Bank/n5941 ), .B(\Reg_Bank/n5926 ), .S(
        rt_index[4]), .Z(reg_target[31]) );
  MUX \Reg_Bank/U6037  ( .A(\Reg_Bank/n5940 ), .B(\Reg_Bank/n5933 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5941 ) );
  MUX \Reg_Bank/U6036  ( .A(\Reg_Bank/n5939 ), .B(\Reg_Bank/n5936 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5940 ) );
  MUX \Reg_Bank/U6035  ( .A(\Reg_Bank/n5938 ), .B(\Reg_Bank/n5937 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5939 ) );
  MUX \Reg_Bank/U6033  ( .A(\Reg_Bank/registers[2][31] ), .B(
        \Reg_Bank/registers[3][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5937 ) );
  MUX \Reg_Bank/U6032  ( .A(\Reg_Bank/n5935 ), .B(\Reg_Bank/n5934 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5936 ) );
  MUX \Reg_Bank/U6031  ( .A(\Reg_Bank/registers[4][31] ), .B(
        \Reg_Bank/registers[5][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5935 ) );
  MUX \Reg_Bank/U6030  ( .A(\Reg_Bank/registers[6][31] ), .B(
        \Reg_Bank/registers[7][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5934 ) );
  MUX \Reg_Bank/U6029  ( .A(\Reg_Bank/n5932 ), .B(\Reg_Bank/n5929 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5933 ) );
  MUX \Reg_Bank/U6028  ( .A(\Reg_Bank/n5931 ), .B(\Reg_Bank/n5930 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5932 ) );
  MUX \Reg_Bank/U6027  ( .A(\Reg_Bank/registers[8][31] ), .B(
        \Reg_Bank/registers[9][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5931 ) );
  MUX \Reg_Bank/U6026  ( .A(\Reg_Bank/registers[10][31] ), .B(
        \Reg_Bank/registers[11][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5930 )
         );
  MUX \Reg_Bank/U6025  ( .A(\Reg_Bank/n5928 ), .B(\Reg_Bank/n5927 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5929 ) );
  MUX \Reg_Bank/U6024  ( .A(\Reg_Bank/registers[12][31] ), .B(
        \Reg_Bank/registers[13][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5928 )
         );
  MUX \Reg_Bank/U6023  ( .A(\Reg_Bank/registers[14][31] ), .B(
        \Reg_Bank/registers[15][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5927 )
         );
  MUX \Reg_Bank/U6022  ( .A(\Reg_Bank/n5925 ), .B(\Reg_Bank/n5918 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5926 ) );
  MUX \Reg_Bank/U6021  ( .A(\Reg_Bank/n5924 ), .B(\Reg_Bank/n5921 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5925 ) );
  MUX \Reg_Bank/U6020  ( .A(\Reg_Bank/n5923 ), .B(\Reg_Bank/n5922 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5924 ) );
  MUX \Reg_Bank/U6019  ( .A(\Reg_Bank/registers[16][31] ), .B(
        \Reg_Bank/registers[17][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5923 )
         );
  MUX \Reg_Bank/U6018  ( .A(\Reg_Bank/registers[18][31] ), .B(
        \Reg_Bank/registers[19][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5922 )
         );
  MUX \Reg_Bank/U6017  ( .A(\Reg_Bank/n5920 ), .B(\Reg_Bank/n5919 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5921 ) );
  MUX \Reg_Bank/U6016  ( .A(\Reg_Bank/registers[20][31] ), .B(
        \Reg_Bank/registers[21][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5920 )
         );
  MUX \Reg_Bank/U6015  ( .A(\Reg_Bank/registers[22][31] ), .B(
        \Reg_Bank/registers[23][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5919 )
         );
  MUX \Reg_Bank/U6014  ( .A(\Reg_Bank/n5917 ), .B(\Reg_Bank/n5914 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5918 ) );
  MUX \Reg_Bank/U6013  ( .A(\Reg_Bank/n5916 ), .B(\Reg_Bank/n5915 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5917 ) );
  MUX \Reg_Bank/U6012  ( .A(\Reg_Bank/registers[24][31] ), .B(
        \Reg_Bank/registers[25][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5916 )
         );
  MUX \Reg_Bank/U6011  ( .A(\Reg_Bank/registers[26][31] ), .B(
        \Reg_Bank/registers[27][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5915 )
         );
  MUX \Reg_Bank/U6010  ( .A(\Reg_Bank/n5913 ), .B(\Reg_Bank/n5912 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5914 ) );
  MUX \Reg_Bank/U6009  ( .A(\Reg_Bank/registers[28][31] ), .B(
        \Reg_Bank/registers[29][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5913 )
         );
  MUX \Reg_Bank/U6008  ( .A(\Reg_Bank/registers[30][31] ), .B(
        \Reg_Bank/registers[31][31] ), .S(rt_index[0]), .Z(\Reg_Bank/n5912 )
         );
  MUX \Reg_Bank/U6007  ( .A(\Reg_Bank/n5911 ), .B(\Reg_Bank/n5896 ), .S(
        rt_index[4]), .Z(reg_target[30]) );
  MUX \Reg_Bank/U6006  ( .A(\Reg_Bank/n5910 ), .B(\Reg_Bank/n5903 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5911 ) );
  MUX \Reg_Bank/U6005  ( .A(\Reg_Bank/n5909 ), .B(\Reg_Bank/n5906 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5910 ) );
  MUX \Reg_Bank/U6004  ( .A(\Reg_Bank/n5908 ), .B(\Reg_Bank/n5907 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5909 ) );
  MUX \Reg_Bank/U6002  ( .A(\Reg_Bank/registers[2][30] ), .B(
        \Reg_Bank/registers[3][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5907 ) );
  MUX \Reg_Bank/U6001  ( .A(\Reg_Bank/n5905 ), .B(\Reg_Bank/n5904 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5906 ) );
  MUX \Reg_Bank/U6000  ( .A(\Reg_Bank/registers[4][30] ), .B(
        \Reg_Bank/registers[5][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5905 ) );
  MUX \Reg_Bank/U5999  ( .A(\Reg_Bank/registers[6][30] ), .B(
        \Reg_Bank/registers[7][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5904 ) );
  MUX \Reg_Bank/U5998  ( .A(\Reg_Bank/n5902 ), .B(\Reg_Bank/n5899 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5903 ) );
  MUX \Reg_Bank/U5997  ( .A(\Reg_Bank/n5901 ), .B(\Reg_Bank/n5900 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5902 ) );
  MUX \Reg_Bank/U5996  ( .A(\Reg_Bank/registers[8][30] ), .B(
        \Reg_Bank/registers[9][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5901 ) );
  MUX \Reg_Bank/U5995  ( .A(\Reg_Bank/registers[10][30] ), .B(
        \Reg_Bank/registers[11][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5900 )
         );
  MUX \Reg_Bank/U5994  ( .A(\Reg_Bank/n5898 ), .B(\Reg_Bank/n5897 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5899 ) );
  MUX \Reg_Bank/U5993  ( .A(\Reg_Bank/registers[12][30] ), .B(
        \Reg_Bank/registers[13][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5898 )
         );
  MUX \Reg_Bank/U5992  ( .A(\Reg_Bank/registers[14][30] ), .B(
        \Reg_Bank/registers[15][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5897 )
         );
  MUX \Reg_Bank/U5991  ( .A(\Reg_Bank/n5895 ), .B(\Reg_Bank/n5888 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5896 ) );
  MUX \Reg_Bank/U5990  ( .A(\Reg_Bank/n5894 ), .B(\Reg_Bank/n5891 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5895 ) );
  MUX \Reg_Bank/U5989  ( .A(\Reg_Bank/n5893 ), .B(\Reg_Bank/n5892 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5894 ) );
  MUX \Reg_Bank/U5988  ( .A(\Reg_Bank/registers[16][30] ), .B(
        \Reg_Bank/registers[17][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5893 )
         );
  MUX \Reg_Bank/U5987  ( .A(\Reg_Bank/registers[18][30] ), .B(
        \Reg_Bank/registers[19][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5892 )
         );
  MUX \Reg_Bank/U5986  ( .A(\Reg_Bank/n5890 ), .B(\Reg_Bank/n5889 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5891 ) );
  MUX \Reg_Bank/U5985  ( .A(\Reg_Bank/registers[20][30] ), .B(
        \Reg_Bank/registers[21][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5890 )
         );
  MUX \Reg_Bank/U5984  ( .A(\Reg_Bank/registers[22][30] ), .B(
        \Reg_Bank/registers[23][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5889 )
         );
  MUX \Reg_Bank/U5983  ( .A(\Reg_Bank/n5887 ), .B(\Reg_Bank/n5884 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5888 ) );
  MUX \Reg_Bank/U5982  ( .A(\Reg_Bank/n5886 ), .B(\Reg_Bank/n5885 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5887 ) );
  MUX \Reg_Bank/U5981  ( .A(\Reg_Bank/registers[24][30] ), .B(
        \Reg_Bank/registers[25][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5886 )
         );
  MUX \Reg_Bank/U5980  ( .A(\Reg_Bank/registers[26][30] ), .B(
        \Reg_Bank/registers[27][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5885 )
         );
  MUX \Reg_Bank/U5979  ( .A(\Reg_Bank/n5883 ), .B(\Reg_Bank/n5882 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5884 ) );
  MUX \Reg_Bank/U5978  ( .A(\Reg_Bank/registers[28][30] ), .B(
        \Reg_Bank/registers[29][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5883 )
         );
  MUX \Reg_Bank/U5977  ( .A(\Reg_Bank/registers[30][30] ), .B(
        \Reg_Bank/registers[31][30] ), .S(rt_index[0]), .Z(\Reg_Bank/n5882 )
         );
  MUX \Reg_Bank/U5976  ( .A(\Reg_Bank/n5881 ), .B(\Reg_Bank/n5866 ), .S(
        rt_index[4]), .Z(reg_target[29]) );
  MUX \Reg_Bank/U5975  ( .A(\Reg_Bank/n5880 ), .B(\Reg_Bank/n5873 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5881 ) );
  MUX \Reg_Bank/U5974  ( .A(\Reg_Bank/n5879 ), .B(\Reg_Bank/n5876 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5880 ) );
  MUX \Reg_Bank/U5973  ( .A(\Reg_Bank/n5878 ), .B(\Reg_Bank/n5877 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5879 ) );
  MUX \Reg_Bank/U5971  ( .A(\Reg_Bank/registers[2][29] ), .B(
        \Reg_Bank/registers[3][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5877 ) );
  MUX \Reg_Bank/U5970  ( .A(\Reg_Bank/n5875 ), .B(\Reg_Bank/n5874 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5876 ) );
  MUX \Reg_Bank/U5969  ( .A(\Reg_Bank/registers[4][29] ), .B(
        \Reg_Bank/registers[5][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5875 ) );
  MUX \Reg_Bank/U5968  ( .A(\Reg_Bank/registers[6][29] ), .B(
        \Reg_Bank/registers[7][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5874 ) );
  MUX \Reg_Bank/U5967  ( .A(\Reg_Bank/n5872 ), .B(\Reg_Bank/n5869 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5873 ) );
  MUX \Reg_Bank/U5966  ( .A(\Reg_Bank/n5871 ), .B(\Reg_Bank/n5870 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5872 ) );
  MUX \Reg_Bank/U5965  ( .A(\Reg_Bank/registers[8][29] ), .B(
        \Reg_Bank/registers[9][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5871 ) );
  MUX \Reg_Bank/U5964  ( .A(\Reg_Bank/registers[10][29] ), .B(
        \Reg_Bank/registers[11][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5870 )
         );
  MUX \Reg_Bank/U5963  ( .A(\Reg_Bank/n5868 ), .B(\Reg_Bank/n5867 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5869 ) );
  MUX \Reg_Bank/U5962  ( .A(\Reg_Bank/registers[12][29] ), .B(
        \Reg_Bank/registers[13][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5868 )
         );
  MUX \Reg_Bank/U5961  ( .A(\Reg_Bank/registers[14][29] ), .B(
        \Reg_Bank/registers[15][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5867 )
         );
  MUX \Reg_Bank/U5960  ( .A(\Reg_Bank/n5865 ), .B(\Reg_Bank/n5858 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5866 ) );
  MUX \Reg_Bank/U5959  ( .A(\Reg_Bank/n5864 ), .B(\Reg_Bank/n5861 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5865 ) );
  MUX \Reg_Bank/U5958  ( .A(\Reg_Bank/n5863 ), .B(\Reg_Bank/n5862 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5864 ) );
  MUX \Reg_Bank/U5957  ( .A(\Reg_Bank/registers[16][29] ), .B(
        \Reg_Bank/registers[17][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5863 )
         );
  MUX \Reg_Bank/U5956  ( .A(\Reg_Bank/registers[18][29] ), .B(
        \Reg_Bank/registers[19][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5862 )
         );
  MUX \Reg_Bank/U5955  ( .A(\Reg_Bank/n5860 ), .B(\Reg_Bank/n5859 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5861 ) );
  MUX \Reg_Bank/U5954  ( .A(\Reg_Bank/registers[20][29] ), .B(
        \Reg_Bank/registers[21][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5860 )
         );
  MUX \Reg_Bank/U5953  ( .A(\Reg_Bank/registers[22][29] ), .B(
        \Reg_Bank/registers[23][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5859 )
         );
  MUX \Reg_Bank/U5952  ( .A(\Reg_Bank/n5857 ), .B(\Reg_Bank/n5854 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5858 ) );
  MUX \Reg_Bank/U5951  ( .A(\Reg_Bank/n5856 ), .B(\Reg_Bank/n5855 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5857 ) );
  MUX \Reg_Bank/U5950  ( .A(\Reg_Bank/registers[24][29] ), .B(
        \Reg_Bank/registers[25][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5856 )
         );
  MUX \Reg_Bank/U5949  ( .A(\Reg_Bank/registers[26][29] ), .B(
        \Reg_Bank/registers[27][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5855 )
         );
  MUX \Reg_Bank/U5948  ( .A(\Reg_Bank/n5853 ), .B(\Reg_Bank/n5852 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5854 ) );
  MUX \Reg_Bank/U5947  ( .A(\Reg_Bank/registers[28][29] ), .B(
        \Reg_Bank/registers[29][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5853 )
         );
  MUX \Reg_Bank/U5946  ( .A(\Reg_Bank/registers[30][29] ), .B(
        \Reg_Bank/registers[31][29] ), .S(rt_index[0]), .Z(\Reg_Bank/n5852 )
         );
  MUX \Reg_Bank/U5945  ( .A(\Reg_Bank/n5851 ), .B(\Reg_Bank/n5836 ), .S(
        rt_index[4]), .Z(reg_target[28]) );
  MUX \Reg_Bank/U5944  ( .A(\Reg_Bank/n5850 ), .B(\Reg_Bank/n5843 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5851 ) );
  MUX \Reg_Bank/U5943  ( .A(\Reg_Bank/n5849 ), .B(\Reg_Bank/n5846 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5850 ) );
  MUX \Reg_Bank/U5942  ( .A(\Reg_Bank/n5848 ), .B(\Reg_Bank/n5847 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5849 ) );
  MUX \Reg_Bank/U5940  ( .A(\Reg_Bank/registers[2][28] ), .B(
        \Reg_Bank/registers[3][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5847 ) );
  MUX \Reg_Bank/U5939  ( .A(\Reg_Bank/n5845 ), .B(\Reg_Bank/n5844 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5846 ) );
  MUX \Reg_Bank/U5938  ( .A(\Reg_Bank/registers[4][28] ), .B(
        \Reg_Bank/registers[5][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5845 ) );
  MUX \Reg_Bank/U5937  ( .A(\Reg_Bank/registers[6][28] ), .B(
        \Reg_Bank/registers[7][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5844 ) );
  MUX \Reg_Bank/U5936  ( .A(\Reg_Bank/n5842 ), .B(\Reg_Bank/n5839 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5843 ) );
  MUX \Reg_Bank/U5935  ( .A(\Reg_Bank/n5841 ), .B(\Reg_Bank/n5840 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5842 ) );
  MUX \Reg_Bank/U5934  ( .A(\Reg_Bank/registers[8][28] ), .B(
        \Reg_Bank/registers[9][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5841 ) );
  MUX \Reg_Bank/U5933  ( .A(\Reg_Bank/registers[10][28] ), .B(
        \Reg_Bank/registers[11][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5840 )
         );
  MUX \Reg_Bank/U5932  ( .A(\Reg_Bank/n5838 ), .B(\Reg_Bank/n5837 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5839 ) );
  MUX \Reg_Bank/U5931  ( .A(\Reg_Bank/registers[12][28] ), .B(
        \Reg_Bank/registers[13][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5838 )
         );
  MUX \Reg_Bank/U5930  ( .A(\Reg_Bank/registers[14][28] ), .B(
        \Reg_Bank/registers[15][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5837 )
         );
  MUX \Reg_Bank/U5929  ( .A(\Reg_Bank/n5835 ), .B(\Reg_Bank/n5828 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5836 ) );
  MUX \Reg_Bank/U5928  ( .A(\Reg_Bank/n5834 ), .B(\Reg_Bank/n5831 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5835 ) );
  MUX \Reg_Bank/U5927  ( .A(\Reg_Bank/n5833 ), .B(\Reg_Bank/n5832 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5834 ) );
  MUX \Reg_Bank/U5926  ( .A(\Reg_Bank/registers[16][28] ), .B(
        \Reg_Bank/registers[17][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5833 )
         );
  MUX \Reg_Bank/U5925  ( .A(\Reg_Bank/registers[18][28] ), .B(
        \Reg_Bank/registers[19][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5832 )
         );
  MUX \Reg_Bank/U5924  ( .A(\Reg_Bank/n5830 ), .B(\Reg_Bank/n5829 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5831 ) );
  MUX \Reg_Bank/U5923  ( .A(\Reg_Bank/registers[20][28] ), .B(
        \Reg_Bank/registers[21][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5830 )
         );
  MUX \Reg_Bank/U5922  ( .A(\Reg_Bank/registers[22][28] ), .B(
        \Reg_Bank/registers[23][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5829 )
         );
  MUX \Reg_Bank/U5921  ( .A(\Reg_Bank/n5827 ), .B(\Reg_Bank/n5824 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5828 ) );
  MUX \Reg_Bank/U5920  ( .A(\Reg_Bank/n5826 ), .B(\Reg_Bank/n5825 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5827 ) );
  MUX \Reg_Bank/U5919  ( .A(\Reg_Bank/registers[24][28] ), .B(
        \Reg_Bank/registers[25][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5826 )
         );
  MUX \Reg_Bank/U5918  ( .A(\Reg_Bank/registers[26][28] ), .B(
        \Reg_Bank/registers[27][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5825 )
         );
  MUX \Reg_Bank/U5917  ( .A(\Reg_Bank/n5823 ), .B(\Reg_Bank/n5822 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5824 ) );
  MUX \Reg_Bank/U5916  ( .A(\Reg_Bank/registers[28][28] ), .B(
        \Reg_Bank/registers[29][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5823 )
         );
  MUX \Reg_Bank/U5915  ( .A(\Reg_Bank/registers[30][28] ), .B(
        \Reg_Bank/registers[31][28] ), .S(rt_index[0]), .Z(\Reg_Bank/n5822 )
         );
  MUX \Reg_Bank/U5914  ( .A(\Reg_Bank/n5821 ), .B(\Reg_Bank/n5806 ), .S(
        rt_index[4]), .Z(reg_target[27]) );
  MUX \Reg_Bank/U5913  ( .A(\Reg_Bank/n5820 ), .B(\Reg_Bank/n5813 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5821 ) );
  MUX \Reg_Bank/U5912  ( .A(\Reg_Bank/n5819 ), .B(\Reg_Bank/n5816 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5820 ) );
  MUX \Reg_Bank/U5911  ( .A(\Reg_Bank/n5818 ), .B(\Reg_Bank/n5817 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5819 ) );
  MUX \Reg_Bank/U5909  ( .A(\Reg_Bank/registers[2][27] ), .B(
        \Reg_Bank/registers[3][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5817 ) );
  MUX \Reg_Bank/U5908  ( .A(\Reg_Bank/n5815 ), .B(\Reg_Bank/n5814 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5816 ) );
  MUX \Reg_Bank/U5907  ( .A(\Reg_Bank/registers[4][27] ), .B(
        \Reg_Bank/registers[5][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5815 ) );
  MUX \Reg_Bank/U5906  ( .A(\Reg_Bank/registers[6][27] ), .B(
        \Reg_Bank/registers[7][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5814 ) );
  MUX \Reg_Bank/U5905  ( .A(\Reg_Bank/n5812 ), .B(\Reg_Bank/n5809 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5813 ) );
  MUX \Reg_Bank/U5904  ( .A(\Reg_Bank/n5811 ), .B(\Reg_Bank/n5810 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5812 ) );
  MUX \Reg_Bank/U5903  ( .A(\Reg_Bank/registers[8][27] ), .B(
        \Reg_Bank/registers[9][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5811 ) );
  MUX \Reg_Bank/U5902  ( .A(\Reg_Bank/registers[10][27] ), .B(
        \Reg_Bank/registers[11][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5810 )
         );
  MUX \Reg_Bank/U5901  ( .A(\Reg_Bank/n5808 ), .B(\Reg_Bank/n5807 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5809 ) );
  MUX \Reg_Bank/U5900  ( .A(\Reg_Bank/registers[12][27] ), .B(
        \Reg_Bank/registers[13][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5808 )
         );
  MUX \Reg_Bank/U5899  ( .A(\Reg_Bank/registers[14][27] ), .B(
        \Reg_Bank/registers[15][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5807 )
         );
  MUX \Reg_Bank/U5898  ( .A(\Reg_Bank/n5805 ), .B(\Reg_Bank/n5798 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5806 ) );
  MUX \Reg_Bank/U5897  ( .A(\Reg_Bank/n5804 ), .B(\Reg_Bank/n5801 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5805 ) );
  MUX \Reg_Bank/U5896  ( .A(\Reg_Bank/n5803 ), .B(\Reg_Bank/n5802 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5804 ) );
  MUX \Reg_Bank/U5895  ( .A(\Reg_Bank/registers[16][27] ), .B(
        \Reg_Bank/registers[17][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5803 )
         );
  MUX \Reg_Bank/U5894  ( .A(\Reg_Bank/registers[18][27] ), .B(
        \Reg_Bank/registers[19][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5802 )
         );
  MUX \Reg_Bank/U5893  ( .A(\Reg_Bank/n5800 ), .B(\Reg_Bank/n5799 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5801 ) );
  MUX \Reg_Bank/U5892  ( .A(\Reg_Bank/registers[20][27] ), .B(
        \Reg_Bank/registers[21][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5800 )
         );
  MUX \Reg_Bank/U5891  ( .A(\Reg_Bank/registers[22][27] ), .B(
        \Reg_Bank/registers[23][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5799 )
         );
  MUX \Reg_Bank/U5890  ( .A(\Reg_Bank/n5797 ), .B(\Reg_Bank/n5794 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5798 ) );
  MUX \Reg_Bank/U5889  ( .A(\Reg_Bank/n5796 ), .B(\Reg_Bank/n5795 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5797 ) );
  MUX \Reg_Bank/U5888  ( .A(\Reg_Bank/registers[24][27] ), .B(
        \Reg_Bank/registers[25][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5796 )
         );
  MUX \Reg_Bank/U5887  ( .A(\Reg_Bank/registers[26][27] ), .B(
        \Reg_Bank/registers[27][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5795 )
         );
  MUX \Reg_Bank/U5886  ( .A(\Reg_Bank/n5793 ), .B(\Reg_Bank/n5792 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5794 ) );
  MUX \Reg_Bank/U5885  ( .A(\Reg_Bank/registers[28][27] ), .B(
        \Reg_Bank/registers[29][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5793 )
         );
  MUX \Reg_Bank/U5884  ( .A(\Reg_Bank/registers[30][27] ), .B(
        \Reg_Bank/registers[31][27] ), .S(rt_index[0]), .Z(\Reg_Bank/n5792 )
         );
  MUX \Reg_Bank/U5883  ( .A(\Reg_Bank/n5791 ), .B(\Reg_Bank/n5776 ), .S(
        rt_index[4]), .Z(reg_target[26]) );
  MUX \Reg_Bank/U5882  ( .A(\Reg_Bank/n5790 ), .B(\Reg_Bank/n5783 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5791 ) );
  MUX \Reg_Bank/U5881  ( .A(\Reg_Bank/n5789 ), .B(\Reg_Bank/n5786 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5790 ) );
  MUX \Reg_Bank/U5880  ( .A(\Reg_Bank/n5788 ), .B(\Reg_Bank/n5787 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5789 ) );
  MUX \Reg_Bank/U5878  ( .A(\Reg_Bank/registers[2][26] ), .B(
        \Reg_Bank/registers[3][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5787 ) );
  MUX \Reg_Bank/U5877  ( .A(\Reg_Bank/n5785 ), .B(\Reg_Bank/n5784 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5786 ) );
  MUX \Reg_Bank/U5876  ( .A(\Reg_Bank/registers[4][26] ), .B(
        \Reg_Bank/registers[5][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5785 ) );
  MUX \Reg_Bank/U5875  ( .A(\Reg_Bank/registers[6][26] ), .B(
        \Reg_Bank/registers[7][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5784 ) );
  MUX \Reg_Bank/U5874  ( .A(\Reg_Bank/n5782 ), .B(\Reg_Bank/n5779 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5783 ) );
  MUX \Reg_Bank/U5873  ( .A(\Reg_Bank/n5781 ), .B(\Reg_Bank/n5780 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5782 ) );
  MUX \Reg_Bank/U5872  ( .A(\Reg_Bank/registers[8][26] ), .B(
        \Reg_Bank/registers[9][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5781 ) );
  MUX \Reg_Bank/U5871  ( .A(\Reg_Bank/registers[10][26] ), .B(
        \Reg_Bank/registers[11][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5780 )
         );
  MUX \Reg_Bank/U5870  ( .A(\Reg_Bank/n5778 ), .B(\Reg_Bank/n5777 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5779 ) );
  MUX \Reg_Bank/U5869  ( .A(\Reg_Bank/registers[12][26] ), .B(
        \Reg_Bank/registers[13][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5778 )
         );
  MUX \Reg_Bank/U5868  ( .A(\Reg_Bank/registers[14][26] ), .B(
        \Reg_Bank/registers[15][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5777 )
         );
  MUX \Reg_Bank/U5867  ( .A(\Reg_Bank/n5775 ), .B(\Reg_Bank/n5768 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5776 ) );
  MUX \Reg_Bank/U5866  ( .A(\Reg_Bank/n5774 ), .B(\Reg_Bank/n5771 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5775 ) );
  MUX \Reg_Bank/U5865  ( .A(\Reg_Bank/n5773 ), .B(\Reg_Bank/n5772 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5774 ) );
  MUX \Reg_Bank/U5864  ( .A(\Reg_Bank/registers[16][26] ), .B(
        \Reg_Bank/registers[17][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5773 )
         );
  MUX \Reg_Bank/U5863  ( .A(\Reg_Bank/registers[18][26] ), .B(
        \Reg_Bank/registers[19][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5772 )
         );
  MUX \Reg_Bank/U5862  ( .A(\Reg_Bank/n5770 ), .B(\Reg_Bank/n5769 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5771 ) );
  MUX \Reg_Bank/U5861  ( .A(\Reg_Bank/registers[20][26] ), .B(
        \Reg_Bank/registers[21][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5770 )
         );
  MUX \Reg_Bank/U5860  ( .A(\Reg_Bank/registers[22][26] ), .B(
        \Reg_Bank/registers[23][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5769 )
         );
  MUX \Reg_Bank/U5859  ( .A(\Reg_Bank/n5767 ), .B(\Reg_Bank/n5764 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5768 ) );
  MUX \Reg_Bank/U5858  ( .A(\Reg_Bank/n5766 ), .B(\Reg_Bank/n5765 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5767 ) );
  MUX \Reg_Bank/U5857  ( .A(\Reg_Bank/registers[24][26] ), .B(
        \Reg_Bank/registers[25][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5766 )
         );
  MUX \Reg_Bank/U5856  ( .A(\Reg_Bank/registers[26][26] ), .B(
        \Reg_Bank/registers[27][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5765 )
         );
  MUX \Reg_Bank/U5855  ( .A(\Reg_Bank/n5763 ), .B(\Reg_Bank/n5762 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5764 ) );
  MUX \Reg_Bank/U5854  ( .A(\Reg_Bank/registers[28][26] ), .B(
        \Reg_Bank/registers[29][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5763 )
         );
  MUX \Reg_Bank/U5853  ( .A(\Reg_Bank/registers[30][26] ), .B(
        \Reg_Bank/registers[31][26] ), .S(rt_index[0]), .Z(\Reg_Bank/n5762 )
         );
  MUX \Reg_Bank/U5852  ( .A(\Reg_Bank/n5761 ), .B(\Reg_Bank/n5746 ), .S(
        rt_index[4]), .Z(reg_target[25]) );
  MUX \Reg_Bank/U5851  ( .A(\Reg_Bank/n5760 ), .B(\Reg_Bank/n5753 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5761 ) );
  MUX \Reg_Bank/U5850  ( .A(\Reg_Bank/n5759 ), .B(\Reg_Bank/n5756 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5760 ) );
  MUX \Reg_Bank/U5849  ( .A(\Reg_Bank/n5758 ), .B(\Reg_Bank/n5757 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5759 ) );
  MUX \Reg_Bank/U5847  ( .A(\Reg_Bank/registers[2][25] ), .B(
        \Reg_Bank/registers[3][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5757 ) );
  MUX \Reg_Bank/U5846  ( .A(\Reg_Bank/n5755 ), .B(\Reg_Bank/n5754 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5756 ) );
  MUX \Reg_Bank/U5845  ( .A(\Reg_Bank/registers[4][25] ), .B(
        \Reg_Bank/registers[5][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5755 ) );
  MUX \Reg_Bank/U5844  ( .A(\Reg_Bank/registers[6][25] ), .B(
        \Reg_Bank/registers[7][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5754 ) );
  MUX \Reg_Bank/U5843  ( .A(\Reg_Bank/n5752 ), .B(\Reg_Bank/n5749 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5753 ) );
  MUX \Reg_Bank/U5842  ( .A(\Reg_Bank/n5751 ), .B(\Reg_Bank/n5750 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5752 ) );
  MUX \Reg_Bank/U5841  ( .A(\Reg_Bank/registers[8][25] ), .B(
        \Reg_Bank/registers[9][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5751 ) );
  MUX \Reg_Bank/U5840  ( .A(\Reg_Bank/registers[10][25] ), .B(
        \Reg_Bank/registers[11][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5750 )
         );
  MUX \Reg_Bank/U5839  ( .A(\Reg_Bank/n5748 ), .B(\Reg_Bank/n5747 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5749 ) );
  MUX \Reg_Bank/U5838  ( .A(\Reg_Bank/registers[12][25] ), .B(
        \Reg_Bank/registers[13][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5748 )
         );
  MUX \Reg_Bank/U5837  ( .A(\Reg_Bank/registers[14][25] ), .B(
        \Reg_Bank/registers[15][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5747 )
         );
  MUX \Reg_Bank/U5836  ( .A(\Reg_Bank/n5745 ), .B(\Reg_Bank/n5738 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5746 ) );
  MUX \Reg_Bank/U5835  ( .A(\Reg_Bank/n5744 ), .B(\Reg_Bank/n5741 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5745 ) );
  MUX \Reg_Bank/U5834  ( .A(\Reg_Bank/n5743 ), .B(\Reg_Bank/n5742 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5744 ) );
  MUX \Reg_Bank/U5833  ( .A(\Reg_Bank/registers[16][25] ), .B(
        \Reg_Bank/registers[17][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5743 )
         );
  MUX \Reg_Bank/U5832  ( .A(\Reg_Bank/registers[18][25] ), .B(
        \Reg_Bank/registers[19][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5742 )
         );
  MUX \Reg_Bank/U5831  ( .A(\Reg_Bank/n5740 ), .B(\Reg_Bank/n5739 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5741 ) );
  MUX \Reg_Bank/U5830  ( .A(\Reg_Bank/registers[20][25] ), .B(
        \Reg_Bank/registers[21][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5740 )
         );
  MUX \Reg_Bank/U5829  ( .A(\Reg_Bank/registers[22][25] ), .B(
        \Reg_Bank/registers[23][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5739 )
         );
  MUX \Reg_Bank/U5828  ( .A(\Reg_Bank/n5737 ), .B(\Reg_Bank/n5734 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5738 ) );
  MUX \Reg_Bank/U5827  ( .A(\Reg_Bank/n5736 ), .B(\Reg_Bank/n5735 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5737 ) );
  MUX \Reg_Bank/U5826  ( .A(\Reg_Bank/registers[24][25] ), .B(
        \Reg_Bank/registers[25][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5736 )
         );
  MUX \Reg_Bank/U5825  ( .A(\Reg_Bank/registers[26][25] ), .B(
        \Reg_Bank/registers[27][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5735 )
         );
  MUX \Reg_Bank/U5824  ( .A(\Reg_Bank/n5733 ), .B(\Reg_Bank/n5732 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5734 ) );
  MUX \Reg_Bank/U5823  ( .A(\Reg_Bank/registers[28][25] ), .B(
        \Reg_Bank/registers[29][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5733 )
         );
  MUX \Reg_Bank/U5822  ( .A(\Reg_Bank/registers[30][25] ), .B(
        \Reg_Bank/registers[31][25] ), .S(rt_index[0]), .Z(\Reg_Bank/n5732 )
         );
  MUX \Reg_Bank/U5821  ( .A(\Reg_Bank/n5731 ), .B(\Reg_Bank/n5716 ), .S(
        rt_index[4]), .Z(reg_target[24]) );
  MUX \Reg_Bank/U5820  ( .A(\Reg_Bank/n5730 ), .B(\Reg_Bank/n5723 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5731 ) );
  MUX \Reg_Bank/U5819  ( .A(\Reg_Bank/n5729 ), .B(\Reg_Bank/n5726 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5730 ) );
  MUX \Reg_Bank/U5818  ( .A(\Reg_Bank/n5728 ), .B(\Reg_Bank/n5727 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5729 ) );
  MUX \Reg_Bank/U5816  ( .A(\Reg_Bank/registers[2][24] ), .B(
        \Reg_Bank/registers[3][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5727 ) );
  MUX \Reg_Bank/U5815  ( .A(\Reg_Bank/n5725 ), .B(\Reg_Bank/n5724 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5726 ) );
  MUX \Reg_Bank/U5814  ( .A(\Reg_Bank/registers[4][24] ), .B(
        \Reg_Bank/registers[5][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5725 ) );
  MUX \Reg_Bank/U5813  ( .A(\Reg_Bank/registers[6][24] ), .B(
        \Reg_Bank/registers[7][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5724 ) );
  MUX \Reg_Bank/U5812  ( .A(\Reg_Bank/n5722 ), .B(\Reg_Bank/n5719 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5723 ) );
  MUX \Reg_Bank/U5811  ( .A(\Reg_Bank/n5721 ), .B(\Reg_Bank/n5720 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5722 ) );
  MUX \Reg_Bank/U5810  ( .A(\Reg_Bank/registers[8][24] ), .B(
        \Reg_Bank/registers[9][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5721 ) );
  MUX \Reg_Bank/U5809  ( .A(\Reg_Bank/registers[10][24] ), .B(
        \Reg_Bank/registers[11][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5720 )
         );
  MUX \Reg_Bank/U5808  ( .A(\Reg_Bank/n5718 ), .B(\Reg_Bank/n5717 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5719 ) );
  MUX \Reg_Bank/U5807  ( .A(\Reg_Bank/registers[12][24] ), .B(
        \Reg_Bank/registers[13][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5718 )
         );
  MUX \Reg_Bank/U5806  ( .A(\Reg_Bank/registers[14][24] ), .B(
        \Reg_Bank/registers[15][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5717 )
         );
  MUX \Reg_Bank/U5805  ( .A(\Reg_Bank/n5715 ), .B(\Reg_Bank/n5708 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5716 ) );
  MUX \Reg_Bank/U5804  ( .A(\Reg_Bank/n5714 ), .B(\Reg_Bank/n5711 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5715 ) );
  MUX \Reg_Bank/U5803  ( .A(\Reg_Bank/n5713 ), .B(\Reg_Bank/n5712 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5714 ) );
  MUX \Reg_Bank/U5802  ( .A(\Reg_Bank/registers[16][24] ), .B(
        \Reg_Bank/registers[17][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5713 )
         );
  MUX \Reg_Bank/U5801  ( .A(\Reg_Bank/registers[18][24] ), .B(
        \Reg_Bank/registers[19][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5712 )
         );
  MUX \Reg_Bank/U5800  ( .A(\Reg_Bank/n5710 ), .B(\Reg_Bank/n5709 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5711 ) );
  MUX \Reg_Bank/U5799  ( .A(\Reg_Bank/registers[20][24] ), .B(
        \Reg_Bank/registers[21][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5710 )
         );
  MUX \Reg_Bank/U5798  ( .A(\Reg_Bank/registers[22][24] ), .B(
        \Reg_Bank/registers[23][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5709 )
         );
  MUX \Reg_Bank/U5797  ( .A(\Reg_Bank/n5707 ), .B(\Reg_Bank/n5704 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5708 ) );
  MUX \Reg_Bank/U5796  ( .A(\Reg_Bank/n5706 ), .B(\Reg_Bank/n5705 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5707 ) );
  MUX \Reg_Bank/U5795  ( .A(\Reg_Bank/registers[24][24] ), .B(
        \Reg_Bank/registers[25][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5706 )
         );
  MUX \Reg_Bank/U5794  ( .A(\Reg_Bank/registers[26][24] ), .B(
        \Reg_Bank/registers[27][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5705 )
         );
  MUX \Reg_Bank/U5793  ( .A(\Reg_Bank/n5703 ), .B(\Reg_Bank/n5702 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5704 ) );
  MUX \Reg_Bank/U5792  ( .A(\Reg_Bank/registers[28][24] ), .B(
        \Reg_Bank/registers[29][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5703 )
         );
  MUX \Reg_Bank/U5791  ( .A(\Reg_Bank/registers[30][24] ), .B(
        \Reg_Bank/registers[31][24] ), .S(rt_index[0]), .Z(\Reg_Bank/n5702 )
         );
  MUX \Reg_Bank/U5790  ( .A(\Reg_Bank/n5701 ), .B(\Reg_Bank/n5686 ), .S(
        rt_index[4]), .Z(reg_target[23]) );
  MUX \Reg_Bank/U5789  ( .A(\Reg_Bank/n5700 ), .B(\Reg_Bank/n5693 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5701 ) );
  MUX \Reg_Bank/U5788  ( .A(\Reg_Bank/n5699 ), .B(\Reg_Bank/n5696 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5700 ) );
  MUX \Reg_Bank/U5787  ( .A(\Reg_Bank/n5698 ), .B(\Reg_Bank/n5697 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5699 ) );
  MUX \Reg_Bank/U5785  ( .A(\Reg_Bank/registers[2][23] ), .B(
        \Reg_Bank/registers[3][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5697 ) );
  MUX \Reg_Bank/U5784  ( .A(\Reg_Bank/n5695 ), .B(\Reg_Bank/n5694 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5696 ) );
  MUX \Reg_Bank/U5783  ( .A(\Reg_Bank/registers[4][23] ), .B(
        \Reg_Bank/registers[5][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5695 ) );
  MUX \Reg_Bank/U5782  ( .A(\Reg_Bank/registers[6][23] ), .B(
        \Reg_Bank/registers[7][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5694 ) );
  MUX \Reg_Bank/U5781  ( .A(\Reg_Bank/n5692 ), .B(\Reg_Bank/n5689 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5693 ) );
  MUX \Reg_Bank/U5780  ( .A(\Reg_Bank/n5691 ), .B(\Reg_Bank/n5690 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5692 ) );
  MUX \Reg_Bank/U5779  ( .A(\Reg_Bank/registers[8][23] ), .B(
        \Reg_Bank/registers[9][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5691 ) );
  MUX \Reg_Bank/U5778  ( .A(\Reg_Bank/registers[10][23] ), .B(
        \Reg_Bank/registers[11][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5690 )
         );
  MUX \Reg_Bank/U5777  ( .A(\Reg_Bank/n5688 ), .B(\Reg_Bank/n5687 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5689 ) );
  MUX \Reg_Bank/U5776  ( .A(\Reg_Bank/registers[12][23] ), .B(
        \Reg_Bank/registers[13][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5688 )
         );
  MUX \Reg_Bank/U5775  ( .A(\Reg_Bank/registers[14][23] ), .B(
        \Reg_Bank/registers[15][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5687 )
         );
  MUX \Reg_Bank/U5774  ( .A(\Reg_Bank/n5685 ), .B(\Reg_Bank/n5678 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5686 ) );
  MUX \Reg_Bank/U5773  ( .A(\Reg_Bank/n5684 ), .B(\Reg_Bank/n5681 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5685 ) );
  MUX \Reg_Bank/U5772  ( .A(\Reg_Bank/n5683 ), .B(\Reg_Bank/n5682 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5684 ) );
  MUX \Reg_Bank/U5771  ( .A(\Reg_Bank/registers[16][23] ), .B(
        \Reg_Bank/registers[17][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5683 )
         );
  MUX \Reg_Bank/U5770  ( .A(\Reg_Bank/registers[18][23] ), .B(
        \Reg_Bank/registers[19][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5682 )
         );
  MUX \Reg_Bank/U5769  ( .A(\Reg_Bank/n5680 ), .B(\Reg_Bank/n5679 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5681 ) );
  MUX \Reg_Bank/U5768  ( .A(\Reg_Bank/registers[20][23] ), .B(
        \Reg_Bank/registers[21][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5680 )
         );
  MUX \Reg_Bank/U5767  ( .A(\Reg_Bank/registers[22][23] ), .B(
        \Reg_Bank/registers[23][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5679 )
         );
  MUX \Reg_Bank/U5766  ( .A(\Reg_Bank/n5677 ), .B(\Reg_Bank/n5674 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5678 ) );
  MUX \Reg_Bank/U5765  ( .A(\Reg_Bank/n5676 ), .B(\Reg_Bank/n5675 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5677 ) );
  MUX \Reg_Bank/U5764  ( .A(\Reg_Bank/registers[24][23] ), .B(
        \Reg_Bank/registers[25][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5676 )
         );
  MUX \Reg_Bank/U5763  ( .A(\Reg_Bank/registers[26][23] ), .B(
        \Reg_Bank/registers[27][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5675 )
         );
  MUX \Reg_Bank/U5762  ( .A(\Reg_Bank/n5673 ), .B(\Reg_Bank/n5672 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5674 ) );
  MUX \Reg_Bank/U5761  ( .A(\Reg_Bank/registers[28][23] ), .B(
        \Reg_Bank/registers[29][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5673 )
         );
  MUX \Reg_Bank/U5760  ( .A(\Reg_Bank/registers[30][23] ), .B(
        \Reg_Bank/registers[31][23] ), .S(rt_index[0]), .Z(\Reg_Bank/n5672 )
         );
  MUX \Reg_Bank/U5759  ( .A(\Reg_Bank/n5671 ), .B(\Reg_Bank/n5656 ), .S(
        rt_index[4]), .Z(reg_target[22]) );
  MUX \Reg_Bank/U5758  ( .A(\Reg_Bank/n5670 ), .B(\Reg_Bank/n5663 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5671 ) );
  MUX \Reg_Bank/U5757  ( .A(\Reg_Bank/n5669 ), .B(\Reg_Bank/n5666 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5670 ) );
  MUX \Reg_Bank/U5756  ( .A(\Reg_Bank/n5668 ), .B(\Reg_Bank/n5667 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5669 ) );
  MUX \Reg_Bank/U5754  ( .A(\Reg_Bank/registers[2][22] ), .B(
        \Reg_Bank/registers[3][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5667 ) );
  MUX \Reg_Bank/U5753  ( .A(\Reg_Bank/n5665 ), .B(\Reg_Bank/n5664 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5666 ) );
  MUX \Reg_Bank/U5752  ( .A(\Reg_Bank/registers[4][22] ), .B(
        \Reg_Bank/registers[5][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5665 ) );
  MUX \Reg_Bank/U5751  ( .A(\Reg_Bank/registers[6][22] ), .B(
        \Reg_Bank/registers[7][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5664 ) );
  MUX \Reg_Bank/U5750  ( .A(\Reg_Bank/n5662 ), .B(\Reg_Bank/n5659 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5663 ) );
  MUX \Reg_Bank/U5749  ( .A(\Reg_Bank/n5661 ), .B(\Reg_Bank/n5660 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5662 ) );
  MUX \Reg_Bank/U5748  ( .A(\Reg_Bank/registers[8][22] ), .B(
        \Reg_Bank/registers[9][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5661 ) );
  MUX \Reg_Bank/U5747  ( .A(\Reg_Bank/registers[10][22] ), .B(
        \Reg_Bank/registers[11][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5660 )
         );
  MUX \Reg_Bank/U5746  ( .A(\Reg_Bank/n5658 ), .B(\Reg_Bank/n5657 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5659 ) );
  MUX \Reg_Bank/U5745  ( .A(\Reg_Bank/registers[12][22] ), .B(
        \Reg_Bank/registers[13][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5658 )
         );
  MUX \Reg_Bank/U5744  ( .A(\Reg_Bank/registers[14][22] ), .B(
        \Reg_Bank/registers[15][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5657 )
         );
  MUX \Reg_Bank/U5743  ( .A(\Reg_Bank/n5655 ), .B(\Reg_Bank/n5648 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5656 ) );
  MUX \Reg_Bank/U5742  ( .A(\Reg_Bank/n5654 ), .B(\Reg_Bank/n5651 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5655 ) );
  MUX \Reg_Bank/U5741  ( .A(\Reg_Bank/n5653 ), .B(\Reg_Bank/n5652 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5654 ) );
  MUX \Reg_Bank/U5740  ( .A(\Reg_Bank/registers[16][22] ), .B(
        \Reg_Bank/registers[17][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5653 )
         );
  MUX \Reg_Bank/U5739  ( .A(\Reg_Bank/registers[18][22] ), .B(
        \Reg_Bank/registers[19][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5652 )
         );
  MUX \Reg_Bank/U5738  ( .A(\Reg_Bank/n5650 ), .B(\Reg_Bank/n5649 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5651 ) );
  MUX \Reg_Bank/U5737  ( .A(\Reg_Bank/registers[20][22] ), .B(
        \Reg_Bank/registers[21][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5650 )
         );
  MUX \Reg_Bank/U5736  ( .A(\Reg_Bank/registers[22][22] ), .B(
        \Reg_Bank/registers[23][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5649 )
         );
  MUX \Reg_Bank/U5735  ( .A(\Reg_Bank/n5647 ), .B(\Reg_Bank/n5644 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5648 ) );
  MUX \Reg_Bank/U5734  ( .A(\Reg_Bank/n5646 ), .B(\Reg_Bank/n5645 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5647 ) );
  MUX \Reg_Bank/U5733  ( .A(\Reg_Bank/registers[24][22] ), .B(
        \Reg_Bank/registers[25][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5646 )
         );
  MUX \Reg_Bank/U5732  ( .A(\Reg_Bank/registers[26][22] ), .B(
        \Reg_Bank/registers[27][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5645 )
         );
  MUX \Reg_Bank/U5731  ( .A(\Reg_Bank/n5643 ), .B(\Reg_Bank/n5642 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5644 ) );
  MUX \Reg_Bank/U5730  ( .A(\Reg_Bank/registers[28][22] ), .B(
        \Reg_Bank/registers[29][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5643 )
         );
  MUX \Reg_Bank/U5729  ( .A(\Reg_Bank/registers[30][22] ), .B(
        \Reg_Bank/registers[31][22] ), .S(rt_index[0]), .Z(\Reg_Bank/n5642 )
         );
  MUX \Reg_Bank/U5728  ( .A(\Reg_Bank/n5641 ), .B(\Reg_Bank/n5626 ), .S(
        rt_index[4]), .Z(reg_target[21]) );
  MUX \Reg_Bank/U5727  ( .A(\Reg_Bank/n5640 ), .B(\Reg_Bank/n5633 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5641 ) );
  MUX \Reg_Bank/U5726  ( .A(\Reg_Bank/n5639 ), .B(\Reg_Bank/n5636 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5640 ) );
  MUX \Reg_Bank/U5725  ( .A(\Reg_Bank/n5638 ), .B(\Reg_Bank/n5637 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5639 ) );
  MUX \Reg_Bank/U5723  ( .A(\Reg_Bank/registers[2][21] ), .B(
        \Reg_Bank/registers[3][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5637 ) );
  MUX \Reg_Bank/U5722  ( .A(\Reg_Bank/n5635 ), .B(\Reg_Bank/n5634 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5636 ) );
  MUX \Reg_Bank/U5721  ( .A(\Reg_Bank/registers[4][21] ), .B(
        \Reg_Bank/registers[5][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5635 ) );
  MUX \Reg_Bank/U5720  ( .A(\Reg_Bank/registers[6][21] ), .B(
        \Reg_Bank/registers[7][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5634 ) );
  MUX \Reg_Bank/U5719  ( .A(\Reg_Bank/n5632 ), .B(\Reg_Bank/n5629 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5633 ) );
  MUX \Reg_Bank/U5718  ( .A(\Reg_Bank/n5631 ), .B(\Reg_Bank/n5630 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5632 ) );
  MUX \Reg_Bank/U5717  ( .A(\Reg_Bank/registers[8][21] ), .B(
        \Reg_Bank/registers[9][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5631 ) );
  MUX \Reg_Bank/U5716  ( .A(\Reg_Bank/registers[10][21] ), .B(
        \Reg_Bank/registers[11][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5630 )
         );
  MUX \Reg_Bank/U5715  ( .A(\Reg_Bank/n5628 ), .B(\Reg_Bank/n5627 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5629 ) );
  MUX \Reg_Bank/U5714  ( .A(\Reg_Bank/registers[12][21] ), .B(
        \Reg_Bank/registers[13][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5628 )
         );
  MUX \Reg_Bank/U5713  ( .A(\Reg_Bank/registers[14][21] ), .B(
        \Reg_Bank/registers[15][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5627 )
         );
  MUX \Reg_Bank/U5712  ( .A(\Reg_Bank/n5625 ), .B(\Reg_Bank/n5618 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5626 ) );
  MUX \Reg_Bank/U5711  ( .A(\Reg_Bank/n5624 ), .B(\Reg_Bank/n5621 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5625 ) );
  MUX \Reg_Bank/U5710  ( .A(\Reg_Bank/n5623 ), .B(\Reg_Bank/n5622 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5624 ) );
  MUX \Reg_Bank/U5709  ( .A(\Reg_Bank/registers[16][21] ), .B(
        \Reg_Bank/registers[17][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5623 )
         );
  MUX \Reg_Bank/U5708  ( .A(\Reg_Bank/registers[18][21] ), .B(
        \Reg_Bank/registers[19][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5622 )
         );
  MUX \Reg_Bank/U5707  ( .A(\Reg_Bank/n5620 ), .B(\Reg_Bank/n5619 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5621 ) );
  MUX \Reg_Bank/U5706  ( .A(\Reg_Bank/registers[20][21] ), .B(
        \Reg_Bank/registers[21][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5620 )
         );
  MUX \Reg_Bank/U5705  ( .A(\Reg_Bank/registers[22][21] ), .B(
        \Reg_Bank/registers[23][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5619 )
         );
  MUX \Reg_Bank/U5704  ( .A(\Reg_Bank/n5617 ), .B(\Reg_Bank/n5614 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5618 ) );
  MUX \Reg_Bank/U5703  ( .A(\Reg_Bank/n5616 ), .B(\Reg_Bank/n5615 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5617 ) );
  MUX \Reg_Bank/U5702  ( .A(\Reg_Bank/registers[24][21] ), .B(
        \Reg_Bank/registers[25][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5616 )
         );
  MUX \Reg_Bank/U5701  ( .A(\Reg_Bank/registers[26][21] ), .B(
        \Reg_Bank/registers[27][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5615 )
         );
  MUX \Reg_Bank/U5700  ( .A(\Reg_Bank/n5613 ), .B(\Reg_Bank/n5612 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5614 ) );
  MUX \Reg_Bank/U5699  ( .A(\Reg_Bank/registers[28][21] ), .B(
        \Reg_Bank/registers[29][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5613 )
         );
  MUX \Reg_Bank/U5698  ( .A(\Reg_Bank/registers[30][21] ), .B(
        \Reg_Bank/registers[31][21] ), .S(rt_index[0]), .Z(\Reg_Bank/n5612 )
         );
  MUX \Reg_Bank/U5697  ( .A(\Reg_Bank/n5611 ), .B(\Reg_Bank/n5596 ), .S(
        rt_index[4]), .Z(reg_target[20]) );
  MUX \Reg_Bank/U5696  ( .A(\Reg_Bank/n5610 ), .B(\Reg_Bank/n5603 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5611 ) );
  MUX \Reg_Bank/U5695  ( .A(\Reg_Bank/n5609 ), .B(\Reg_Bank/n5606 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5610 ) );
  MUX \Reg_Bank/U5694  ( .A(\Reg_Bank/n5608 ), .B(\Reg_Bank/n5607 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5609 ) );
  MUX \Reg_Bank/U5692  ( .A(\Reg_Bank/registers[2][20] ), .B(
        \Reg_Bank/registers[3][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5607 ) );
  MUX \Reg_Bank/U5691  ( .A(\Reg_Bank/n5605 ), .B(\Reg_Bank/n5604 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5606 ) );
  MUX \Reg_Bank/U5690  ( .A(\Reg_Bank/registers[4][20] ), .B(
        \Reg_Bank/registers[5][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5605 ) );
  MUX \Reg_Bank/U5689  ( .A(\Reg_Bank/registers[6][20] ), .B(
        \Reg_Bank/registers[7][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5604 ) );
  MUX \Reg_Bank/U5688  ( .A(\Reg_Bank/n5602 ), .B(\Reg_Bank/n5599 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5603 ) );
  MUX \Reg_Bank/U5687  ( .A(\Reg_Bank/n5601 ), .B(\Reg_Bank/n5600 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5602 ) );
  MUX \Reg_Bank/U5686  ( .A(\Reg_Bank/registers[8][20] ), .B(
        \Reg_Bank/registers[9][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5601 ) );
  MUX \Reg_Bank/U5685  ( .A(\Reg_Bank/registers[10][20] ), .B(
        \Reg_Bank/registers[11][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5600 )
         );
  MUX \Reg_Bank/U5684  ( .A(\Reg_Bank/n5598 ), .B(\Reg_Bank/n5597 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5599 ) );
  MUX \Reg_Bank/U5683  ( .A(\Reg_Bank/registers[12][20] ), .B(
        \Reg_Bank/registers[13][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5598 )
         );
  MUX \Reg_Bank/U5682  ( .A(\Reg_Bank/registers[14][20] ), .B(
        \Reg_Bank/registers[15][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5597 )
         );
  MUX \Reg_Bank/U5681  ( .A(\Reg_Bank/n5595 ), .B(\Reg_Bank/n5588 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5596 ) );
  MUX \Reg_Bank/U5680  ( .A(\Reg_Bank/n5594 ), .B(\Reg_Bank/n5591 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5595 ) );
  MUX \Reg_Bank/U5679  ( .A(\Reg_Bank/n5593 ), .B(\Reg_Bank/n5592 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5594 ) );
  MUX \Reg_Bank/U5678  ( .A(\Reg_Bank/registers[16][20] ), .B(
        \Reg_Bank/registers[17][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5593 )
         );
  MUX \Reg_Bank/U5677  ( .A(\Reg_Bank/registers[18][20] ), .B(
        \Reg_Bank/registers[19][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5592 )
         );
  MUX \Reg_Bank/U5676  ( .A(\Reg_Bank/n5590 ), .B(\Reg_Bank/n5589 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5591 ) );
  MUX \Reg_Bank/U5675  ( .A(\Reg_Bank/registers[20][20] ), .B(
        \Reg_Bank/registers[21][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5590 )
         );
  MUX \Reg_Bank/U5674  ( .A(\Reg_Bank/registers[22][20] ), .B(
        \Reg_Bank/registers[23][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5589 )
         );
  MUX \Reg_Bank/U5673  ( .A(\Reg_Bank/n5587 ), .B(\Reg_Bank/n5584 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5588 ) );
  MUX \Reg_Bank/U5672  ( .A(\Reg_Bank/n5586 ), .B(\Reg_Bank/n5585 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5587 ) );
  MUX \Reg_Bank/U5671  ( .A(\Reg_Bank/registers[24][20] ), .B(
        \Reg_Bank/registers[25][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5586 )
         );
  MUX \Reg_Bank/U5670  ( .A(\Reg_Bank/registers[26][20] ), .B(
        \Reg_Bank/registers[27][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5585 )
         );
  MUX \Reg_Bank/U5669  ( .A(\Reg_Bank/n5583 ), .B(\Reg_Bank/n5582 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5584 ) );
  MUX \Reg_Bank/U5668  ( .A(\Reg_Bank/registers[28][20] ), .B(
        \Reg_Bank/registers[29][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5583 )
         );
  MUX \Reg_Bank/U5667  ( .A(\Reg_Bank/registers[30][20] ), .B(
        \Reg_Bank/registers[31][20] ), .S(rt_index[0]), .Z(\Reg_Bank/n5582 )
         );
  MUX \Reg_Bank/U5666  ( .A(\Reg_Bank/n5581 ), .B(\Reg_Bank/n5566 ), .S(
        rt_index[4]), .Z(reg_target[19]) );
  MUX \Reg_Bank/U5665  ( .A(\Reg_Bank/n5580 ), .B(\Reg_Bank/n5573 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5581 ) );
  MUX \Reg_Bank/U5664  ( .A(\Reg_Bank/n5579 ), .B(\Reg_Bank/n5576 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5580 ) );
  MUX \Reg_Bank/U5663  ( .A(\Reg_Bank/n5578 ), .B(\Reg_Bank/n5577 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5579 ) );
  MUX \Reg_Bank/U5661  ( .A(\Reg_Bank/registers[2][19] ), .B(
        \Reg_Bank/registers[3][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5577 ) );
  MUX \Reg_Bank/U5660  ( .A(\Reg_Bank/n5575 ), .B(\Reg_Bank/n5574 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5576 ) );
  MUX \Reg_Bank/U5659  ( .A(\Reg_Bank/registers[4][19] ), .B(
        \Reg_Bank/registers[5][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5575 ) );
  MUX \Reg_Bank/U5658  ( .A(\Reg_Bank/registers[6][19] ), .B(
        \Reg_Bank/registers[7][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5574 ) );
  MUX \Reg_Bank/U5657  ( .A(\Reg_Bank/n5572 ), .B(\Reg_Bank/n5569 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5573 ) );
  MUX \Reg_Bank/U5656  ( .A(\Reg_Bank/n5571 ), .B(\Reg_Bank/n5570 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5572 ) );
  MUX \Reg_Bank/U5655  ( .A(\Reg_Bank/registers[8][19] ), .B(
        \Reg_Bank/registers[9][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5571 ) );
  MUX \Reg_Bank/U5654  ( .A(\Reg_Bank/registers[10][19] ), .B(
        \Reg_Bank/registers[11][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5570 )
         );
  MUX \Reg_Bank/U5653  ( .A(\Reg_Bank/n5568 ), .B(\Reg_Bank/n5567 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5569 ) );
  MUX \Reg_Bank/U5652  ( .A(\Reg_Bank/registers[12][19] ), .B(
        \Reg_Bank/registers[13][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5568 )
         );
  MUX \Reg_Bank/U5651  ( .A(\Reg_Bank/registers[14][19] ), .B(
        \Reg_Bank/registers[15][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5567 )
         );
  MUX \Reg_Bank/U5650  ( .A(\Reg_Bank/n5565 ), .B(\Reg_Bank/n5558 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5566 ) );
  MUX \Reg_Bank/U5649  ( .A(\Reg_Bank/n5564 ), .B(\Reg_Bank/n5561 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5565 ) );
  MUX \Reg_Bank/U5648  ( .A(\Reg_Bank/n5563 ), .B(\Reg_Bank/n5562 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5564 ) );
  MUX \Reg_Bank/U5647  ( .A(\Reg_Bank/registers[16][19] ), .B(
        \Reg_Bank/registers[17][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5563 )
         );
  MUX \Reg_Bank/U5646  ( .A(\Reg_Bank/registers[18][19] ), .B(
        \Reg_Bank/registers[19][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5562 )
         );
  MUX \Reg_Bank/U5645  ( .A(\Reg_Bank/n5560 ), .B(\Reg_Bank/n5559 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5561 ) );
  MUX \Reg_Bank/U5644  ( .A(\Reg_Bank/registers[20][19] ), .B(
        \Reg_Bank/registers[21][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5560 )
         );
  MUX \Reg_Bank/U5643  ( .A(\Reg_Bank/registers[22][19] ), .B(
        \Reg_Bank/registers[23][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5559 )
         );
  MUX \Reg_Bank/U5642  ( .A(\Reg_Bank/n5557 ), .B(\Reg_Bank/n5554 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5558 ) );
  MUX \Reg_Bank/U5641  ( .A(\Reg_Bank/n5556 ), .B(\Reg_Bank/n5555 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5557 ) );
  MUX \Reg_Bank/U5640  ( .A(\Reg_Bank/registers[24][19] ), .B(
        \Reg_Bank/registers[25][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5556 )
         );
  MUX \Reg_Bank/U5639  ( .A(\Reg_Bank/registers[26][19] ), .B(
        \Reg_Bank/registers[27][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5555 )
         );
  MUX \Reg_Bank/U5638  ( .A(\Reg_Bank/n5553 ), .B(\Reg_Bank/n5552 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5554 ) );
  MUX \Reg_Bank/U5637  ( .A(\Reg_Bank/registers[28][19] ), .B(
        \Reg_Bank/registers[29][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5553 )
         );
  MUX \Reg_Bank/U5636  ( .A(\Reg_Bank/registers[30][19] ), .B(
        \Reg_Bank/registers[31][19] ), .S(rt_index[0]), .Z(\Reg_Bank/n5552 )
         );
  MUX \Reg_Bank/U5635  ( .A(\Reg_Bank/n5551 ), .B(\Reg_Bank/n5536 ), .S(
        rt_index[4]), .Z(reg_target[18]) );
  MUX \Reg_Bank/U5634  ( .A(\Reg_Bank/n5550 ), .B(\Reg_Bank/n5543 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5551 ) );
  MUX \Reg_Bank/U5633  ( .A(\Reg_Bank/n5549 ), .B(\Reg_Bank/n5546 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5550 ) );
  MUX \Reg_Bank/U5632  ( .A(\Reg_Bank/n5548 ), .B(\Reg_Bank/n5547 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5549 ) );
  MUX \Reg_Bank/U5630  ( .A(\Reg_Bank/registers[2][18] ), .B(
        \Reg_Bank/registers[3][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5547 ) );
  MUX \Reg_Bank/U5629  ( .A(\Reg_Bank/n5545 ), .B(\Reg_Bank/n5544 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5546 ) );
  MUX \Reg_Bank/U5628  ( .A(\Reg_Bank/registers[4][18] ), .B(
        \Reg_Bank/registers[5][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5545 ) );
  MUX \Reg_Bank/U5627  ( .A(\Reg_Bank/registers[6][18] ), .B(
        \Reg_Bank/registers[7][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5544 ) );
  MUX \Reg_Bank/U5626  ( .A(\Reg_Bank/n5542 ), .B(\Reg_Bank/n5539 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5543 ) );
  MUX \Reg_Bank/U5625  ( .A(\Reg_Bank/n5541 ), .B(\Reg_Bank/n5540 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5542 ) );
  MUX \Reg_Bank/U5624  ( .A(\Reg_Bank/registers[8][18] ), .B(
        \Reg_Bank/registers[9][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5541 ) );
  MUX \Reg_Bank/U5623  ( .A(\Reg_Bank/registers[10][18] ), .B(
        \Reg_Bank/registers[11][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5540 )
         );
  MUX \Reg_Bank/U5622  ( .A(\Reg_Bank/n5538 ), .B(\Reg_Bank/n5537 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5539 ) );
  MUX \Reg_Bank/U5621  ( .A(\Reg_Bank/registers[12][18] ), .B(
        \Reg_Bank/registers[13][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5538 )
         );
  MUX \Reg_Bank/U5620  ( .A(\Reg_Bank/registers[14][18] ), .B(
        \Reg_Bank/registers[15][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5537 )
         );
  MUX \Reg_Bank/U5619  ( .A(\Reg_Bank/n5535 ), .B(\Reg_Bank/n5528 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5536 ) );
  MUX \Reg_Bank/U5618  ( .A(\Reg_Bank/n5534 ), .B(\Reg_Bank/n5531 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5535 ) );
  MUX \Reg_Bank/U5617  ( .A(\Reg_Bank/n5533 ), .B(\Reg_Bank/n5532 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5534 ) );
  MUX \Reg_Bank/U5616  ( .A(\Reg_Bank/registers[16][18] ), .B(
        \Reg_Bank/registers[17][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5533 )
         );
  MUX \Reg_Bank/U5615  ( .A(\Reg_Bank/registers[18][18] ), .B(
        \Reg_Bank/registers[19][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5532 )
         );
  MUX \Reg_Bank/U5614  ( .A(\Reg_Bank/n5530 ), .B(\Reg_Bank/n5529 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5531 ) );
  MUX \Reg_Bank/U5613  ( .A(\Reg_Bank/registers[20][18] ), .B(
        \Reg_Bank/registers[21][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5530 )
         );
  MUX \Reg_Bank/U5612  ( .A(\Reg_Bank/registers[22][18] ), .B(
        \Reg_Bank/registers[23][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5529 )
         );
  MUX \Reg_Bank/U5611  ( .A(\Reg_Bank/n5527 ), .B(\Reg_Bank/n5524 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5528 ) );
  MUX \Reg_Bank/U5610  ( .A(\Reg_Bank/n5526 ), .B(\Reg_Bank/n5525 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5527 ) );
  MUX \Reg_Bank/U5609  ( .A(\Reg_Bank/registers[24][18] ), .B(
        \Reg_Bank/registers[25][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5526 )
         );
  MUX \Reg_Bank/U5608  ( .A(\Reg_Bank/registers[26][18] ), .B(
        \Reg_Bank/registers[27][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5525 )
         );
  MUX \Reg_Bank/U5607  ( .A(\Reg_Bank/n5523 ), .B(\Reg_Bank/n5522 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5524 ) );
  MUX \Reg_Bank/U5606  ( .A(\Reg_Bank/registers[28][18] ), .B(
        \Reg_Bank/registers[29][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5523 )
         );
  MUX \Reg_Bank/U5605  ( .A(\Reg_Bank/registers[30][18] ), .B(
        \Reg_Bank/registers[31][18] ), .S(rt_index[0]), .Z(\Reg_Bank/n5522 )
         );
  MUX \Reg_Bank/U5604  ( .A(\Reg_Bank/n5521 ), .B(\Reg_Bank/n5506 ), .S(
        rt_index[4]), .Z(reg_target[17]) );
  MUX \Reg_Bank/U5603  ( .A(\Reg_Bank/n5520 ), .B(\Reg_Bank/n5513 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5521 ) );
  MUX \Reg_Bank/U5602  ( .A(\Reg_Bank/n5519 ), .B(\Reg_Bank/n5516 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5520 ) );
  MUX \Reg_Bank/U5601  ( .A(\Reg_Bank/n5518 ), .B(\Reg_Bank/n5517 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5519 ) );
  MUX \Reg_Bank/U5599  ( .A(\Reg_Bank/registers[2][17] ), .B(
        \Reg_Bank/registers[3][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5517 ) );
  MUX \Reg_Bank/U5598  ( .A(\Reg_Bank/n5515 ), .B(\Reg_Bank/n5514 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5516 ) );
  MUX \Reg_Bank/U5597  ( .A(\Reg_Bank/registers[4][17] ), .B(
        \Reg_Bank/registers[5][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5515 ) );
  MUX \Reg_Bank/U5596  ( .A(\Reg_Bank/registers[6][17] ), .B(
        \Reg_Bank/registers[7][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5514 ) );
  MUX \Reg_Bank/U5595  ( .A(\Reg_Bank/n5512 ), .B(\Reg_Bank/n5509 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5513 ) );
  MUX \Reg_Bank/U5594  ( .A(\Reg_Bank/n5511 ), .B(\Reg_Bank/n5510 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5512 ) );
  MUX \Reg_Bank/U5593  ( .A(\Reg_Bank/registers[8][17] ), .B(
        \Reg_Bank/registers[9][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5511 ) );
  MUX \Reg_Bank/U5592  ( .A(\Reg_Bank/registers[10][17] ), .B(
        \Reg_Bank/registers[11][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5510 )
         );
  MUX \Reg_Bank/U5591  ( .A(\Reg_Bank/n5508 ), .B(\Reg_Bank/n5507 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5509 ) );
  MUX \Reg_Bank/U5590  ( .A(\Reg_Bank/registers[12][17] ), .B(
        \Reg_Bank/registers[13][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5508 )
         );
  MUX \Reg_Bank/U5589  ( .A(\Reg_Bank/registers[14][17] ), .B(
        \Reg_Bank/registers[15][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5507 )
         );
  MUX \Reg_Bank/U5588  ( .A(\Reg_Bank/n5505 ), .B(\Reg_Bank/n5498 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5506 ) );
  MUX \Reg_Bank/U5587  ( .A(\Reg_Bank/n5504 ), .B(\Reg_Bank/n5501 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5505 ) );
  MUX \Reg_Bank/U5586  ( .A(\Reg_Bank/n5503 ), .B(\Reg_Bank/n5502 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5504 ) );
  MUX \Reg_Bank/U5585  ( .A(\Reg_Bank/registers[16][17] ), .B(
        \Reg_Bank/registers[17][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5503 )
         );
  MUX \Reg_Bank/U5584  ( .A(\Reg_Bank/registers[18][17] ), .B(
        \Reg_Bank/registers[19][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5502 )
         );
  MUX \Reg_Bank/U5583  ( .A(\Reg_Bank/n5500 ), .B(\Reg_Bank/n5499 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5501 ) );
  MUX \Reg_Bank/U5582  ( .A(\Reg_Bank/registers[20][17] ), .B(
        \Reg_Bank/registers[21][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5500 )
         );
  MUX \Reg_Bank/U5581  ( .A(\Reg_Bank/registers[22][17] ), .B(
        \Reg_Bank/registers[23][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5499 )
         );
  MUX \Reg_Bank/U5580  ( .A(\Reg_Bank/n5497 ), .B(\Reg_Bank/n5494 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5498 ) );
  MUX \Reg_Bank/U5579  ( .A(\Reg_Bank/n5496 ), .B(\Reg_Bank/n5495 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5497 ) );
  MUX \Reg_Bank/U5578  ( .A(\Reg_Bank/registers[24][17] ), .B(
        \Reg_Bank/registers[25][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5496 )
         );
  MUX \Reg_Bank/U5577  ( .A(\Reg_Bank/registers[26][17] ), .B(
        \Reg_Bank/registers[27][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5495 )
         );
  MUX \Reg_Bank/U5576  ( .A(\Reg_Bank/n5493 ), .B(\Reg_Bank/n5492 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5494 ) );
  MUX \Reg_Bank/U5575  ( .A(\Reg_Bank/registers[28][17] ), .B(
        \Reg_Bank/registers[29][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5493 )
         );
  MUX \Reg_Bank/U5574  ( .A(\Reg_Bank/registers[30][17] ), .B(
        \Reg_Bank/registers[31][17] ), .S(rt_index[0]), .Z(\Reg_Bank/n5492 )
         );
  MUX \Reg_Bank/U5573  ( .A(\Reg_Bank/n5491 ), .B(\Reg_Bank/n5476 ), .S(
        rt_index[4]), .Z(reg_target[16]) );
  MUX \Reg_Bank/U5572  ( .A(\Reg_Bank/n5490 ), .B(\Reg_Bank/n5483 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5491 ) );
  MUX \Reg_Bank/U5571  ( .A(\Reg_Bank/n5489 ), .B(\Reg_Bank/n5486 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5490 ) );
  MUX \Reg_Bank/U5570  ( .A(\Reg_Bank/n5488 ), .B(\Reg_Bank/n5487 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5489 ) );
  MUX \Reg_Bank/U5568  ( .A(\Reg_Bank/registers[2][16] ), .B(
        \Reg_Bank/registers[3][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5487 ) );
  MUX \Reg_Bank/U5567  ( .A(\Reg_Bank/n5485 ), .B(\Reg_Bank/n5484 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5486 ) );
  MUX \Reg_Bank/U5566  ( .A(\Reg_Bank/registers[4][16] ), .B(
        \Reg_Bank/registers[5][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5485 ) );
  MUX \Reg_Bank/U5565  ( .A(\Reg_Bank/registers[6][16] ), .B(
        \Reg_Bank/registers[7][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5484 ) );
  MUX \Reg_Bank/U5564  ( .A(\Reg_Bank/n5482 ), .B(\Reg_Bank/n5479 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5483 ) );
  MUX \Reg_Bank/U5563  ( .A(\Reg_Bank/n5481 ), .B(\Reg_Bank/n5480 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5482 ) );
  MUX \Reg_Bank/U5562  ( .A(\Reg_Bank/registers[8][16] ), .B(
        \Reg_Bank/registers[9][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5481 ) );
  MUX \Reg_Bank/U5561  ( .A(\Reg_Bank/registers[10][16] ), .B(
        \Reg_Bank/registers[11][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5480 )
         );
  MUX \Reg_Bank/U5560  ( .A(\Reg_Bank/n5478 ), .B(\Reg_Bank/n5477 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5479 ) );
  MUX \Reg_Bank/U5559  ( .A(\Reg_Bank/registers[12][16] ), .B(
        \Reg_Bank/registers[13][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5478 )
         );
  MUX \Reg_Bank/U5558  ( .A(\Reg_Bank/registers[14][16] ), .B(
        \Reg_Bank/registers[15][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5477 )
         );
  MUX \Reg_Bank/U5557  ( .A(\Reg_Bank/n5475 ), .B(\Reg_Bank/n5468 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5476 ) );
  MUX \Reg_Bank/U5556  ( .A(\Reg_Bank/n5474 ), .B(\Reg_Bank/n5471 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5475 ) );
  MUX \Reg_Bank/U5555  ( .A(\Reg_Bank/n5473 ), .B(\Reg_Bank/n5472 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5474 ) );
  MUX \Reg_Bank/U5554  ( .A(\Reg_Bank/registers[16][16] ), .B(
        \Reg_Bank/registers[17][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5473 )
         );
  MUX \Reg_Bank/U5553  ( .A(\Reg_Bank/registers[18][16] ), .B(
        \Reg_Bank/registers[19][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5472 )
         );
  MUX \Reg_Bank/U5552  ( .A(\Reg_Bank/n5470 ), .B(\Reg_Bank/n5469 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5471 ) );
  MUX \Reg_Bank/U5551  ( .A(\Reg_Bank/registers[20][16] ), .B(
        \Reg_Bank/registers[21][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5470 )
         );
  MUX \Reg_Bank/U5550  ( .A(\Reg_Bank/registers[22][16] ), .B(
        \Reg_Bank/registers[23][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5469 )
         );
  MUX \Reg_Bank/U5549  ( .A(\Reg_Bank/n5467 ), .B(\Reg_Bank/n5464 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5468 ) );
  MUX \Reg_Bank/U5548  ( .A(\Reg_Bank/n5466 ), .B(\Reg_Bank/n5465 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5467 ) );
  MUX \Reg_Bank/U5547  ( .A(\Reg_Bank/registers[24][16] ), .B(
        \Reg_Bank/registers[25][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5466 )
         );
  MUX \Reg_Bank/U5546  ( .A(\Reg_Bank/registers[26][16] ), .B(
        \Reg_Bank/registers[27][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5465 )
         );
  MUX \Reg_Bank/U5545  ( .A(\Reg_Bank/n5463 ), .B(\Reg_Bank/n5462 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5464 ) );
  MUX \Reg_Bank/U5544  ( .A(\Reg_Bank/registers[28][16] ), .B(
        \Reg_Bank/registers[29][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5463 )
         );
  MUX \Reg_Bank/U5543  ( .A(\Reg_Bank/registers[30][16] ), .B(
        \Reg_Bank/registers[31][16] ), .S(rt_index[0]), .Z(\Reg_Bank/n5462 )
         );
  MUX \Reg_Bank/U5542  ( .A(\Reg_Bank/n5461 ), .B(\Reg_Bank/n5446 ), .S(
        rt_index[4]), .Z(reg_target[15]) );
  MUX \Reg_Bank/U5541  ( .A(\Reg_Bank/n5460 ), .B(\Reg_Bank/n5453 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5461 ) );
  MUX \Reg_Bank/U5540  ( .A(\Reg_Bank/n5459 ), .B(\Reg_Bank/n5456 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5460 ) );
  MUX \Reg_Bank/U5539  ( .A(\Reg_Bank/n5458 ), .B(\Reg_Bank/n5457 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5459 ) );
  MUX \Reg_Bank/U5537  ( .A(\Reg_Bank/registers[2][15] ), .B(
        \Reg_Bank/registers[3][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5457 ) );
  MUX \Reg_Bank/U5536  ( .A(\Reg_Bank/n5455 ), .B(\Reg_Bank/n5454 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5456 ) );
  MUX \Reg_Bank/U5535  ( .A(\Reg_Bank/registers[4][15] ), .B(
        \Reg_Bank/registers[5][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5455 ) );
  MUX \Reg_Bank/U5534  ( .A(\Reg_Bank/registers[6][15] ), .B(
        \Reg_Bank/registers[7][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5454 ) );
  MUX \Reg_Bank/U5533  ( .A(\Reg_Bank/n5452 ), .B(\Reg_Bank/n5449 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5453 ) );
  MUX \Reg_Bank/U5532  ( .A(\Reg_Bank/n5451 ), .B(\Reg_Bank/n5450 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5452 ) );
  MUX \Reg_Bank/U5531  ( .A(\Reg_Bank/registers[8][15] ), .B(
        \Reg_Bank/registers[9][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5451 ) );
  MUX \Reg_Bank/U5530  ( .A(\Reg_Bank/registers[10][15] ), .B(
        \Reg_Bank/registers[11][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5450 )
         );
  MUX \Reg_Bank/U5529  ( .A(\Reg_Bank/n5448 ), .B(\Reg_Bank/n5447 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5449 ) );
  MUX \Reg_Bank/U5528  ( .A(\Reg_Bank/registers[12][15] ), .B(
        \Reg_Bank/registers[13][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5448 )
         );
  MUX \Reg_Bank/U5527  ( .A(\Reg_Bank/registers[14][15] ), .B(
        \Reg_Bank/registers[15][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5447 )
         );
  MUX \Reg_Bank/U5526  ( .A(\Reg_Bank/n5445 ), .B(\Reg_Bank/n5438 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5446 ) );
  MUX \Reg_Bank/U5525  ( .A(\Reg_Bank/n5444 ), .B(\Reg_Bank/n5441 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5445 ) );
  MUX \Reg_Bank/U5524  ( .A(\Reg_Bank/n5443 ), .B(\Reg_Bank/n5442 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5444 ) );
  MUX \Reg_Bank/U5523  ( .A(\Reg_Bank/registers[16][15] ), .B(
        \Reg_Bank/registers[17][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5443 )
         );
  MUX \Reg_Bank/U5522  ( .A(\Reg_Bank/registers[18][15] ), .B(
        \Reg_Bank/registers[19][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5442 )
         );
  MUX \Reg_Bank/U5521  ( .A(\Reg_Bank/n5440 ), .B(\Reg_Bank/n5439 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5441 ) );
  MUX \Reg_Bank/U5520  ( .A(\Reg_Bank/registers[20][15] ), .B(
        \Reg_Bank/registers[21][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5440 )
         );
  MUX \Reg_Bank/U5519  ( .A(\Reg_Bank/registers[22][15] ), .B(
        \Reg_Bank/registers[23][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5439 )
         );
  MUX \Reg_Bank/U5518  ( .A(\Reg_Bank/n5437 ), .B(\Reg_Bank/n5434 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5438 ) );
  MUX \Reg_Bank/U5517  ( .A(\Reg_Bank/n5436 ), .B(\Reg_Bank/n5435 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5437 ) );
  MUX \Reg_Bank/U5516  ( .A(\Reg_Bank/registers[24][15] ), .B(
        \Reg_Bank/registers[25][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5436 )
         );
  MUX \Reg_Bank/U5515  ( .A(\Reg_Bank/registers[26][15] ), .B(
        \Reg_Bank/registers[27][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5435 )
         );
  MUX \Reg_Bank/U5514  ( .A(\Reg_Bank/n5433 ), .B(\Reg_Bank/n5432 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5434 ) );
  MUX \Reg_Bank/U5513  ( .A(\Reg_Bank/registers[28][15] ), .B(
        \Reg_Bank/registers[29][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5433 )
         );
  MUX \Reg_Bank/U5512  ( .A(\Reg_Bank/registers[30][15] ), .B(
        \Reg_Bank/registers[31][15] ), .S(rt_index[0]), .Z(\Reg_Bank/n5432 )
         );
  MUX \Reg_Bank/U5511  ( .A(\Reg_Bank/n5431 ), .B(\Reg_Bank/n5416 ), .S(
        rt_index[4]), .Z(reg_target[14]) );
  MUX \Reg_Bank/U5510  ( .A(\Reg_Bank/n5430 ), .B(\Reg_Bank/n5423 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5431 ) );
  MUX \Reg_Bank/U5509  ( .A(\Reg_Bank/n5429 ), .B(\Reg_Bank/n5426 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5430 ) );
  MUX \Reg_Bank/U5508  ( .A(\Reg_Bank/n5428 ), .B(\Reg_Bank/n5427 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5429 ) );
  MUX \Reg_Bank/U5506  ( .A(\Reg_Bank/registers[2][14] ), .B(
        \Reg_Bank/registers[3][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5427 ) );
  MUX \Reg_Bank/U5505  ( .A(\Reg_Bank/n5425 ), .B(\Reg_Bank/n5424 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5426 ) );
  MUX \Reg_Bank/U5504  ( .A(\Reg_Bank/registers[4][14] ), .B(
        \Reg_Bank/registers[5][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5425 ) );
  MUX \Reg_Bank/U5503  ( .A(\Reg_Bank/registers[6][14] ), .B(
        \Reg_Bank/registers[7][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5424 ) );
  MUX \Reg_Bank/U5502  ( .A(\Reg_Bank/n5422 ), .B(\Reg_Bank/n5419 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5423 ) );
  MUX \Reg_Bank/U5501  ( .A(\Reg_Bank/n5421 ), .B(\Reg_Bank/n5420 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5422 ) );
  MUX \Reg_Bank/U5500  ( .A(\Reg_Bank/registers[8][14] ), .B(
        \Reg_Bank/registers[9][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5421 ) );
  MUX \Reg_Bank/U5499  ( .A(\Reg_Bank/registers[10][14] ), .B(
        \Reg_Bank/registers[11][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5420 )
         );
  MUX \Reg_Bank/U5498  ( .A(\Reg_Bank/n5418 ), .B(\Reg_Bank/n5417 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5419 ) );
  MUX \Reg_Bank/U5497  ( .A(\Reg_Bank/registers[12][14] ), .B(
        \Reg_Bank/registers[13][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5418 )
         );
  MUX \Reg_Bank/U5496  ( .A(\Reg_Bank/registers[14][14] ), .B(
        \Reg_Bank/registers[15][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5417 )
         );
  MUX \Reg_Bank/U5495  ( .A(\Reg_Bank/n5415 ), .B(\Reg_Bank/n5408 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5416 ) );
  MUX \Reg_Bank/U5494  ( .A(\Reg_Bank/n5414 ), .B(\Reg_Bank/n5411 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5415 ) );
  MUX \Reg_Bank/U5493  ( .A(\Reg_Bank/n5413 ), .B(\Reg_Bank/n5412 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5414 ) );
  MUX \Reg_Bank/U5492  ( .A(\Reg_Bank/registers[16][14] ), .B(
        \Reg_Bank/registers[17][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5413 )
         );
  MUX \Reg_Bank/U5491  ( .A(\Reg_Bank/registers[18][14] ), .B(
        \Reg_Bank/registers[19][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5412 )
         );
  MUX \Reg_Bank/U5490  ( .A(\Reg_Bank/n5410 ), .B(\Reg_Bank/n5409 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5411 ) );
  MUX \Reg_Bank/U5489  ( .A(\Reg_Bank/registers[20][14] ), .B(
        \Reg_Bank/registers[21][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5410 )
         );
  MUX \Reg_Bank/U5488  ( .A(\Reg_Bank/registers[22][14] ), .B(
        \Reg_Bank/registers[23][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5409 )
         );
  MUX \Reg_Bank/U5487  ( .A(\Reg_Bank/n5407 ), .B(\Reg_Bank/n5404 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5408 ) );
  MUX \Reg_Bank/U5486  ( .A(\Reg_Bank/n5406 ), .B(\Reg_Bank/n5405 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5407 ) );
  MUX \Reg_Bank/U5485  ( .A(\Reg_Bank/registers[24][14] ), .B(
        \Reg_Bank/registers[25][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5406 )
         );
  MUX \Reg_Bank/U5484  ( .A(\Reg_Bank/registers[26][14] ), .B(
        \Reg_Bank/registers[27][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5405 )
         );
  MUX \Reg_Bank/U5483  ( .A(\Reg_Bank/n5403 ), .B(\Reg_Bank/n5402 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5404 ) );
  MUX \Reg_Bank/U5482  ( .A(\Reg_Bank/registers[28][14] ), .B(
        \Reg_Bank/registers[29][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5403 )
         );
  MUX \Reg_Bank/U5481  ( .A(\Reg_Bank/registers[30][14] ), .B(
        \Reg_Bank/registers[31][14] ), .S(rt_index[0]), .Z(\Reg_Bank/n5402 )
         );
  MUX \Reg_Bank/U5480  ( .A(\Reg_Bank/n5401 ), .B(\Reg_Bank/n5386 ), .S(
        rt_index[4]), .Z(reg_target[13]) );
  MUX \Reg_Bank/U5479  ( .A(\Reg_Bank/n5400 ), .B(\Reg_Bank/n5393 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5401 ) );
  MUX \Reg_Bank/U5478  ( .A(\Reg_Bank/n5399 ), .B(\Reg_Bank/n5396 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5400 ) );
  MUX \Reg_Bank/U5477  ( .A(\Reg_Bank/n5398 ), .B(\Reg_Bank/n5397 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5399 ) );
  MUX \Reg_Bank/U5475  ( .A(\Reg_Bank/registers[2][13] ), .B(
        \Reg_Bank/registers[3][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5397 ) );
  MUX \Reg_Bank/U5474  ( .A(\Reg_Bank/n5395 ), .B(\Reg_Bank/n5394 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5396 ) );
  MUX \Reg_Bank/U5473  ( .A(\Reg_Bank/registers[4][13] ), .B(
        \Reg_Bank/registers[5][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5395 ) );
  MUX \Reg_Bank/U5472  ( .A(\Reg_Bank/registers[6][13] ), .B(
        \Reg_Bank/registers[7][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5394 ) );
  MUX \Reg_Bank/U5471  ( .A(\Reg_Bank/n5392 ), .B(\Reg_Bank/n5389 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5393 ) );
  MUX \Reg_Bank/U5470  ( .A(\Reg_Bank/n5391 ), .B(\Reg_Bank/n5390 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5392 ) );
  MUX \Reg_Bank/U5469  ( .A(\Reg_Bank/registers[8][13] ), .B(
        \Reg_Bank/registers[9][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5391 ) );
  MUX \Reg_Bank/U5468  ( .A(\Reg_Bank/registers[10][13] ), .B(
        \Reg_Bank/registers[11][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5390 )
         );
  MUX \Reg_Bank/U5467  ( .A(\Reg_Bank/n5388 ), .B(\Reg_Bank/n5387 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5389 ) );
  MUX \Reg_Bank/U5466  ( .A(\Reg_Bank/registers[12][13] ), .B(
        \Reg_Bank/registers[13][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5388 )
         );
  MUX \Reg_Bank/U5465  ( .A(\Reg_Bank/registers[14][13] ), .B(
        \Reg_Bank/registers[15][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5387 )
         );
  MUX \Reg_Bank/U5464  ( .A(\Reg_Bank/n5385 ), .B(\Reg_Bank/n5378 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5386 ) );
  MUX \Reg_Bank/U5463  ( .A(\Reg_Bank/n5384 ), .B(\Reg_Bank/n5381 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5385 ) );
  MUX \Reg_Bank/U5462  ( .A(\Reg_Bank/n5383 ), .B(\Reg_Bank/n5382 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5384 ) );
  MUX \Reg_Bank/U5461  ( .A(\Reg_Bank/registers[16][13] ), .B(
        \Reg_Bank/registers[17][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5383 )
         );
  MUX \Reg_Bank/U5460  ( .A(\Reg_Bank/registers[18][13] ), .B(
        \Reg_Bank/registers[19][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5382 )
         );
  MUX \Reg_Bank/U5459  ( .A(\Reg_Bank/n5380 ), .B(\Reg_Bank/n5379 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5381 ) );
  MUX \Reg_Bank/U5458  ( .A(\Reg_Bank/registers[20][13] ), .B(
        \Reg_Bank/registers[21][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5380 )
         );
  MUX \Reg_Bank/U5457  ( .A(\Reg_Bank/registers[22][13] ), .B(
        \Reg_Bank/registers[23][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5379 )
         );
  MUX \Reg_Bank/U5456  ( .A(\Reg_Bank/n5377 ), .B(\Reg_Bank/n5374 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5378 ) );
  MUX \Reg_Bank/U5455  ( .A(\Reg_Bank/n5376 ), .B(\Reg_Bank/n5375 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5377 ) );
  MUX \Reg_Bank/U5454  ( .A(\Reg_Bank/registers[24][13] ), .B(
        \Reg_Bank/registers[25][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5376 )
         );
  MUX \Reg_Bank/U5453  ( .A(\Reg_Bank/registers[26][13] ), .B(
        \Reg_Bank/registers[27][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5375 )
         );
  MUX \Reg_Bank/U5452  ( .A(\Reg_Bank/n5373 ), .B(\Reg_Bank/n5372 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5374 ) );
  MUX \Reg_Bank/U5451  ( .A(\Reg_Bank/registers[28][13] ), .B(
        \Reg_Bank/registers[29][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5373 )
         );
  MUX \Reg_Bank/U5450  ( .A(\Reg_Bank/registers[30][13] ), .B(
        \Reg_Bank/registers[31][13] ), .S(rt_index[0]), .Z(\Reg_Bank/n5372 )
         );
  MUX \Reg_Bank/U5449  ( .A(\Reg_Bank/n5371 ), .B(\Reg_Bank/n5356 ), .S(
        rt_index[4]), .Z(reg_target[12]) );
  MUX \Reg_Bank/U5448  ( .A(\Reg_Bank/n5370 ), .B(\Reg_Bank/n5363 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5371 ) );
  MUX \Reg_Bank/U5447  ( .A(\Reg_Bank/n5369 ), .B(\Reg_Bank/n5366 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5370 ) );
  MUX \Reg_Bank/U5446  ( .A(\Reg_Bank/n5368 ), .B(\Reg_Bank/n5367 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5369 ) );
  MUX \Reg_Bank/U5444  ( .A(\Reg_Bank/registers[2][12] ), .B(
        \Reg_Bank/registers[3][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5367 ) );
  MUX \Reg_Bank/U5443  ( .A(\Reg_Bank/n5365 ), .B(\Reg_Bank/n5364 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5366 ) );
  MUX \Reg_Bank/U5442  ( .A(\Reg_Bank/registers[4][12] ), .B(
        \Reg_Bank/registers[5][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5365 ) );
  MUX \Reg_Bank/U5441  ( .A(\Reg_Bank/registers[6][12] ), .B(
        \Reg_Bank/registers[7][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5364 ) );
  MUX \Reg_Bank/U5440  ( .A(\Reg_Bank/n5362 ), .B(\Reg_Bank/n5359 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5363 ) );
  MUX \Reg_Bank/U5439  ( .A(\Reg_Bank/n5361 ), .B(\Reg_Bank/n5360 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5362 ) );
  MUX \Reg_Bank/U5438  ( .A(\Reg_Bank/registers[8][12] ), .B(
        \Reg_Bank/registers[9][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5361 ) );
  MUX \Reg_Bank/U5437  ( .A(\Reg_Bank/registers[10][12] ), .B(
        \Reg_Bank/registers[11][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5360 )
         );
  MUX \Reg_Bank/U5436  ( .A(\Reg_Bank/n5358 ), .B(\Reg_Bank/n5357 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5359 ) );
  MUX \Reg_Bank/U5435  ( .A(\Reg_Bank/registers[12][12] ), .B(
        \Reg_Bank/registers[13][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5358 )
         );
  MUX \Reg_Bank/U5434  ( .A(\Reg_Bank/registers[14][12] ), .B(
        \Reg_Bank/registers[15][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5357 )
         );
  MUX \Reg_Bank/U5433  ( .A(\Reg_Bank/n5355 ), .B(\Reg_Bank/n5348 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5356 ) );
  MUX \Reg_Bank/U5432  ( .A(\Reg_Bank/n5354 ), .B(\Reg_Bank/n5351 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5355 ) );
  MUX \Reg_Bank/U5431  ( .A(\Reg_Bank/n5353 ), .B(\Reg_Bank/n5352 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5354 ) );
  MUX \Reg_Bank/U5430  ( .A(\Reg_Bank/registers[16][12] ), .B(
        \Reg_Bank/registers[17][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5353 )
         );
  MUX \Reg_Bank/U5429  ( .A(\Reg_Bank/registers[18][12] ), .B(
        \Reg_Bank/registers[19][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5352 )
         );
  MUX \Reg_Bank/U5428  ( .A(\Reg_Bank/n5350 ), .B(\Reg_Bank/n5349 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5351 ) );
  MUX \Reg_Bank/U5427  ( .A(\Reg_Bank/registers[20][12] ), .B(
        \Reg_Bank/registers[21][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5350 )
         );
  MUX \Reg_Bank/U5426  ( .A(\Reg_Bank/registers[22][12] ), .B(
        \Reg_Bank/registers[23][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5349 )
         );
  MUX \Reg_Bank/U5425  ( .A(\Reg_Bank/n5347 ), .B(\Reg_Bank/n5344 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5348 ) );
  MUX \Reg_Bank/U5424  ( .A(\Reg_Bank/n5346 ), .B(\Reg_Bank/n5345 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5347 ) );
  MUX \Reg_Bank/U5423  ( .A(\Reg_Bank/registers[24][12] ), .B(
        \Reg_Bank/registers[25][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5346 )
         );
  MUX \Reg_Bank/U5422  ( .A(\Reg_Bank/registers[26][12] ), .B(
        \Reg_Bank/registers[27][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5345 )
         );
  MUX \Reg_Bank/U5421  ( .A(\Reg_Bank/n5343 ), .B(\Reg_Bank/n5342 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5344 ) );
  MUX \Reg_Bank/U5420  ( .A(\Reg_Bank/registers[28][12] ), .B(
        \Reg_Bank/registers[29][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5343 )
         );
  MUX \Reg_Bank/U5419  ( .A(\Reg_Bank/registers[30][12] ), .B(
        \Reg_Bank/registers[31][12] ), .S(rt_index[0]), .Z(\Reg_Bank/n5342 )
         );
  MUX \Reg_Bank/U5418  ( .A(\Reg_Bank/n5341 ), .B(\Reg_Bank/n5326 ), .S(
        rt_index[4]), .Z(reg_target[11]) );
  MUX \Reg_Bank/U5417  ( .A(\Reg_Bank/n5340 ), .B(\Reg_Bank/n5333 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5341 ) );
  MUX \Reg_Bank/U5416  ( .A(\Reg_Bank/n5339 ), .B(\Reg_Bank/n5336 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5340 ) );
  MUX \Reg_Bank/U5415  ( .A(\Reg_Bank/n5338 ), .B(\Reg_Bank/n5337 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5339 ) );
  MUX \Reg_Bank/U5413  ( .A(\Reg_Bank/registers[2][11] ), .B(
        \Reg_Bank/registers[3][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5337 ) );
  MUX \Reg_Bank/U5412  ( .A(\Reg_Bank/n5335 ), .B(\Reg_Bank/n5334 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5336 ) );
  MUX \Reg_Bank/U5411  ( .A(\Reg_Bank/registers[4][11] ), .B(
        \Reg_Bank/registers[5][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5335 ) );
  MUX \Reg_Bank/U5410  ( .A(\Reg_Bank/registers[6][11] ), .B(
        \Reg_Bank/registers[7][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5334 ) );
  MUX \Reg_Bank/U5409  ( .A(\Reg_Bank/n5332 ), .B(\Reg_Bank/n5329 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5333 ) );
  MUX \Reg_Bank/U5408  ( .A(\Reg_Bank/n5331 ), .B(\Reg_Bank/n5330 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5332 ) );
  MUX \Reg_Bank/U5407  ( .A(\Reg_Bank/registers[8][11] ), .B(
        \Reg_Bank/registers[9][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5331 ) );
  MUX \Reg_Bank/U5406  ( .A(\Reg_Bank/registers[10][11] ), .B(
        \Reg_Bank/registers[11][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5330 )
         );
  MUX \Reg_Bank/U5405  ( .A(\Reg_Bank/n5328 ), .B(\Reg_Bank/n5327 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5329 ) );
  MUX \Reg_Bank/U5404  ( .A(\Reg_Bank/registers[12][11] ), .B(
        \Reg_Bank/registers[13][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5328 )
         );
  MUX \Reg_Bank/U5403  ( .A(\Reg_Bank/registers[14][11] ), .B(
        \Reg_Bank/registers[15][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5327 )
         );
  MUX \Reg_Bank/U5402  ( .A(\Reg_Bank/n5325 ), .B(\Reg_Bank/n5318 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5326 ) );
  MUX \Reg_Bank/U5401  ( .A(\Reg_Bank/n5324 ), .B(\Reg_Bank/n5321 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5325 ) );
  MUX \Reg_Bank/U5400  ( .A(\Reg_Bank/n5323 ), .B(\Reg_Bank/n5322 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5324 ) );
  MUX \Reg_Bank/U5399  ( .A(\Reg_Bank/registers[16][11] ), .B(
        \Reg_Bank/registers[17][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5323 )
         );
  MUX \Reg_Bank/U5398  ( .A(\Reg_Bank/registers[18][11] ), .B(
        \Reg_Bank/registers[19][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5322 )
         );
  MUX \Reg_Bank/U5397  ( .A(\Reg_Bank/n5320 ), .B(\Reg_Bank/n5319 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5321 ) );
  MUX \Reg_Bank/U5396  ( .A(\Reg_Bank/registers[20][11] ), .B(
        \Reg_Bank/registers[21][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5320 )
         );
  MUX \Reg_Bank/U5395  ( .A(\Reg_Bank/registers[22][11] ), .B(
        \Reg_Bank/registers[23][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5319 )
         );
  MUX \Reg_Bank/U5394  ( .A(\Reg_Bank/n5317 ), .B(\Reg_Bank/n5314 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5318 ) );
  MUX \Reg_Bank/U5393  ( .A(\Reg_Bank/n5316 ), .B(\Reg_Bank/n5315 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5317 ) );
  MUX \Reg_Bank/U5392  ( .A(\Reg_Bank/registers[24][11] ), .B(
        \Reg_Bank/registers[25][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5316 )
         );
  MUX \Reg_Bank/U5391  ( .A(\Reg_Bank/registers[26][11] ), .B(
        \Reg_Bank/registers[27][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5315 )
         );
  MUX \Reg_Bank/U5390  ( .A(\Reg_Bank/n5313 ), .B(\Reg_Bank/n5312 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5314 ) );
  MUX \Reg_Bank/U5389  ( .A(\Reg_Bank/registers[28][11] ), .B(
        \Reg_Bank/registers[29][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5313 )
         );
  MUX \Reg_Bank/U5388  ( .A(\Reg_Bank/registers[30][11] ), .B(
        \Reg_Bank/registers[31][11] ), .S(rt_index[0]), .Z(\Reg_Bank/n5312 )
         );
  MUX \Reg_Bank/U5387  ( .A(\Reg_Bank/n5311 ), .B(\Reg_Bank/n5296 ), .S(
        rt_index[4]), .Z(reg_target[10]) );
  MUX \Reg_Bank/U5386  ( .A(\Reg_Bank/n5310 ), .B(\Reg_Bank/n5303 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5311 ) );
  MUX \Reg_Bank/U5385  ( .A(\Reg_Bank/n5309 ), .B(\Reg_Bank/n5306 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5310 ) );
  MUX \Reg_Bank/U5384  ( .A(\Reg_Bank/n5308 ), .B(\Reg_Bank/n5307 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5309 ) );
  MUX \Reg_Bank/U5382  ( .A(\Reg_Bank/registers[2][10] ), .B(
        \Reg_Bank/registers[3][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5307 ) );
  MUX \Reg_Bank/U5381  ( .A(\Reg_Bank/n5305 ), .B(\Reg_Bank/n5304 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5306 ) );
  MUX \Reg_Bank/U5380  ( .A(\Reg_Bank/registers[4][10] ), .B(
        \Reg_Bank/registers[5][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5305 ) );
  MUX \Reg_Bank/U5379  ( .A(\Reg_Bank/registers[6][10] ), .B(
        \Reg_Bank/registers[7][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5304 ) );
  MUX \Reg_Bank/U5378  ( .A(\Reg_Bank/n5302 ), .B(\Reg_Bank/n5299 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5303 ) );
  MUX \Reg_Bank/U5377  ( .A(\Reg_Bank/n5301 ), .B(\Reg_Bank/n5300 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5302 ) );
  MUX \Reg_Bank/U5376  ( .A(\Reg_Bank/registers[8][10] ), .B(
        \Reg_Bank/registers[9][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5301 ) );
  MUX \Reg_Bank/U5375  ( .A(\Reg_Bank/registers[10][10] ), .B(
        \Reg_Bank/registers[11][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5300 )
         );
  MUX \Reg_Bank/U5374  ( .A(\Reg_Bank/n5298 ), .B(\Reg_Bank/n5297 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5299 ) );
  MUX \Reg_Bank/U5373  ( .A(\Reg_Bank/registers[12][10] ), .B(
        \Reg_Bank/registers[13][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5298 )
         );
  MUX \Reg_Bank/U5372  ( .A(\Reg_Bank/registers[14][10] ), .B(
        \Reg_Bank/registers[15][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5297 )
         );
  MUX \Reg_Bank/U5371  ( .A(\Reg_Bank/n5295 ), .B(\Reg_Bank/n5288 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5296 ) );
  MUX \Reg_Bank/U5370  ( .A(\Reg_Bank/n5294 ), .B(\Reg_Bank/n5291 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5295 ) );
  MUX \Reg_Bank/U5369  ( .A(\Reg_Bank/n5293 ), .B(\Reg_Bank/n5292 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5294 ) );
  MUX \Reg_Bank/U5368  ( .A(\Reg_Bank/registers[16][10] ), .B(
        \Reg_Bank/registers[17][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5293 )
         );
  MUX \Reg_Bank/U5367  ( .A(\Reg_Bank/registers[18][10] ), .B(
        \Reg_Bank/registers[19][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5292 )
         );
  MUX \Reg_Bank/U5366  ( .A(\Reg_Bank/n5290 ), .B(\Reg_Bank/n5289 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5291 ) );
  MUX \Reg_Bank/U5365  ( .A(\Reg_Bank/registers[20][10] ), .B(
        \Reg_Bank/registers[21][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5290 )
         );
  MUX \Reg_Bank/U5364  ( .A(\Reg_Bank/registers[22][10] ), .B(
        \Reg_Bank/registers[23][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5289 )
         );
  MUX \Reg_Bank/U5363  ( .A(\Reg_Bank/n5287 ), .B(\Reg_Bank/n5284 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5288 ) );
  MUX \Reg_Bank/U5362  ( .A(\Reg_Bank/n5286 ), .B(\Reg_Bank/n5285 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5287 ) );
  MUX \Reg_Bank/U5361  ( .A(\Reg_Bank/registers[24][10] ), .B(
        \Reg_Bank/registers[25][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5286 )
         );
  MUX \Reg_Bank/U5360  ( .A(\Reg_Bank/registers[26][10] ), .B(
        \Reg_Bank/registers[27][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5285 )
         );
  MUX \Reg_Bank/U5359  ( .A(\Reg_Bank/n5283 ), .B(\Reg_Bank/n5282 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5284 ) );
  MUX \Reg_Bank/U5358  ( .A(\Reg_Bank/registers[28][10] ), .B(
        \Reg_Bank/registers[29][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5283 )
         );
  MUX \Reg_Bank/U5357  ( .A(\Reg_Bank/registers[30][10] ), .B(
        \Reg_Bank/registers[31][10] ), .S(rt_index[0]), .Z(\Reg_Bank/n5282 )
         );
  MUX \Reg_Bank/U5356  ( .A(\Reg_Bank/n5281 ), .B(\Reg_Bank/n5266 ), .S(
        rt_index[4]), .Z(reg_target[9]) );
  MUX \Reg_Bank/U5355  ( .A(\Reg_Bank/n5280 ), .B(\Reg_Bank/n5273 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5281 ) );
  MUX \Reg_Bank/U5354  ( .A(\Reg_Bank/n5279 ), .B(\Reg_Bank/n5276 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5280 ) );
  MUX \Reg_Bank/U5353  ( .A(\Reg_Bank/n5278 ), .B(\Reg_Bank/n5277 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5279 ) );
  MUX \Reg_Bank/U5351  ( .A(\Reg_Bank/registers[2][9] ), .B(
        \Reg_Bank/registers[3][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5277 ) );
  MUX \Reg_Bank/U5350  ( .A(\Reg_Bank/n5275 ), .B(\Reg_Bank/n5274 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5276 ) );
  MUX \Reg_Bank/U5349  ( .A(\Reg_Bank/registers[4][9] ), .B(
        \Reg_Bank/registers[5][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5275 ) );
  MUX \Reg_Bank/U5348  ( .A(\Reg_Bank/registers[6][9] ), .B(
        \Reg_Bank/registers[7][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5274 ) );
  MUX \Reg_Bank/U5347  ( .A(\Reg_Bank/n5272 ), .B(\Reg_Bank/n5269 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5273 ) );
  MUX \Reg_Bank/U5346  ( .A(\Reg_Bank/n5271 ), .B(\Reg_Bank/n5270 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5272 ) );
  MUX \Reg_Bank/U5345  ( .A(\Reg_Bank/registers[8][9] ), .B(
        \Reg_Bank/registers[9][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5271 ) );
  MUX \Reg_Bank/U5344  ( .A(\Reg_Bank/registers[10][9] ), .B(
        \Reg_Bank/registers[11][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5270 ) );
  MUX \Reg_Bank/U5343  ( .A(\Reg_Bank/n5268 ), .B(\Reg_Bank/n5267 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5269 ) );
  MUX \Reg_Bank/U5342  ( .A(\Reg_Bank/registers[12][9] ), .B(
        \Reg_Bank/registers[13][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5268 ) );
  MUX \Reg_Bank/U5341  ( .A(\Reg_Bank/registers[14][9] ), .B(
        \Reg_Bank/registers[15][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5267 ) );
  MUX \Reg_Bank/U5340  ( .A(\Reg_Bank/n5265 ), .B(\Reg_Bank/n5258 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5266 ) );
  MUX \Reg_Bank/U5339  ( .A(\Reg_Bank/n5264 ), .B(\Reg_Bank/n5261 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5265 ) );
  MUX \Reg_Bank/U5338  ( .A(\Reg_Bank/n5263 ), .B(\Reg_Bank/n5262 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5264 ) );
  MUX \Reg_Bank/U5337  ( .A(\Reg_Bank/registers[16][9] ), .B(
        \Reg_Bank/registers[17][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5263 ) );
  MUX \Reg_Bank/U5336  ( .A(\Reg_Bank/registers[18][9] ), .B(
        \Reg_Bank/registers[19][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5262 ) );
  MUX \Reg_Bank/U5335  ( .A(\Reg_Bank/n5260 ), .B(\Reg_Bank/n5259 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5261 ) );
  MUX \Reg_Bank/U5334  ( .A(\Reg_Bank/registers[20][9] ), .B(
        \Reg_Bank/registers[21][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5260 ) );
  MUX \Reg_Bank/U5333  ( .A(\Reg_Bank/registers[22][9] ), .B(
        \Reg_Bank/registers[23][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5259 ) );
  MUX \Reg_Bank/U5332  ( .A(\Reg_Bank/n5257 ), .B(\Reg_Bank/n5254 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5258 ) );
  MUX \Reg_Bank/U5331  ( .A(\Reg_Bank/n5256 ), .B(\Reg_Bank/n5255 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5257 ) );
  MUX \Reg_Bank/U5330  ( .A(\Reg_Bank/registers[24][9] ), .B(
        \Reg_Bank/registers[25][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5256 ) );
  MUX \Reg_Bank/U5329  ( .A(\Reg_Bank/registers[26][9] ), .B(
        \Reg_Bank/registers[27][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5255 ) );
  MUX \Reg_Bank/U5328  ( .A(\Reg_Bank/n5253 ), .B(\Reg_Bank/n5252 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5254 ) );
  MUX \Reg_Bank/U5327  ( .A(\Reg_Bank/registers[28][9] ), .B(
        \Reg_Bank/registers[29][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5253 ) );
  MUX \Reg_Bank/U5326  ( .A(\Reg_Bank/registers[30][9] ), .B(
        \Reg_Bank/registers[31][9] ), .S(rt_index[0]), .Z(\Reg_Bank/n5252 ) );
  MUX \Reg_Bank/U5325  ( .A(\Reg_Bank/n5251 ), .B(\Reg_Bank/n5236 ), .S(
        rt_index[4]), .Z(reg_target[8]) );
  MUX \Reg_Bank/U5324  ( .A(\Reg_Bank/n5250 ), .B(\Reg_Bank/n5243 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5251 ) );
  MUX \Reg_Bank/U5323  ( .A(\Reg_Bank/n5249 ), .B(\Reg_Bank/n5246 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5250 ) );
  MUX \Reg_Bank/U5322  ( .A(\Reg_Bank/n5248 ), .B(\Reg_Bank/n5247 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5249 ) );
  MUX \Reg_Bank/U5320  ( .A(\Reg_Bank/registers[2][8] ), .B(
        \Reg_Bank/registers[3][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5247 ) );
  MUX \Reg_Bank/U5319  ( .A(\Reg_Bank/n5245 ), .B(\Reg_Bank/n5244 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5246 ) );
  MUX \Reg_Bank/U5318  ( .A(\Reg_Bank/registers[4][8] ), .B(
        \Reg_Bank/registers[5][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5245 ) );
  MUX \Reg_Bank/U5317  ( .A(\Reg_Bank/registers[6][8] ), .B(
        \Reg_Bank/registers[7][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5244 ) );
  MUX \Reg_Bank/U5316  ( .A(\Reg_Bank/n5242 ), .B(\Reg_Bank/n5239 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5243 ) );
  MUX \Reg_Bank/U5315  ( .A(\Reg_Bank/n5241 ), .B(\Reg_Bank/n5240 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5242 ) );
  MUX \Reg_Bank/U5314  ( .A(\Reg_Bank/registers[8][8] ), .B(
        \Reg_Bank/registers[9][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5241 ) );
  MUX \Reg_Bank/U5313  ( .A(\Reg_Bank/registers[10][8] ), .B(
        \Reg_Bank/registers[11][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5240 ) );
  MUX \Reg_Bank/U5312  ( .A(\Reg_Bank/n5238 ), .B(\Reg_Bank/n5237 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5239 ) );
  MUX \Reg_Bank/U5311  ( .A(\Reg_Bank/registers[12][8] ), .B(
        \Reg_Bank/registers[13][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5238 ) );
  MUX \Reg_Bank/U5310  ( .A(\Reg_Bank/registers[14][8] ), .B(
        \Reg_Bank/registers[15][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5237 ) );
  MUX \Reg_Bank/U5309  ( .A(\Reg_Bank/n5235 ), .B(\Reg_Bank/n5228 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5236 ) );
  MUX \Reg_Bank/U5308  ( .A(\Reg_Bank/n5234 ), .B(\Reg_Bank/n5231 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5235 ) );
  MUX \Reg_Bank/U5307  ( .A(\Reg_Bank/n5233 ), .B(\Reg_Bank/n5232 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5234 ) );
  MUX \Reg_Bank/U5306  ( .A(\Reg_Bank/registers[16][8] ), .B(
        \Reg_Bank/registers[17][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5233 ) );
  MUX \Reg_Bank/U5305  ( .A(\Reg_Bank/registers[18][8] ), .B(
        \Reg_Bank/registers[19][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5232 ) );
  MUX \Reg_Bank/U5304  ( .A(\Reg_Bank/n5230 ), .B(\Reg_Bank/n5229 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5231 ) );
  MUX \Reg_Bank/U5303  ( .A(\Reg_Bank/registers[20][8] ), .B(
        \Reg_Bank/registers[21][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5230 ) );
  MUX \Reg_Bank/U5302  ( .A(\Reg_Bank/registers[22][8] ), .B(
        \Reg_Bank/registers[23][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5229 ) );
  MUX \Reg_Bank/U5301  ( .A(\Reg_Bank/n5227 ), .B(\Reg_Bank/n5224 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5228 ) );
  MUX \Reg_Bank/U5300  ( .A(\Reg_Bank/n5226 ), .B(\Reg_Bank/n5225 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5227 ) );
  MUX \Reg_Bank/U5299  ( .A(\Reg_Bank/registers[24][8] ), .B(
        \Reg_Bank/registers[25][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5226 ) );
  MUX \Reg_Bank/U5298  ( .A(\Reg_Bank/registers[26][8] ), .B(
        \Reg_Bank/registers[27][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5225 ) );
  MUX \Reg_Bank/U5297  ( .A(\Reg_Bank/n5223 ), .B(\Reg_Bank/n5222 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5224 ) );
  MUX \Reg_Bank/U5296  ( .A(\Reg_Bank/registers[28][8] ), .B(
        \Reg_Bank/registers[29][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5223 ) );
  MUX \Reg_Bank/U5295  ( .A(\Reg_Bank/registers[30][8] ), .B(
        \Reg_Bank/registers[31][8] ), .S(rt_index[0]), .Z(\Reg_Bank/n5222 ) );
  MUX \Reg_Bank/U5294  ( .A(\Reg_Bank/n5221 ), .B(\Reg_Bank/n5206 ), .S(
        rt_index[4]), .Z(reg_target[7]) );
  MUX \Reg_Bank/U5293  ( .A(\Reg_Bank/n5220 ), .B(\Reg_Bank/n5213 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5221 ) );
  MUX \Reg_Bank/U5292  ( .A(\Reg_Bank/n5219 ), .B(\Reg_Bank/n5216 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5220 ) );
  MUX \Reg_Bank/U5291  ( .A(\Reg_Bank/n5218 ), .B(\Reg_Bank/n5217 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5219 ) );
  MUX \Reg_Bank/U5289  ( .A(\Reg_Bank/registers[2][7] ), .B(
        \Reg_Bank/registers[3][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5217 ) );
  MUX \Reg_Bank/U5288  ( .A(\Reg_Bank/n5215 ), .B(\Reg_Bank/n5214 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5216 ) );
  MUX \Reg_Bank/U5287  ( .A(\Reg_Bank/registers[4][7] ), .B(
        \Reg_Bank/registers[5][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5215 ) );
  MUX \Reg_Bank/U5286  ( .A(\Reg_Bank/registers[6][7] ), .B(
        \Reg_Bank/registers[7][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5214 ) );
  MUX \Reg_Bank/U5285  ( .A(\Reg_Bank/n5212 ), .B(\Reg_Bank/n5209 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5213 ) );
  MUX \Reg_Bank/U5284  ( .A(\Reg_Bank/n5211 ), .B(\Reg_Bank/n5210 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5212 ) );
  MUX \Reg_Bank/U5283  ( .A(\Reg_Bank/registers[8][7] ), .B(
        \Reg_Bank/registers[9][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5211 ) );
  MUX \Reg_Bank/U5282  ( .A(\Reg_Bank/registers[10][7] ), .B(
        \Reg_Bank/registers[11][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5210 ) );
  MUX \Reg_Bank/U5281  ( .A(\Reg_Bank/n5208 ), .B(\Reg_Bank/n5207 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5209 ) );
  MUX \Reg_Bank/U5280  ( .A(\Reg_Bank/registers[12][7] ), .B(
        \Reg_Bank/registers[13][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5208 ) );
  MUX \Reg_Bank/U5279  ( .A(\Reg_Bank/registers[14][7] ), .B(
        \Reg_Bank/registers[15][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5207 ) );
  MUX \Reg_Bank/U5278  ( .A(\Reg_Bank/n5205 ), .B(\Reg_Bank/n5198 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5206 ) );
  MUX \Reg_Bank/U5277  ( .A(\Reg_Bank/n5204 ), .B(\Reg_Bank/n5201 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5205 ) );
  MUX \Reg_Bank/U5276  ( .A(\Reg_Bank/n5203 ), .B(\Reg_Bank/n5202 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5204 ) );
  MUX \Reg_Bank/U5275  ( .A(\Reg_Bank/registers[16][7] ), .B(
        \Reg_Bank/registers[17][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5203 ) );
  MUX \Reg_Bank/U5274  ( .A(\Reg_Bank/registers[18][7] ), .B(
        \Reg_Bank/registers[19][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5202 ) );
  MUX \Reg_Bank/U5273  ( .A(\Reg_Bank/n5200 ), .B(\Reg_Bank/n5199 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5201 ) );
  MUX \Reg_Bank/U5272  ( .A(\Reg_Bank/registers[20][7] ), .B(
        \Reg_Bank/registers[21][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5200 ) );
  MUX \Reg_Bank/U5271  ( .A(\Reg_Bank/registers[22][7] ), .B(
        \Reg_Bank/registers[23][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5199 ) );
  MUX \Reg_Bank/U5270  ( .A(\Reg_Bank/n5197 ), .B(\Reg_Bank/n5194 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5198 ) );
  MUX \Reg_Bank/U5269  ( .A(\Reg_Bank/n5196 ), .B(\Reg_Bank/n5195 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5197 ) );
  MUX \Reg_Bank/U5268  ( .A(\Reg_Bank/registers[24][7] ), .B(
        \Reg_Bank/registers[25][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5196 ) );
  MUX \Reg_Bank/U5267  ( .A(\Reg_Bank/registers[26][7] ), .B(
        \Reg_Bank/registers[27][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5195 ) );
  MUX \Reg_Bank/U5266  ( .A(\Reg_Bank/n5193 ), .B(\Reg_Bank/n5192 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5194 ) );
  MUX \Reg_Bank/U5265  ( .A(\Reg_Bank/registers[28][7] ), .B(
        \Reg_Bank/registers[29][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5193 ) );
  MUX \Reg_Bank/U5264  ( .A(\Reg_Bank/registers[30][7] ), .B(
        \Reg_Bank/registers[31][7] ), .S(rt_index[0]), .Z(\Reg_Bank/n5192 ) );
  MUX \Reg_Bank/U5263  ( .A(\Reg_Bank/n5191 ), .B(\Reg_Bank/n5176 ), .S(
        rt_index[4]), .Z(reg_target[6]) );
  MUX \Reg_Bank/U5262  ( .A(\Reg_Bank/n5190 ), .B(\Reg_Bank/n5183 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5191 ) );
  MUX \Reg_Bank/U5261  ( .A(\Reg_Bank/n5189 ), .B(\Reg_Bank/n5186 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5190 ) );
  MUX \Reg_Bank/U5260  ( .A(\Reg_Bank/n5188 ), .B(\Reg_Bank/n5187 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5189 ) );
  MUX \Reg_Bank/U5258  ( .A(\Reg_Bank/registers[2][6] ), .B(
        \Reg_Bank/registers[3][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5187 ) );
  MUX \Reg_Bank/U5257  ( .A(\Reg_Bank/n5185 ), .B(\Reg_Bank/n5184 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5186 ) );
  MUX \Reg_Bank/U5256  ( .A(\Reg_Bank/registers[4][6] ), .B(
        \Reg_Bank/registers[5][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5185 ) );
  MUX \Reg_Bank/U5255  ( .A(\Reg_Bank/registers[6][6] ), .B(
        \Reg_Bank/registers[7][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5184 ) );
  MUX \Reg_Bank/U5254  ( .A(\Reg_Bank/n5182 ), .B(\Reg_Bank/n5179 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5183 ) );
  MUX \Reg_Bank/U5253  ( .A(\Reg_Bank/n5181 ), .B(\Reg_Bank/n5180 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5182 ) );
  MUX \Reg_Bank/U5252  ( .A(\Reg_Bank/registers[8][6] ), .B(
        \Reg_Bank/registers[9][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5181 ) );
  MUX \Reg_Bank/U5251  ( .A(\Reg_Bank/registers[10][6] ), .B(
        \Reg_Bank/registers[11][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5180 ) );
  MUX \Reg_Bank/U5250  ( .A(\Reg_Bank/n5178 ), .B(\Reg_Bank/n5177 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5179 ) );
  MUX \Reg_Bank/U5249  ( .A(\Reg_Bank/registers[12][6] ), .B(
        \Reg_Bank/registers[13][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5178 ) );
  MUX \Reg_Bank/U5248  ( .A(\Reg_Bank/registers[14][6] ), .B(
        \Reg_Bank/registers[15][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5177 ) );
  MUX \Reg_Bank/U5247  ( .A(\Reg_Bank/n5175 ), .B(\Reg_Bank/n5168 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5176 ) );
  MUX \Reg_Bank/U5246  ( .A(\Reg_Bank/n5174 ), .B(\Reg_Bank/n5171 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5175 ) );
  MUX \Reg_Bank/U5245  ( .A(\Reg_Bank/n5173 ), .B(\Reg_Bank/n5172 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5174 ) );
  MUX \Reg_Bank/U5244  ( .A(\Reg_Bank/registers[16][6] ), .B(
        \Reg_Bank/registers[17][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5173 ) );
  MUX \Reg_Bank/U5243  ( .A(\Reg_Bank/registers[18][6] ), .B(
        \Reg_Bank/registers[19][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5172 ) );
  MUX \Reg_Bank/U5242  ( .A(\Reg_Bank/n5170 ), .B(\Reg_Bank/n5169 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5171 ) );
  MUX \Reg_Bank/U5241  ( .A(\Reg_Bank/registers[20][6] ), .B(
        \Reg_Bank/registers[21][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5170 ) );
  MUX \Reg_Bank/U5240  ( .A(\Reg_Bank/registers[22][6] ), .B(
        \Reg_Bank/registers[23][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5169 ) );
  MUX \Reg_Bank/U5239  ( .A(\Reg_Bank/n5167 ), .B(\Reg_Bank/n5164 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5168 ) );
  MUX \Reg_Bank/U5238  ( .A(\Reg_Bank/n5166 ), .B(\Reg_Bank/n5165 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5167 ) );
  MUX \Reg_Bank/U5237  ( .A(\Reg_Bank/registers[24][6] ), .B(
        \Reg_Bank/registers[25][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5166 ) );
  MUX \Reg_Bank/U5236  ( .A(\Reg_Bank/registers[26][6] ), .B(
        \Reg_Bank/registers[27][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5165 ) );
  MUX \Reg_Bank/U5235  ( .A(\Reg_Bank/n5163 ), .B(\Reg_Bank/n5162 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5164 ) );
  MUX \Reg_Bank/U5234  ( .A(\Reg_Bank/registers[28][6] ), .B(
        \Reg_Bank/registers[29][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5163 ) );
  MUX \Reg_Bank/U5233  ( .A(\Reg_Bank/registers[30][6] ), .B(
        \Reg_Bank/registers[31][6] ), .S(rt_index[0]), .Z(\Reg_Bank/n5162 ) );
  MUX \Reg_Bank/U5232  ( .A(\Reg_Bank/n5161 ), .B(\Reg_Bank/n5146 ), .S(
        rt_index[4]), .Z(reg_target[5]) );
  MUX \Reg_Bank/U5231  ( .A(\Reg_Bank/n5160 ), .B(\Reg_Bank/n5153 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5161 ) );
  MUX \Reg_Bank/U5230  ( .A(\Reg_Bank/n5159 ), .B(\Reg_Bank/n5156 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5160 ) );
  MUX \Reg_Bank/U5229  ( .A(\Reg_Bank/n5158 ), .B(\Reg_Bank/n5157 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5159 ) );
  MUX \Reg_Bank/U5227  ( .A(\Reg_Bank/registers[2][5] ), .B(
        \Reg_Bank/registers[3][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5157 ) );
  MUX \Reg_Bank/U5226  ( .A(\Reg_Bank/n5155 ), .B(\Reg_Bank/n5154 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5156 ) );
  MUX \Reg_Bank/U5225  ( .A(\Reg_Bank/registers[4][5] ), .B(
        \Reg_Bank/registers[5][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5155 ) );
  MUX \Reg_Bank/U5224  ( .A(\Reg_Bank/registers[6][5] ), .B(
        \Reg_Bank/registers[7][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5154 ) );
  MUX \Reg_Bank/U5223  ( .A(\Reg_Bank/n5152 ), .B(\Reg_Bank/n5149 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5153 ) );
  MUX \Reg_Bank/U5222  ( .A(\Reg_Bank/n5151 ), .B(\Reg_Bank/n5150 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5152 ) );
  MUX \Reg_Bank/U5221  ( .A(\Reg_Bank/registers[8][5] ), .B(
        \Reg_Bank/registers[9][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5151 ) );
  MUX \Reg_Bank/U5220  ( .A(\Reg_Bank/registers[10][5] ), .B(
        \Reg_Bank/registers[11][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5150 ) );
  MUX \Reg_Bank/U5219  ( .A(\Reg_Bank/n5148 ), .B(\Reg_Bank/n5147 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5149 ) );
  MUX \Reg_Bank/U5218  ( .A(\Reg_Bank/registers[12][5] ), .B(
        \Reg_Bank/registers[13][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5148 ) );
  MUX \Reg_Bank/U5217  ( .A(\Reg_Bank/registers[14][5] ), .B(
        \Reg_Bank/registers[15][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5147 ) );
  MUX \Reg_Bank/U5216  ( .A(\Reg_Bank/n5145 ), .B(\Reg_Bank/n5138 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5146 ) );
  MUX \Reg_Bank/U5215  ( .A(\Reg_Bank/n5144 ), .B(\Reg_Bank/n5141 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5145 ) );
  MUX \Reg_Bank/U5214  ( .A(\Reg_Bank/n5143 ), .B(\Reg_Bank/n5142 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5144 ) );
  MUX \Reg_Bank/U5213  ( .A(\Reg_Bank/registers[16][5] ), .B(
        \Reg_Bank/registers[17][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5143 ) );
  MUX \Reg_Bank/U5212  ( .A(\Reg_Bank/registers[18][5] ), .B(
        \Reg_Bank/registers[19][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5142 ) );
  MUX \Reg_Bank/U5211  ( .A(\Reg_Bank/n5140 ), .B(\Reg_Bank/n5139 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5141 ) );
  MUX \Reg_Bank/U5210  ( .A(\Reg_Bank/registers[20][5] ), .B(
        \Reg_Bank/registers[21][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5140 ) );
  MUX \Reg_Bank/U5209  ( .A(\Reg_Bank/registers[22][5] ), .B(
        \Reg_Bank/registers[23][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5139 ) );
  MUX \Reg_Bank/U5208  ( .A(\Reg_Bank/n5137 ), .B(\Reg_Bank/n5134 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5138 ) );
  MUX \Reg_Bank/U5207  ( .A(\Reg_Bank/n5136 ), .B(\Reg_Bank/n5135 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5137 ) );
  MUX \Reg_Bank/U5206  ( .A(\Reg_Bank/registers[24][5] ), .B(
        \Reg_Bank/registers[25][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5136 ) );
  MUX \Reg_Bank/U5205  ( .A(\Reg_Bank/registers[26][5] ), .B(
        \Reg_Bank/registers[27][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5135 ) );
  MUX \Reg_Bank/U5204  ( .A(\Reg_Bank/n5133 ), .B(\Reg_Bank/n5132 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5134 ) );
  MUX \Reg_Bank/U5203  ( .A(\Reg_Bank/registers[28][5] ), .B(
        \Reg_Bank/registers[29][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5133 ) );
  MUX \Reg_Bank/U5202  ( .A(\Reg_Bank/registers[30][5] ), .B(
        \Reg_Bank/registers[31][5] ), .S(rt_index[0]), .Z(\Reg_Bank/n5132 ) );
  MUX \Reg_Bank/U5201  ( .A(\Reg_Bank/n5131 ), .B(\Reg_Bank/n5116 ), .S(
        rt_index[4]), .Z(reg_target[4]) );
  MUX \Reg_Bank/U5200  ( .A(\Reg_Bank/n5130 ), .B(\Reg_Bank/n5123 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5131 ) );
  MUX \Reg_Bank/U5199  ( .A(\Reg_Bank/n5129 ), .B(\Reg_Bank/n5126 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5130 ) );
  MUX \Reg_Bank/U5198  ( .A(\Reg_Bank/n5128 ), .B(\Reg_Bank/n5127 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5129 ) );
  MUX \Reg_Bank/U5196  ( .A(\Reg_Bank/registers[2][4] ), .B(
        \Reg_Bank/registers[3][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5127 ) );
  MUX \Reg_Bank/U5195  ( .A(\Reg_Bank/n5125 ), .B(\Reg_Bank/n5124 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5126 ) );
  MUX \Reg_Bank/U5194  ( .A(\Reg_Bank/registers[4][4] ), .B(
        \Reg_Bank/registers[5][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5125 ) );
  MUX \Reg_Bank/U5193  ( .A(\Reg_Bank/registers[6][4] ), .B(
        \Reg_Bank/registers[7][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5124 ) );
  MUX \Reg_Bank/U5192  ( .A(\Reg_Bank/n5122 ), .B(\Reg_Bank/n5119 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5123 ) );
  MUX \Reg_Bank/U5191  ( .A(\Reg_Bank/n5121 ), .B(\Reg_Bank/n5120 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5122 ) );
  MUX \Reg_Bank/U5190  ( .A(\Reg_Bank/registers[8][4] ), .B(
        \Reg_Bank/registers[9][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5121 ) );
  MUX \Reg_Bank/U5189  ( .A(\Reg_Bank/registers[10][4] ), .B(
        \Reg_Bank/registers[11][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5120 ) );
  MUX \Reg_Bank/U5188  ( .A(\Reg_Bank/n5118 ), .B(\Reg_Bank/n5117 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5119 ) );
  MUX \Reg_Bank/U5187  ( .A(\Reg_Bank/registers[12][4] ), .B(
        \Reg_Bank/registers[13][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5118 ) );
  MUX \Reg_Bank/U5186  ( .A(\Reg_Bank/registers[14][4] ), .B(
        \Reg_Bank/registers[15][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5117 ) );
  MUX \Reg_Bank/U5185  ( .A(\Reg_Bank/n5115 ), .B(\Reg_Bank/n5108 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5116 ) );
  MUX \Reg_Bank/U5184  ( .A(\Reg_Bank/n5114 ), .B(\Reg_Bank/n5111 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5115 ) );
  MUX \Reg_Bank/U5183  ( .A(\Reg_Bank/n5113 ), .B(\Reg_Bank/n5112 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5114 ) );
  MUX \Reg_Bank/U5182  ( .A(\Reg_Bank/registers[16][4] ), .B(
        \Reg_Bank/registers[17][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5113 ) );
  MUX \Reg_Bank/U5181  ( .A(\Reg_Bank/registers[18][4] ), .B(
        \Reg_Bank/registers[19][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5112 ) );
  MUX \Reg_Bank/U5180  ( .A(\Reg_Bank/n5110 ), .B(\Reg_Bank/n5109 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5111 ) );
  MUX \Reg_Bank/U5179  ( .A(\Reg_Bank/registers[20][4] ), .B(
        \Reg_Bank/registers[21][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5110 ) );
  MUX \Reg_Bank/U5178  ( .A(\Reg_Bank/registers[22][4] ), .B(
        \Reg_Bank/registers[23][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5109 ) );
  MUX \Reg_Bank/U5177  ( .A(\Reg_Bank/n5107 ), .B(\Reg_Bank/n5104 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5108 ) );
  MUX \Reg_Bank/U5176  ( .A(\Reg_Bank/n5106 ), .B(\Reg_Bank/n5105 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5107 ) );
  MUX \Reg_Bank/U5175  ( .A(\Reg_Bank/registers[24][4] ), .B(
        \Reg_Bank/registers[25][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5106 ) );
  MUX \Reg_Bank/U5174  ( .A(\Reg_Bank/registers[26][4] ), .B(
        \Reg_Bank/registers[27][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5105 ) );
  MUX \Reg_Bank/U5173  ( .A(\Reg_Bank/n5103 ), .B(\Reg_Bank/n5102 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5104 ) );
  MUX \Reg_Bank/U5172  ( .A(\Reg_Bank/registers[28][4] ), .B(
        \Reg_Bank/registers[29][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5103 ) );
  MUX \Reg_Bank/U5171  ( .A(\Reg_Bank/registers[30][4] ), .B(
        \Reg_Bank/registers[31][4] ), .S(rt_index[0]), .Z(\Reg_Bank/n5102 ) );
  MUX \Reg_Bank/U5170  ( .A(\Reg_Bank/n5101 ), .B(\Reg_Bank/n5086 ), .S(
        rt_index[4]), .Z(reg_target[3]) );
  MUX \Reg_Bank/U5169  ( .A(\Reg_Bank/n5100 ), .B(\Reg_Bank/n5093 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5101 ) );
  MUX \Reg_Bank/U5168  ( .A(\Reg_Bank/n5099 ), .B(\Reg_Bank/n5096 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5100 ) );
  MUX \Reg_Bank/U5167  ( .A(\Reg_Bank/n5098 ), .B(\Reg_Bank/n5097 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5099 ) );
  MUX \Reg_Bank/U5165  ( .A(\Reg_Bank/registers[2][3] ), .B(
        \Reg_Bank/registers[3][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5097 ) );
  MUX \Reg_Bank/U5164  ( .A(\Reg_Bank/n5095 ), .B(\Reg_Bank/n5094 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5096 ) );
  MUX \Reg_Bank/U5163  ( .A(\Reg_Bank/registers[4][3] ), .B(
        \Reg_Bank/registers[5][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5095 ) );
  MUX \Reg_Bank/U5162  ( .A(\Reg_Bank/registers[6][3] ), .B(
        \Reg_Bank/registers[7][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5094 ) );
  MUX \Reg_Bank/U5161  ( .A(\Reg_Bank/n5092 ), .B(\Reg_Bank/n5089 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5093 ) );
  MUX \Reg_Bank/U5160  ( .A(\Reg_Bank/n5091 ), .B(\Reg_Bank/n5090 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5092 ) );
  MUX \Reg_Bank/U5159  ( .A(\Reg_Bank/registers[8][3] ), .B(
        \Reg_Bank/registers[9][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5091 ) );
  MUX \Reg_Bank/U5158  ( .A(\Reg_Bank/registers[10][3] ), .B(
        \Reg_Bank/registers[11][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5090 ) );
  MUX \Reg_Bank/U5157  ( .A(\Reg_Bank/n5088 ), .B(\Reg_Bank/n5087 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5089 ) );
  MUX \Reg_Bank/U5156  ( .A(\Reg_Bank/registers[12][3] ), .B(
        \Reg_Bank/registers[13][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5088 ) );
  MUX \Reg_Bank/U5155  ( .A(\Reg_Bank/registers[14][3] ), .B(
        \Reg_Bank/registers[15][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5087 ) );
  MUX \Reg_Bank/U5154  ( .A(\Reg_Bank/n5085 ), .B(\Reg_Bank/n5078 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5086 ) );
  MUX \Reg_Bank/U5153  ( .A(\Reg_Bank/n5084 ), .B(\Reg_Bank/n5081 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5085 ) );
  MUX \Reg_Bank/U5152  ( .A(\Reg_Bank/n5083 ), .B(\Reg_Bank/n5082 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5084 ) );
  MUX \Reg_Bank/U5151  ( .A(\Reg_Bank/registers[16][3] ), .B(
        \Reg_Bank/registers[17][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5083 ) );
  MUX \Reg_Bank/U5150  ( .A(\Reg_Bank/registers[18][3] ), .B(
        \Reg_Bank/registers[19][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5082 ) );
  MUX \Reg_Bank/U5149  ( .A(\Reg_Bank/n5080 ), .B(\Reg_Bank/n5079 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5081 ) );
  MUX \Reg_Bank/U5148  ( .A(\Reg_Bank/registers[20][3] ), .B(
        \Reg_Bank/registers[21][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5080 ) );
  MUX \Reg_Bank/U5147  ( .A(\Reg_Bank/registers[22][3] ), .B(
        \Reg_Bank/registers[23][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5079 ) );
  MUX \Reg_Bank/U5146  ( .A(\Reg_Bank/n5077 ), .B(\Reg_Bank/n5074 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5078 ) );
  MUX \Reg_Bank/U5145  ( .A(\Reg_Bank/n5076 ), .B(\Reg_Bank/n5075 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5077 ) );
  MUX \Reg_Bank/U5144  ( .A(\Reg_Bank/registers[24][3] ), .B(
        \Reg_Bank/registers[25][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5076 ) );
  MUX \Reg_Bank/U5143  ( .A(\Reg_Bank/registers[26][3] ), .B(
        \Reg_Bank/registers[27][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5075 ) );
  MUX \Reg_Bank/U5142  ( .A(\Reg_Bank/n5073 ), .B(\Reg_Bank/n5072 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5074 ) );
  MUX \Reg_Bank/U5141  ( .A(\Reg_Bank/registers[28][3] ), .B(
        \Reg_Bank/registers[29][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5073 ) );
  MUX \Reg_Bank/U5140  ( .A(\Reg_Bank/registers[30][3] ), .B(
        \Reg_Bank/registers[31][3] ), .S(rt_index[0]), .Z(\Reg_Bank/n5072 ) );
  MUX \Reg_Bank/U5139  ( .A(\Reg_Bank/n5071 ), .B(\Reg_Bank/n5056 ), .S(
        rt_index[4]), .Z(reg_target[2]) );
  MUX \Reg_Bank/U5138  ( .A(\Reg_Bank/n5070 ), .B(\Reg_Bank/n5063 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5071 ) );
  MUX \Reg_Bank/U5137  ( .A(\Reg_Bank/n5069 ), .B(\Reg_Bank/n5066 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5070 ) );
  MUX \Reg_Bank/U5136  ( .A(\Reg_Bank/n5068 ), .B(\Reg_Bank/n5067 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5069 ) );
  MUX \Reg_Bank/U5134  ( .A(\Reg_Bank/registers[2][2] ), .B(
        \Reg_Bank/registers[3][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5067 ) );
  MUX \Reg_Bank/U5133  ( .A(\Reg_Bank/n5065 ), .B(\Reg_Bank/n5064 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5066 ) );
  MUX \Reg_Bank/U5132  ( .A(\Reg_Bank/registers[4][2] ), .B(
        \Reg_Bank/registers[5][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5065 ) );
  MUX \Reg_Bank/U5131  ( .A(\Reg_Bank/registers[6][2] ), .B(
        \Reg_Bank/registers[7][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5064 ) );
  MUX \Reg_Bank/U5130  ( .A(\Reg_Bank/n5062 ), .B(\Reg_Bank/n5059 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5063 ) );
  MUX \Reg_Bank/U5129  ( .A(\Reg_Bank/n5061 ), .B(\Reg_Bank/n5060 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5062 ) );
  MUX \Reg_Bank/U5128  ( .A(\Reg_Bank/registers[8][2] ), .B(
        \Reg_Bank/registers[9][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5061 ) );
  MUX \Reg_Bank/U5127  ( .A(\Reg_Bank/registers[10][2] ), .B(
        \Reg_Bank/registers[11][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5060 ) );
  MUX \Reg_Bank/U5126  ( .A(\Reg_Bank/n5058 ), .B(\Reg_Bank/n5057 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5059 ) );
  MUX \Reg_Bank/U5125  ( .A(\Reg_Bank/registers[12][2] ), .B(
        \Reg_Bank/registers[13][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5058 ) );
  MUX \Reg_Bank/U5124  ( .A(\Reg_Bank/registers[14][2] ), .B(
        \Reg_Bank/registers[15][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5057 ) );
  MUX \Reg_Bank/U5123  ( .A(\Reg_Bank/n5055 ), .B(\Reg_Bank/n5048 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5056 ) );
  MUX \Reg_Bank/U5122  ( .A(\Reg_Bank/n5054 ), .B(\Reg_Bank/n5051 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5055 ) );
  MUX \Reg_Bank/U5121  ( .A(\Reg_Bank/n5053 ), .B(\Reg_Bank/n5052 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5054 ) );
  MUX \Reg_Bank/U5120  ( .A(\Reg_Bank/registers[16][2] ), .B(
        \Reg_Bank/registers[17][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5053 ) );
  MUX \Reg_Bank/U5119  ( .A(\Reg_Bank/registers[18][2] ), .B(
        \Reg_Bank/registers[19][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5052 ) );
  MUX \Reg_Bank/U5118  ( .A(\Reg_Bank/n5050 ), .B(\Reg_Bank/n5049 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5051 ) );
  MUX \Reg_Bank/U5117  ( .A(\Reg_Bank/registers[20][2] ), .B(
        \Reg_Bank/registers[21][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5050 ) );
  MUX \Reg_Bank/U5116  ( .A(\Reg_Bank/registers[22][2] ), .B(
        \Reg_Bank/registers[23][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5049 ) );
  MUX \Reg_Bank/U5115  ( .A(\Reg_Bank/n5047 ), .B(\Reg_Bank/n5044 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5048 ) );
  MUX \Reg_Bank/U5114  ( .A(\Reg_Bank/n5046 ), .B(\Reg_Bank/n5045 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5047 ) );
  MUX \Reg_Bank/U5113  ( .A(\Reg_Bank/registers[24][2] ), .B(
        \Reg_Bank/registers[25][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5046 ) );
  MUX \Reg_Bank/U5112  ( .A(\Reg_Bank/registers[26][2] ), .B(
        \Reg_Bank/registers[27][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5045 ) );
  MUX \Reg_Bank/U5111  ( .A(\Reg_Bank/n5043 ), .B(\Reg_Bank/n5042 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5044 ) );
  MUX \Reg_Bank/U5110  ( .A(\Reg_Bank/registers[28][2] ), .B(
        \Reg_Bank/registers[29][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5043 ) );
  MUX \Reg_Bank/U5109  ( .A(\Reg_Bank/registers[30][2] ), .B(
        \Reg_Bank/registers[31][2] ), .S(rt_index[0]), .Z(\Reg_Bank/n5042 ) );
  MUX \Reg_Bank/U5108  ( .A(\Reg_Bank/n5041 ), .B(\Reg_Bank/n5026 ), .S(
        rt_index[4]), .Z(reg_target[1]) );
  MUX \Reg_Bank/U5107  ( .A(\Reg_Bank/n5040 ), .B(\Reg_Bank/n5033 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5041 ) );
  MUX \Reg_Bank/U5106  ( .A(\Reg_Bank/n5039 ), .B(\Reg_Bank/n5036 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5040 ) );
  MUX \Reg_Bank/U5105  ( .A(\Reg_Bank/n5038 ), .B(\Reg_Bank/n5037 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5039 ) );
  MUX \Reg_Bank/U5103  ( .A(\Reg_Bank/registers[2][1] ), .B(
        \Reg_Bank/registers[3][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5037 ) );
  MUX \Reg_Bank/U5102  ( .A(\Reg_Bank/n5035 ), .B(\Reg_Bank/n5034 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5036 ) );
  MUX \Reg_Bank/U5101  ( .A(\Reg_Bank/registers[4][1] ), .B(
        \Reg_Bank/registers[5][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5035 ) );
  MUX \Reg_Bank/U5100  ( .A(\Reg_Bank/registers[6][1] ), .B(
        \Reg_Bank/registers[7][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5034 ) );
  MUX \Reg_Bank/U5099  ( .A(\Reg_Bank/n5032 ), .B(\Reg_Bank/n5029 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5033 ) );
  MUX \Reg_Bank/U5098  ( .A(\Reg_Bank/n5031 ), .B(\Reg_Bank/n5030 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5032 ) );
  MUX \Reg_Bank/U5097  ( .A(\Reg_Bank/registers[8][1] ), .B(
        \Reg_Bank/registers[9][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5031 ) );
  MUX \Reg_Bank/U5096  ( .A(\Reg_Bank/registers[10][1] ), .B(
        \Reg_Bank/registers[11][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5030 ) );
  MUX \Reg_Bank/U5095  ( .A(\Reg_Bank/n5028 ), .B(\Reg_Bank/n5027 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5029 ) );
  MUX \Reg_Bank/U5094  ( .A(\Reg_Bank/registers[12][1] ), .B(
        \Reg_Bank/registers[13][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5028 ) );
  MUX \Reg_Bank/U5093  ( .A(\Reg_Bank/registers[14][1] ), .B(
        \Reg_Bank/registers[15][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5027 ) );
  MUX \Reg_Bank/U5092  ( .A(\Reg_Bank/n5025 ), .B(\Reg_Bank/n5018 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5026 ) );
  MUX \Reg_Bank/U5091  ( .A(\Reg_Bank/n5024 ), .B(\Reg_Bank/n5021 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5025 ) );
  MUX \Reg_Bank/U5090  ( .A(\Reg_Bank/n5023 ), .B(\Reg_Bank/n5022 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5024 ) );
  MUX \Reg_Bank/U5089  ( .A(\Reg_Bank/registers[16][1] ), .B(
        \Reg_Bank/registers[17][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5023 ) );
  MUX \Reg_Bank/U5088  ( .A(\Reg_Bank/registers[18][1] ), .B(
        \Reg_Bank/registers[19][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5022 ) );
  MUX \Reg_Bank/U5087  ( .A(\Reg_Bank/n5020 ), .B(\Reg_Bank/n5019 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5021 ) );
  MUX \Reg_Bank/U5086  ( .A(\Reg_Bank/registers[20][1] ), .B(
        \Reg_Bank/registers[21][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5020 ) );
  MUX \Reg_Bank/U5085  ( .A(\Reg_Bank/registers[22][1] ), .B(
        \Reg_Bank/registers[23][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5019 ) );
  MUX \Reg_Bank/U5084  ( .A(\Reg_Bank/n5017 ), .B(\Reg_Bank/n5014 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5018 ) );
  MUX \Reg_Bank/U5083  ( .A(\Reg_Bank/n5016 ), .B(\Reg_Bank/n5015 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5017 ) );
  MUX \Reg_Bank/U5082  ( .A(\Reg_Bank/registers[24][1] ), .B(
        \Reg_Bank/registers[25][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5016 ) );
  MUX \Reg_Bank/U5081  ( .A(\Reg_Bank/registers[26][1] ), .B(
        \Reg_Bank/registers[27][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5015 ) );
  MUX \Reg_Bank/U5080  ( .A(\Reg_Bank/n5013 ), .B(\Reg_Bank/n5012 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5014 ) );
  MUX \Reg_Bank/U5079  ( .A(\Reg_Bank/registers[28][1] ), .B(
        \Reg_Bank/registers[29][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5013 ) );
  MUX \Reg_Bank/U5078  ( .A(\Reg_Bank/registers[30][1] ), .B(
        \Reg_Bank/registers[31][1] ), .S(rt_index[0]), .Z(\Reg_Bank/n5012 ) );
  MUX \Reg_Bank/U5077  ( .A(\Reg_Bank/n5011 ), .B(\Reg_Bank/n4996 ), .S(
        rt_index[4]), .Z(reg_target[0]) );
  MUX \Reg_Bank/U5076  ( .A(\Reg_Bank/n5010 ), .B(\Reg_Bank/n5003 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n5011 ) );
  MUX \Reg_Bank/U5075  ( .A(\Reg_Bank/n5009 ), .B(\Reg_Bank/n5006 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5010 ) );
  MUX \Reg_Bank/U5074  ( .A(\Reg_Bank/n5008 ), .B(\Reg_Bank/n5007 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5009 ) );
  MUX \Reg_Bank/U5072  ( .A(\Reg_Bank/registers[2][0] ), .B(
        \Reg_Bank/registers[3][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n5007 ) );
  MUX \Reg_Bank/U5071  ( .A(\Reg_Bank/n5005 ), .B(\Reg_Bank/n5004 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5006 ) );
  MUX \Reg_Bank/U5070  ( .A(\Reg_Bank/registers[4][0] ), .B(
        \Reg_Bank/registers[5][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n5005 ) );
  MUX \Reg_Bank/U5069  ( .A(\Reg_Bank/registers[6][0] ), .B(
        \Reg_Bank/registers[7][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n5004 ) );
  MUX \Reg_Bank/U5068  ( .A(\Reg_Bank/n5002 ), .B(\Reg_Bank/n4999 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n5003 ) );
  MUX \Reg_Bank/U5067  ( .A(\Reg_Bank/n5001 ), .B(\Reg_Bank/n5000 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n5002 ) );
  MUX \Reg_Bank/U5066  ( .A(\Reg_Bank/registers[8][0] ), .B(
        \Reg_Bank/registers[9][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n5001 ) );
  MUX \Reg_Bank/U5065  ( .A(\Reg_Bank/registers[10][0] ), .B(
        \Reg_Bank/registers[11][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n5000 ) );
  MUX \Reg_Bank/U5064  ( .A(\Reg_Bank/n4998 ), .B(\Reg_Bank/n4997 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n4999 ) );
  MUX \Reg_Bank/U5063  ( .A(\Reg_Bank/registers[12][0] ), .B(
        \Reg_Bank/registers[13][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4998 ) );
  MUX \Reg_Bank/U5062  ( .A(\Reg_Bank/registers[14][0] ), .B(
        \Reg_Bank/registers[15][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4997 ) );
  MUX \Reg_Bank/U5061  ( .A(\Reg_Bank/n4995 ), .B(\Reg_Bank/n4988 ), .S(
        rt_index[3]), .Z(\Reg_Bank/n4996 ) );
  MUX \Reg_Bank/U5060  ( .A(\Reg_Bank/n4994 ), .B(\Reg_Bank/n4991 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n4995 ) );
  MUX \Reg_Bank/U5059  ( .A(\Reg_Bank/n4993 ), .B(\Reg_Bank/n4992 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n4994 ) );
  MUX \Reg_Bank/U5058  ( .A(\Reg_Bank/registers[16][0] ), .B(
        \Reg_Bank/registers[17][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4993 ) );
  MUX \Reg_Bank/U5057  ( .A(\Reg_Bank/registers[18][0] ), .B(
        \Reg_Bank/registers[19][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4992 ) );
  MUX \Reg_Bank/U5056  ( .A(\Reg_Bank/n4990 ), .B(\Reg_Bank/n4989 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n4991 ) );
  MUX \Reg_Bank/U5055  ( .A(\Reg_Bank/registers[20][0] ), .B(
        \Reg_Bank/registers[21][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4990 ) );
  MUX \Reg_Bank/U5054  ( .A(\Reg_Bank/registers[22][0] ), .B(
        \Reg_Bank/registers[23][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4989 ) );
  MUX \Reg_Bank/U5053  ( .A(\Reg_Bank/n4987 ), .B(\Reg_Bank/n4984 ), .S(
        rt_index[2]), .Z(\Reg_Bank/n4988 ) );
  MUX \Reg_Bank/U5052  ( .A(\Reg_Bank/n4986 ), .B(\Reg_Bank/n4985 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n4987 ) );
  MUX \Reg_Bank/U5051  ( .A(\Reg_Bank/registers[24][0] ), .B(
        \Reg_Bank/registers[25][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4986 ) );
  MUX \Reg_Bank/U5050  ( .A(\Reg_Bank/registers[26][0] ), .B(
        \Reg_Bank/registers[27][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4985 ) );
  MUX \Reg_Bank/U5049  ( .A(\Reg_Bank/n4983 ), .B(\Reg_Bank/n4982 ), .S(
        rt_index[1]), .Z(\Reg_Bank/n4984 ) );
  MUX \Reg_Bank/U5048  ( .A(\Reg_Bank/registers[28][0] ), .B(
        \Reg_Bank/registers[29][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4983 ) );
  MUX \Reg_Bank/U5047  ( .A(\Reg_Bank/registers[30][0] ), .B(
        \Reg_Bank/registers[31][0] ), .S(rt_index[0]), .Z(\Reg_Bank/n4982 ) );
  MUX \Reg_Bank/U5046  ( .A(\Reg_Bank/n4981 ), .B(\Reg_Bank/n4966 ), .S(
        rs_index[4]), .Z(reg_source[31]) );
  MUX \Reg_Bank/U5045  ( .A(\Reg_Bank/n4980 ), .B(\Reg_Bank/n4973 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4981 ) );
  MUX \Reg_Bank/U5044  ( .A(\Reg_Bank/n4979 ), .B(\Reg_Bank/n4976 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4980 ) );
  MUX \Reg_Bank/U5043  ( .A(\Reg_Bank/n4978 ), .B(\Reg_Bank/n4977 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4979 ) );
  MUX \Reg_Bank/U5041  ( .A(\Reg_Bank/registers[2][31] ), .B(
        \Reg_Bank/registers[3][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4977 ) );
  MUX \Reg_Bank/U5040  ( .A(\Reg_Bank/n4975 ), .B(\Reg_Bank/n4974 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4976 ) );
  MUX \Reg_Bank/U5039  ( .A(\Reg_Bank/registers[4][31] ), .B(
        \Reg_Bank/registers[5][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4975 ) );
  MUX \Reg_Bank/U5038  ( .A(\Reg_Bank/registers[6][31] ), .B(
        \Reg_Bank/registers[7][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4974 ) );
  MUX \Reg_Bank/U5037  ( .A(\Reg_Bank/n4972 ), .B(\Reg_Bank/n4969 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4973 ) );
  MUX \Reg_Bank/U5036  ( .A(\Reg_Bank/n4971 ), .B(\Reg_Bank/n4970 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4972 ) );
  MUX \Reg_Bank/U5035  ( .A(\Reg_Bank/registers[8][31] ), .B(
        \Reg_Bank/registers[9][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4971 ) );
  MUX \Reg_Bank/U5034  ( .A(\Reg_Bank/registers[10][31] ), .B(
        \Reg_Bank/registers[11][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4970 )
         );
  MUX \Reg_Bank/U5033  ( .A(\Reg_Bank/n4968 ), .B(\Reg_Bank/n4967 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4969 ) );
  MUX \Reg_Bank/U5032  ( .A(\Reg_Bank/registers[12][31] ), .B(
        \Reg_Bank/registers[13][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4968 )
         );
  MUX \Reg_Bank/U5031  ( .A(\Reg_Bank/registers[14][31] ), .B(
        \Reg_Bank/registers[15][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4967 )
         );
  MUX \Reg_Bank/U5030  ( .A(\Reg_Bank/n4965 ), .B(\Reg_Bank/n4958 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4966 ) );
  MUX \Reg_Bank/U5029  ( .A(\Reg_Bank/n4964 ), .B(\Reg_Bank/n4961 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4965 ) );
  MUX \Reg_Bank/U5028  ( .A(\Reg_Bank/n4963 ), .B(\Reg_Bank/n4962 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4964 ) );
  MUX \Reg_Bank/U5027  ( .A(\Reg_Bank/registers[16][31] ), .B(
        \Reg_Bank/registers[17][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4963 )
         );
  MUX \Reg_Bank/U5026  ( .A(\Reg_Bank/registers[18][31] ), .B(
        \Reg_Bank/registers[19][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4962 )
         );
  MUX \Reg_Bank/U5025  ( .A(\Reg_Bank/n4960 ), .B(\Reg_Bank/n4959 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4961 ) );
  MUX \Reg_Bank/U5024  ( .A(\Reg_Bank/registers[20][31] ), .B(
        \Reg_Bank/registers[21][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4960 )
         );
  MUX \Reg_Bank/U5023  ( .A(\Reg_Bank/registers[22][31] ), .B(
        \Reg_Bank/registers[23][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4959 )
         );
  MUX \Reg_Bank/U5022  ( .A(\Reg_Bank/n4957 ), .B(\Reg_Bank/n4954 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4958 ) );
  MUX \Reg_Bank/U5021  ( .A(\Reg_Bank/n4956 ), .B(\Reg_Bank/n4955 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4957 ) );
  MUX \Reg_Bank/U5020  ( .A(\Reg_Bank/registers[24][31] ), .B(
        \Reg_Bank/registers[25][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4956 )
         );
  MUX \Reg_Bank/U5019  ( .A(\Reg_Bank/registers[26][31] ), .B(
        \Reg_Bank/registers[27][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4955 )
         );
  MUX \Reg_Bank/U5018  ( .A(\Reg_Bank/n4953 ), .B(\Reg_Bank/n4952 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4954 ) );
  MUX \Reg_Bank/U5017  ( .A(\Reg_Bank/registers[28][31] ), .B(
        \Reg_Bank/registers[29][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4953 )
         );
  MUX \Reg_Bank/U5016  ( .A(\Reg_Bank/registers[30][31] ), .B(
        \Reg_Bank/registers[31][31] ), .S(rs_index[0]), .Z(\Reg_Bank/n4952 )
         );
  MUX \Reg_Bank/U5015  ( .A(\Reg_Bank/n4951 ), .B(\Reg_Bank/n4936 ), .S(
        rs_index[4]), .Z(reg_source[30]) );
  MUX \Reg_Bank/U5014  ( .A(\Reg_Bank/n4950 ), .B(\Reg_Bank/n4943 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4951 ) );
  MUX \Reg_Bank/U5013  ( .A(\Reg_Bank/n4949 ), .B(\Reg_Bank/n4946 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4950 ) );
  MUX \Reg_Bank/U5012  ( .A(\Reg_Bank/n4948 ), .B(\Reg_Bank/n4947 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4949 ) );
  MUX \Reg_Bank/U5010  ( .A(\Reg_Bank/registers[2][30] ), .B(
        \Reg_Bank/registers[3][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4947 ) );
  MUX \Reg_Bank/U5009  ( .A(\Reg_Bank/n4945 ), .B(\Reg_Bank/n4944 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4946 ) );
  MUX \Reg_Bank/U5008  ( .A(\Reg_Bank/registers[4][30] ), .B(
        \Reg_Bank/registers[5][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4945 ) );
  MUX \Reg_Bank/U5007  ( .A(\Reg_Bank/registers[6][30] ), .B(
        \Reg_Bank/registers[7][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4944 ) );
  MUX \Reg_Bank/U5006  ( .A(\Reg_Bank/n4942 ), .B(\Reg_Bank/n4939 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4943 ) );
  MUX \Reg_Bank/U5005  ( .A(\Reg_Bank/n4941 ), .B(\Reg_Bank/n4940 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4942 ) );
  MUX \Reg_Bank/U5004  ( .A(\Reg_Bank/registers[8][30] ), .B(
        \Reg_Bank/registers[9][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4941 ) );
  MUX \Reg_Bank/U5003  ( .A(\Reg_Bank/registers[10][30] ), .B(
        \Reg_Bank/registers[11][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4940 )
         );
  MUX \Reg_Bank/U5002  ( .A(\Reg_Bank/n4938 ), .B(\Reg_Bank/n4937 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4939 ) );
  MUX \Reg_Bank/U5001  ( .A(\Reg_Bank/registers[12][30] ), .B(
        \Reg_Bank/registers[13][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4938 )
         );
  MUX \Reg_Bank/U5000  ( .A(\Reg_Bank/registers[14][30] ), .B(
        \Reg_Bank/registers[15][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4937 )
         );
  MUX \Reg_Bank/U4999  ( .A(\Reg_Bank/n4935 ), .B(\Reg_Bank/n4928 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4936 ) );
  MUX \Reg_Bank/U4998  ( .A(\Reg_Bank/n4934 ), .B(\Reg_Bank/n4931 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4935 ) );
  MUX \Reg_Bank/U4997  ( .A(\Reg_Bank/n4933 ), .B(\Reg_Bank/n4932 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4934 ) );
  MUX \Reg_Bank/U4996  ( .A(\Reg_Bank/registers[16][30] ), .B(
        \Reg_Bank/registers[17][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4933 )
         );
  MUX \Reg_Bank/U4995  ( .A(\Reg_Bank/registers[18][30] ), .B(
        \Reg_Bank/registers[19][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4932 )
         );
  MUX \Reg_Bank/U4994  ( .A(\Reg_Bank/n4930 ), .B(\Reg_Bank/n4929 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4931 ) );
  MUX \Reg_Bank/U4993  ( .A(\Reg_Bank/registers[20][30] ), .B(
        \Reg_Bank/registers[21][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4930 )
         );
  MUX \Reg_Bank/U4992  ( .A(\Reg_Bank/registers[22][30] ), .B(
        \Reg_Bank/registers[23][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4929 )
         );
  MUX \Reg_Bank/U4991  ( .A(\Reg_Bank/n4927 ), .B(\Reg_Bank/n4924 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4928 ) );
  MUX \Reg_Bank/U4990  ( .A(\Reg_Bank/n4926 ), .B(\Reg_Bank/n4925 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4927 ) );
  MUX \Reg_Bank/U4989  ( .A(\Reg_Bank/registers[24][30] ), .B(
        \Reg_Bank/registers[25][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4926 )
         );
  MUX \Reg_Bank/U4988  ( .A(\Reg_Bank/registers[26][30] ), .B(
        \Reg_Bank/registers[27][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4925 )
         );
  MUX \Reg_Bank/U4987  ( .A(\Reg_Bank/n4923 ), .B(\Reg_Bank/n4922 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4924 ) );
  MUX \Reg_Bank/U4986  ( .A(\Reg_Bank/registers[28][30] ), .B(
        \Reg_Bank/registers[29][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4923 )
         );
  MUX \Reg_Bank/U4985  ( .A(\Reg_Bank/registers[30][30] ), .B(
        \Reg_Bank/registers[31][30] ), .S(rs_index[0]), .Z(\Reg_Bank/n4922 )
         );
  MUX \Reg_Bank/U4984  ( .A(\Reg_Bank/n4921 ), .B(\Reg_Bank/n4906 ), .S(
        rs_index[4]), .Z(reg_source[29]) );
  MUX \Reg_Bank/U4983  ( .A(\Reg_Bank/n4920 ), .B(\Reg_Bank/n4913 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4921 ) );
  MUX \Reg_Bank/U4982  ( .A(\Reg_Bank/n4919 ), .B(\Reg_Bank/n4916 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4920 ) );
  MUX \Reg_Bank/U4981  ( .A(\Reg_Bank/n4918 ), .B(\Reg_Bank/n4917 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4919 ) );
  MUX \Reg_Bank/U4979  ( .A(\Reg_Bank/registers[2][29] ), .B(
        \Reg_Bank/registers[3][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4917 ) );
  MUX \Reg_Bank/U4978  ( .A(\Reg_Bank/n4915 ), .B(\Reg_Bank/n4914 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4916 ) );
  MUX \Reg_Bank/U4977  ( .A(\Reg_Bank/registers[4][29] ), .B(
        \Reg_Bank/registers[5][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4915 ) );
  MUX \Reg_Bank/U4976  ( .A(\Reg_Bank/registers[6][29] ), .B(
        \Reg_Bank/registers[7][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4914 ) );
  MUX \Reg_Bank/U4975  ( .A(\Reg_Bank/n4912 ), .B(\Reg_Bank/n4909 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4913 ) );
  MUX \Reg_Bank/U4974  ( .A(\Reg_Bank/n4911 ), .B(\Reg_Bank/n4910 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4912 ) );
  MUX \Reg_Bank/U4973  ( .A(\Reg_Bank/registers[8][29] ), .B(
        \Reg_Bank/registers[9][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4911 ) );
  MUX \Reg_Bank/U4972  ( .A(\Reg_Bank/registers[10][29] ), .B(
        \Reg_Bank/registers[11][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4910 )
         );
  MUX \Reg_Bank/U4971  ( .A(\Reg_Bank/n4908 ), .B(\Reg_Bank/n4907 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4909 ) );
  MUX \Reg_Bank/U4970  ( .A(\Reg_Bank/registers[12][29] ), .B(
        \Reg_Bank/registers[13][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4908 )
         );
  MUX \Reg_Bank/U4969  ( .A(\Reg_Bank/registers[14][29] ), .B(
        \Reg_Bank/registers[15][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4907 )
         );
  MUX \Reg_Bank/U4968  ( .A(\Reg_Bank/n4905 ), .B(\Reg_Bank/n4898 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4906 ) );
  MUX \Reg_Bank/U4967  ( .A(\Reg_Bank/n4904 ), .B(\Reg_Bank/n4901 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4905 ) );
  MUX \Reg_Bank/U4966  ( .A(\Reg_Bank/n4903 ), .B(\Reg_Bank/n4902 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4904 ) );
  MUX \Reg_Bank/U4965  ( .A(\Reg_Bank/registers[16][29] ), .B(
        \Reg_Bank/registers[17][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4903 )
         );
  MUX \Reg_Bank/U4964  ( .A(\Reg_Bank/registers[18][29] ), .B(
        \Reg_Bank/registers[19][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4902 )
         );
  MUX \Reg_Bank/U4963  ( .A(\Reg_Bank/n4900 ), .B(\Reg_Bank/n4899 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4901 ) );
  MUX \Reg_Bank/U4962  ( .A(\Reg_Bank/registers[20][29] ), .B(
        \Reg_Bank/registers[21][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4900 )
         );
  MUX \Reg_Bank/U4961  ( .A(\Reg_Bank/registers[22][29] ), .B(
        \Reg_Bank/registers[23][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4899 )
         );
  MUX \Reg_Bank/U4960  ( .A(\Reg_Bank/n4897 ), .B(\Reg_Bank/n4894 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4898 ) );
  MUX \Reg_Bank/U4959  ( .A(\Reg_Bank/n4896 ), .B(\Reg_Bank/n4895 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4897 ) );
  MUX \Reg_Bank/U4958  ( .A(\Reg_Bank/registers[24][29] ), .B(
        \Reg_Bank/registers[25][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4896 )
         );
  MUX \Reg_Bank/U4957  ( .A(\Reg_Bank/registers[26][29] ), .B(
        \Reg_Bank/registers[27][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4895 )
         );
  MUX \Reg_Bank/U4956  ( .A(\Reg_Bank/n4893 ), .B(\Reg_Bank/n4892 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4894 ) );
  MUX \Reg_Bank/U4955  ( .A(\Reg_Bank/registers[28][29] ), .B(
        \Reg_Bank/registers[29][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4893 )
         );
  MUX \Reg_Bank/U4954  ( .A(\Reg_Bank/registers[30][29] ), .B(
        \Reg_Bank/registers[31][29] ), .S(rs_index[0]), .Z(\Reg_Bank/n4892 )
         );
  MUX \Reg_Bank/U4953  ( .A(\Reg_Bank/n4891 ), .B(\Reg_Bank/n4876 ), .S(
        rs_index[4]), .Z(reg_source[28]) );
  MUX \Reg_Bank/U4952  ( .A(\Reg_Bank/n4890 ), .B(\Reg_Bank/n4883 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4891 ) );
  MUX \Reg_Bank/U4951  ( .A(\Reg_Bank/n4889 ), .B(\Reg_Bank/n4886 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4890 ) );
  MUX \Reg_Bank/U4950  ( .A(\Reg_Bank/n4888 ), .B(\Reg_Bank/n4887 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4889 ) );
  MUX \Reg_Bank/U4948  ( .A(\Reg_Bank/registers[2][28] ), .B(
        \Reg_Bank/registers[3][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4887 ) );
  MUX \Reg_Bank/U4947  ( .A(\Reg_Bank/n4885 ), .B(\Reg_Bank/n4884 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4886 ) );
  MUX \Reg_Bank/U4946  ( .A(\Reg_Bank/registers[4][28] ), .B(
        \Reg_Bank/registers[5][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4885 ) );
  MUX \Reg_Bank/U4945  ( .A(\Reg_Bank/registers[6][28] ), .B(
        \Reg_Bank/registers[7][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4884 ) );
  MUX \Reg_Bank/U4944  ( .A(\Reg_Bank/n4882 ), .B(\Reg_Bank/n4879 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4883 ) );
  MUX \Reg_Bank/U4943  ( .A(\Reg_Bank/n4881 ), .B(\Reg_Bank/n4880 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4882 ) );
  MUX \Reg_Bank/U4942  ( .A(\Reg_Bank/registers[8][28] ), .B(
        \Reg_Bank/registers[9][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4881 ) );
  MUX \Reg_Bank/U4941  ( .A(\Reg_Bank/registers[10][28] ), .B(
        \Reg_Bank/registers[11][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4880 )
         );
  MUX \Reg_Bank/U4940  ( .A(\Reg_Bank/n4878 ), .B(\Reg_Bank/n4877 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4879 ) );
  MUX \Reg_Bank/U4939  ( .A(\Reg_Bank/registers[12][28] ), .B(
        \Reg_Bank/registers[13][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4878 )
         );
  MUX \Reg_Bank/U4938  ( .A(\Reg_Bank/registers[14][28] ), .B(
        \Reg_Bank/registers[15][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4877 )
         );
  MUX \Reg_Bank/U4937  ( .A(\Reg_Bank/n4875 ), .B(\Reg_Bank/n4868 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4876 ) );
  MUX \Reg_Bank/U4936  ( .A(\Reg_Bank/n4874 ), .B(\Reg_Bank/n4871 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4875 ) );
  MUX \Reg_Bank/U4935  ( .A(\Reg_Bank/n4873 ), .B(\Reg_Bank/n4872 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4874 ) );
  MUX \Reg_Bank/U4934  ( .A(\Reg_Bank/registers[16][28] ), .B(
        \Reg_Bank/registers[17][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4873 )
         );
  MUX \Reg_Bank/U4933  ( .A(\Reg_Bank/registers[18][28] ), .B(
        \Reg_Bank/registers[19][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4872 )
         );
  MUX \Reg_Bank/U4932  ( .A(\Reg_Bank/n4870 ), .B(\Reg_Bank/n4869 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4871 ) );
  MUX \Reg_Bank/U4931  ( .A(\Reg_Bank/registers[20][28] ), .B(
        \Reg_Bank/registers[21][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4870 )
         );
  MUX \Reg_Bank/U4930  ( .A(\Reg_Bank/registers[22][28] ), .B(
        \Reg_Bank/registers[23][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4869 )
         );
  MUX \Reg_Bank/U4929  ( .A(\Reg_Bank/n4867 ), .B(\Reg_Bank/n4864 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4868 ) );
  MUX \Reg_Bank/U4928  ( .A(\Reg_Bank/n4866 ), .B(\Reg_Bank/n4865 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4867 ) );
  MUX \Reg_Bank/U4927  ( .A(\Reg_Bank/registers[24][28] ), .B(
        \Reg_Bank/registers[25][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4866 )
         );
  MUX \Reg_Bank/U4926  ( .A(\Reg_Bank/registers[26][28] ), .B(
        \Reg_Bank/registers[27][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4865 )
         );
  MUX \Reg_Bank/U4925  ( .A(\Reg_Bank/n4863 ), .B(\Reg_Bank/n4862 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4864 ) );
  MUX \Reg_Bank/U4924  ( .A(\Reg_Bank/registers[28][28] ), .B(
        \Reg_Bank/registers[29][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4863 )
         );
  MUX \Reg_Bank/U4923  ( .A(\Reg_Bank/registers[30][28] ), .B(
        \Reg_Bank/registers[31][28] ), .S(rs_index[0]), .Z(\Reg_Bank/n4862 )
         );
  MUX \Reg_Bank/U4922  ( .A(\Reg_Bank/n4861 ), .B(\Reg_Bank/n4846 ), .S(
        rs_index[4]), .Z(reg_source[27]) );
  MUX \Reg_Bank/U4921  ( .A(\Reg_Bank/n4860 ), .B(\Reg_Bank/n4853 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4861 ) );
  MUX \Reg_Bank/U4920  ( .A(\Reg_Bank/n4859 ), .B(\Reg_Bank/n4856 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4860 ) );
  MUX \Reg_Bank/U4919  ( .A(\Reg_Bank/n4858 ), .B(\Reg_Bank/n4857 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4859 ) );
  MUX \Reg_Bank/U4917  ( .A(\Reg_Bank/registers[2][27] ), .B(
        \Reg_Bank/registers[3][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4857 ) );
  MUX \Reg_Bank/U4916  ( .A(\Reg_Bank/n4855 ), .B(\Reg_Bank/n4854 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4856 ) );
  MUX \Reg_Bank/U4915  ( .A(\Reg_Bank/registers[4][27] ), .B(
        \Reg_Bank/registers[5][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4855 ) );
  MUX \Reg_Bank/U4914  ( .A(\Reg_Bank/registers[6][27] ), .B(
        \Reg_Bank/registers[7][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4854 ) );
  MUX \Reg_Bank/U4913  ( .A(\Reg_Bank/n4852 ), .B(\Reg_Bank/n4849 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4853 ) );
  MUX \Reg_Bank/U4912  ( .A(\Reg_Bank/n4851 ), .B(\Reg_Bank/n4850 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4852 ) );
  MUX \Reg_Bank/U4911  ( .A(\Reg_Bank/registers[8][27] ), .B(
        \Reg_Bank/registers[9][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4851 ) );
  MUX \Reg_Bank/U4910  ( .A(\Reg_Bank/registers[10][27] ), .B(
        \Reg_Bank/registers[11][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4850 )
         );
  MUX \Reg_Bank/U4909  ( .A(\Reg_Bank/n4848 ), .B(\Reg_Bank/n4847 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4849 ) );
  MUX \Reg_Bank/U4908  ( .A(\Reg_Bank/registers[12][27] ), .B(
        \Reg_Bank/registers[13][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4848 )
         );
  MUX \Reg_Bank/U4907  ( .A(\Reg_Bank/registers[14][27] ), .B(
        \Reg_Bank/registers[15][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4847 )
         );
  MUX \Reg_Bank/U4906  ( .A(\Reg_Bank/n4845 ), .B(\Reg_Bank/n4838 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4846 ) );
  MUX \Reg_Bank/U4905  ( .A(\Reg_Bank/n4844 ), .B(\Reg_Bank/n4841 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4845 ) );
  MUX \Reg_Bank/U4904  ( .A(\Reg_Bank/n4843 ), .B(\Reg_Bank/n4842 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4844 ) );
  MUX \Reg_Bank/U4903  ( .A(\Reg_Bank/registers[16][27] ), .B(
        \Reg_Bank/registers[17][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4843 )
         );
  MUX \Reg_Bank/U4902  ( .A(\Reg_Bank/registers[18][27] ), .B(
        \Reg_Bank/registers[19][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4842 )
         );
  MUX \Reg_Bank/U4901  ( .A(\Reg_Bank/n4840 ), .B(\Reg_Bank/n4839 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4841 ) );
  MUX \Reg_Bank/U4900  ( .A(\Reg_Bank/registers[20][27] ), .B(
        \Reg_Bank/registers[21][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4840 )
         );
  MUX \Reg_Bank/U4899  ( .A(\Reg_Bank/registers[22][27] ), .B(
        \Reg_Bank/registers[23][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4839 )
         );
  MUX \Reg_Bank/U4898  ( .A(\Reg_Bank/n4837 ), .B(\Reg_Bank/n4834 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4838 ) );
  MUX \Reg_Bank/U4897  ( .A(\Reg_Bank/n4836 ), .B(\Reg_Bank/n4835 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4837 ) );
  MUX \Reg_Bank/U4896  ( .A(\Reg_Bank/registers[24][27] ), .B(
        \Reg_Bank/registers[25][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4836 )
         );
  MUX \Reg_Bank/U4895  ( .A(\Reg_Bank/registers[26][27] ), .B(
        \Reg_Bank/registers[27][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4835 )
         );
  MUX \Reg_Bank/U4894  ( .A(\Reg_Bank/n4833 ), .B(\Reg_Bank/n4832 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4834 ) );
  MUX \Reg_Bank/U4893  ( .A(\Reg_Bank/registers[28][27] ), .B(
        \Reg_Bank/registers[29][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4833 )
         );
  MUX \Reg_Bank/U4892  ( .A(\Reg_Bank/registers[30][27] ), .B(
        \Reg_Bank/registers[31][27] ), .S(rs_index[0]), .Z(\Reg_Bank/n4832 )
         );
  MUX \Reg_Bank/U4891  ( .A(\Reg_Bank/n4831 ), .B(\Reg_Bank/n4816 ), .S(
        rs_index[4]), .Z(reg_source[26]) );
  MUX \Reg_Bank/U4890  ( .A(\Reg_Bank/n4830 ), .B(\Reg_Bank/n4823 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4831 ) );
  MUX \Reg_Bank/U4889  ( .A(\Reg_Bank/n4829 ), .B(\Reg_Bank/n4826 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4830 ) );
  MUX \Reg_Bank/U4888  ( .A(\Reg_Bank/n4828 ), .B(\Reg_Bank/n4827 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4829 ) );
  MUX \Reg_Bank/U4886  ( .A(\Reg_Bank/registers[2][26] ), .B(
        \Reg_Bank/registers[3][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4827 ) );
  MUX \Reg_Bank/U4885  ( .A(\Reg_Bank/n4825 ), .B(\Reg_Bank/n4824 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4826 ) );
  MUX \Reg_Bank/U4884  ( .A(\Reg_Bank/registers[4][26] ), .B(
        \Reg_Bank/registers[5][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4825 ) );
  MUX \Reg_Bank/U4883  ( .A(\Reg_Bank/registers[6][26] ), .B(
        \Reg_Bank/registers[7][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4824 ) );
  MUX \Reg_Bank/U4882  ( .A(\Reg_Bank/n4822 ), .B(\Reg_Bank/n4819 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4823 ) );
  MUX \Reg_Bank/U4881  ( .A(\Reg_Bank/n4821 ), .B(\Reg_Bank/n4820 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4822 ) );
  MUX \Reg_Bank/U4880  ( .A(\Reg_Bank/registers[8][26] ), .B(
        \Reg_Bank/registers[9][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4821 ) );
  MUX \Reg_Bank/U4879  ( .A(\Reg_Bank/registers[10][26] ), .B(
        \Reg_Bank/registers[11][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4820 )
         );
  MUX \Reg_Bank/U4878  ( .A(\Reg_Bank/n4818 ), .B(\Reg_Bank/n4817 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4819 ) );
  MUX \Reg_Bank/U4877  ( .A(\Reg_Bank/registers[12][26] ), .B(
        \Reg_Bank/registers[13][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4818 )
         );
  MUX \Reg_Bank/U4876  ( .A(\Reg_Bank/registers[14][26] ), .B(
        \Reg_Bank/registers[15][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4817 )
         );
  MUX \Reg_Bank/U4875  ( .A(\Reg_Bank/n4815 ), .B(\Reg_Bank/n4808 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4816 ) );
  MUX \Reg_Bank/U4874  ( .A(\Reg_Bank/n4814 ), .B(\Reg_Bank/n4811 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4815 ) );
  MUX \Reg_Bank/U4873  ( .A(\Reg_Bank/n4813 ), .B(\Reg_Bank/n4812 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4814 ) );
  MUX \Reg_Bank/U4872  ( .A(\Reg_Bank/registers[16][26] ), .B(
        \Reg_Bank/registers[17][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4813 )
         );
  MUX \Reg_Bank/U4871  ( .A(\Reg_Bank/registers[18][26] ), .B(
        \Reg_Bank/registers[19][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4812 )
         );
  MUX \Reg_Bank/U4870  ( .A(\Reg_Bank/n4810 ), .B(\Reg_Bank/n4809 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4811 ) );
  MUX \Reg_Bank/U4869  ( .A(\Reg_Bank/registers[20][26] ), .B(
        \Reg_Bank/registers[21][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4810 )
         );
  MUX \Reg_Bank/U4868  ( .A(\Reg_Bank/registers[22][26] ), .B(
        \Reg_Bank/registers[23][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4809 )
         );
  MUX \Reg_Bank/U4867  ( .A(\Reg_Bank/n4807 ), .B(\Reg_Bank/n4804 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4808 ) );
  MUX \Reg_Bank/U4866  ( .A(\Reg_Bank/n4806 ), .B(\Reg_Bank/n4805 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4807 ) );
  MUX \Reg_Bank/U4865  ( .A(\Reg_Bank/registers[24][26] ), .B(
        \Reg_Bank/registers[25][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4806 )
         );
  MUX \Reg_Bank/U4864  ( .A(\Reg_Bank/registers[26][26] ), .B(
        \Reg_Bank/registers[27][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4805 )
         );
  MUX \Reg_Bank/U4863  ( .A(\Reg_Bank/n4803 ), .B(\Reg_Bank/n4802 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4804 ) );
  MUX \Reg_Bank/U4862  ( .A(\Reg_Bank/registers[28][26] ), .B(
        \Reg_Bank/registers[29][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4803 )
         );
  MUX \Reg_Bank/U4861  ( .A(\Reg_Bank/registers[30][26] ), .B(
        \Reg_Bank/registers[31][26] ), .S(rs_index[0]), .Z(\Reg_Bank/n4802 )
         );
  MUX \Reg_Bank/U4860  ( .A(\Reg_Bank/n4801 ), .B(\Reg_Bank/n4786 ), .S(
        rs_index[4]), .Z(reg_source[25]) );
  MUX \Reg_Bank/U4859  ( .A(\Reg_Bank/n4800 ), .B(\Reg_Bank/n4793 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4801 ) );
  MUX \Reg_Bank/U4858  ( .A(\Reg_Bank/n4799 ), .B(\Reg_Bank/n4796 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4800 ) );
  MUX \Reg_Bank/U4857  ( .A(\Reg_Bank/n4798 ), .B(\Reg_Bank/n4797 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4799 ) );
  MUX \Reg_Bank/U4855  ( .A(\Reg_Bank/registers[2][25] ), .B(
        \Reg_Bank/registers[3][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4797 ) );
  MUX \Reg_Bank/U4854  ( .A(\Reg_Bank/n4795 ), .B(\Reg_Bank/n4794 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4796 ) );
  MUX \Reg_Bank/U4853  ( .A(\Reg_Bank/registers[4][25] ), .B(
        \Reg_Bank/registers[5][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4795 ) );
  MUX \Reg_Bank/U4852  ( .A(\Reg_Bank/registers[6][25] ), .B(
        \Reg_Bank/registers[7][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4794 ) );
  MUX \Reg_Bank/U4851  ( .A(\Reg_Bank/n4792 ), .B(\Reg_Bank/n4789 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4793 ) );
  MUX \Reg_Bank/U4850  ( .A(\Reg_Bank/n4791 ), .B(\Reg_Bank/n4790 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4792 ) );
  MUX \Reg_Bank/U4849  ( .A(\Reg_Bank/registers[8][25] ), .B(
        \Reg_Bank/registers[9][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4791 ) );
  MUX \Reg_Bank/U4848  ( .A(\Reg_Bank/registers[10][25] ), .B(
        \Reg_Bank/registers[11][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4790 )
         );
  MUX \Reg_Bank/U4847  ( .A(\Reg_Bank/n4788 ), .B(\Reg_Bank/n4787 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4789 ) );
  MUX \Reg_Bank/U4846  ( .A(\Reg_Bank/registers[12][25] ), .B(
        \Reg_Bank/registers[13][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4788 )
         );
  MUX \Reg_Bank/U4845  ( .A(\Reg_Bank/registers[14][25] ), .B(
        \Reg_Bank/registers[15][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4787 )
         );
  MUX \Reg_Bank/U4844  ( .A(\Reg_Bank/n4785 ), .B(\Reg_Bank/n4778 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4786 ) );
  MUX \Reg_Bank/U4843  ( .A(\Reg_Bank/n4784 ), .B(\Reg_Bank/n4781 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4785 ) );
  MUX \Reg_Bank/U4842  ( .A(\Reg_Bank/n4783 ), .B(\Reg_Bank/n4782 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4784 ) );
  MUX \Reg_Bank/U4841  ( .A(\Reg_Bank/registers[16][25] ), .B(
        \Reg_Bank/registers[17][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4783 )
         );
  MUX \Reg_Bank/U4840  ( .A(\Reg_Bank/registers[18][25] ), .B(
        \Reg_Bank/registers[19][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4782 )
         );
  MUX \Reg_Bank/U4839  ( .A(\Reg_Bank/n4780 ), .B(\Reg_Bank/n4779 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4781 ) );
  MUX \Reg_Bank/U4838  ( .A(\Reg_Bank/registers[20][25] ), .B(
        \Reg_Bank/registers[21][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4780 )
         );
  MUX \Reg_Bank/U4837  ( .A(\Reg_Bank/registers[22][25] ), .B(
        \Reg_Bank/registers[23][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4779 )
         );
  MUX \Reg_Bank/U4836  ( .A(\Reg_Bank/n4777 ), .B(\Reg_Bank/n4774 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4778 ) );
  MUX \Reg_Bank/U4835  ( .A(\Reg_Bank/n4776 ), .B(\Reg_Bank/n4775 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4777 ) );
  MUX \Reg_Bank/U4834  ( .A(\Reg_Bank/registers[24][25] ), .B(
        \Reg_Bank/registers[25][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4776 )
         );
  MUX \Reg_Bank/U4833  ( .A(\Reg_Bank/registers[26][25] ), .B(
        \Reg_Bank/registers[27][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4775 )
         );
  MUX \Reg_Bank/U4832  ( .A(\Reg_Bank/n4773 ), .B(\Reg_Bank/n4772 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4774 ) );
  MUX \Reg_Bank/U4831  ( .A(\Reg_Bank/registers[28][25] ), .B(
        \Reg_Bank/registers[29][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4773 )
         );
  MUX \Reg_Bank/U4830  ( .A(\Reg_Bank/registers[30][25] ), .B(
        \Reg_Bank/registers[31][25] ), .S(rs_index[0]), .Z(\Reg_Bank/n4772 )
         );
  MUX \Reg_Bank/U4829  ( .A(\Reg_Bank/n4771 ), .B(\Reg_Bank/n4756 ), .S(
        rs_index[4]), .Z(reg_source[24]) );
  MUX \Reg_Bank/U4828  ( .A(\Reg_Bank/n4770 ), .B(\Reg_Bank/n4763 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4771 ) );
  MUX \Reg_Bank/U4827  ( .A(\Reg_Bank/n4769 ), .B(\Reg_Bank/n4766 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4770 ) );
  MUX \Reg_Bank/U4826  ( .A(\Reg_Bank/n4768 ), .B(\Reg_Bank/n4767 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4769 ) );
  MUX \Reg_Bank/U4824  ( .A(\Reg_Bank/registers[2][24] ), .B(
        \Reg_Bank/registers[3][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4767 ) );
  MUX \Reg_Bank/U4823  ( .A(\Reg_Bank/n4765 ), .B(\Reg_Bank/n4764 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4766 ) );
  MUX \Reg_Bank/U4822  ( .A(\Reg_Bank/registers[4][24] ), .B(
        \Reg_Bank/registers[5][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4765 ) );
  MUX \Reg_Bank/U4821  ( .A(\Reg_Bank/registers[6][24] ), .B(
        \Reg_Bank/registers[7][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4764 ) );
  MUX \Reg_Bank/U4820  ( .A(\Reg_Bank/n4762 ), .B(\Reg_Bank/n4759 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4763 ) );
  MUX \Reg_Bank/U4819  ( .A(\Reg_Bank/n4761 ), .B(\Reg_Bank/n4760 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4762 ) );
  MUX \Reg_Bank/U4818  ( .A(\Reg_Bank/registers[8][24] ), .B(
        \Reg_Bank/registers[9][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4761 ) );
  MUX \Reg_Bank/U4817  ( .A(\Reg_Bank/registers[10][24] ), .B(
        \Reg_Bank/registers[11][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4760 )
         );
  MUX \Reg_Bank/U4816  ( .A(\Reg_Bank/n4758 ), .B(\Reg_Bank/n4757 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4759 ) );
  MUX \Reg_Bank/U4815  ( .A(\Reg_Bank/registers[12][24] ), .B(
        \Reg_Bank/registers[13][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4758 )
         );
  MUX \Reg_Bank/U4814  ( .A(\Reg_Bank/registers[14][24] ), .B(
        \Reg_Bank/registers[15][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4757 )
         );
  MUX \Reg_Bank/U4813  ( .A(\Reg_Bank/n4755 ), .B(\Reg_Bank/n4748 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4756 ) );
  MUX \Reg_Bank/U4812  ( .A(\Reg_Bank/n4754 ), .B(\Reg_Bank/n4751 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4755 ) );
  MUX \Reg_Bank/U4811  ( .A(\Reg_Bank/n4753 ), .B(\Reg_Bank/n4752 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4754 ) );
  MUX \Reg_Bank/U4810  ( .A(\Reg_Bank/registers[16][24] ), .B(
        \Reg_Bank/registers[17][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4753 )
         );
  MUX \Reg_Bank/U4809  ( .A(\Reg_Bank/registers[18][24] ), .B(
        \Reg_Bank/registers[19][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4752 )
         );
  MUX \Reg_Bank/U4808  ( .A(\Reg_Bank/n4750 ), .B(\Reg_Bank/n4749 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4751 ) );
  MUX \Reg_Bank/U4807  ( .A(\Reg_Bank/registers[20][24] ), .B(
        \Reg_Bank/registers[21][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4750 )
         );
  MUX \Reg_Bank/U4806  ( .A(\Reg_Bank/registers[22][24] ), .B(
        \Reg_Bank/registers[23][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4749 )
         );
  MUX \Reg_Bank/U4805  ( .A(\Reg_Bank/n4747 ), .B(\Reg_Bank/n4744 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4748 ) );
  MUX \Reg_Bank/U4804  ( .A(\Reg_Bank/n4746 ), .B(\Reg_Bank/n4745 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4747 ) );
  MUX \Reg_Bank/U4803  ( .A(\Reg_Bank/registers[24][24] ), .B(
        \Reg_Bank/registers[25][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4746 )
         );
  MUX \Reg_Bank/U4802  ( .A(\Reg_Bank/registers[26][24] ), .B(
        \Reg_Bank/registers[27][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4745 )
         );
  MUX \Reg_Bank/U4801  ( .A(\Reg_Bank/n4743 ), .B(\Reg_Bank/n4742 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4744 ) );
  MUX \Reg_Bank/U4800  ( .A(\Reg_Bank/registers[28][24] ), .B(
        \Reg_Bank/registers[29][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4743 )
         );
  MUX \Reg_Bank/U4799  ( .A(\Reg_Bank/registers[30][24] ), .B(
        \Reg_Bank/registers[31][24] ), .S(rs_index[0]), .Z(\Reg_Bank/n4742 )
         );
  MUX \Reg_Bank/U4798  ( .A(\Reg_Bank/n4741 ), .B(\Reg_Bank/n4726 ), .S(
        rs_index[4]), .Z(reg_source[23]) );
  MUX \Reg_Bank/U4797  ( .A(\Reg_Bank/n4740 ), .B(\Reg_Bank/n4733 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4741 ) );
  MUX \Reg_Bank/U4796  ( .A(\Reg_Bank/n4739 ), .B(\Reg_Bank/n4736 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4740 ) );
  MUX \Reg_Bank/U4795  ( .A(\Reg_Bank/n4738 ), .B(\Reg_Bank/n4737 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4739 ) );
  MUX \Reg_Bank/U4793  ( .A(\Reg_Bank/registers[2][23] ), .B(
        \Reg_Bank/registers[3][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4737 ) );
  MUX \Reg_Bank/U4792  ( .A(\Reg_Bank/n4735 ), .B(\Reg_Bank/n4734 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4736 ) );
  MUX \Reg_Bank/U4791  ( .A(\Reg_Bank/registers[4][23] ), .B(
        \Reg_Bank/registers[5][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4735 ) );
  MUX \Reg_Bank/U4790  ( .A(\Reg_Bank/registers[6][23] ), .B(
        \Reg_Bank/registers[7][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4734 ) );
  MUX \Reg_Bank/U4789  ( .A(\Reg_Bank/n4732 ), .B(\Reg_Bank/n4729 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4733 ) );
  MUX \Reg_Bank/U4788  ( .A(\Reg_Bank/n4731 ), .B(\Reg_Bank/n4730 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4732 ) );
  MUX \Reg_Bank/U4787  ( .A(\Reg_Bank/registers[8][23] ), .B(
        \Reg_Bank/registers[9][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4731 ) );
  MUX \Reg_Bank/U4786  ( .A(\Reg_Bank/registers[10][23] ), .B(
        \Reg_Bank/registers[11][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4730 )
         );
  MUX \Reg_Bank/U4785  ( .A(\Reg_Bank/n4728 ), .B(\Reg_Bank/n4727 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4729 ) );
  MUX \Reg_Bank/U4784  ( .A(\Reg_Bank/registers[12][23] ), .B(
        \Reg_Bank/registers[13][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4728 )
         );
  MUX \Reg_Bank/U4783  ( .A(\Reg_Bank/registers[14][23] ), .B(
        \Reg_Bank/registers[15][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4727 )
         );
  MUX \Reg_Bank/U4782  ( .A(\Reg_Bank/n4725 ), .B(\Reg_Bank/n4718 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4726 ) );
  MUX \Reg_Bank/U4781  ( .A(\Reg_Bank/n4724 ), .B(\Reg_Bank/n4721 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4725 ) );
  MUX \Reg_Bank/U4780  ( .A(\Reg_Bank/n4723 ), .B(\Reg_Bank/n4722 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4724 ) );
  MUX \Reg_Bank/U4779  ( .A(\Reg_Bank/registers[16][23] ), .B(
        \Reg_Bank/registers[17][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4723 )
         );
  MUX \Reg_Bank/U4778  ( .A(\Reg_Bank/registers[18][23] ), .B(
        \Reg_Bank/registers[19][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4722 )
         );
  MUX \Reg_Bank/U4777  ( .A(\Reg_Bank/n4720 ), .B(\Reg_Bank/n4719 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4721 ) );
  MUX \Reg_Bank/U4776  ( .A(\Reg_Bank/registers[20][23] ), .B(
        \Reg_Bank/registers[21][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4720 )
         );
  MUX \Reg_Bank/U4775  ( .A(\Reg_Bank/registers[22][23] ), .B(
        \Reg_Bank/registers[23][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4719 )
         );
  MUX \Reg_Bank/U4774  ( .A(\Reg_Bank/n4717 ), .B(\Reg_Bank/n4714 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4718 ) );
  MUX \Reg_Bank/U4773  ( .A(\Reg_Bank/n4716 ), .B(\Reg_Bank/n4715 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4717 ) );
  MUX \Reg_Bank/U4772  ( .A(\Reg_Bank/registers[24][23] ), .B(
        \Reg_Bank/registers[25][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4716 )
         );
  MUX \Reg_Bank/U4771  ( .A(\Reg_Bank/registers[26][23] ), .B(
        \Reg_Bank/registers[27][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4715 )
         );
  MUX \Reg_Bank/U4770  ( .A(\Reg_Bank/n4713 ), .B(\Reg_Bank/n4712 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4714 ) );
  MUX \Reg_Bank/U4769  ( .A(\Reg_Bank/registers[28][23] ), .B(
        \Reg_Bank/registers[29][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4713 )
         );
  MUX \Reg_Bank/U4768  ( .A(\Reg_Bank/registers[30][23] ), .B(
        \Reg_Bank/registers[31][23] ), .S(rs_index[0]), .Z(\Reg_Bank/n4712 )
         );
  MUX \Reg_Bank/U4767  ( .A(\Reg_Bank/n4711 ), .B(\Reg_Bank/n4696 ), .S(
        rs_index[4]), .Z(reg_source[22]) );
  MUX \Reg_Bank/U4766  ( .A(\Reg_Bank/n4710 ), .B(\Reg_Bank/n4703 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4711 ) );
  MUX \Reg_Bank/U4765  ( .A(\Reg_Bank/n4709 ), .B(\Reg_Bank/n4706 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4710 ) );
  MUX \Reg_Bank/U4764  ( .A(\Reg_Bank/n4708 ), .B(\Reg_Bank/n4707 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4709 ) );
  MUX \Reg_Bank/U4762  ( .A(\Reg_Bank/registers[2][22] ), .B(
        \Reg_Bank/registers[3][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4707 ) );
  MUX \Reg_Bank/U4761  ( .A(\Reg_Bank/n4705 ), .B(\Reg_Bank/n4704 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4706 ) );
  MUX \Reg_Bank/U4760  ( .A(\Reg_Bank/registers[4][22] ), .B(
        \Reg_Bank/registers[5][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4705 ) );
  MUX \Reg_Bank/U4759  ( .A(\Reg_Bank/registers[6][22] ), .B(
        \Reg_Bank/registers[7][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4704 ) );
  MUX \Reg_Bank/U4758  ( .A(\Reg_Bank/n4702 ), .B(\Reg_Bank/n4699 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4703 ) );
  MUX \Reg_Bank/U4757  ( .A(\Reg_Bank/n4701 ), .B(\Reg_Bank/n4700 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4702 ) );
  MUX \Reg_Bank/U4756  ( .A(\Reg_Bank/registers[8][22] ), .B(
        \Reg_Bank/registers[9][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4701 ) );
  MUX \Reg_Bank/U4755  ( .A(\Reg_Bank/registers[10][22] ), .B(
        \Reg_Bank/registers[11][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4700 )
         );
  MUX \Reg_Bank/U4754  ( .A(\Reg_Bank/n4698 ), .B(\Reg_Bank/n4697 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4699 ) );
  MUX \Reg_Bank/U4753  ( .A(\Reg_Bank/registers[12][22] ), .B(
        \Reg_Bank/registers[13][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4698 )
         );
  MUX \Reg_Bank/U4752  ( .A(\Reg_Bank/registers[14][22] ), .B(
        \Reg_Bank/registers[15][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4697 )
         );
  MUX \Reg_Bank/U4751  ( .A(\Reg_Bank/n4695 ), .B(\Reg_Bank/n4688 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4696 ) );
  MUX \Reg_Bank/U4750  ( .A(\Reg_Bank/n4694 ), .B(\Reg_Bank/n4691 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4695 ) );
  MUX \Reg_Bank/U4749  ( .A(\Reg_Bank/n4693 ), .B(\Reg_Bank/n4692 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4694 ) );
  MUX \Reg_Bank/U4748  ( .A(\Reg_Bank/registers[16][22] ), .B(
        \Reg_Bank/registers[17][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4693 )
         );
  MUX \Reg_Bank/U4747  ( .A(\Reg_Bank/registers[18][22] ), .B(
        \Reg_Bank/registers[19][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4692 )
         );
  MUX \Reg_Bank/U4746  ( .A(\Reg_Bank/n4690 ), .B(\Reg_Bank/n4689 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4691 ) );
  MUX \Reg_Bank/U4745  ( .A(\Reg_Bank/registers[20][22] ), .B(
        \Reg_Bank/registers[21][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4690 )
         );
  MUX \Reg_Bank/U4744  ( .A(\Reg_Bank/registers[22][22] ), .B(
        \Reg_Bank/registers[23][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4689 )
         );
  MUX \Reg_Bank/U4743  ( .A(\Reg_Bank/n4687 ), .B(\Reg_Bank/n4684 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4688 ) );
  MUX \Reg_Bank/U4742  ( .A(\Reg_Bank/n4686 ), .B(\Reg_Bank/n4685 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4687 ) );
  MUX \Reg_Bank/U4741  ( .A(\Reg_Bank/registers[24][22] ), .B(
        \Reg_Bank/registers[25][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4686 )
         );
  MUX \Reg_Bank/U4740  ( .A(\Reg_Bank/registers[26][22] ), .B(
        \Reg_Bank/registers[27][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4685 )
         );
  MUX \Reg_Bank/U4739  ( .A(\Reg_Bank/n4683 ), .B(\Reg_Bank/n4682 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4684 ) );
  MUX \Reg_Bank/U4738  ( .A(\Reg_Bank/registers[28][22] ), .B(
        \Reg_Bank/registers[29][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4683 )
         );
  MUX \Reg_Bank/U4737  ( .A(\Reg_Bank/registers[30][22] ), .B(
        \Reg_Bank/registers[31][22] ), .S(rs_index[0]), .Z(\Reg_Bank/n4682 )
         );
  MUX \Reg_Bank/U4736  ( .A(\Reg_Bank/n4681 ), .B(\Reg_Bank/n4666 ), .S(
        rs_index[4]), .Z(reg_source[21]) );
  MUX \Reg_Bank/U4735  ( .A(\Reg_Bank/n4680 ), .B(\Reg_Bank/n4673 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4681 ) );
  MUX \Reg_Bank/U4734  ( .A(\Reg_Bank/n4679 ), .B(\Reg_Bank/n4676 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4680 ) );
  MUX \Reg_Bank/U4733  ( .A(\Reg_Bank/n4678 ), .B(\Reg_Bank/n4677 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4679 ) );
  MUX \Reg_Bank/U4731  ( .A(\Reg_Bank/registers[2][21] ), .B(
        \Reg_Bank/registers[3][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4677 ) );
  MUX \Reg_Bank/U4730  ( .A(\Reg_Bank/n4675 ), .B(\Reg_Bank/n4674 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4676 ) );
  MUX \Reg_Bank/U4729  ( .A(\Reg_Bank/registers[4][21] ), .B(
        \Reg_Bank/registers[5][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4675 ) );
  MUX \Reg_Bank/U4728  ( .A(\Reg_Bank/registers[6][21] ), .B(
        \Reg_Bank/registers[7][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4674 ) );
  MUX \Reg_Bank/U4727  ( .A(\Reg_Bank/n4672 ), .B(\Reg_Bank/n4669 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4673 ) );
  MUX \Reg_Bank/U4726  ( .A(\Reg_Bank/n4671 ), .B(\Reg_Bank/n4670 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4672 ) );
  MUX \Reg_Bank/U4725  ( .A(\Reg_Bank/registers[8][21] ), .B(
        \Reg_Bank/registers[9][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4671 ) );
  MUX \Reg_Bank/U4724  ( .A(\Reg_Bank/registers[10][21] ), .B(
        \Reg_Bank/registers[11][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4670 )
         );
  MUX \Reg_Bank/U4723  ( .A(\Reg_Bank/n4668 ), .B(\Reg_Bank/n4667 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4669 ) );
  MUX \Reg_Bank/U4722  ( .A(\Reg_Bank/registers[12][21] ), .B(
        \Reg_Bank/registers[13][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4668 )
         );
  MUX \Reg_Bank/U4721  ( .A(\Reg_Bank/registers[14][21] ), .B(
        \Reg_Bank/registers[15][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4667 )
         );
  MUX \Reg_Bank/U4720  ( .A(\Reg_Bank/n4665 ), .B(\Reg_Bank/n4658 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4666 ) );
  MUX \Reg_Bank/U4719  ( .A(\Reg_Bank/n4664 ), .B(\Reg_Bank/n4661 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4665 ) );
  MUX \Reg_Bank/U4718  ( .A(\Reg_Bank/n4663 ), .B(\Reg_Bank/n4662 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4664 ) );
  MUX \Reg_Bank/U4717  ( .A(\Reg_Bank/registers[16][21] ), .B(
        \Reg_Bank/registers[17][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4663 )
         );
  MUX \Reg_Bank/U4716  ( .A(\Reg_Bank/registers[18][21] ), .B(
        \Reg_Bank/registers[19][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4662 )
         );
  MUX \Reg_Bank/U4715  ( .A(\Reg_Bank/n4660 ), .B(\Reg_Bank/n4659 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4661 ) );
  MUX \Reg_Bank/U4714  ( .A(\Reg_Bank/registers[20][21] ), .B(
        \Reg_Bank/registers[21][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4660 )
         );
  MUX \Reg_Bank/U4713  ( .A(\Reg_Bank/registers[22][21] ), .B(
        \Reg_Bank/registers[23][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4659 )
         );
  MUX \Reg_Bank/U4712  ( .A(\Reg_Bank/n4657 ), .B(\Reg_Bank/n4654 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4658 ) );
  MUX \Reg_Bank/U4711  ( .A(\Reg_Bank/n4656 ), .B(\Reg_Bank/n4655 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4657 ) );
  MUX \Reg_Bank/U4710  ( .A(\Reg_Bank/registers[24][21] ), .B(
        \Reg_Bank/registers[25][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4656 )
         );
  MUX \Reg_Bank/U4709  ( .A(\Reg_Bank/registers[26][21] ), .B(
        \Reg_Bank/registers[27][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4655 )
         );
  MUX \Reg_Bank/U4708  ( .A(\Reg_Bank/n4653 ), .B(\Reg_Bank/n4652 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4654 ) );
  MUX \Reg_Bank/U4707  ( .A(\Reg_Bank/registers[28][21] ), .B(
        \Reg_Bank/registers[29][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4653 )
         );
  MUX \Reg_Bank/U4706  ( .A(\Reg_Bank/registers[30][21] ), .B(
        \Reg_Bank/registers[31][21] ), .S(rs_index[0]), .Z(\Reg_Bank/n4652 )
         );
  MUX \Reg_Bank/U4705  ( .A(\Reg_Bank/n4651 ), .B(\Reg_Bank/n4636 ), .S(
        rs_index[4]), .Z(reg_source[20]) );
  MUX \Reg_Bank/U4704  ( .A(\Reg_Bank/n4650 ), .B(\Reg_Bank/n4643 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4651 ) );
  MUX \Reg_Bank/U4703  ( .A(\Reg_Bank/n4649 ), .B(\Reg_Bank/n4646 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4650 ) );
  MUX \Reg_Bank/U4702  ( .A(\Reg_Bank/n4648 ), .B(\Reg_Bank/n4647 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4649 ) );
  MUX \Reg_Bank/U4700  ( .A(\Reg_Bank/registers[2][20] ), .B(
        \Reg_Bank/registers[3][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4647 ) );
  MUX \Reg_Bank/U4699  ( .A(\Reg_Bank/n4645 ), .B(\Reg_Bank/n4644 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4646 ) );
  MUX \Reg_Bank/U4698  ( .A(\Reg_Bank/registers[4][20] ), .B(
        \Reg_Bank/registers[5][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4645 ) );
  MUX \Reg_Bank/U4697  ( .A(\Reg_Bank/registers[6][20] ), .B(
        \Reg_Bank/registers[7][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4644 ) );
  MUX \Reg_Bank/U4696  ( .A(\Reg_Bank/n4642 ), .B(\Reg_Bank/n4639 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4643 ) );
  MUX \Reg_Bank/U4695  ( .A(\Reg_Bank/n4641 ), .B(\Reg_Bank/n4640 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4642 ) );
  MUX \Reg_Bank/U4694  ( .A(\Reg_Bank/registers[8][20] ), .B(
        \Reg_Bank/registers[9][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4641 ) );
  MUX \Reg_Bank/U4693  ( .A(\Reg_Bank/registers[10][20] ), .B(
        \Reg_Bank/registers[11][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4640 )
         );
  MUX \Reg_Bank/U4692  ( .A(\Reg_Bank/n4638 ), .B(\Reg_Bank/n4637 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4639 ) );
  MUX \Reg_Bank/U4691  ( .A(\Reg_Bank/registers[12][20] ), .B(
        \Reg_Bank/registers[13][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4638 )
         );
  MUX \Reg_Bank/U4690  ( .A(\Reg_Bank/registers[14][20] ), .B(
        \Reg_Bank/registers[15][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4637 )
         );
  MUX \Reg_Bank/U4689  ( .A(\Reg_Bank/n4635 ), .B(\Reg_Bank/n4628 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4636 ) );
  MUX \Reg_Bank/U4688  ( .A(\Reg_Bank/n4634 ), .B(\Reg_Bank/n4631 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4635 ) );
  MUX \Reg_Bank/U4687  ( .A(\Reg_Bank/n4633 ), .B(\Reg_Bank/n4632 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4634 ) );
  MUX \Reg_Bank/U4686  ( .A(\Reg_Bank/registers[16][20] ), .B(
        \Reg_Bank/registers[17][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4633 )
         );
  MUX \Reg_Bank/U4685  ( .A(\Reg_Bank/registers[18][20] ), .B(
        \Reg_Bank/registers[19][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4632 )
         );
  MUX \Reg_Bank/U4684  ( .A(\Reg_Bank/n4630 ), .B(\Reg_Bank/n4629 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4631 ) );
  MUX \Reg_Bank/U4683  ( .A(\Reg_Bank/registers[20][20] ), .B(
        \Reg_Bank/registers[21][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4630 )
         );
  MUX \Reg_Bank/U4682  ( .A(\Reg_Bank/registers[22][20] ), .B(
        \Reg_Bank/registers[23][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4629 )
         );
  MUX \Reg_Bank/U4681  ( .A(\Reg_Bank/n4627 ), .B(\Reg_Bank/n4624 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4628 ) );
  MUX \Reg_Bank/U4680  ( .A(\Reg_Bank/n4626 ), .B(\Reg_Bank/n4625 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4627 ) );
  MUX \Reg_Bank/U4679  ( .A(\Reg_Bank/registers[24][20] ), .B(
        \Reg_Bank/registers[25][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4626 )
         );
  MUX \Reg_Bank/U4678  ( .A(\Reg_Bank/registers[26][20] ), .B(
        \Reg_Bank/registers[27][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4625 )
         );
  MUX \Reg_Bank/U4677  ( .A(\Reg_Bank/n4623 ), .B(\Reg_Bank/n4622 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4624 ) );
  MUX \Reg_Bank/U4676  ( .A(\Reg_Bank/registers[28][20] ), .B(
        \Reg_Bank/registers[29][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4623 )
         );
  MUX \Reg_Bank/U4675  ( .A(\Reg_Bank/registers[30][20] ), .B(
        \Reg_Bank/registers[31][20] ), .S(rs_index[0]), .Z(\Reg_Bank/n4622 )
         );
  MUX \Reg_Bank/U4674  ( .A(\Reg_Bank/n4621 ), .B(\Reg_Bank/n4606 ), .S(
        rs_index[4]), .Z(reg_source[19]) );
  MUX \Reg_Bank/U4673  ( .A(\Reg_Bank/n4620 ), .B(\Reg_Bank/n4613 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4621 ) );
  MUX \Reg_Bank/U4672  ( .A(\Reg_Bank/n4619 ), .B(\Reg_Bank/n4616 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4620 ) );
  MUX \Reg_Bank/U4671  ( .A(\Reg_Bank/n4618 ), .B(\Reg_Bank/n4617 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4619 ) );
  MUX \Reg_Bank/U4669  ( .A(\Reg_Bank/registers[2][19] ), .B(
        \Reg_Bank/registers[3][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4617 ) );
  MUX \Reg_Bank/U4668  ( .A(\Reg_Bank/n4615 ), .B(\Reg_Bank/n4614 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4616 ) );
  MUX \Reg_Bank/U4667  ( .A(\Reg_Bank/registers[4][19] ), .B(
        \Reg_Bank/registers[5][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4615 ) );
  MUX \Reg_Bank/U4666  ( .A(\Reg_Bank/registers[6][19] ), .B(
        \Reg_Bank/registers[7][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4614 ) );
  MUX \Reg_Bank/U4665  ( .A(\Reg_Bank/n4612 ), .B(\Reg_Bank/n4609 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4613 ) );
  MUX \Reg_Bank/U4664  ( .A(\Reg_Bank/n4611 ), .B(\Reg_Bank/n4610 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4612 ) );
  MUX \Reg_Bank/U4663  ( .A(\Reg_Bank/registers[8][19] ), .B(
        \Reg_Bank/registers[9][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4611 ) );
  MUX \Reg_Bank/U4662  ( .A(\Reg_Bank/registers[10][19] ), .B(
        \Reg_Bank/registers[11][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4610 )
         );
  MUX \Reg_Bank/U4661  ( .A(\Reg_Bank/n4608 ), .B(\Reg_Bank/n4607 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4609 ) );
  MUX \Reg_Bank/U4660  ( .A(\Reg_Bank/registers[12][19] ), .B(
        \Reg_Bank/registers[13][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4608 )
         );
  MUX \Reg_Bank/U4659  ( .A(\Reg_Bank/registers[14][19] ), .B(
        \Reg_Bank/registers[15][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4607 )
         );
  MUX \Reg_Bank/U4658  ( .A(\Reg_Bank/n4605 ), .B(\Reg_Bank/n4598 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4606 ) );
  MUX \Reg_Bank/U4657  ( .A(\Reg_Bank/n4604 ), .B(\Reg_Bank/n4601 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4605 ) );
  MUX \Reg_Bank/U4656  ( .A(\Reg_Bank/n4603 ), .B(\Reg_Bank/n4602 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4604 ) );
  MUX \Reg_Bank/U4655  ( .A(\Reg_Bank/registers[16][19] ), .B(
        \Reg_Bank/registers[17][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4603 )
         );
  MUX \Reg_Bank/U4654  ( .A(\Reg_Bank/registers[18][19] ), .B(
        \Reg_Bank/registers[19][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4602 )
         );
  MUX \Reg_Bank/U4653  ( .A(\Reg_Bank/n4600 ), .B(\Reg_Bank/n4599 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4601 ) );
  MUX \Reg_Bank/U4652  ( .A(\Reg_Bank/registers[20][19] ), .B(
        \Reg_Bank/registers[21][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4600 )
         );
  MUX \Reg_Bank/U4651  ( .A(\Reg_Bank/registers[22][19] ), .B(
        \Reg_Bank/registers[23][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4599 )
         );
  MUX \Reg_Bank/U4650  ( .A(\Reg_Bank/n4597 ), .B(\Reg_Bank/n4594 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4598 ) );
  MUX \Reg_Bank/U4649  ( .A(\Reg_Bank/n4596 ), .B(\Reg_Bank/n4595 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4597 ) );
  MUX \Reg_Bank/U4648  ( .A(\Reg_Bank/registers[24][19] ), .B(
        \Reg_Bank/registers[25][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4596 )
         );
  MUX \Reg_Bank/U4647  ( .A(\Reg_Bank/registers[26][19] ), .B(
        \Reg_Bank/registers[27][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4595 )
         );
  MUX \Reg_Bank/U4646  ( .A(\Reg_Bank/n4593 ), .B(\Reg_Bank/n4592 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4594 ) );
  MUX \Reg_Bank/U4645  ( .A(\Reg_Bank/registers[28][19] ), .B(
        \Reg_Bank/registers[29][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4593 )
         );
  MUX \Reg_Bank/U4644  ( .A(\Reg_Bank/registers[30][19] ), .B(
        \Reg_Bank/registers[31][19] ), .S(rs_index[0]), .Z(\Reg_Bank/n4592 )
         );
  MUX \Reg_Bank/U4643  ( .A(\Reg_Bank/n4591 ), .B(\Reg_Bank/n4576 ), .S(
        rs_index[4]), .Z(reg_source[18]) );
  MUX \Reg_Bank/U4642  ( .A(\Reg_Bank/n4590 ), .B(\Reg_Bank/n4583 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4591 ) );
  MUX \Reg_Bank/U4641  ( .A(\Reg_Bank/n4589 ), .B(\Reg_Bank/n4586 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4590 ) );
  MUX \Reg_Bank/U4640  ( .A(\Reg_Bank/n4588 ), .B(\Reg_Bank/n4587 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4589 ) );
  MUX \Reg_Bank/U4638  ( .A(\Reg_Bank/registers[2][18] ), .B(
        \Reg_Bank/registers[3][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4587 ) );
  MUX \Reg_Bank/U4637  ( .A(\Reg_Bank/n4585 ), .B(\Reg_Bank/n4584 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4586 ) );
  MUX \Reg_Bank/U4636  ( .A(\Reg_Bank/registers[4][18] ), .B(
        \Reg_Bank/registers[5][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4585 ) );
  MUX \Reg_Bank/U4635  ( .A(\Reg_Bank/registers[6][18] ), .B(
        \Reg_Bank/registers[7][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4584 ) );
  MUX \Reg_Bank/U4634  ( .A(\Reg_Bank/n4582 ), .B(\Reg_Bank/n4579 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4583 ) );
  MUX \Reg_Bank/U4633  ( .A(\Reg_Bank/n4581 ), .B(\Reg_Bank/n4580 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4582 ) );
  MUX \Reg_Bank/U4632  ( .A(\Reg_Bank/registers[8][18] ), .B(
        \Reg_Bank/registers[9][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4581 ) );
  MUX \Reg_Bank/U4631  ( .A(\Reg_Bank/registers[10][18] ), .B(
        \Reg_Bank/registers[11][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4580 )
         );
  MUX \Reg_Bank/U4630  ( .A(\Reg_Bank/n4578 ), .B(\Reg_Bank/n4577 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4579 ) );
  MUX \Reg_Bank/U4629  ( .A(\Reg_Bank/registers[12][18] ), .B(
        \Reg_Bank/registers[13][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4578 )
         );
  MUX \Reg_Bank/U4628  ( .A(\Reg_Bank/registers[14][18] ), .B(
        \Reg_Bank/registers[15][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4577 )
         );
  MUX \Reg_Bank/U4627  ( .A(\Reg_Bank/n4575 ), .B(\Reg_Bank/n4568 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4576 ) );
  MUX \Reg_Bank/U4626  ( .A(\Reg_Bank/n4574 ), .B(\Reg_Bank/n4571 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4575 ) );
  MUX \Reg_Bank/U4625  ( .A(\Reg_Bank/n4573 ), .B(\Reg_Bank/n4572 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4574 ) );
  MUX \Reg_Bank/U4624  ( .A(\Reg_Bank/registers[16][18] ), .B(
        \Reg_Bank/registers[17][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4573 )
         );
  MUX \Reg_Bank/U4623  ( .A(\Reg_Bank/registers[18][18] ), .B(
        \Reg_Bank/registers[19][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4572 )
         );
  MUX \Reg_Bank/U4622  ( .A(\Reg_Bank/n4570 ), .B(\Reg_Bank/n4569 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4571 ) );
  MUX \Reg_Bank/U4621  ( .A(\Reg_Bank/registers[20][18] ), .B(
        \Reg_Bank/registers[21][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4570 )
         );
  MUX \Reg_Bank/U4620  ( .A(\Reg_Bank/registers[22][18] ), .B(
        \Reg_Bank/registers[23][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4569 )
         );
  MUX \Reg_Bank/U4619  ( .A(\Reg_Bank/n4567 ), .B(\Reg_Bank/n4564 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4568 ) );
  MUX \Reg_Bank/U4618  ( .A(\Reg_Bank/n4566 ), .B(\Reg_Bank/n4565 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4567 ) );
  MUX \Reg_Bank/U4617  ( .A(\Reg_Bank/registers[24][18] ), .B(
        \Reg_Bank/registers[25][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4566 )
         );
  MUX \Reg_Bank/U4616  ( .A(\Reg_Bank/registers[26][18] ), .B(
        \Reg_Bank/registers[27][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4565 )
         );
  MUX \Reg_Bank/U4615  ( .A(\Reg_Bank/n4563 ), .B(\Reg_Bank/n4562 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4564 ) );
  MUX \Reg_Bank/U4614  ( .A(\Reg_Bank/registers[28][18] ), .B(
        \Reg_Bank/registers[29][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4563 )
         );
  MUX \Reg_Bank/U4613  ( .A(\Reg_Bank/registers[30][18] ), .B(
        \Reg_Bank/registers[31][18] ), .S(rs_index[0]), .Z(\Reg_Bank/n4562 )
         );
  MUX \Reg_Bank/U4612  ( .A(\Reg_Bank/n4561 ), .B(\Reg_Bank/n4546 ), .S(
        rs_index[4]), .Z(reg_source[17]) );
  MUX \Reg_Bank/U4611  ( .A(\Reg_Bank/n4560 ), .B(\Reg_Bank/n4553 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4561 ) );
  MUX \Reg_Bank/U4610  ( .A(\Reg_Bank/n4559 ), .B(\Reg_Bank/n4556 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4560 ) );
  MUX \Reg_Bank/U4609  ( .A(\Reg_Bank/n4558 ), .B(\Reg_Bank/n4557 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4559 ) );
  MUX \Reg_Bank/U4607  ( .A(\Reg_Bank/registers[2][17] ), .B(
        \Reg_Bank/registers[3][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4557 ) );
  MUX \Reg_Bank/U4606  ( .A(\Reg_Bank/n4555 ), .B(\Reg_Bank/n4554 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4556 ) );
  MUX \Reg_Bank/U4605  ( .A(\Reg_Bank/registers[4][17] ), .B(
        \Reg_Bank/registers[5][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4555 ) );
  MUX \Reg_Bank/U4604  ( .A(\Reg_Bank/registers[6][17] ), .B(
        \Reg_Bank/registers[7][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4554 ) );
  MUX \Reg_Bank/U4603  ( .A(\Reg_Bank/n4552 ), .B(\Reg_Bank/n4549 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4553 ) );
  MUX \Reg_Bank/U4602  ( .A(\Reg_Bank/n4551 ), .B(\Reg_Bank/n4550 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4552 ) );
  MUX \Reg_Bank/U4601  ( .A(\Reg_Bank/registers[8][17] ), .B(
        \Reg_Bank/registers[9][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4551 ) );
  MUX \Reg_Bank/U4600  ( .A(\Reg_Bank/registers[10][17] ), .B(
        \Reg_Bank/registers[11][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4550 )
         );
  MUX \Reg_Bank/U4599  ( .A(\Reg_Bank/n4548 ), .B(\Reg_Bank/n4547 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4549 ) );
  MUX \Reg_Bank/U4598  ( .A(\Reg_Bank/registers[12][17] ), .B(
        \Reg_Bank/registers[13][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4548 )
         );
  MUX \Reg_Bank/U4597  ( .A(\Reg_Bank/registers[14][17] ), .B(
        \Reg_Bank/registers[15][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4547 )
         );
  MUX \Reg_Bank/U4596  ( .A(\Reg_Bank/n4545 ), .B(\Reg_Bank/n4538 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4546 ) );
  MUX \Reg_Bank/U4595  ( .A(\Reg_Bank/n4544 ), .B(\Reg_Bank/n4541 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4545 ) );
  MUX \Reg_Bank/U4594  ( .A(\Reg_Bank/n4543 ), .B(\Reg_Bank/n4542 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4544 ) );
  MUX \Reg_Bank/U4593  ( .A(\Reg_Bank/registers[16][17] ), .B(
        \Reg_Bank/registers[17][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4543 )
         );
  MUX \Reg_Bank/U4592  ( .A(\Reg_Bank/registers[18][17] ), .B(
        \Reg_Bank/registers[19][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4542 )
         );
  MUX \Reg_Bank/U4591  ( .A(\Reg_Bank/n4540 ), .B(\Reg_Bank/n4539 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4541 ) );
  MUX \Reg_Bank/U4590  ( .A(\Reg_Bank/registers[20][17] ), .B(
        \Reg_Bank/registers[21][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4540 )
         );
  MUX \Reg_Bank/U4589  ( .A(\Reg_Bank/registers[22][17] ), .B(
        \Reg_Bank/registers[23][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4539 )
         );
  MUX \Reg_Bank/U4588  ( .A(\Reg_Bank/n4537 ), .B(\Reg_Bank/n4534 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4538 ) );
  MUX \Reg_Bank/U4587  ( .A(\Reg_Bank/n4536 ), .B(\Reg_Bank/n4535 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4537 ) );
  MUX \Reg_Bank/U4586  ( .A(\Reg_Bank/registers[24][17] ), .B(
        \Reg_Bank/registers[25][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4536 )
         );
  MUX \Reg_Bank/U4585  ( .A(\Reg_Bank/registers[26][17] ), .B(
        \Reg_Bank/registers[27][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4535 )
         );
  MUX \Reg_Bank/U4584  ( .A(\Reg_Bank/n4533 ), .B(\Reg_Bank/n4532 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4534 ) );
  MUX \Reg_Bank/U4583  ( .A(\Reg_Bank/registers[28][17] ), .B(
        \Reg_Bank/registers[29][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4533 )
         );
  MUX \Reg_Bank/U4582  ( .A(\Reg_Bank/registers[30][17] ), .B(
        \Reg_Bank/registers[31][17] ), .S(rs_index[0]), .Z(\Reg_Bank/n4532 )
         );
  MUX \Reg_Bank/U4581  ( .A(\Reg_Bank/n4531 ), .B(\Reg_Bank/n4516 ), .S(
        rs_index[4]), .Z(reg_source[16]) );
  MUX \Reg_Bank/U4580  ( .A(\Reg_Bank/n4530 ), .B(\Reg_Bank/n4523 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4531 ) );
  MUX \Reg_Bank/U4579  ( .A(\Reg_Bank/n4529 ), .B(\Reg_Bank/n4526 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4530 ) );
  MUX \Reg_Bank/U4578  ( .A(\Reg_Bank/n4528 ), .B(\Reg_Bank/n4527 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4529 ) );
  MUX \Reg_Bank/U4576  ( .A(\Reg_Bank/registers[2][16] ), .B(
        \Reg_Bank/registers[3][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4527 ) );
  MUX \Reg_Bank/U4575  ( .A(\Reg_Bank/n4525 ), .B(\Reg_Bank/n4524 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4526 ) );
  MUX \Reg_Bank/U4574  ( .A(\Reg_Bank/registers[4][16] ), .B(
        \Reg_Bank/registers[5][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4525 ) );
  MUX \Reg_Bank/U4573  ( .A(\Reg_Bank/registers[6][16] ), .B(
        \Reg_Bank/registers[7][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4524 ) );
  MUX \Reg_Bank/U4572  ( .A(\Reg_Bank/n4522 ), .B(\Reg_Bank/n4519 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4523 ) );
  MUX \Reg_Bank/U4571  ( .A(\Reg_Bank/n4521 ), .B(\Reg_Bank/n4520 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4522 ) );
  MUX \Reg_Bank/U4570  ( .A(\Reg_Bank/registers[8][16] ), .B(
        \Reg_Bank/registers[9][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4521 ) );
  MUX \Reg_Bank/U4569  ( .A(\Reg_Bank/registers[10][16] ), .B(
        \Reg_Bank/registers[11][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4520 )
         );
  MUX \Reg_Bank/U4568  ( .A(\Reg_Bank/n4518 ), .B(\Reg_Bank/n4517 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4519 ) );
  MUX \Reg_Bank/U4567  ( .A(\Reg_Bank/registers[12][16] ), .B(
        \Reg_Bank/registers[13][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4518 )
         );
  MUX \Reg_Bank/U4566  ( .A(\Reg_Bank/registers[14][16] ), .B(
        \Reg_Bank/registers[15][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4517 )
         );
  MUX \Reg_Bank/U4565  ( .A(\Reg_Bank/n4515 ), .B(\Reg_Bank/n4508 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4516 ) );
  MUX \Reg_Bank/U4564  ( .A(\Reg_Bank/n4514 ), .B(\Reg_Bank/n4511 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4515 ) );
  MUX \Reg_Bank/U4563  ( .A(\Reg_Bank/n4513 ), .B(\Reg_Bank/n4512 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4514 ) );
  MUX \Reg_Bank/U4562  ( .A(\Reg_Bank/registers[16][16] ), .B(
        \Reg_Bank/registers[17][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4513 )
         );
  MUX \Reg_Bank/U4561  ( .A(\Reg_Bank/registers[18][16] ), .B(
        \Reg_Bank/registers[19][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4512 )
         );
  MUX \Reg_Bank/U4560  ( .A(\Reg_Bank/n4510 ), .B(\Reg_Bank/n4509 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4511 ) );
  MUX \Reg_Bank/U4559  ( .A(\Reg_Bank/registers[20][16] ), .B(
        \Reg_Bank/registers[21][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4510 )
         );
  MUX \Reg_Bank/U4558  ( .A(\Reg_Bank/registers[22][16] ), .B(
        \Reg_Bank/registers[23][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4509 )
         );
  MUX \Reg_Bank/U4557  ( .A(\Reg_Bank/n4507 ), .B(\Reg_Bank/n4504 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4508 ) );
  MUX \Reg_Bank/U4556  ( .A(\Reg_Bank/n4506 ), .B(\Reg_Bank/n4505 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4507 ) );
  MUX \Reg_Bank/U4555  ( .A(\Reg_Bank/registers[24][16] ), .B(
        \Reg_Bank/registers[25][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4506 )
         );
  MUX \Reg_Bank/U4554  ( .A(\Reg_Bank/registers[26][16] ), .B(
        \Reg_Bank/registers[27][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4505 )
         );
  MUX \Reg_Bank/U4553  ( .A(\Reg_Bank/n4503 ), .B(\Reg_Bank/n4502 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4504 ) );
  MUX \Reg_Bank/U4552  ( .A(\Reg_Bank/registers[28][16] ), .B(
        \Reg_Bank/registers[29][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4503 )
         );
  MUX \Reg_Bank/U4551  ( .A(\Reg_Bank/registers[30][16] ), .B(
        \Reg_Bank/registers[31][16] ), .S(rs_index[0]), .Z(\Reg_Bank/n4502 )
         );
  MUX \Reg_Bank/U4550  ( .A(\Reg_Bank/n4501 ), .B(\Reg_Bank/n4486 ), .S(
        rs_index[4]), .Z(reg_source[15]) );
  MUX \Reg_Bank/U4549  ( .A(\Reg_Bank/n4500 ), .B(\Reg_Bank/n4493 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4501 ) );
  MUX \Reg_Bank/U4548  ( .A(\Reg_Bank/n4499 ), .B(\Reg_Bank/n4496 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4500 ) );
  MUX \Reg_Bank/U4547  ( .A(\Reg_Bank/n4498 ), .B(\Reg_Bank/n4497 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4499 ) );
  MUX \Reg_Bank/U4545  ( .A(\Reg_Bank/registers[2][15] ), .B(
        \Reg_Bank/registers[3][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4497 ) );
  MUX \Reg_Bank/U4544  ( .A(\Reg_Bank/n4495 ), .B(\Reg_Bank/n4494 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4496 ) );
  MUX \Reg_Bank/U4543  ( .A(\Reg_Bank/registers[4][15] ), .B(
        \Reg_Bank/registers[5][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4495 ) );
  MUX \Reg_Bank/U4542  ( .A(\Reg_Bank/registers[6][15] ), .B(
        \Reg_Bank/registers[7][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4494 ) );
  MUX \Reg_Bank/U4541  ( .A(\Reg_Bank/n4492 ), .B(\Reg_Bank/n4489 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4493 ) );
  MUX \Reg_Bank/U4540  ( .A(\Reg_Bank/n4491 ), .B(\Reg_Bank/n4490 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4492 ) );
  MUX \Reg_Bank/U4539  ( .A(\Reg_Bank/registers[8][15] ), .B(
        \Reg_Bank/registers[9][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4491 ) );
  MUX \Reg_Bank/U4538  ( .A(\Reg_Bank/registers[10][15] ), .B(
        \Reg_Bank/registers[11][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4490 )
         );
  MUX \Reg_Bank/U4537  ( .A(\Reg_Bank/n4488 ), .B(\Reg_Bank/n4487 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4489 ) );
  MUX \Reg_Bank/U4536  ( .A(\Reg_Bank/registers[12][15] ), .B(
        \Reg_Bank/registers[13][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4488 )
         );
  MUX \Reg_Bank/U4535  ( .A(\Reg_Bank/registers[14][15] ), .B(
        \Reg_Bank/registers[15][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4487 )
         );
  MUX \Reg_Bank/U4534  ( .A(\Reg_Bank/n4485 ), .B(\Reg_Bank/n4478 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4486 ) );
  MUX \Reg_Bank/U4533  ( .A(\Reg_Bank/n4484 ), .B(\Reg_Bank/n4481 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4485 ) );
  MUX \Reg_Bank/U4532  ( .A(\Reg_Bank/n4483 ), .B(\Reg_Bank/n4482 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4484 ) );
  MUX \Reg_Bank/U4531  ( .A(\Reg_Bank/registers[16][15] ), .B(
        \Reg_Bank/registers[17][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4483 )
         );
  MUX \Reg_Bank/U4530  ( .A(\Reg_Bank/registers[18][15] ), .B(
        \Reg_Bank/registers[19][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4482 )
         );
  MUX \Reg_Bank/U4529  ( .A(\Reg_Bank/n4480 ), .B(\Reg_Bank/n4479 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4481 ) );
  MUX \Reg_Bank/U4528  ( .A(\Reg_Bank/registers[20][15] ), .B(
        \Reg_Bank/registers[21][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4480 )
         );
  MUX \Reg_Bank/U4527  ( .A(\Reg_Bank/registers[22][15] ), .B(
        \Reg_Bank/registers[23][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4479 )
         );
  MUX \Reg_Bank/U4526  ( .A(\Reg_Bank/n4477 ), .B(\Reg_Bank/n4474 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4478 ) );
  MUX \Reg_Bank/U4525  ( .A(\Reg_Bank/n4476 ), .B(\Reg_Bank/n4475 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4477 ) );
  MUX \Reg_Bank/U4524  ( .A(\Reg_Bank/registers[24][15] ), .B(
        \Reg_Bank/registers[25][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4476 )
         );
  MUX \Reg_Bank/U4523  ( .A(\Reg_Bank/registers[26][15] ), .B(
        \Reg_Bank/registers[27][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4475 )
         );
  MUX \Reg_Bank/U4522  ( .A(\Reg_Bank/n4473 ), .B(\Reg_Bank/n4472 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4474 ) );
  MUX \Reg_Bank/U4521  ( .A(\Reg_Bank/registers[28][15] ), .B(
        \Reg_Bank/registers[29][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4473 )
         );
  MUX \Reg_Bank/U4520  ( .A(\Reg_Bank/registers[30][15] ), .B(
        \Reg_Bank/registers[31][15] ), .S(rs_index[0]), .Z(\Reg_Bank/n4472 )
         );
  MUX \Reg_Bank/U4519  ( .A(\Reg_Bank/n4471 ), .B(\Reg_Bank/n4456 ), .S(
        rs_index[4]), .Z(reg_source[14]) );
  MUX \Reg_Bank/U4518  ( .A(\Reg_Bank/n4470 ), .B(\Reg_Bank/n4463 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4471 ) );
  MUX \Reg_Bank/U4517  ( .A(\Reg_Bank/n4469 ), .B(\Reg_Bank/n4466 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4470 ) );
  MUX \Reg_Bank/U4516  ( .A(\Reg_Bank/n4468 ), .B(\Reg_Bank/n4467 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4469 ) );
  MUX \Reg_Bank/U4514  ( .A(\Reg_Bank/registers[2][14] ), .B(
        \Reg_Bank/registers[3][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4467 ) );
  MUX \Reg_Bank/U4513  ( .A(\Reg_Bank/n4465 ), .B(\Reg_Bank/n4464 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4466 ) );
  MUX \Reg_Bank/U4512  ( .A(\Reg_Bank/registers[4][14] ), .B(
        \Reg_Bank/registers[5][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4465 ) );
  MUX \Reg_Bank/U4511  ( .A(\Reg_Bank/registers[6][14] ), .B(
        \Reg_Bank/registers[7][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4464 ) );
  MUX \Reg_Bank/U4510  ( .A(\Reg_Bank/n4462 ), .B(\Reg_Bank/n4459 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4463 ) );
  MUX \Reg_Bank/U4509  ( .A(\Reg_Bank/n4461 ), .B(\Reg_Bank/n4460 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4462 ) );
  MUX \Reg_Bank/U4508  ( .A(\Reg_Bank/registers[8][14] ), .B(
        \Reg_Bank/registers[9][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4461 ) );
  MUX \Reg_Bank/U4507  ( .A(\Reg_Bank/registers[10][14] ), .B(
        \Reg_Bank/registers[11][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4460 )
         );
  MUX \Reg_Bank/U4506  ( .A(\Reg_Bank/n4458 ), .B(\Reg_Bank/n4457 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4459 ) );
  MUX \Reg_Bank/U4505  ( .A(\Reg_Bank/registers[12][14] ), .B(
        \Reg_Bank/registers[13][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4458 )
         );
  MUX \Reg_Bank/U4504  ( .A(\Reg_Bank/registers[14][14] ), .B(
        \Reg_Bank/registers[15][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4457 )
         );
  MUX \Reg_Bank/U4503  ( .A(\Reg_Bank/n4455 ), .B(\Reg_Bank/n4448 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4456 ) );
  MUX \Reg_Bank/U4502  ( .A(\Reg_Bank/n4454 ), .B(\Reg_Bank/n4451 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4455 ) );
  MUX \Reg_Bank/U4501  ( .A(\Reg_Bank/n4453 ), .B(\Reg_Bank/n4452 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4454 ) );
  MUX \Reg_Bank/U4500  ( .A(\Reg_Bank/registers[16][14] ), .B(
        \Reg_Bank/registers[17][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4453 )
         );
  MUX \Reg_Bank/U4499  ( .A(\Reg_Bank/registers[18][14] ), .B(
        \Reg_Bank/registers[19][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4452 )
         );
  MUX \Reg_Bank/U4498  ( .A(\Reg_Bank/n4450 ), .B(\Reg_Bank/n4449 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4451 ) );
  MUX \Reg_Bank/U4497  ( .A(\Reg_Bank/registers[20][14] ), .B(
        \Reg_Bank/registers[21][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4450 )
         );
  MUX \Reg_Bank/U4496  ( .A(\Reg_Bank/registers[22][14] ), .B(
        \Reg_Bank/registers[23][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4449 )
         );
  MUX \Reg_Bank/U4495  ( .A(\Reg_Bank/n4447 ), .B(\Reg_Bank/n4444 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4448 ) );
  MUX \Reg_Bank/U4494  ( .A(\Reg_Bank/n4446 ), .B(\Reg_Bank/n4445 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4447 ) );
  MUX \Reg_Bank/U4493  ( .A(\Reg_Bank/registers[24][14] ), .B(
        \Reg_Bank/registers[25][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4446 )
         );
  MUX \Reg_Bank/U4492  ( .A(\Reg_Bank/registers[26][14] ), .B(
        \Reg_Bank/registers[27][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4445 )
         );
  MUX \Reg_Bank/U4491  ( .A(\Reg_Bank/n4443 ), .B(\Reg_Bank/n4442 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4444 ) );
  MUX \Reg_Bank/U4490  ( .A(\Reg_Bank/registers[28][14] ), .B(
        \Reg_Bank/registers[29][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4443 )
         );
  MUX \Reg_Bank/U4489  ( .A(\Reg_Bank/registers[30][14] ), .B(
        \Reg_Bank/registers[31][14] ), .S(rs_index[0]), .Z(\Reg_Bank/n4442 )
         );
  MUX \Reg_Bank/U4488  ( .A(\Reg_Bank/n4441 ), .B(\Reg_Bank/n4426 ), .S(
        rs_index[4]), .Z(reg_source[13]) );
  MUX \Reg_Bank/U4487  ( .A(\Reg_Bank/n4440 ), .B(\Reg_Bank/n4433 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4441 ) );
  MUX \Reg_Bank/U4486  ( .A(\Reg_Bank/n4439 ), .B(\Reg_Bank/n4436 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4440 ) );
  MUX \Reg_Bank/U4485  ( .A(\Reg_Bank/n4438 ), .B(\Reg_Bank/n4437 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4439 ) );
  MUX \Reg_Bank/U4483  ( .A(\Reg_Bank/registers[2][13] ), .B(
        \Reg_Bank/registers[3][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4437 ) );
  MUX \Reg_Bank/U4482  ( .A(\Reg_Bank/n4435 ), .B(\Reg_Bank/n4434 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4436 ) );
  MUX \Reg_Bank/U4481  ( .A(\Reg_Bank/registers[4][13] ), .B(
        \Reg_Bank/registers[5][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4435 ) );
  MUX \Reg_Bank/U4480  ( .A(\Reg_Bank/registers[6][13] ), .B(
        \Reg_Bank/registers[7][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4434 ) );
  MUX \Reg_Bank/U4479  ( .A(\Reg_Bank/n4432 ), .B(\Reg_Bank/n4429 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4433 ) );
  MUX \Reg_Bank/U4478  ( .A(\Reg_Bank/n4431 ), .B(\Reg_Bank/n4430 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4432 ) );
  MUX \Reg_Bank/U4477  ( .A(\Reg_Bank/registers[8][13] ), .B(
        \Reg_Bank/registers[9][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4431 ) );
  MUX \Reg_Bank/U4476  ( .A(\Reg_Bank/registers[10][13] ), .B(
        \Reg_Bank/registers[11][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4430 )
         );
  MUX \Reg_Bank/U4475  ( .A(\Reg_Bank/n4428 ), .B(\Reg_Bank/n4427 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4429 ) );
  MUX \Reg_Bank/U4474  ( .A(\Reg_Bank/registers[12][13] ), .B(
        \Reg_Bank/registers[13][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4428 )
         );
  MUX \Reg_Bank/U4473  ( .A(\Reg_Bank/registers[14][13] ), .B(
        \Reg_Bank/registers[15][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4427 )
         );
  MUX \Reg_Bank/U4472  ( .A(\Reg_Bank/n4425 ), .B(\Reg_Bank/n4418 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4426 ) );
  MUX \Reg_Bank/U4471  ( .A(\Reg_Bank/n4424 ), .B(\Reg_Bank/n4421 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4425 ) );
  MUX \Reg_Bank/U4470  ( .A(\Reg_Bank/n4423 ), .B(\Reg_Bank/n4422 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4424 ) );
  MUX \Reg_Bank/U4469  ( .A(\Reg_Bank/registers[16][13] ), .B(
        \Reg_Bank/registers[17][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4423 )
         );
  MUX \Reg_Bank/U4468  ( .A(\Reg_Bank/registers[18][13] ), .B(
        \Reg_Bank/registers[19][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4422 )
         );
  MUX \Reg_Bank/U4467  ( .A(\Reg_Bank/n4420 ), .B(\Reg_Bank/n4419 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4421 ) );
  MUX \Reg_Bank/U4466  ( .A(\Reg_Bank/registers[20][13] ), .B(
        \Reg_Bank/registers[21][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4420 )
         );
  MUX \Reg_Bank/U4465  ( .A(\Reg_Bank/registers[22][13] ), .B(
        \Reg_Bank/registers[23][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4419 )
         );
  MUX \Reg_Bank/U4464  ( .A(\Reg_Bank/n4417 ), .B(\Reg_Bank/n4414 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4418 ) );
  MUX \Reg_Bank/U4463  ( .A(\Reg_Bank/n4416 ), .B(\Reg_Bank/n4415 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4417 ) );
  MUX \Reg_Bank/U4462  ( .A(\Reg_Bank/registers[24][13] ), .B(
        \Reg_Bank/registers[25][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4416 )
         );
  MUX \Reg_Bank/U4461  ( .A(\Reg_Bank/registers[26][13] ), .B(
        \Reg_Bank/registers[27][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4415 )
         );
  MUX \Reg_Bank/U4460  ( .A(\Reg_Bank/n4413 ), .B(\Reg_Bank/n4412 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4414 ) );
  MUX \Reg_Bank/U4459  ( .A(\Reg_Bank/registers[28][13] ), .B(
        \Reg_Bank/registers[29][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4413 )
         );
  MUX \Reg_Bank/U4458  ( .A(\Reg_Bank/registers[30][13] ), .B(
        \Reg_Bank/registers[31][13] ), .S(rs_index[0]), .Z(\Reg_Bank/n4412 )
         );
  MUX \Reg_Bank/U4457  ( .A(\Reg_Bank/n4411 ), .B(\Reg_Bank/n4396 ), .S(
        rs_index[4]), .Z(reg_source[12]) );
  MUX \Reg_Bank/U4456  ( .A(\Reg_Bank/n4410 ), .B(\Reg_Bank/n4403 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4411 ) );
  MUX \Reg_Bank/U4455  ( .A(\Reg_Bank/n4409 ), .B(\Reg_Bank/n4406 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4410 ) );
  MUX \Reg_Bank/U4454  ( .A(\Reg_Bank/n4408 ), .B(\Reg_Bank/n4407 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4409 ) );
  MUX \Reg_Bank/U4452  ( .A(\Reg_Bank/registers[2][12] ), .B(
        \Reg_Bank/registers[3][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4407 ) );
  MUX \Reg_Bank/U4451  ( .A(\Reg_Bank/n4405 ), .B(\Reg_Bank/n4404 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4406 ) );
  MUX \Reg_Bank/U4450  ( .A(\Reg_Bank/registers[4][12] ), .B(
        \Reg_Bank/registers[5][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4405 ) );
  MUX \Reg_Bank/U4449  ( .A(\Reg_Bank/registers[6][12] ), .B(
        \Reg_Bank/registers[7][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4404 ) );
  MUX \Reg_Bank/U4448  ( .A(\Reg_Bank/n4402 ), .B(\Reg_Bank/n4399 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4403 ) );
  MUX \Reg_Bank/U4447  ( .A(\Reg_Bank/n4401 ), .B(\Reg_Bank/n4400 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4402 ) );
  MUX \Reg_Bank/U4446  ( .A(\Reg_Bank/registers[8][12] ), .B(
        \Reg_Bank/registers[9][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4401 ) );
  MUX \Reg_Bank/U4445  ( .A(\Reg_Bank/registers[10][12] ), .B(
        \Reg_Bank/registers[11][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4400 )
         );
  MUX \Reg_Bank/U4444  ( .A(\Reg_Bank/n4398 ), .B(\Reg_Bank/n4397 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4399 ) );
  MUX \Reg_Bank/U4443  ( .A(\Reg_Bank/registers[12][12] ), .B(
        \Reg_Bank/registers[13][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4398 )
         );
  MUX \Reg_Bank/U4442  ( .A(\Reg_Bank/registers[14][12] ), .B(
        \Reg_Bank/registers[15][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4397 )
         );
  MUX \Reg_Bank/U4441  ( .A(\Reg_Bank/n4395 ), .B(\Reg_Bank/n4388 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4396 ) );
  MUX \Reg_Bank/U4440  ( .A(\Reg_Bank/n4394 ), .B(\Reg_Bank/n4391 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4395 ) );
  MUX \Reg_Bank/U4439  ( .A(\Reg_Bank/n4393 ), .B(\Reg_Bank/n4392 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4394 ) );
  MUX \Reg_Bank/U4438  ( .A(\Reg_Bank/registers[16][12] ), .B(
        \Reg_Bank/registers[17][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4393 )
         );
  MUX \Reg_Bank/U4437  ( .A(\Reg_Bank/registers[18][12] ), .B(
        \Reg_Bank/registers[19][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4392 )
         );
  MUX \Reg_Bank/U4436  ( .A(\Reg_Bank/n4390 ), .B(\Reg_Bank/n4389 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4391 ) );
  MUX \Reg_Bank/U4435  ( .A(\Reg_Bank/registers[20][12] ), .B(
        \Reg_Bank/registers[21][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4390 )
         );
  MUX \Reg_Bank/U4434  ( .A(\Reg_Bank/registers[22][12] ), .B(
        \Reg_Bank/registers[23][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4389 )
         );
  MUX \Reg_Bank/U4433  ( .A(\Reg_Bank/n4387 ), .B(\Reg_Bank/n4384 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4388 ) );
  MUX \Reg_Bank/U4432  ( .A(\Reg_Bank/n4386 ), .B(\Reg_Bank/n4385 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4387 ) );
  MUX \Reg_Bank/U4431  ( .A(\Reg_Bank/registers[24][12] ), .B(
        \Reg_Bank/registers[25][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4386 )
         );
  MUX \Reg_Bank/U4430  ( .A(\Reg_Bank/registers[26][12] ), .B(
        \Reg_Bank/registers[27][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4385 )
         );
  MUX \Reg_Bank/U4429  ( .A(\Reg_Bank/n4383 ), .B(\Reg_Bank/n4382 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4384 ) );
  MUX \Reg_Bank/U4428  ( .A(\Reg_Bank/registers[28][12] ), .B(
        \Reg_Bank/registers[29][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4383 )
         );
  MUX \Reg_Bank/U4427  ( .A(\Reg_Bank/registers[30][12] ), .B(
        \Reg_Bank/registers[31][12] ), .S(rs_index[0]), .Z(\Reg_Bank/n4382 )
         );
  MUX \Reg_Bank/U4426  ( .A(\Reg_Bank/n4381 ), .B(\Reg_Bank/n4366 ), .S(
        rs_index[4]), .Z(reg_source[11]) );
  MUX \Reg_Bank/U4425  ( .A(\Reg_Bank/n4380 ), .B(\Reg_Bank/n4373 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4381 ) );
  MUX \Reg_Bank/U4424  ( .A(\Reg_Bank/n4379 ), .B(\Reg_Bank/n4376 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4380 ) );
  MUX \Reg_Bank/U4423  ( .A(\Reg_Bank/n4378 ), .B(\Reg_Bank/n4377 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4379 ) );
  MUX \Reg_Bank/U4421  ( .A(\Reg_Bank/registers[2][11] ), .B(
        \Reg_Bank/registers[3][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4377 ) );
  MUX \Reg_Bank/U4420  ( .A(\Reg_Bank/n4375 ), .B(\Reg_Bank/n4374 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4376 ) );
  MUX \Reg_Bank/U4419  ( .A(\Reg_Bank/registers[4][11] ), .B(
        \Reg_Bank/registers[5][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4375 ) );
  MUX \Reg_Bank/U4418  ( .A(\Reg_Bank/registers[6][11] ), .B(
        \Reg_Bank/registers[7][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4374 ) );
  MUX \Reg_Bank/U4417  ( .A(\Reg_Bank/n4372 ), .B(\Reg_Bank/n4369 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4373 ) );
  MUX \Reg_Bank/U4416  ( .A(\Reg_Bank/n4371 ), .B(\Reg_Bank/n4370 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4372 ) );
  MUX \Reg_Bank/U4415  ( .A(\Reg_Bank/registers[8][11] ), .B(
        \Reg_Bank/registers[9][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4371 ) );
  MUX \Reg_Bank/U4414  ( .A(\Reg_Bank/registers[10][11] ), .B(
        \Reg_Bank/registers[11][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4370 )
         );
  MUX \Reg_Bank/U4413  ( .A(\Reg_Bank/n4368 ), .B(\Reg_Bank/n4367 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4369 ) );
  MUX \Reg_Bank/U4412  ( .A(\Reg_Bank/registers[12][11] ), .B(
        \Reg_Bank/registers[13][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4368 )
         );
  MUX \Reg_Bank/U4411  ( .A(\Reg_Bank/registers[14][11] ), .B(
        \Reg_Bank/registers[15][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4367 )
         );
  MUX \Reg_Bank/U4410  ( .A(\Reg_Bank/n4365 ), .B(\Reg_Bank/n4358 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4366 ) );
  MUX \Reg_Bank/U4409  ( .A(\Reg_Bank/n4364 ), .B(\Reg_Bank/n4361 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4365 ) );
  MUX \Reg_Bank/U4408  ( .A(\Reg_Bank/n4363 ), .B(\Reg_Bank/n4362 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4364 ) );
  MUX \Reg_Bank/U4407  ( .A(\Reg_Bank/registers[16][11] ), .B(
        \Reg_Bank/registers[17][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4363 )
         );
  MUX \Reg_Bank/U4406  ( .A(\Reg_Bank/registers[18][11] ), .B(
        \Reg_Bank/registers[19][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4362 )
         );
  MUX \Reg_Bank/U4405  ( .A(\Reg_Bank/n4360 ), .B(\Reg_Bank/n4359 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4361 ) );
  MUX \Reg_Bank/U4404  ( .A(\Reg_Bank/registers[20][11] ), .B(
        \Reg_Bank/registers[21][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4360 )
         );
  MUX \Reg_Bank/U4403  ( .A(\Reg_Bank/registers[22][11] ), .B(
        \Reg_Bank/registers[23][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4359 )
         );
  MUX \Reg_Bank/U4402  ( .A(\Reg_Bank/n4357 ), .B(\Reg_Bank/n4354 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4358 ) );
  MUX \Reg_Bank/U4401  ( .A(\Reg_Bank/n4356 ), .B(\Reg_Bank/n4355 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4357 ) );
  MUX \Reg_Bank/U4400  ( .A(\Reg_Bank/registers[24][11] ), .B(
        \Reg_Bank/registers[25][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4356 )
         );
  MUX \Reg_Bank/U4399  ( .A(\Reg_Bank/registers[26][11] ), .B(
        \Reg_Bank/registers[27][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4355 )
         );
  MUX \Reg_Bank/U4398  ( .A(\Reg_Bank/n4353 ), .B(\Reg_Bank/n4352 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4354 ) );
  MUX \Reg_Bank/U4397  ( .A(\Reg_Bank/registers[28][11] ), .B(
        \Reg_Bank/registers[29][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4353 )
         );
  MUX \Reg_Bank/U4396  ( .A(\Reg_Bank/registers[30][11] ), .B(
        \Reg_Bank/registers[31][11] ), .S(rs_index[0]), .Z(\Reg_Bank/n4352 )
         );
  MUX \Reg_Bank/U4395  ( .A(\Reg_Bank/n4351 ), .B(\Reg_Bank/n4336 ), .S(
        rs_index[4]), .Z(reg_source[10]) );
  MUX \Reg_Bank/U4394  ( .A(\Reg_Bank/n4350 ), .B(\Reg_Bank/n4343 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4351 ) );
  MUX \Reg_Bank/U4393  ( .A(\Reg_Bank/n4349 ), .B(\Reg_Bank/n4346 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4350 ) );
  MUX \Reg_Bank/U4392  ( .A(\Reg_Bank/n4348 ), .B(\Reg_Bank/n4347 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4349 ) );
  MUX \Reg_Bank/U4390  ( .A(\Reg_Bank/registers[2][10] ), .B(
        \Reg_Bank/registers[3][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4347 ) );
  MUX \Reg_Bank/U4389  ( .A(\Reg_Bank/n4345 ), .B(\Reg_Bank/n4344 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4346 ) );
  MUX \Reg_Bank/U4388  ( .A(\Reg_Bank/registers[4][10] ), .B(
        \Reg_Bank/registers[5][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4345 ) );
  MUX \Reg_Bank/U4387  ( .A(\Reg_Bank/registers[6][10] ), .B(
        \Reg_Bank/registers[7][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4344 ) );
  MUX \Reg_Bank/U4386  ( .A(\Reg_Bank/n4342 ), .B(\Reg_Bank/n4339 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4343 ) );
  MUX \Reg_Bank/U4385  ( .A(\Reg_Bank/n4341 ), .B(\Reg_Bank/n4340 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4342 ) );
  MUX \Reg_Bank/U4384  ( .A(\Reg_Bank/registers[8][10] ), .B(
        \Reg_Bank/registers[9][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4341 ) );
  MUX \Reg_Bank/U4383  ( .A(\Reg_Bank/registers[10][10] ), .B(
        \Reg_Bank/registers[11][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4340 )
         );
  MUX \Reg_Bank/U4382  ( .A(\Reg_Bank/n4338 ), .B(\Reg_Bank/n4337 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4339 ) );
  MUX \Reg_Bank/U4381  ( .A(\Reg_Bank/registers[12][10] ), .B(
        \Reg_Bank/registers[13][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4338 )
         );
  MUX \Reg_Bank/U4380  ( .A(\Reg_Bank/registers[14][10] ), .B(
        \Reg_Bank/registers[15][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4337 )
         );
  MUX \Reg_Bank/U4379  ( .A(\Reg_Bank/n4335 ), .B(\Reg_Bank/n4328 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4336 ) );
  MUX \Reg_Bank/U4378  ( .A(\Reg_Bank/n4334 ), .B(\Reg_Bank/n4331 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4335 ) );
  MUX \Reg_Bank/U4377  ( .A(\Reg_Bank/n4333 ), .B(\Reg_Bank/n4332 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4334 ) );
  MUX \Reg_Bank/U4376  ( .A(\Reg_Bank/registers[16][10] ), .B(
        \Reg_Bank/registers[17][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4333 )
         );
  MUX \Reg_Bank/U4375  ( .A(\Reg_Bank/registers[18][10] ), .B(
        \Reg_Bank/registers[19][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4332 )
         );
  MUX \Reg_Bank/U4374  ( .A(\Reg_Bank/n4330 ), .B(\Reg_Bank/n4329 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4331 ) );
  MUX \Reg_Bank/U4373  ( .A(\Reg_Bank/registers[20][10] ), .B(
        \Reg_Bank/registers[21][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4330 )
         );
  MUX \Reg_Bank/U4372  ( .A(\Reg_Bank/registers[22][10] ), .B(
        \Reg_Bank/registers[23][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4329 )
         );
  MUX \Reg_Bank/U4371  ( .A(\Reg_Bank/n4327 ), .B(\Reg_Bank/n4324 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4328 ) );
  MUX \Reg_Bank/U4370  ( .A(\Reg_Bank/n4326 ), .B(\Reg_Bank/n4325 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4327 ) );
  MUX \Reg_Bank/U4369  ( .A(\Reg_Bank/registers[24][10] ), .B(
        \Reg_Bank/registers[25][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4326 )
         );
  MUX \Reg_Bank/U4368  ( .A(\Reg_Bank/registers[26][10] ), .B(
        \Reg_Bank/registers[27][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4325 )
         );
  MUX \Reg_Bank/U4367  ( .A(\Reg_Bank/n4323 ), .B(\Reg_Bank/n4322 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4324 ) );
  MUX \Reg_Bank/U4366  ( .A(\Reg_Bank/registers[28][10] ), .B(
        \Reg_Bank/registers[29][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4323 )
         );
  MUX \Reg_Bank/U4365  ( .A(\Reg_Bank/registers[30][10] ), .B(
        \Reg_Bank/registers[31][10] ), .S(rs_index[0]), .Z(\Reg_Bank/n4322 )
         );
  MUX \Reg_Bank/U4364  ( .A(\Reg_Bank/n4321 ), .B(\Reg_Bank/n4306 ), .S(
        rs_index[4]), .Z(reg_source[9]) );
  MUX \Reg_Bank/U4363  ( .A(\Reg_Bank/n4320 ), .B(\Reg_Bank/n4313 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4321 ) );
  MUX \Reg_Bank/U4362  ( .A(\Reg_Bank/n4319 ), .B(\Reg_Bank/n4316 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4320 ) );
  MUX \Reg_Bank/U4361  ( .A(\Reg_Bank/n4318 ), .B(\Reg_Bank/n4317 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4319 ) );
  MUX \Reg_Bank/U4359  ( .A(\Reg_Bank/registers[2][9] ), .B(
        \Reg_Bank/registers[3][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4317 ) );
  MUX \Reg_Bank/U4358  ( .A(\Reg_Bank/n4315 ), .B(\Reg_Bank/n4314 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4316 ) );
  MUX \Reg_Bank/U4357  ( .A(\Reg_Bank/registers[4][9] ), .B(
        \Reg_Bank/registers[5][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4315 ) );
  MUX \Reg_Bank/U4356  ( .A(\Reg_Bank/registers[6][9] ), .B(
        \Reg_Bank/registers[7][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4314 ) );
  MUX \Reg_Bank/U4355  ( .A(\Reg_Bank/n4312 ), .B(\Reg_Bank/n4309 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4313 ) );
  MUX \Reg_Bank/U4354  ( .A(\Reg_Bank/n4311 ), .B(\Reg_Bank/n4310 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4312 ) );
  MUX \Reg_Bank/U4353  ( .A(\Reg_Bank/registers[8][9] ), .B(
        \Reg_Bank/registers[9][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4311 ) );
  MUX \Reg_Bank/U4352  ( .A(\Reg_Bank/registers[10][9] ), .B(
        \Reg_Bank/registers[11][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4310 ) );
  MUX \Reg_Bank/U4351  ( .A(\Reg_Bank/n4308 ), .B(\Reg_Bank/n4307 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4309 ) );
  MUX \Reg_Bank/U4350  ( .A(\Reg_Bank/registers[12][9] ), .B(
        \Reg_Bank/registers[13][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4308 ) );
  MUX \Reg_Bank/U4349  ( .A(\Reg_Bank/registers[14][9] ), .B(
        \Reg_Bank/registers[15][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4307 ) );
  MUX \Reg_Bank/U4348  ( .A(\Reg_Bank/n4305 ), .B(\Reg_Bank/n4298 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4306 ) );
  MUX \Reg_Bank/U4347  ( .A(\Reg_Bank/n4304 ), .B(\Reg_Bank/n4301 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4305 ) );
  MUX \Reg_Bank/U4346  ( .A(\Reg_Bank/n4303 ), .B(\Reg_Bank/n4302 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4304 ) );
  MUX \Reg_Bank/U4345  ( .A(\Reg_Bank/registers[16][9] ), .B(
        \Reg_Bank/registers[17][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4303 ) );
  MUX \Reg_Bank/U4344  ( .A(\Reg_Bank/registers[18][9] ), .B(
        \Reg_Bank/registers[19][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4302 ) );
  MUX \Reg_Bank/U4343  ( .A(\Reg_Bank/n4300 ), .B(\Reg_Bank/n4299 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4301 ) );
  MUX \Reg_Bank/U4342  ( .A(\Reg_Bank/registers[20][9] ), .B(
        \Reg_Bank/registers[21][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4300 ) );
  MUX \Reg_Bank/U4341  ( .A(\Reg_Bank/registers[22][9] ), .B(
        \Reg_Bank/registers[23][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4299 ) );
  MUX \Reg_Bank/U4340  ( .A(\Reg_Bank/n4297 ), .B(\Reg_Bank/n4294 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4298 ) );
  MUX \Reg_Bank/U4339  ( .A(\Reg_Bank/n4296 ), .B(\Reg_Bank/n4295 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4297 ) );
  MUX \Reg_Bank/U4338  ( .A(\Reg_Bank/registers[24][9] ), .B(
        \Reg_Bank/registers[25][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4296 ) );
  MUX \Reg_Bank/U4337  ( .A(\Reg_Bank/registers[26][9] ), .B(
        \Reg_Bank/registers[27][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4295 ) );
  MUX \Reg_Bank/U4336  ( .A(\Reg_Bank/n4293 ), .B(\Reg_Bank/n4292 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4294 ) );
  MUX \Reg_Bank/U4335  ( .A(\Reg_Bank/registers[28][9] ), .B(
        \Reg_Bank/registers[29][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4293 ) );
  MUX \Reg_Bank/U4334  ( .A(\Reg_Bank/registers[30][9] ), .B(
        \Reg_Bank/registers[31][9] ), .S(rs_index[0]), .Z(\Reg_Bank/n4292 ) );
  MUX \Reg_Bank/U4333  ( .A(\Reg_Bank/n4291 ), .B(\Reg_Bank/n4276 ), .S(
        rs_index[4]), .Z(reg_source[8]) );
  MUX \Reg_Bank/U4332  ( .A(\Reg_Bank/n4290 ), .B(\Reg_Bank/n4283 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4291 ) );
  MUX \Reg_Bank/U4331  ( .A(\Reg_Bank/n4289 ), .B(\Reg_Bank/n4286 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4290 ) );
  MUX \Reg_Bank/U4330  ( .A(\Reg_Bank/n4288 ), .B(\Reg_Bank/n4287 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4289 ) );
  MUX \Reg_Bank/U4328  ( .A(\Reg_Bank/registers[2][8] ), .B(
        \Reg_Bank/registers[3][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4287 ) );
  MUX \Reg_Bank/U4327  ( .A(\Reg_Bank/n4285 ), .B(\Reg_Bank/n4284 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4286 ) );
  MUX \Reg_Bank/U4326  ( .A(\Reg_Bank/registers[4][8] ), .B(
        \Reg_Bank/registers[5][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4285 ) );
  MUX \Reg_Bank/U4325  ( .A(\Reg_Bank/registers[6][8] ), .B(
        \Reg_Bank/registers[7][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4284 ) );
  MUX \Reg_Bank/U4324  ( .A(\Reg_Bank/n4282 ), .B(\Reg_Bank/n4279 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4283 ) );
  MUX \Reg_Bank/U4323  ( .A(\Reg_Bank/n4281 ), .B(\Reg_Bank/n4280 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4282 ) );
  MUX \Reg_Bank/U4322  ( .A(\Reg_Bank/registers[8][8] ), .B(
        \Reg_Bank/registers[9][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4281 ) );
  MUX \Reg_Bank/U4321  ( .A(\Reg_Bank/registers[10][8] ), .B(
        \Reg_Bank/registers[11][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4280 ) );
  MUX \Reg_Bank/U4320  ( .A(\Reg_Bank/n4278 ), .B(\Reg_Bank/n4277 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4279 ) );
  MUX \Reg_Bank/U4319  ( .A(\Reg_Bank/registers[12][8] ), .B(
        \Reg_Bank/registers[13][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4278 ) );
  MUX \Reg_Bank/U4318  ( .A(\Reg_Bank/registers[14][8] ), .B(
        \Reg_Bank/registers[15][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4277 ) );
  MUX \Reg_Bank/U4317  ( .A(\Reg_Bank/n4275 ), .B(\Reg_Bank/n4268 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4276 ) );
  MUX \Reg_Bank/U4316  ( .A(\Reg_Bank/n4274 ), .B(\Reg_Bank/n4271 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4275 ) );
  MUX \Reg_Bank/U4315  ( .A(\Reg_Bank/n4273 ), .B(\Reg_Bank/n4272 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4274 ) );
  MUX \Reg_Bank/U4314  ( .A(\Reg_Bank/registers[16][8] ), .B(
        \Reg_Bank/registers[17][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4273 ) );
  MUX \Reg_Bank/U4313  ( .A(\Reg_Bank/registers[18][8] ), .B(
        \Reg_Bank/registers[19][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4272 ) );
  MUX \Reg_Bank/U4312  ( .A(\Reg_Bank/n4270 ), .B(\Reg_Bank/n4269 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4271 ) );
  MUX \Reg_Bank/U4311  ( .A(\Reg_Bank/registers[20][8] ), .B(
        \Reg_Bank/registers[21][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4270 ) );
  MUX \Reg_Bank/U4310  ( .A(\Reg_Bank/registers[22][8] ), .B(
        \Reg_Bank/registers[23][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4269 ) );
  MUX \Reg_Bank/U4309  ( .A(\Reg_Bank/n4267 ), .B(\Reg_Bank/n4264 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4268 ) );
  MUX \Reg_Bank/U4308  ( .A(\Reg_Bank/n4266 ), .B(\Reg_Bank/n4265 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4267 ) );
  MUX \Reg_Bank/U4307  ( .A(\Reg_Bank/registers[24][8] ), .B(
        \Reg_Bank/registers[25][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4266 ) );
  MUX \Reg_Bank/U4306  ( .A(\Reg_Bank/registers[26][8] ), .B(
        \Reg_Bank/registers[27][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4265 ) );
  MUX \Reg_Bank/U4305  ( .A(\Reg_Bank/n4263 ), .B(\Reg_Bank/n4262 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4264 ) );
  MUX \Reg_Bank/U4304  ( .A(\Reg_Bank/registers[28][8] ), .B(
        \Reg_Bank/registers[29][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4263 ) );
  MUX \Reg_Bank/U4303  ( .A(\Reg_Bank/registers[30][8] ), .B(
        \Reg_Bank/registers[31][8] ), .S(rs_index[0]), .Z(\Reg_Bank/n4262 ) );
  MUX \Reg_Bank/U4302  ( .A(\Reg_Bank/n4261 ), .B(\Reg_Bank/n4246 ), .S(
        rs_index[4]), .Z(reg_source[7]) );
  MUX \Reg_Bank/U4301  ( .A(\Reg_Bank/n4260 ), .B(\Reg_Bank/n4253 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4261 ) );
  MUX \Reg_Bank/U4300  ( .A(\Reg_Bank/n4259 ), .B(\Reg_Bank/n4256 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4260 ) );
  MUX \Reg_Bank/U4299  ( .A(\Reg_Bank/n4258 ), .B(\Reg_Bank/n4257 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4259 ) );
  MUX \Reg_Bank/U4297  ( .A(\Reg_Bank/registers[2][7] ), .B(
        \Reg_Bank/registers[3][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4257 ) );
  MUX \Reg_Bank/U4296  ( .A(\Reg_Bank/n4255 ), .B(\Reg_Bank/n4254 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4256 ) );
  MUX \Reg_Bank/U4295  ( .A(\Reg_Bank/registers[4][7] ), .B(
        \Reg_Bank/registers[5][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4255 ) );
  MUX \Reg_Bank/U4294  ( .A(\Reg_Bank/registers[6][7] ), .B(
        \Reg_Bank/registers[7][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4254 ) );
  MUX \Reg_Bank/U4293  ( .A(\Reg_Bank/n4252 ), .B(\Reg_Bank/n4249 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4253 ) );
  MUX \Reg_Bank/U4292  ( .A(\Reg_Bank/n4251 ), .B(\Reg_Bank/n4250 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4252 ) );
  MUX \Reg_Bank/U4291  ( .A(\Reg_Bank/registers[8][7] ), .B(
        \Reg_Bank/registers[9][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4251 ) );
  MUX \Reg_Bank/U4290  ( .A(\Reg_Bank/registers[10][7] ), .B(
        \Reg_Bank/registers[11][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4250 ) );
  MUX \Reg_Bank/U4289  ( .A(\Reg_Bank/n4248 ), .B(\Reg_Bank/n4247 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4249 ) );
  MUX \Reg_Bank/U4288  ( .A(\Reg_Bank/registers[12][7] ), .B(
        \Reg_Bank/registers[13][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4248 ) );
  MUX \Reg_Bank/U4287  ( .A(\Reg_Bank/registers[14][7] ), .B(
        \Reg_Bank/registers[15][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4247 ) );
  MUX \Reg_Bank/U4286  ( .A(\Reg_Bank/n4245 ), .B(\Reg_Bank/n4238 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4246 ) );
  MUX \Reg_Bank/U4285  ( .A(\Reg_Bank/n4244 ), .B(\Reg_Bank/n4241 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4245 ) );
  MUX \Reg_Bank/U4284  ( .A(\Reg_Bank/n4243 ), .B(\Reg_Bank/n4242 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4244 ) );
  MUX \Reg_Bank/U4283  ( .A(\Reg_Bank/registers[16][7] ), .B(
        \Reg_Bank/registers[17][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4243 ) );
  MUX \Reg_Bank/U4282  ( .A(\Reg_Bank/registers[18][7] ), .B(
        \Reg_Bank/registers[19][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4242 ) );
  MUX \Reg_Bank/U4281  ( .A(\Reg_Bank/n4240 ), .B(\Reg_Bank/n4239 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4241 ) );
  MUX \Reg_Bank/U4280  ( .A(\Reg_Bank/registers[20][7] ), .B(
        \Reg_Bank/registers[21][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4240 ) );
  MUX \Reg_Bank/U4279  ( .A(\Reg_Bank/registers[22][7] ), .B(
        \Reg_Bank/registers[23][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4239 ) );
  MUX \Reg_Bank/U4278  ( .A(\Reg_Bank/n4237 ), .B(\Reg_Bank/n4234 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4238 ) );
  MUX \Reg_Bank/U4277  ( .A(\Reg_Bank/n4236 ), .B(\Reg_Bank/n4235 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4237 ) );
  MUX \Reg_Bank/U4276  ( .A(\Reg_Bank/registers[24][7] ), .B(
        \Reg_Bank/registers[25][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4236 ) );
  MUX \Reg_Bank/U4275  ( .A(\Reg_Bank/registers[26][7] ), .B(
        \Reg_Bank/registers[27][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4235 ) );
  MUX \Reg_Bank/U4274  ( .A(\Reg_Bank/n4233 ), .B(\Reg_Bank/n4232 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4234 ) );
  MUX \Reg_Bank/U4273  ( .A(\Reg_Bank/registers[28][7] ), .B(
        \Reg_Bank/registers[29][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4233 ) );
  MUX \Reg_Bank/U4272  ( .A(\Reg_Bank/registers[30][7] ), .B(
        \Reg_Bank/registers[31][7] ), .S(rs_index[0]), .Z(\Reg_Bank/n4232 ) );
  MUX \Reg_Bank/U4271  ( .A(\Reg_Bank/n4231 ), .B(\Reg_Bank/n4216 ), .S(
        rs_index[4]), .Z(reg_source[6]) );
  MUX \Reg_Bank/U4270  ( .A(\Reg_Bank/n4230 ), .B(\Reg_Bank/n4223 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4231 ) );
  MUX \Reg_Bank/U4269  ( .A(\Reg_Bank/n4229 ), .B(\Reg_Bank/n4226 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4230 ) );
  MUX \Reg_Bank/U4268  ( .A(\Reg_Bank/n4228 ), .B(\Reg_Bank/n4227 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4229 ) );
  MUX \Reg_Bank/U4266  ( .A(\Reg_Bank/registers[2][6] ), .B(
        \Reg_Bank/registers[3][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4227 ) );
  MUX \Reg_Bank/U4265  ( .A(\Reg_Bank/n4225 ), .B(\Reg_Bank/n4224 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4226 ) );
  MUX \Reg_Bank/U4264  ( .A(\Reg_Bank/registers[4][6] ), .B(
        \Reg_Bank/registers[5][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4225 ) );
  MUX \Reg_Bank/U4263  ( .A(\Reg_Bank/registers[6][6] ), .B(
        \Reg_Bank/registers[7][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4224 ) );
  MUX \Reg_Bank/U4262  ( .A(\Reg_Bank/n4222 ), .B(\Reg_Bank/n4219 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4223 ) );
  MUX \Reg_Bank/U4261  ( .A(\Reg_Bank/n4221 ), .B(\Reg_Bank/n4220 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4222 ) );
  MUX \Reg_Bank/U4260  ( .A(\Reg_Bank/registers[8][6] ), .B(
        \Reg_Bank/registers[9][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4221 ) );
  MUX \Reg_Bank/U4259  ( .A(\Reg_Bank/registers[10][6] ), .B(
        \Reg_Bank/registers[11][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4220 ) );
  MUX \Reg_Bank/U4258  ( .A(\Reg_Bank/n4218 ), .B(\Reg_Bank/n4217 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4219 ) );
  MUX \Reg_Bank/U4257  ( .A(\Reg_Bank/registers[12][6] ), .B(
        \Reg_Bank/registers[13][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4218 ) );
  MUX \Reg_Bank/U4256  ( .A(\Reg_Bank/registers[14][6] ), .B(
        \Reg_Bank/registers[15][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4217 ) );
  MUX \Reg_Bank/U4255  ( .A(\Reg_Bank/n4215 ), .B(\Reg_Bank/n4208 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4216 ) );
  MUX \Reg_Bank/U4254  ( .A(\Reg_Bank/n4214 ), .B(\Reg_Bank/n4211 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4215 ) );
  MUX \Reg_Bank/U4253  ( .A(\Reg_Bank/n4213 ), .B(\Reg_Bank/n4212 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4214 ) );
  MUX \Reg_Bank/U4252  ( .A(\Reg_Bank/registers[16][6] ), .B(
        \Reg_Bank/registers[17][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4213 ) );
  MUX \Reg_Bank/U4251  ( .A(\Reg_Bank/registers[18][6] ), .B(
        \Reg_Bank/registers[19][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4212 ) );
  MUX \Reg_Bank/U4250  ( .A(\Reg_Bank/n4210 ), .B(\Reg_Bank/n4209 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4211 ) );
  MUX \Reg_Bank/U4249  ( .A(\Reg_Bank/registers[20][6] ), .B(
        \Reg_Bank/registers[21][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4210 ) );
  MUX \Reg_Bank/U4248  ( .A(\Reg_Bank/registers[22][6] ), .B(
        \Reg_Bank/registers[23][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4209 ) );
  MUX \Reg_Bank/U4247  ( .A(\Reg_Bank/n4207 ), .B(\Reg_Bank/n4204 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4208 ) );
  MUX \Reg_Bank/U4246  ( .A(\Reg_Bank/n4206 ), .B(\Reg_Bank/n4205 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4207 ) );
  MUX \Reg_Bank/U4245  ( .A(\Reg_Bank/registers[24][6] ), .B(
        \Reg_Bank/registers[25][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4206 ) );
  MUX \Reg_Bank/U4244  ( .A(\Reg_Bank/registers[26][6] ), .B(
        \Reg_Bank/registers[27][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4205 ) );
  MUX \Reg_Bank/U4243  ( .A(\Reg_Bank/n4203 ), .B(\Reg_Bank/n4202 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4204 ) );
  MUX \Reg_Bank/U4242  ( .A(\Reg_Bank/registers[28][6] ), .B(
        \Reg_Bank/registers[29][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4203 ) );
  MUX \Reg_Bank/U4241  ( .A(\Reg_Bank/registers[30][6] ), .B(
        \Reg_Bank/registers[31][6] ), .S(rs_index[0]), .Z(\Reg_Bank/n4202 ) );
  MUX \Reg_Bank/U4240  ( .A(\Reg_Bank/n4201 ), .B(\Reg_Bank/n4186 ), .S(
        rs_index[4]), .Z(reg_source[5]) );
  MUX \Reg_Bank/U4239  ( .A(\Reg_Bank/n4200 ), .B(\Reg_Bank/n4193 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4201 ) );
  MUX \Reg_Bank/U4238  ( .A(\Reg_Bank/n4199 ), .B(\Reg_Bank/n4196 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4200 ) );
  MUX \Reg_Bank/U4237  ( .A(\Reg_Bank/n4198 ), .B(\Reg_Bank/n4197 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4199 ) );
  MUX \Reg_Bank/U4235  ( .A(\Reg_Bank/registers[2][5] ), .B(
        \Reg_Bank/registers[3][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4197 ) );
  MUX \Reg_Bank/U4234  ( .A(\Reg_Bank/n4195 ), .B(\Reg_Bank/n4194 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4196 ) );
  MUX \Reg_Bank/U4233  ( .A(\Reg_Bank/registers[4][5] ), .B(
        \Reg_Bank/registers[5][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4195 ) );
  MUX \Reg_Bank/U4232  ( .A(\Reg_Bank/registers[6][5] ), .B(
        \Reg_Bank/registers[7][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4194 ) );
  MUX \Reg_Bank/U4231  ( .A(\Reg_Bank/n4192 ), .B(\Reg_Bank/n4189 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4193 ) );
  MUX \Reg_Bank/U4230  ( .A(\Reg_Bank/n4191 ), .B(\Reg_Bank/n4190 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4192 ) );
  MUX \Reg_Bank/U4229  ( .A(\Reg_Bank/registers[8][5] ), .B(
        \Reg_Bank/registers[9][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4191 ) );
  MUX \Reg_Bank/U4228  ( .A(\Reg_Bank/registers[10][5] ), .B(
        \Reg_Bank/registers[11][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4190 ) );
  MUX \Reg_Bank/U4227  ( .A(\Reg_Bank/n4188 ), .B(\Reg_Bank/n4187 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4189 ) );
  MUX \Reg_Bank/U4226  ( .A(\Reg_Bank/registers[12][5] ), .B(
        \Reg_Bank/registers[13][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4188 ) );
  MUX \Reg_Bank/U4225  ( .A(\Reg_Bank/registers[14][5] ), .B(
        \Reg_Bank/registers[15][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4187 ) );
  MUX \Reg_Bank/U4224  ( .A(\Reg_Bank/n4185 ), .B(\Reg_Bank/n4178 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4186 ) );
  MUX \Reg_Bank/U4223  ( .A(\Reg_Bank/n4184 ), .B(\Reg_Bank/n4181 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4185 ) );
  MUX \Reg_Bank/U4222  ( .A(\Reg_Bank/n4183 ), .B(\Reg_Bank/n4182 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4184 ) );
  MUX \Reg_Bank/U4221  ( .A(\Reg_Bank/registers[16][5] ), .B(
        \Reg_Bank/registers[17][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4183 ) );
  MUX \Reg_Bank/U4220  ( .A(\Reg_Bank/registers[18][5] ), .B(
        \Reg_Bank/registers[19][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4182 ) );
  MUX \Reg_Bank/U4219  ( .A(\Reg_Bank/n4180 ), .B(\Reg_Bank/n4179 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4181 ) );
  MUX \Reg_Bank/U4218  ( .A(\Reg_Bank/registers[20][5] ), .B(
        \Reg_Bank/registers[21][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4180 ) );
  MUX \Reg_Bank/U4217  ( .A(\Reg_Bank/registers[22][5] ), .B(
        \Reg_Bank/registers[23][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4179 ) );
  MUX \Reg_Bank/U4216  ( .A(\Reg_Bank/n4177 ), .B(\Reg_Bank/n4174 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4178 ) );
  MUX \Reg_Bank/U4215  ( .A(\Reg_Bank/n4176 ), .B(\Reg_Bank/n4175 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4177 ) );
  MUX \Reg_Bank/U4214  ( .A(\Reg_Bank/registers[24][5] ), .B(
        \Reg_Bank/registers[25][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4176 ) );
  MUX \Reg_Bank/U4213  ( .A(\Reg_Bank/registers[26][5] ), .B(
        \Reg_Bank/registers[27][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4175 ) );
  MUX \Reg_Bank/U4212  ( .A(\Reg_Bank/n4173 ), .B(\Reg_Bank/n4172 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4174 ) );
  MUX \Reg_Bank/U4211  ( .A(\Reg_Bank/registers[28][5] ), .B(
        \Reg_Bank/registers[29][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4173 ) );
  MUX \Reg_Bank/U4210  ( .A(\Reg_Bank/registers[30][5] ), .B(
        \Reg_Bank/registers[31][5] ), .S(rs_index[0]), .Z(\Reg_Bank/n4172 ) );
  MUX \Reg_Bank/U4209  ( .A(\Reg_Bank/n4171 ), .B(\Reg_Bank/n4156 ), .S(
        rs_index[4]), .Z(reg_source[4]) );
  MUX \Reg_Bank/U4208  ( .A(\Reg_Bank/n4170 ), .B(\Reg_Bank/n4163 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4171 ) );
  MUX \Reg_Bank/U4207  ( .A(\Reg_Bank/n4169 ), .B(\Reg_Bank/n4166 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4170 ) );
  MUX \Reg_Bank/U4206  ( .A(\Reg_Bank/n4168 ), .B(\Reg_Bank/n4167 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4169 ) );
  MUX \Reg_Bank/U4204  ( .A(\Reg_Bank/registers[2][4] ), .B(
        \Reg_Bank/registers[3][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4167 ) );
  MUX \Reg_Bank/U4203  ( .A(\Reg_Bank/n4165 ), .B(\Reg_Bank/n4164 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4166 ) );
  MUX \Reg_Bank/U4202  ( .A(\Reg_Bank/registers[4][4] ), .B(
        \Reg_Bank/registers[5][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4165 ) );
  MUX \Reg_Bank/U4201  ( .A(\Reg_Bank/registers[6][4] ), .B(
        \Reg_Bank/registers[7][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4164 ) );
  MUX \Reg_Bank/U4200  ( .A(\Reg_Bank/n4162 ), .B(\Reg_Bank/n4159 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4163 ) );
  MUX \Reg_Bank/U4199  ( .A(\Reg_Bank/n4161 ), .B(\Reg_Bank/n4160 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4162 ) );
  MUX \Reg_Bank/U4198  ( .A(\Reg_Bank/registers[8][4] ), .B(
        \Reg_Bank/registers[9][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4161 ) );
  MUX \Reg_Bank/U4197  ( .A(\Reg_Bank/registers[10][4] ), .B(
        \Reg_Bank/registers[11][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4160 ) );
  MUX \Reg_Bank/U4196  ( .A(\Reg_Bank/n4158 ), .B(\Reg_Bank/n4157 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4159 ) );
  MUX \Reg_Bank/U4195  ( .A(\Reg_Bank/registers[12][4] ), .B(
        \Reg_Bank/registers[13][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4158 ) );
  MUX \Reg_Bank/U4194  ( .A(\Reg_Bank/registers[14][4] ), .B(
        \Reg_Bank/registers[15][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4157 ) );
  MUX \Reg_Bank/U4193  ( .A(\Reg_Bank/n4155 ), .B(\Reg_Bank/n4148 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4156 ) );
  MUX \Reg_Bank/U4192  ( .A(\Reg_Bank/n4154 ), .B(\Reg_Bank/n4151 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4155 ) );
  MUX \Reg_Bank/U4191  ( .A(\Reg_Bank/n4153 ), .B(\Reg_Bank/n4152 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4154 ) );
  MUX \Reg_Bank/U4190  ( .A(\Reg_Bank/registers[16][4] ), .B(
        \Reg_Bank/registers[17][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4153 ) );
  MUX \Reg_Bank/U4189  ( .A(\Reg_Bank/registers[18][4] ), .B(
        \Reg_Bank/registers[19][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4152 ) );
  MUX \Reg_Bank/U4188  ( .A(\Reg_Bank/n4150 ), .B(\Reg_Bank/n4149 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4151 ) );
  MUX \Reg_Bank/U4187  ( .A(\Reg_Bank/registers[20][4] ), .B(
        \Reg_Bank/registers[21][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4150 ) );
  MUX \Reg_Bank/U4186  ( .A(\Reg_Bank/registers[22][4] ), .B(
        \Reg_Bank/registers[23][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4149 ) );
  MUX \Reg_Bank/U4185  ( .A(\Reg_Bank/n4147 ), .B(\Reg_Bank/n4144 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4148 ) );
  MUX \Reg_Bank/U4184  ( .A(\Reg_Bank/n4146 ), .B(\Reg_Bank/n4145 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4147 ) );
  MUX \Reg_Bank/U4183  ( .A(\Reg_Bank/registers[24][4] ), .B(
        \Reg_Bank/registers[25][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4146 ) );
  MUX \Reg_Bank/U4182  ( .A(\Reg_Bank/registers[26][4] ), .B(
        \Reg_Bank/registers[27][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4145 ) );
  MUX \Reg_Bank/U4181  ( .A(\Reg_Bank/n4143 ), .B(\Reg_Bank/n4142 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4144 ) );
  MUX \Reg_Bank/U4180  ( .A(\Reg_Bank/registers[28][4] ), .B(
        \Reg_Bank/registers[29][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4143 ) );
  MUX \Reg_Bank/U4179  ( .A(\Reg_Bank/registers[30][4] ), .B(
        \Reg_Bank/registers[31][4] ), .S(rs_index[0]), .Z(\Reg_Bank/n4142 ) );
  MUX \Reg_Bank/U4178  ( .A(\Reg_Bank/n4141 ), .B(\Reg_Bank/n4126 ), .S(
        rs_index[4]), .Z(reg_source[3]) );
  MUX \Reg_Bank/U4177  ( .A(\Reg_Bank/n4140 ), .B(\Reg_Bank/n4133 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4141 ) );
  MUX \Reg_Bank/U4176  ( .A(\Reg_Bank/n4139 ), .B(\Reg_Bank/n4136 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4140 ) );
  MUX \Reg_Bank/U4175  ( .A(\Reg_Bank/n4138 ), .B(\Reg_Bank/n4137 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4139 ) );
  MUX \Reg_Bank/U4173  ( .A(\Reg_Bank/registers[2][3] ), .B(
        \Reg_Bank/registers[3][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4137 ) );
  MUX \Reg_Bank/U4172  ( .A(\Reg_Bank/n4135 ), .B(\Reg_Bank/n4134 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4136 ) );
  MUX \Reg_Bank/U4171  ( .A(\Reg_Bank/registers[4][3] ), .B(
        \Reg_Bank/registers[5][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4135 ) );
  MUX \Reg_Bank/U4170  ( .A(\Reg_Bank/registers[6][3] ), .B(
        \Reg_Bank/registers[7][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4134 ) );
  MUX \Reg_Bank/U4169  ( .A(\Reg_Bank/n4132 ), .B(\Reg_Bank/n4129 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4133 ) );
  MUX \Reg_Bank/U4168  ( .A(\Reg_Bank/n4131 ), .B(\Reg_Bank/n4130 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4132 ) );
  MUX \Reg_Bank/U4167  ( .A(\Reg_Bank/registers[8][3] ), .B(
        \Reg_Bank/registers[9][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4131 ) );
  MUX \Reg_Bank/U4166  ( .A(\Reg_Bank/registers[10][3] ), .B(
        \Reg_Bank/registers[11][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4130 ) );
  MUX \Reg_Bank/U4165  ( .A(\Reg_Bank/n4128 ), .B(\Reg_Bank/n4127 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4129 ) );
  MUX \Reg_Bank/U4164  ( .A(\Reg_Bank/registers[12][3] ), .B(
        \Reg_Bank/registers[13][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4128 ) );
  MUX \Reg_Bank/U4163  ( .A(\Reg_Bank/registers[14][3] ), .B(
        \Reg_Bank/registers[15][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4127 ) );
  MUX \Reg_Bank/U4162  ( .A(\Reg_Bank/n4125 ), .B(\Reg_Bank/n4118 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4126 ) );
  MUX \Reg_Bank/U4161  ( .A(\Reg_Bank/n4124 ), .B(\Reg_Bank/n4121 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4125 ) );
  MUX \Reg_Bank/U4160  ( .A(\Reg_Bank/n4123 ), .B(\Reg_Bank/n4122 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4124 ) );
  MUX \Reg_Bank/U4159  ( .A(\Reg_Bank/registers[16][3] ), .B(
        \Reg_Bank/registers[17][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4123 ) );
  MUX \Reg_Bank/U4158  ( .A(\Reg_Bank/registers[18][3] ), .B(
        \Reg_Bank/registers[19][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4122 ) );
  MUX \Reg_Bank/U4157  ( .A(\Reg_Bank/n4120 ), .B(\Reg_Bank/n4119 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4121 ) );
  MUX \Reg_Bank/U4156  ( .A(\Reg_Bank/registers[20][3] ), .B(
        \Reg_Bank/registers[21][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4120 ) );
  MUX \Reg_Bank/U4155  ( .A(\Reg_Bank/registers[22][3] ), .B(
        \Reg_Bank/registers[23][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4119 ) );
  MUX \Reg_Bank/U4154  ( .A(\Reg_Bank/n4117 ), .B(\Reg_Bank/n4114 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4118 ) );
  MUX \Reg_Bank/U4153  ( .A(\Reg_Bank/n4116 ), .B(\Reg_Bank/n4115 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4117 ) );
  MUX \Reg_Bank/U4152  ( .A(\Reg_Bank/registers[24][3] ), .B(
        \Reg_Bank/registers[25][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4116 ) );
  MUX \Reg_Bank/U4151  ( .A(\Reg_Bank/registers[26][3] ), .B(
        \Reg_Bank/registers[27][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4115 ) );
  MUX \Reg_Bank/U4150  ( .A(\Reg_Bank/n4113 ), .B(\Reg_Bank/n4112 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4114 ) );
  MUX \Reg_Bank/U4149  ( .A(\Reg_Bank/registers[28][3] ), .B(
        \Reg_Bank/registers[29][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4113 ) );
  MUX \Reg_Bank/U4148  ( .A(\Reg_Bank/registers[30][3] ), .B(
        \Reg_Bank/registers[31][3] ), .S(rs_index[0]), .Z(\Reg_Bank/n4112 ) );
  MUX \Reg_Bank/U4147  ( .A(\Reg_Bank/n4111 ), .B(\Reg_Bank/n4096 ), .S(
        rs_index[4]), .Z(reg_source[2]) );
  MUX \Reg_Bank/U4146  ( .A(\Reg_Bank/n4110 ), .B(\Reg_Bank/n4103 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4111 ) );
  MUX \Reg_Bank/U4145  ( .A(\Reg_Bank/n4109 ), .B(\Reg_Bank/n4106 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4110 ) );
  MUX \Reg_Bank/U4144  ( .A(\Reg_Bank/n4108 ), .B(\Reg_Bank/n4107 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4109 ) );
  MUX \Reg_Bank/U4142  ( .A(\Reg_Bank/registers[2][2] ), .B(
        \Reg_Bank/registers[3][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4107 ) );
  MUX \Reg_Bank/U4141  ( .A(\Reg_Bank/n4105 ), .B(\Reg_Bank/n4104 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4106 ) );
  MUX \Reg_Bank/U4140  ( .A(\Reg_Bank/registers[4][2] ), .B(
        \Reg_Bank/registers[5][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4105 ) );
  MUX \Reg_Bank/U4139  ( .A(\Reg_Bank/registers[6][2] ), .B(
        \Reg_Bank/registers[7][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4104 ) );
  MUX \Reg_Bank/U4138  ( .A(\Reg_Bank/n4102 ), .B(\Reg_Bank/n4099 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4103 ) );
  MUX \Reg_Bank/U4137  ( .A(\Reg_Bank/n4101 ), .B(\Reg_Bank/n4100 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4102 ) );
  MUX \Reg_Bank/U4136  ( .A(\Reg_Bank/registers[8][2] ), .B(
        \Reg_Bank/registers[9][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4101 ) );
  MUX \Reg_Bank/U4135  ( .A(\Reg_Bank/registers[10][2] ), .B(
        \Reg_Bank/registers[11][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4100 ) );
  MUX \Reg_Bank/U4134  ( .A(\Reg_Bank/n4098 ), .B(\Reg_Bank/n4097 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4099 ) );
  MUX \Reg_Bank/U4133  ( .A(\Reg_Bank/registers[12][2] ), .B(
        \Reg_Bank/registers[13][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4098 ) );
  MUX \Reg_Bank/U4132  ( .A(\Reg_Bank/registers[14][2] ), .B(
        \Reg_Bank/registers[15][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4097 ) );
  MUX \Reg_Bank/U4131  ( .A(\Reg_Bank/n4095 ), .B(\Reg_Bank/n4088 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4096 ) );
  MUX \Reg_Bank/U4130  ( .A(\Reg_Bank/n4094 ), .B(\Reg_Bank/n4091 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4095 ) );
  MUX \Reg_Bank/U4129  ( .A(\Reg_Bank/n4093 ), .B(\Reg_Bank/n4092 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4094 ) );
  MUX \Reg_Bank/U4128  ( .A(\Reg_Bank/registers[16][2] ), .B(
        \Reg_Bank/registers[17][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4093 ) );
  MUX \Reg_Bank/U4127  ( .A(\Reg_Bank/registers[18][2] ), .B(
        \Reg_Bank/registers[19][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4092 ) );
  MUX \Reg_Bank/U4126  ( .A(\Reg_Bank/n4090 ), .B(\Reg_Bank/n4089 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4091 ) );
  MUX \Reg_Bank/U4125  ( .A(\Reg_Bank/registers[20][2] ), .B(
        \Reg_Bank/registers[21][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4090 ) );
  MUX \Reg_Bank/U4124  ( .A(\Reg_Bank/registers[22][2] ), .B(
        \Reg_Bank/registers[23][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4089 ) );
  MUX \Reg_Bank/U4123  ( .A(\Reg_Bank/n4087 ), .B(\Reg_Bank/n4084 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4088 ) );
  MUX \Reg_Bank/U4122  ( .A(\Reg_Bank/n4086 ), .B(\Reg_Bank/n4085 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4087 ) );
  MUX \Reg_Bank/U4121  ( .A(\Reg_Bank/registers[24][2] ), .B(
        \Reg_Bank/registers[25][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4086 ) );
  MUX \Reg_Bank/U4120  ( .A(\Reg_Bank/registers[26][2] ), .B(
        \Reg_Bank/registers[27][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4085 ) );
  MUX \Reg_Bank/U4119  ( .A(\Reg_Bank/n4083 ), .B(\Reg_Bank/n4082 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4084 ) );
  MUX \Reg_Bank/U4118  ( .A(\Reg_Bank/registers[28][2] ), .B(
        \Reg_Bank/registers[29][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4083 ) );
  MUX \Reg_Bank/U4117  ( .A(\Reg_Bank/registers[30][2] ), .B(
        \Reg_Bank/registers[31][2] ), .S(rs_index[0]), .Z(\Reg_Bank/n4082 ) );
  MUX \Reg_Bank/U4116  ( .A(\Reg_Bank/n4081 ), .B(\Reg_Bank/n4066 ), .S(
        rs_index[4]), .Z(reg_source[1]) );
  MUX \Reg_Bank/U4115  ( .A(\Reg_Bank/n4080 ), .B(\Reg_Bank/n4073 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4081 ) );
  MUX \Reg_Bank/U4114  ( .A(\Reg_Bank/n4079 ), .B(\Reg_Bank/n4076 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4080 ) );
  MUX \Reg_Bank/U4113  ( .A(\Reg_Bank/n4078 ), .B(\Reg_Bank/n4077 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4079 ) );
  MUX \Reg_Bank/U4111  ( .A(\Reg_Bank/registers[2][1] ), .B(
        \Reg_Bank/registers[3][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4077 ) );
  MUX \Reg_Bank/U4110  ( .A(\Reg_Bank/n4075 ), .B(\Reg_Bank/n4074 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4076 ) );
  MUX \Reg_Bank/U4109  ( .A(\Reg_Bank/registers[4][1] ), .B(
        \Reg_Bank/registers[5][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4075 ) );
  MUX \Reg_Bank/U4108  ( .A(\Reg_Bank/registers[6][1] ), .B(
        \Reg_Bank/registers[7][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4074 ) );
  MUX \Reg_Bank/U4107  ( .A(\Reg_Bank/n4072 ), .B(\Reg_Bank/n4069 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4073 ) );
  MUX \Reg_Bank/U4106  ( .A(\Reg_Bank/n4071 ), .B(\Reg_Bank/n4070 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4072 ) );
  MUX \Reg_Bank/U4105  ( .A(\Reg_Bank/registers[8][1] ), .B(
        \Reg_Bank/registers[9][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4071 ) );
  MUX \Reg_Bank/U4104  ( .A(\Reg_Bank/registers[10][1] ), .B(
        \Reg_Bank/registers[11][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4070 ) );
  MUX \Reg_Bank/U4103  ( .A(\Reg_Bank/n4068 ), .B(\Reg_Bank/n4067 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4069 ) );
  MUX \Reg_Bank/U4102  ( .A(\Reg_Bank/registers[12][1] ), .B(
        \Reg_Bank/registers[13][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4068 ) );
  MUX \Reg_Bank/U4101  ( .A(\Reg_Bank/registers[14][1] ), .B(
        \Reg_Bank/registers[15][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4067 ) );
  MUX \Reg_Bank/U4100  ( .A(\Reg_Bank/n4065 ), .B(\Reg_Bank/n4058 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4066 ) );
  MUX \Reg_Bank/U4099  ( .A(\Reg_Bank/n4064 ), .B(\Reg_Bank/n4061 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4065 ) );
  MUX \Reg_Bank/U4098  ( .A(\Reg_Bank/n4063 ), .B(\Reg_Bank/n4062 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4064 ) );
  MUX \Reg_Bank/U4097  ( .A(\Reg_Bank/registers[16][1] ), .B(
        \Reg_Bank/registers[17][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4063 ) );
  MUX \Reg_Bank/U4096  ( .A(\Reg_Bank/registers[18][1] ), .B(
        \Reg_Bank/registers[19][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4062 ) );
  MUX \Reg_Bank/U4095  ( .A(\Reg_Bank/n4060 ), .B(\Reg_Bank/n4059 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4061 ) );
  MUX \Reg_Bank/U4094  ( .A(\Reg_Bank/registers[20][1] ), .B(
        \Reg_Bank/registers[21][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4060 ) );
  MUX \Reg_Bank/U4093  ( .A(\Reg_Bank/registers[22][1] ), .B(
        \Reg_Bank/registers[23][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4059 ) );
  MUX \Reg_Bank/U4092  ( .A(\Reg_Bank/n4057 ), .B(\Reg_Bank/n4054 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4058 ) );
  MUX \Reg_Bank/U4091  ( .A(\Reg_Bank/n4056 ), .B(\Reg_Bank/n4055 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4057 ) );
  MUX \Reg_Bank/U4090  ( .A(\Reg_Bank/registers[24][1] ), .B(
        \Reg_Bank/registers[25][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4056 ) );
  MUX \Reg_Bank/U4089  ( .A(\Reg_Bank/registers[26][1] ), .B(
        \Reg_Bank/registers[27][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4055 ) );
  MUX \Reg_Bank/U4088  ( .A(\Reg_Bank/n4053 ), .B(\Reg_Bank/n4052 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4054 ) );
  MUX \Reg_Bank/U4087  ( .A(\Reg_Bank/registers[28][1] ), .B(
        \Reg_Bank/registers[29][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4053 ) );
  MUX \Reg_Bank/U4086  ( .A(\Reg_Bank/registers[30][1] ), .B(
        \Reg_Bank/registers[31][1] ), .S(rs_index[0]), .Z(\Reg_Bank/n4052 ) );
  MUX \Reg_Bank/U4085  ( .A(\Reg_Bank/n4051 ), .B(\Reg_Bank/n4036 ), .S(
        rs_index[4]), .Z(reg_source[0]) );
  MUX \Reg_Bank/U4084  ( .A(\Reg_Bank/n4050 ), .B(\Reg_Bank/n4043 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4051 ) );
  MUX \Reg_Bank/U4083  ( .A(\Reg_Bank/n4049 ), .B(\Reg_Bank/n4046 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4050 ) );
  MUX \Reg_Bank/U4082  ( .A(\Reg_Bank/n4048 ), .B(\Reg_Bank/n4047 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4049 ) );
  MUX \Reg_Bank/U4080  ( .A(\Reg_Bank/registers[2][0] ), .B(
        \Reg_Bank/registers[3][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4047 ) );
  MUX \Reg_Bank/U4079  ( .A(\Reg_Bank/n4045 ), .B(\Reg_Bank/n4044 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4046 ) );
  MUX \Reg_Bank/U4078  ( .A(\Reg_Bank/registers[4][0] ), .B(
        \Reg_Bank/registers[5][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4045 ) );
  MUX \Reg_Bank/U4077  ( .A(\Reg_Bank/registers[6][0] ), .B(
        \Reg_Bank/registers[7][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4044 ) );
  MUX \Reg_Bank/U4076  ( .A(\Reg_Bank/n4042 ), .B(\Reg_Bank/n4039 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4043 ) );
  MUX \Reg_Bank/U4075  ( .A(\Reg_Bank/n4041 ), .B(\Reg_Bank/n4040 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4042 ) );
  MUX \Reg_Bank/U4074  ( .A(\Reg_Bank/registers[8][0] ), .B(
        \Reg_Bank/registers[9][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4041 ) );
  MUX \Reg_Bank/U4073  ( .A(\Reg_Bank/registers[10][0] ), .B(
        \Reg_Bank/registers[11][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4040 ) );
  MUX \Reg_Bank/U4072  ( .A(\Reg_Bank/n4038 ), .B(\Reg_Bank/n4037 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4039 ) );
  MUX \Reg_Bank/U4071  ( .A(\Reg_Bank/registers[12][0] ), .B(
        \Reg_Bank/registers[13][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4038 ) );
  MUX \Reg_Bank/U4070  ( .A(\Reg_Bank/registers[14][0] ), .B(
        \Reg_Bank/registers[15][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4037 ) );
  MUX \Reg_Bank/U4069  ( .A(\Reg_Bank/n4035 ), .B(\Reg_Bank/n4028 ), .S(
        rs_index[3]), .Z(\Reg_Bank/n4036 ) );
  MUX \Reg_Bank/U4068  ( .A(\Reg_Bank/n4034 ), .B(\Reg_Bank/n4031 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4035 ) );
  MUX \Reg_Bank/U4067  ( .A(\Reg_Bank/n4033 ), .B(\Reg_Bank/n4032 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4034 ) );
  MUX \Reg_Bank/U4066  ( .A(\Reg_Bank/registers[16][0] ), .B(
        \Reg_Bank/registers[17][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4033 ) );
  MUX \Reg_Bank/U4065  ( .A(\Reg_Bank/registers[18][0] ), .B(
        \Reg_Bank/registers[19][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4032 ) );
  MUX \Reg_Bank/U4064  ( .A(\Reg_Bank/n4030 ), .B(\Reg_Bank/n4029 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4031 ) );
  MUX \Reg_Bank/U4063  ( .A(\Reg_Bank/registers[20][0] ), .B(
        \Reg_Bank/registers[21][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4030 ) );
  MUX \Reg_Bank/U4062  ( .A(\Reg_Bank/registers[22][0] ), .B(
        \Reg_Bank/registers[23][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4029 ) );
  MUX \Reg_Bank/U4061  ( .A(\Reg_Bank/n4027 ), .B(\Reg_Bank/n4024 ), .S(
        rs_index[2]), .Z(\Reg_Bank/n4028 ) );
  MUX \Reg_Bank/U4060  ( .A(\Reg_Bank/n4026 ), .B(\Reg_Bank/n4025 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4027 ) );
  MUX \Reg_Bank/U4059  ( .A(\Reg_Bank/registers[24][0] ), .B(
        \Reg_Bank/registers[25][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4026 ) );
  MUX \Reg_Bank/U4058  ( .A(\Reg_Bank/registers[26][0] ), .B(
        \Reg_Bank/registers[27][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4025 ) );
  MUX \Reg_Bank/U4057  ( .A(\Reg_Bank/n4023 ), .B(\Reg_Bank/n4022 ), .S(
        rs_index[1]), .Z(\Reg_Bank/n4024 ) );
  MUX \Reg_Bank/U4056  ( .A(\Reg_Bank/registers[28][0] ), .B(
        \Reg_Bank/registers[29][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4023 ) );
  MUX \Reg_Bank/U4055  ( .A(\Reg_Bank/registers[30][0] ), .B(
        \Reg_Bank/registers[31][0] ), .S(rs_index[0]), .Z(\Reg_Bank/n4022 ) );
  DFF \Reg_Bank/registers_reg[1][0]  ( .D(\Reg_Bank/n3030 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][0] ) );
  DFF \Reg_Bank/registers_reg[1][1]  ( .D(\Reg_Bank/n3031 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][1] ) );
  DFF \Reg_Bank/registers_reg[1][2]  ( .D(\Reg_Bank/n3032 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][2] ) );
  DFF \Reg_Bank/registers_reg[1][3]  ( .D(\Reg_Bank/n3033 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][3] ) );
  DFF \Reg_Bank/registers_reg[1][4]  ( .D(\Reg_Bank/n3034 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][4] ) );
  DFF \Reg_Bank/registers_reg[1][5]  ( .D(\Reg_Bank/n3035 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][5] ) );
  DFF \Reg_Bank/registers_reg[1][6]  ( .D(\Reg_Bank/n3036 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][6] ) );
  DFF \Reg_Bank/registers_reg[1][7]  ( .D(\Reg_Bank/n3037 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][7] ) );
  DFF \Reg_Bank/registers_reg[1][8]  ( .D(\Reg_Bank/n3038 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][8] ) );
  DFF \Reg_Bank/registers_reg[1][9]  ( .D(\Reg_Bank/n3039 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][9] ) );
  DFF \Reg_Bank/registers_reg[1][10]  ( .D(\Reg_Bank/n3040 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][10] ) );
  DFF \Reg_Bank/registers_reg[1][11]  ( .D(\Reg_Bank/n3041 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][11] ) );
  DFF \Reg_Bank/registers_reg[1][12]  ( .D(\Reg_Bank/n3042 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][12] ) );
  DFF \Reg_Bank/registers_reg[1][13]  ( .D(\Reg_Bank/n3043 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][13] ) );
  DFF \Reg_Bank/registers_reg[1][14]  ( .D(\Reg_Bank/n3044 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][14] ) );
  DFF \Reg_Bank/registers_reg[1][15]  ( .D(\Reg_Bank/n3045 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][15] ) );
  DFF \Reg_Bank/registers_reg[1][16]  ( .D(\Reg_Bank/n3046 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][16] ) );
  DFF \Reg_Bank/registers_reg[1][17]  ( .D(\Reg_Bank/n3047 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][17] ) );
  DFF \Reg_Bank/registers_reg[1][18]  ( .D(\Reg_Bank/n3048 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][18] ) );
  DFF \Reg_Bank/registers_reg[1][19]  ( .D(\Reg_Bank/n3049 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][19] ) );
  DFF \Reg_Bank/registers_reg[1][20]  ( .D(\Reg_Bank/n3050 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][20] ) );
  DFF \Reg_Bank/registers_reg[1][21]  ( .D(\Reg_Bank/n3051 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][21] ) );
  DFF \Reg_Bank/registers_reg[1][22]  ( .D(\Reg_Bank/n3052 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][22] ) );
  DFF \Reg_Bank/registers_reg[1][23]  ( .D(\Reg_Bank/n3053 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][23] ) );
  DFF \Reg_Bank/registers_reg[1][24]  ( .D(\Reg_Bank/n3054 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][24] ) );
  DFF \Reg_Bank/registers_reg[1][25]  ( .D(\Reg_Bank/n3055 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][25] ) );
  DFF \Reg_Bank/registers_reg[1][26]  ( .D(\Reg_Bank/n3056 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][26] ) );
  DFF \Reg_Bank/registers_reg[1][27]  ( .D(\Reg_Bank/n3057 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][27] ) );
  DFF \Reg_Bank/registers_reg[1][28]  ( .D(\Reg_Bank/n3058 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][28] ) );
  DFF \Reg_Bank/registers_reg[1][29]  ( .D(\Reg_Bank/n3059 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][29] ) );
  DFF \Reg_Bank/registers_reg[1][30]  ( .D(\Reg_Bank/n3060 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][30] ) );
  DFF \Reg_Bank/registers_reg[1][31]  ( .D(\Reg_Bank/n3061 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][31] ) );
  DFF \Reg_Bank/registers_reg[2][0]  ( .D(\Reg_Bank/n3062 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][0] ) );
  DFF \Reg_Bank/registers_reg[2][1]  ( .D(\Reg_Bank/n3063 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][1] ) );
  DFF \Reg_Bank/registers_reg[2][2]  ( .D(\Reg_Bank/n3064 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][2] ) );
  DFF \Reg_Bank/registers_reg[2][3]  ( .D(\Reg_Bank/n3065 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][3] ) );
  DFF \Reg_Bank/registers_reg[2][4]  ( .D(\Reg_Bank/n3066 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][4] ) );
  DFF \Reg_Bank/registers_reg[2][5]  ( .D(\Reg_Bank/n3067 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][5] ) );
  DFF \Reg_Bank/registers_reg[2][6]  ( .D(\Reg_Bank/n3068 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][6] ) );
  DFF \Reg_Bank/registers_reg[2][7]  ( .D(\Reg_Bank/n3069 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][7] ) );
  DFF \Reg_Bank/registers_reg[2][8]  ( .D(\Reg_Bank/n3070 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][8] ) );
  DFF \Reg_Bank/registers_reg[2][9]  ( .D(\Reg_Bank/n3071 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][9] ) );
  DFF \Reg_Bank/registers_reg[2][10]  ( .D(\Reg_Bank/n3072 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][10] ) );
  DFF \Reg_Bank/registers_reg[2][11]  ( .D(\Reg_Bank/n3073 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][11] ) );
  DFF \Reg_Bank/registers_reg[2][12]  ( .D(\Reg_Bank/n3074 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][12] ) );
  DFF \Reg_Bank/registers_reg[2][13]  ( .D(\Reg_Bank/n3075 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][13] ) );
  DFF \Reg_Bank/registers_reg[2][14]  ( .D(\Reg_Bank/n3076 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][14] ) );
  DFF \Reg_Bank/registers_reg[2][15]  ( .D(\Reg_Bank/n3077 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][15] ) );
  DFF \Reg_Bank/registers_reg[2][16]  ( .D(\Reg_Bank/n3078 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][16] ) );
  DFF \Reg_Bank/registers_reg[2][17]  ( .D(\Reg_Bank/n3079 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][17] ) );
  DFF \Reg_Bank/registers_reg[2][18]  ( .D(\Reg_Bank/n3080 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][18] ) );
  DFF \Reg_Bank/registers_reg[2][19]  ( .D(\Reg_Bank/n3081 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][19] ) );
  DFF \Reg_Bank/registers_reg[2][20]  ( .D(\Reg_Bank/n3082 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][20] ) );
  DFF \Reg_Bank/registers_reg[2][21]  ( .D(\Reg_Bank/n3083 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][21] ) );
  DFF \Reg_Bank/registers_reg[2][22]  ( .D(\Reg_Bank/n3084 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][22] ) );
  DFF \Reg_Bank/registers_reg[2][23]  ( .D(\Reg_Bank/n3085 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][23] ) );
  DFF \Reg_Bank/registers_reg[2][24]  ( .D(\Reg_Bank/n3086 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][24] ) );
  DFF \Reg_Bank/registers_reg[2][25]  ( .D(\Reg_Bank/n3087 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][25] ) );
  DFF \Reg_Bank/registers_reg[2][26]  ( .D(\Reg_Bank/n3088 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][26] ) );
  DFF \Reg_Bank/registers_reg[2][27]  ( .D(\Reg_Bank/n3089 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][27] ) );
  DFF \Reg_Bank/registers_reg[2][28]  ( .D(\Reg_Bank/n3090 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][28] ) );
  DFF \Reg_Bank/registers_reg[2][29]  ( .D(\Reg_Bank/n3091 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][29] ) );
  DFF \Reg_Bank/registers_reg[2][30]  ( .D(\Reg_Bank/n3092 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][30] ) );
  DFF \Reg_Bank/registers_reg[2][31]  ( .D(\Reg_Bank/n3093 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][31] ) );
  DFF \Reg_Bank/registers_reg[3][0]  ( .D(\Reg_Bank/n3094 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][0] ) );
  DFF \Reg_Bank/registers_reg[3][1]  ( .D(\Reg_Bank/n3095 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][1] ) );
  DFF \Reg_Bank/registers_reg[3][2]  ( .D(\Reg_Bank/n3096 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][2] ) );
  DFF \Reg_Bank/registers_reg[3][3]  ( .D(\Reg_Bank/n3097 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][3] ) );
  DFF \Reg_Bank/registers_reg[3][4]  ( .D(\Reg_Bank/n3098 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][4] ) );
  DFF \Reg_Bank/registers_reg[3][5]  ( .D(\Reg_Bank/n3099 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][5] ) );
  DFF \Reg_Bank/registers_reg[3][6]  ( .D(\Reg_Bank/n3100 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][6] ) );
  DFF \Reg_Bank/registers_reg[3][7]  ( .D(\Reg_Bank/n3101 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][7] ) );
  DFF \Reg_Bank/registers_reg[3][8]  ( .D(\Reg_Bank/n3102 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][8] ) );
  DFF \Reg_Bank/registers_reg[3][9]  ( .D(\Reg_Bank/n3103 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][9] ) );
  DFF \Reg_Bank/registers_reg[3][10]  ( .D(\Reg_Bank/n3104 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][10] ) );
  DFF \Reg_Bank/registers_reg[3][11]  ( .D(\Reg_Bank/n3105 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][11] ) );
  DFF \Reg_Bank/registers_reg[3][12]  ( .D(\Reg_Bank/n3106 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][12] ) );
  DFF \Reg_Bank/registers_reg[3][13]  ( .D(\Reg_Bank/n3107 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][13] ) );
  DFF \Reg_Bank/registers_reg[3][14]  ( .D(\Reg_Bank/n3108 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][14] ) );
  DFF \Reg_Bank/registers_reg[3][15]  ( .D(\Reg_Bank/n3109 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][15] ) );
  DFF \Reg_Bank/registers_reg[3][16]  ( .D(\Reg_Bank/n3110 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][16] ) );
  DFF \Reg_Bank/registers_reg[3][17]  ( .D(\Reg_Bank/n3111 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][17] ) );
  DFF \Reg_Bank/registers_reg[3][18]  ( .D(\Reg_Bank/n3112 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][18] ) );
  DFF \Reg_Bank/registers_reg[3][19]  ( .D(\Reg_Bank/n3113 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][19] ) );
  DFF \Reg_Bank/registers_reg[3][20]  ( .D(\Reg_Bank/n3114 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][20] ) );
  DFF \Reg_Bank/registers_reg[3][21]  ( .D(\Reg_Bank/n3115 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][21] ) );
  DFF \Reg_Bank/registers_reg[3][22]  ( .D(\Reg_Bank/n3116 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][22] ) );
  DFF \Reg_Bank/registers_reg[3][23]  ( .D(\Reg_Bank/n3117 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][23] ) );
  DFF \Reg_Bank/registers_reg[3][24]  ( .D(\Reg_Bank/n3118 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][24] ) );
  DFF \Reg_Bank/registers_reg[3][25]  ( .D(\Reg_Bank/n3119 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][25] ) );
  DFF \Reg_Bank/registers_reg[3][26]  ( .D(\Reg_Bank/n3120 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][26] ) );
  DFF \Reg_Bank/registers_reg[3][27]  ( .D(\Reg_Bank/n3121 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][27] ) );
  DFF \Reg_Bank/registers_reg[3][28]  ( .D(\Reg_Bank/n3122 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][28] ) );
  DFF \Reg_Bank/registers_reg[3][29]  ( .D(\Reg_Bank/n3123 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][29] ) );
  DFF \Reg_Bank/registers_reg[3][30]  ( .D(\Reg_Bank/n3124 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][30] ) );
  DFF \Reg_Bank/registers_reg[3][31]  ( .D(\Reg_Bank/n3125 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][31] ) );
  DFF \Reg_Bank/registers_reg[4][0]  ( .D(\Reg_Bank/n3126 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][0] ) );
  DFF \Reg_Bank/registers_reg[4][1]  ( .D(\Reg_Bank/n3127 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][1] ) );
  DFF \Reg_Bank/registers_reg[4][2]  ( .D(\Reg_Bank/n3128 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][2] ) );
  DFF \Reg_Bank/registers_reg[4][3]  ( .D(\Reg_Bank/n3129 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][3] ) );
  DFF \Reg_Bank/registers_reg[4][4]  ( .D(\Reg_Bank/n3130 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][4] ) );
  DFF \Reg_Bank/registers_reg[4][5]  ( .D(\Reg_Bank/n3131 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][5] ) );
  DFF \Reg_Bank/registers_reg[4][6]  ( .D(\Reg_Bank/n3132 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][6] ) );
  DFF \Reg_Bank/registers_reg[4][7]  ( .D(\Reg_Bank/n3133 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][7] ) );
  DFF \Reg_Bank/registers_reg[4][8]  ( .D(\Reg_Bank/n3134 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][8] ) );
  DFF \Reg_Bank/registers_reg[4][9]  ( .D(\Reg_Bank/n3135 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][9] ) );
  DFF \Reg_Bank/registers_reg[4][10]  ( .D(\Reg_Bank/n3136 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][10] ) );
  DFF \Reg_Bank/registers_reg[4][11]  ( .D(\Reg_Bank/n3137 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][11] ) );
  DFF \Reg_Bank/registers_reg[4][12]  ( .D(\Reg_Bank/n3138 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][12] ) );
  DFF \Reg_Bank/registers_reg[4][13]  ( .D(\Reg_Bank/n3139 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][13] ) );
  DFF \Reg_Bank/registers_reg[4][14]  ( .D(\Reg_Bank/n3140 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][14] ) );
  DFF \Reg_Bank/registers_reg[4][15]  ( .D(\Reg_Bank/n3141 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][15] ) );
  DFF \Reg_Bank/registers_reg[4][16]  ( .D(\Reg_Bank/n3142 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][16] ) );
  DFF \Reg_Bank/registers_reg[4][17]  ( .D(\Reg_Bank/n3143 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][17] ) );
  DFF \Reg_Bank/registers_reg[4][18]  ( .D(\Reg_Bank/n3144 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][18] ) );
  DFF \Reg_Bank/registers_reg[4][19]  ( .D(\Reg_Bank/n3145 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][19] ) );
  DFF \Reg_Bank/registers_reg[4][20]  ( .D(\Reg_Bank/n3146 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][20] ) );
  DFF \Reg_Bank/registers_reg[4][21]  ( .D(\Reg_Bank/n3147 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][21] ) );
  DFF \Reg_Bank/registers_reg[4][22]  ( .D(\Reg_Bank/n3148 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][22] ) );
  DFF \Reg_Bank/registers_reg[4][23]  ( .D(\Reg_Bank/n3149 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][23] ) );
  DFF \Reg_Bank/registers_reg[4][24]  ( .D(\Reg_Bank/n3150 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][24] ) );
  DFF \Reg_Bank/registers_reg[4][25]  ( .D(\Reg_Bank/n3151 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][25] ) );
  DFF \Reg_Bank/registers_reg[4][26]  ( .D(\Reg_Bank/n3152 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][26] ) );
  DFF \Reg_Bank/registers_reg[4][27]  ( .D(\Reg_Bank/n3153 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][27] ) );
  DFF \Reg_Bank/registers_reg[4][28]  ( .D(\Reg_Bank/n3154 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][28] ) );
  DFF \Reg_Bank/registers_reg[4][29]  ( .D(\Reg_Bank/n3155 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][29] ) );
  DFF \Reg_Bank/registers_reg[4][30]  ( .D(\Reg_Bank/n3156 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][30] ) );
  DFF \Reg_Bank/registers_reg[4][31]  ( .D(\Reg_Bank/n3157 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][31] ) );
  DFF \Reg_Bank/registers_reg[5][0]  ( .D(\Reg_Bank/n3158 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][0] ) );
  DFF \Reg_Bank/registers_reg[5][1]  ( .D(\Reg_Bank/n3159 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][1] ) );
  DFF \Reg_Bank/registers_reg[5][2]  ( .D(\Reg_Bank/n3160 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][2] ) );
  DFF \Reg_Bank/registers_reg[5][3]  ( .D(\Reg_Bank/n3161 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][3] ) );
  DFF \Reg_Bank/registers_reg[5][4]  ( .D(\Reg_Bank/n3162 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][4] ) );
  DFF \Reg_Bank/registers_reg[5][5]  ( .D(\Reg_Bank/n3163 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][5] ) );
  DFF \Reg_Bank/registers_reg[5][6]  ( .D(\Reg_Bank/n3164 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][6] ) );
  DFF \Reg_Bank/registers_reg[5][7]  ( .D(\Reg_Bank/n3165 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][7] ) );
  DFF \Reg_Bank/registers_reg[5][8]  ( .D(\Reg_Bank/n3166 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][8] ) );
  DFF \Reg_Bank/registers_reg[5][9]  ( .D(\Reg_Bank/n3167 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][9] ) );
  DFF \Reg_Bank/registers_reg[5][10]  ( .D(\Reg_Bank/n3168 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][10] ) );
  DFF \Reg_Bank/registers_reg[5][11]  ( .D(\Reg_Bank/n3169 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][11] ) );
  DFF \Reg_Bank/registers_reg[5][12]  ( .D(\Reg_Bank/n3170 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][12] ) );
  DFF \Reg_Bank/registers_reg[5][13]  ( .D(\Reg_Bank/n3171 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][13] ) );
  DFF \Reg_Bank/registers_reg[5][14]  ( .D(\Reg_Bank/n3172 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][14] ) );
  DFF \Reg_Bank/registers_reg[5][15]  ( .D(\Reg_Bank/n3173 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][15] ) );
  DFF \Reg_Bank/registers_reg[5][16]  ( .D(\Reg_Bank/n3174 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][16] ) );
  DFF \Reg_Bank/registers_reg[5][17]  ( .D(\Reg_Bank/n3175 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][17] ) );
  DFF \Reg_Bank/registers_reg[5][18]  ( .D(\Reg_Bank/n3176 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][18] ) );
  DFF \Reg_Bank/registers_reg[5][19]  ( .D(\Reg_Bank/n3177 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][19] ) );
  DFF \Reg_Bank/registers_reg[5][20]  ( .D(\Reg_Bank/n3178 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][20] ) );
  DFF \Reg_Bank/registers_reg[5][21]  ( .D(\Reg_Bank/n3179 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][21] ) );
  DFF \Reg_Bank/registers_reg[5][22]  ( .D(\Reg_Bank/n3180 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][22] ) );
  DFF \Reg_Bank/registers_reg[5][23]  ( .D(\Reg_Bank/n3181 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][23] ) );
  DFF \Reg_Bank/registers_reg[5][24]  ( .D(\Reg_Bank/n3182 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][24] ) );
  DFF \Reg_Bank/registers_reg[5][25]  ( .D(\Reg_Bank/n3183 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][25] ) );
  DFF \Reg_Bank/registers_reg[5][26]  ( .D(\Reg_Bank/n3184 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][26] ) );
  DFF \Reg_Bank/registers_reg[5][27]  ( .D(\Reg_Bank/n3185 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][27] ) );
  DFF \Reg_Bank/registers_reg[5][28]  ( .D(\Reg_Bank/n3186 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][28] ) );
  DFF \Reg_Bank/registers_reg[5][29]  ( .D(\Reg_Bank/n3187 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][29] ) );
  DFF \Reg_Bank/registers_reg[5][30]  ( .D(\Reg_Bank/n3188 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][30] ) );
  DFF \Reg_Bank/registers_reg[5][31]  ( .D(\Reg_Bank/n3189 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][31] ) );
  DFF \Reg_Bank/registers_reg[6][0]  ( .D(\Reg_Bank/n3190 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][0] ) );
  DFF \Reg_Bank/registers_reg[6][1]  ( .D(\Reg_Bank/n3191 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][1] ) );
  DFF \Reg_Bank/registers_reg[6][2]  ( .D(\Reg_Bank/n3192 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][2] ) );
  DFF \Reg_Bank/registers_reg[6][3]  ( .D(\Reg_Bank/n3193 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][3] ) );
  DFF \Reg_Bank/registers_reg[6][4]  ( .D(\Reg_Bank/n3194 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][4] ) );
  DFF \Reg_Bank/registers_reg[6][5]  ( .D(\Reg_Bank/n3195 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][5] ) );
  DFF \Reg_Bank/registers_reg[6][6]  ( .D(\Reg_Bank/n3196 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][6] ) );
  DFF \Reg_Bank/registers_reg[6][7]  ( .D(\Reg_Bank/n3197 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][7] ) );
  DFF \Reg_Bank/registers_reg[6][8]  ( .D(\Reg_Bank/n3198 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][8] ) );
  DFF \Reg_Bank/registers_reg[6][9]  ( .D(\Reg_Bank/n3199 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][9] ) );
  DFF \Reg_Bank/registers_reg[6][10]  ( .D(\Reg_Bank/n3200 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][10] ) );
  DFF \Reg_Bank/registers_reg[6][11]  ( .D(\Reg_Bank/n3201 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][11] ) );
  DFF \Reg_Bank/registers_reg[6][12]  ( .D(\Reg_Bank/n3202 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][12] ) );
  DFF \Reg_Bank/registers_reg[6][13]  ( .D(\Reg_Bank/n3203 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][13] ) );
  DFF \Reg_Bank/registers_reg[6][14]  ( .D(\Reg_Bank/n3204 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][14] ) );
  DFF \Reg_Bank/registers_reg[6][15]  ( .D(\Reg_Bank/n3205 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][15] ) );
  DFF \Reg_Bank/registers_reg[6][16]  ( .D(\Reg_Bank/n3206 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][16] ) );
  DFF \Reg_Bank/registers_reg[6][17]  ( .D(\Reg_Bank/n3207 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][17] ) );
  DFF \Reg_Bank/registers_reg[6][18]  ( .D(\Reg_Bank/n3208 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][18] ) );
  DFF \Reg_Bank/registers_reg[6][19]  ( .D(\Reg_Bank/n3209 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][19] ) );
  DFF \Reg_Bank/registers_reg[6][20]  ( .D(\Reg_Bank/n3210 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][20] ) );
  DFF \Reg_Bank/registers_reg[6][21]  ( .D(\Reg_Bank/n3211 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][21] ) );
  DFF \Reg_Bank/registers_reg[6][22]  ( .D(\Reg_Bank/n3212 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][22] ) );
  DFF \Reg_Bank/registers_reg[6][23]  ( .D(\Reg_Bank/n3213 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][23] ) );
  DFF \Reg_Bank/registers_reg[6][24]  ( .D(\Reg_Bank/n3214 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][24] ) );
  DFF \Reg_Bank/registers_reg[6][25]  ( .D(\Reg_Bank/n3215 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][25] ) );
  DFF \Reg_Bank/registers_reg[6][26]  ( .D(\Reg_Bank/n3216 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][26] ) );
  DFF \Reg_Bank/registers_reg[6][27]  ( .D(\Reg_Bank/n3217 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][27] ) );
  DFF \Reg_Bank/registers_reg[6][28]  ( .D(\Reg_Bank/n3218 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][28] ) );
  DFF \Reg_Bank/registers_reg[6][29]  ( .D(\Reg_Bank/n3219 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][29] ) );
  DFF \Reg_Bank/registers_reg[6][30]  ( .D(\Reg_Bank/n3220 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][30] ) );
  DFF \Reg_Bank/registers_reg[6][31]  ( .D(\Reg_Bank/n3221 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][31] ) );
  DFF \Reg_Bank/registers_reg[7][0]  ( .D(\Reg_Bank/n3222 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][0] ) );
  DFF \Reg_Bank/registers_reg[7][1]  ( .D(\Reg_Bank/n3223 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][1] ) );
  DFF \Reg_Bank/registers_reg[7][2]  ( .D(\Reg_Bank/n3224 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][2] ) );
  DFF \Reg_Bank/registers_reg[7][3]  ( .D(\Reg_Bank/n3225 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][3] ) );
  DFF \Reg_Bank/registers_reg[7][4]  ( .D(\Reg_Bank/n3226 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][4] ) );
  DFF \Reg_Bank/registers_reg[7][5]  ( .D(\Reg_Bank/n3227 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][5] ) );
  DFF \Reg_Bank/registers_reg[7][6]  ( .D(\Reg_Bank/n3228 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][6] ) );
  DFF \Reg_Bank/registers_reg[7][7]  ( .D(\Reg_Bank/n3229 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][7] ) );
  DFF \Reg_Bank/registers_reg[7][8]  ( .D(\Reg_Bank/n3230 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][8] ) );
  DFF \Reg_Bank/registers_reg[7][9]  ( .D(\Reg_Bank/n3231 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][9] ) );
  DFF \Reg_Bank/registers_reg[7][10]  ( .D(\Reg_Bank/n3232 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][10] ) );
  DFF \Reg_Bank/registers_reg[7][11]  ( .D(\Reg_Bank/n3233 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][11] ) );
  DFF \Reg_Bank/registers_reg[7][12]  ( .D(\Reg_Bank/n3234 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][12] ) );
  DFF \Reg_Bank/registers_reg[7][13]  ( .D(\Reg_Bank/n3235 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][13] ) );
  DFF \Reg_Bank/registers_reg[7][14]  ( .D(\Reg_Bank/n3236 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][14] ) );
  DFF \Reg_Bank/registers_reg[7][15]  ( .D(\Reg_Bank/n3237 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][15] ) );
  DFF \Reg_Bank/registers_reg[7][16]  ( .D(\Reg_Bank/n3238 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][16] ) );
  DFF \Reg_Bank/registers_reg[7][17]  ( .D(\Reg_Bank/n3239 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][17] ) );
  DFF \Reg_Bank/registers_reg[7][18]  ( .D(\Reg_Bank/n3240 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][18] ) );
  DFF \Reg_Bank/registers_reg[7][19]  ( .D(\Reg_Bank/n3241 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][19] ) );
  DFF \Reg_Bank/registers_reg[7][20]  ( .D(\Reg_Bank/n3242 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][20] ) );
  DFF \Reg_Bank/registers_reg[7][21]  ( .D(\Reg_Bank/n3243 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][21] ) );
  DFF \Reg_Bank/registers_reg[7][22]  ( .D(\Reg_Bank/n3244 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][22] ) );
  DFF \Reg_Bank/registers_reg[7][23]  ( .D(\Reg_Bank/n3245 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][23] ) );
  DFF \Reg_Bank/registers_reg[7][24]  ( .D(\Reg_Bank/n3246 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][24] ) );
  DFF \Reg_Bank/registers_reg[7][25]  ( .D(\Reg_Bank/n3247 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][25] ) );
  DFF \Reg_Bank/registers_reg[7][26]  ( .D(\Reg_Bank/n3248 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][26] ) );
  DFF \Reg_Bank/registers_reg[7][27]  ( .D(\Reg_Bank/n3249 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][27] ) );
  DFF \Reg_Bank/registers_reg[7][28]  ( .D(\Reg_Bank/n3250 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][28] ) );
  DFF \Reg_Bank/registers_reg[7][29]  ( .D(\Reg_Bank/n3251 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][29] ) );
  DFF \Reg_Bank/registers_reg[7][30]  ( .D(\Reg_Bank/n3252 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][30] ) );
  DFF \Reg_Bank/registers_reg[7][31]  ( .D(\Reg_Bank/n3253 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][31] ) );
  DFF \Reg_Bank/registers_reg[8][0]  ( .D(\Reg_Bank/n3254 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][0] ) );
  DFF \Reg_Bank/registers_reg[8][1]  ( .D(\Reg_Bank/n3255 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][1] ) );
  DFF \Reg_Bank/registers_reg[8][2]  ( .D(\Reg_Bank/n3256 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][2] ) );
  DFF \Reg_Bank/registers_reg[8][3]  ( .D(\Reg_Bank/n3257 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][3] ) );
  DFF \Reg_Bank/registers_reg[8][4]  ( .D(\Reg_Bank/n3258 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][4] ) );
  DFF \Reg_Bank/registers_reg[8][5]  ( .D(\Reg_Bank/n3259 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][5] ) );
  DFF \Reg_Bank/registers_reg[8][6]  ( .D(\Reg_Bank/n3260 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][6] ) );
  DFF \Reg_Bank/registers_reg[8][7]  ( .D(\Reg_Bank/n3261 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][7] ) );
  DFF \Reg_Bank/registers_reg[8][8]  ( .D(\Reg_Bank/n3262 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][8] ) );
  DFF \Reg_Bank/registers_reg[8][9]  ( .D(\Reg_Bank/n3263 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][9] ) );
  DFF \Reg_Bank/registers_reg[8][10]  ( .D(\Reg_Bank/n3264 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][10] ) );
  DFF \Reg_Bank/registers_reg[8][11]  ( .D(\Reg_Bank/n3265 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][11] ) );
  DFF \Reg_Bank/registers_reg[8][12]  ( .D(\Reg_Bank/n3266 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][12] ) );
  DFF \Reg_Bank/registers_reg[8][13]  ( .D(\Reg_Bank/n3267 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][13] ) );
  DFF \Reg_Bank/registers_reg[8][14]  ( .D(\Reg_Bank/n3268 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][14] ) );
  DFF \Reg_Bank/registers_reg[8][15]  ( .D(\Reg_Bank/n3269 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][15] ) );
  DFF \Reg_Bank/registers_reg[8][16]  ( .D(\Reg_Bank/n3270 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][16] ) );
  DFF \Reg_Bank/registers_reg[8][17]  ( .D(\Reg_Bank/n3271 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][17] ) );
  DFF \Reg_Bank/registers_reg[8][18]  ( .D(\Reg_Bank/n3272 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][18] ) );
  DFF \Reg_Bank/registers_reg[8][19]  ( .D(\Reg_Bank/n3273 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][19] ) );
  DFF \Reg_Bank/registers_reg[8][20]  ( .D(\Reg_Bank/n3274 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][20] ) );
  DFF \Reg_Bank/registers_reg[8][21]  ( .D(\Reg_Bank/n3275 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][21] ) );
  DFF \Reg_Bank/registers_reg[8][22]  ( .D(\Reg_Bank/n3276 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][22] ) );
  DFF \Reg_Bank/registers_reg[8][23]  ( .D(\Reg_Bank/n3277 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][23] ) );
  DFF \Reg_Bank/registers_reg[8][24]  ( .D(\Reg_Bank/n3278 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][24] ) );
  DFF \Reg_Bank/registers_reg[8][25]  ( .D(\Reg_Bank/n3279 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][25] ) );
  DFF \Reg_Bank/registers_reg[8][26]  ( .D(\Reg_Bank/n3280 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][26] ) );
  DFF \Reg_Bank/registers_reg[8][27]  ( .D(\Reg_Bank/n3281 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][27] ) );
  DFF \Reg_Bank/registers_reg[8][28]  ( .D(\Reg_Bank/n3282 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][28] ) );
  DFF \Reg_Bank/registers_reg[8][29]  ( .D(\Reg_Bank/n3283 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][29] ) );
  DFF \Reg_Bank/registers_reg[8][30]  ( .D(\Reg_Bank/n3284 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][30] ) );
  DFF \Reg_Bank/registers_reg[8][31]  ( .D(\Reg_Bank/n3285 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][31] ) );
  DFF \Reg_Bank/registers_reg[9][0]  ( .D(\Reg_Bank/n3286 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][0] ) );
  DFF \Reg_Bank/registers_reg[9][1]  ( .D(\Reg_Bank/n3287 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][1] ) );
  DFF \Reg_Bank/registers_reg[9][2]  ( .D(\Reg_Bank/n3288 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][2] ) );
  DFF \Reg_Bank/registers_reg[9][3]  ( .D(\Reg_Bank/n3289 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][3] ) );
  DFF \Reg_Bank/registers_reg[9][4]  ( .D(\Reg_Bank/n3290 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][4] ) );
  DFF \Reg_Bank/registers_reg[9][5]  ( .D(\Reg_Bank/n3291 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][5] ) );
  DFF \Reg_Bank/registers_reg[9][6]  ( .D(\Reg_Bank/n3292 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][6] ) );
  DFF \Reg_Bank/registers_reg[9][7]  ( .D(\Reg_Bank/n3293 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][7] ) );
  DFF \Reg_Bank/registers_reg[9][8]  ( .D(\Reg_Bank/n3294 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][8] ) );
  DFF \Reg_Bank/registers_reg[9][9]  ( .D(\Reg_Bank/n3295 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][9] ) );
  DFF \Reg_Bank/registers_reg[9][10]  ( .D(\Reg_Bank/n3296 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][10] ) );
  DFF \Reg_Bank/registers_reg[9][11]  ( .D(\Reg_Bank/n3297 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][11] ) );
  DFF \Reg_Bank/registers_reg[9][12]  ( .D(\Reg_Bank/n3298 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][12] ) );
  DFF \Reg_Bank/registers_reg[9][13]  ( .D(\Reg_Bank/n3299 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][13] ) );
  DFF \Reg_Bank/registers_reg[9][14]  ( .D(\Reg_Bank/n3300 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][14] ) );
  DFF \Reg_Bank/registers_reg[9][15]  ( .D(\Reg_Bank/n3301 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][15] ) );
  DFF \Reg_Bank/registers_reg[9][16]  ( .D(\Reg_Bank/n3302 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][16] ) );
  DFF \Reg_Bank/registers_reg[9][17]  ( .D(\Reg_Bank/n3303 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][17] ) );
  DFF \Reg_Bank/registers_reg[9][18]  ( .D(\Reg_Bank/n3304 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][18] ) );
  DFF \Reg_Bank/registers_reg[9][19]  ( .D(\Reg_Bank/n3305 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][19] ) );
  DFF \Reg_Bank/registers_reg[9][20]  ( .D(\Reg_Bank/n3306 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][20] ) );
  DFF \Reg_Bank/registers_reg[9][21]  ( .D(\Reg_Bank/n3307 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][21] ) );
  DFF \Reg_Bank/registers_reg[9][22]  ( .D(\Reg_Bank/n3308 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][22] ) );
  DFF \Reg_Bank/registers_reg[9][23]  ( .D(\Reg_Bank/n3309 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][23] ) );
  DFF \Reg_Bank/registers_reg[9][24]  ( .D(\Reg_Bank/n3310 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][24] ) );
  DFF \Reg_Bank/registers_reg[9][25]  ( .D(\Reg_Bank/n3311 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][25] ) );
  DFF \Reg_Bank/registers_reg[9][26]  ( .D(\Reg_Bank/n3312 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][26] ) );
  DFF \Reg_Bank/registers_reg[9][27]  ( .D(\Reg_Bank/n3313 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][27] ) );
  DFF \Reg_Bank/registers_reg[9][28]  ( .D(\Reg_Bank/n3314 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][28] ) );
  DFF \Reg_Bank/registers_reg[9][29]  ( .D(\Reg_Bank/n3315 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][29] ) );
  DFF \Reg_Bank/registers_reg[9][30]  ( .D(\Reg_Bank/n3316 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][30] ) );
  DFF \Reg_Bank/registers_reg[9][31]  ( .D(\Reg_Bank/n3317 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][31] ) );
  DFF \Reg_Bank/registers_reg[10][0]  ( .D(\Reg_Bank/n3318 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][0] ) );
  DFF \Reg_Bank/registers_reg[10][1]  ( .D(\Reg_Bank/n3319 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][1] ) );
  DFF \Reg_Bank/registers_reg[10][2]  ( .D(\Reg_Bank/n3320 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][2] ) );
  DFF \Reg_Bank/registers_reg[10][3]  ( .D(\Reg_Bank/n3321 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][3] ) );
  DFF \Reg_Bank/registers_reg[10][4]  ( .D(\Reg_Bank/n3322 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][4] ) );
  DFF \Reg_Bank/registers_reg[10][5]  ( .D(\Reg_Bank/n3323 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][5] ) );
  DFF \Reg_Bank/registers_reg[10][6]  ( .D(\Reg_Bank/n3324 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][6] ) );
  DFF \Reg_Bank/registers_reg[10][7]  ( .D(\Reg_Bank/n3325 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][7] ) );
  DFF \Reg_Bank/registers_reg[10][8]  ( .D(\Reg_Bank/n3326 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][8] ) );
  DFF \Reg_Bank/registers_reg[10][9]  ( .D(\Reg_Bank/n3327 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][9] ) );
  DFF \Reg_Bank/registers_reg[10][10]  ( .D(\Reg_Bank/n3328 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][10] ) );
  DFF \Reg_Bank/registers_reg[10][11]  ( .D(\Reg_Bank/n3329 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][11] ) );
  DFF \Reg_Bank/registers_reg[10][12]  ( .D(\Reg_Bank/n3330 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][12] ) );
  DFF \Reg_Bank/registers_reg[10][13]  ( .D(\Reg_Bank/n3331 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][13] ) );
  DFF \Reg_Bank/registers_reg[10][14]  ( .D(\Reg_Bank/n3332 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][14] ) );
  DFF \Reg_Bank/registers_reg[10][15]  ( .D(\Reg_Bank/n3333 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][15] ) );
  DFF \Reg_Bank/registers_reg[10][16]  ( .D(\Reg_Bank/n3334 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][16] ) );
  DFF \Reg_Bank/registers_reg[10][17]  ( .D(\Reg_Bank/n3335 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][17] ) );
  DFF \Reg_Bank/registers_reg[10][18]  ( .D(\Reg_Bank/n3336 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][18] ) );
  DFF \Reg_Bank/registers_reg[10][19]  ( .D(\Reg_Bank/n3337 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][19] ) );
  DFF \Reg_Bank/registers_reg[10][20]  ( .D(\Reg_Bank/n3338 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][20] ) );
  DFF \Reg_Bank/registers_reg[10][21]  ( .D(\Reg_Bank/n3339 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][21] ) );
  DFF \Reg_Bank/registers_reg[10][22]  ( .D(\Reg_Bank/n3340 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][22] ) );
  DFF \Reg_Bank/registers_reg[10][23]  ( .D(\Reg_Bank/n3341 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][23] ) );
  DFF \Reg_Bank/registers_reg[10][24]  ( .D(\Reg_Bank/n3342 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][24] ) );
  DFF \Reg_Bank/registers_reg[10][25]  ( .D(\Reg_Bank/n3343 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][25] ) );
  DFF \Reg_Bank/registers_reg[10][26]  ( .D(\Reg_Bank/n3344 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][26] ) );
  DFF \Reg_Bank/registers_reg[10][27]  ( .D(\Reg_Bank/n3345 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][27] ) );
  DFF \Reg_Bank/registers_reg[10][28]  ( .D(\Reg_Bank/n3346 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][28] ) );
  DFF \Reg_Bank/registers_reg[10][29]  ( .D(\Reg_Bank/n3347 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][29] ) );
  DFF \Reg_Bank/registers_reg[10][30]  ( .D(\Reg_Bank/n3348 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][30] ) );
  DFF \Reg_Bank/registers_reg[10][31]  ( .D(\Reg_Bank/n3349 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][31] ) );
  DFF \Reg_Bank/registers_reg[11][0]  ( .D(\Reg_Bank/n3350 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][0] ) );
  DFF \Reg_Bank/registers_reg[11][1]  ( .D(\Reg_Bank/n3351 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][1] ) );
  DFF \Reg_Bank/registers_reg[11][2]  ( .D(\Reg_Bank/n3352 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][2] ) );
  DFF \Reg_Bank/registers_reg[11][3]  ( .D(\Reg_Bank/n3353 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][3] ) );
  DFF \Reg_Bank/registers_reg[11][4]  ( .D(\Reg_Bank/n3354 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][4] ) );
  DFF \Reg_Bank/registers_reg[11][5]  ( .D(\Reg_Bank/n3355 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][5] ) );
  DFF \Reg_Bank/registers_reg[11][6]  ( .D(\Reg_Bank/n3356 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][6] ) );
  DFF \Reg_Bank/registers_reg[11][7]  ( .D(\Reg_Bank/n3357 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][7] ) );
  DFF \Reg_Bank/registers_reg[11][8]  ( .D(\Reg_Bank/n3358 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][8] ) );
  DFF \Reg_Bank/registers_reg[11][9]  ( .D(\Reg_Bank/n3359 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][9] ) );
  DFF \Reg_Bank/registers_reg[11][10]  ( .D(\Reg_Bank/n3360 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][10] ) );
  DFF \Reg_Bank/registers_reg[11][11]  ( .D(\Reg_Bank/n3361 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][11] ) );
  DFF \Reg_Bank/registers_reg[11][12]  ( .D(\Reg_Bank/n3362 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][12] ) );
  DFF \Reg_Bank/registers_reg[11][13]  ( .D(\Reg_Bank/n3363 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][13] ) );
  DFF \Reg_Bank/registers_reg[11][14]  ( .D(\Reg_Bank/n3364 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][14] ) );
  DFF \Reg_Bank/registers_reg[11][15]  ( .D(\Reg_Bank/n3365 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][15] ) );
  DFF \Reg_Bank/registers_reg[11][16]  ( .D(\Reg_Bank/n3366 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][16] ) );
  DFF \Reg_Bank/registers_reg[11][17]  ( .D(\Reg_Bank/n3367 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][17] ) );
  DFF \Reg_Bank/registers_reg[11][18]  ( .D(\Reg_Bank/n3368 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][18] ) );
  DFF \Reg_Bank/registers_reg[11][19]  ( .D(\Reg_Bank/n3369 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][19] ) );
  DFF \Reg_Bank/registers_reg[11][20]  ( .D(\Reg_Bank/n3370 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][20] ) );
  DFF \Reg_Bank/registers_reg[11][21]  ( .D(\Reg_Bank/n3371 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][21] ) );
  DFF \Reg_Bank/registers_reg[11][22]  ( .D(\Reg_Bank/n3372 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][22] ) );
  DFF \Reg_Bank/registers_reg[11][23]  ( .D(\Reg_Bank/n3373 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][23] ) );
  DFF \Reg_Bank/registers_reg[11][24]  ( .D(\Reg_Bank/n3374 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][24] ) );
  DFF \Reg_Bank/registers_reg[11][25]  ( .D(\Reg_Bank/n3375 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][25] ) );
  DFF \Reg_Bank/registers_reg[11][26]  ( .D(\Reg_Bank/n3376 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][26] ) );
  DFF \Reg_Bank/registers_reg[11][27]  ( .D(\Reg_Bank/n3377 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][27] ) );
  DFF \Reg_Bank/registers_reg[11][28]  ( .D(\Reg_Bank/n3378 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][28] ) );
  DFF \Reg_Bank/registers_reg[11][29]  ( .D(\Reg_Bank/n3379 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][29] ) );
  DFF \Reg_Bank/registers_reg[11][30]  ( .D(\Reg_Bank/n3380 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][30] ) );
  DFF \Reg_Bank/registers_reg[11][31]  ( .D(\Reg_Bank/n3381 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][31] ) );
  DFF \Reg_Bank/registers_reg[12][0]  ( .D(\Reg_Bank/n3382 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][0] ) );
  DFF \Reg_Bank/registers_reg[12][1]  ( .D(\Reg_Bank/n3383 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][1] ) );
  DFF \Reg_Bank/registers_reg[12][2]  ( .D(\Reg_Bank/n3384 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][2] ) );
  DFF \Reg_Bank/registers_reg[12][3]  ( .D(\Reg_Bank/n3385 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][3] ) );
  DFF \Reg_Bank/registers_reg[12][4]  ( .D(\Reg_Bank/n3386 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][4] ) );
  DFF \Reg_Bank/registers_reg[12][5]  ( .D(\Reg_Bank/n3387 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][5] ) );
  DFF \Reg_Bank/registers_reg[12][6]  ( .D(\Reg_Bank/n3388 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][6] ) );
  DFF \Reg_Bank/registers_reg[12][7]  ( .D(\Reg_Bank/n3389 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][7] ) );
  DFF \Reg_Bank/registers_reg[12][8]  ( .D(\Reg_Bank/n3390 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][8] ) );
  DFF \Reg_Bank/registers_reg[12][9]  ( .D(\Reg_Bank/n3391 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][9] ) );
  DFF \Reg_Bank/registers_reg[12][10]  ( .D(\Reg_Bank/n3392 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][10] ) );
  DFF \Reg_Bank/registers_reg[12][11]  ( .D(\Reg_Bank/n3393 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][11] ) );
  DFF \Reg_Bank/registers_reg[12][12]  ( .D(\Reg_Bank/n3394 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][12] ) );
  DFF \Reg_Bank/registers_reg[12][13]  ( .D(\Reg_Bank/n3395 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][13] ) );
  DFF \Reg_Bank/registers_reg[12][14]  ( .D(\Reg_Bank/n3396 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][14] ) );
  DFF \Reg_Bank/registers_reg[12][15]  ( .D(\Reg_Bank/n3397 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][15] ) );
  DFF \Reg_Bank/registers_reg[12][16]  ( .D(\Reg_Bank/n3398 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][16] ) );
  DFF \Reg_Bank/registers_reg[12][17]  ( .D(\Reg_Bank/n3399 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][17] ) );
  DFF \Reg_Bank/registers_reg[12][18]  ( .D(\Reg_Bank/n3400 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][18] ) );
  DFF \Reg_Bank/registers_reg[12][19]  ( .D(\Reg_Bank/n3401 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][19] ) );
  DFF \Reg_Bank/registers_reg[12][20]  ( .D(\Reg_Bank/n3402 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][20] ) );
  DFF \Reg_Bank/registers_reg[12][21]  ( .D(\Reg_Bank/n3403 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][21] ) );
  DFF \Reg_Bank/registers_reg[12][22]  ( .D(\Reg_Bank/n3404 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][22] ) );
  DFF \Reg_Bank/registers_reg[12][23]  ( .D(\Reg_Bank/n3405 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][23] ) );
  DFF \Reg_Bank/registers_reg[12][24]  ( .D(\Reg_Bank/n3406 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][24] ) );
  DFF \Reg_Bank/registers_reg[12][25]  ( .D(\Reg_Bank/n3407 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][25] ) );
  DFF \Reg_Bank/registers_reg[12][26]  ( .D(\Reg_Bank/n3408 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][26] ) );
  DFF \Reg_Bank/registers_reg[12][27]  ( .D(\Reg_Bank/n3409 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][27] ) );
  DFF \Reg_Bank/registers_reg[12][28]  ( .D(\Reg_Bank/n3410 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][28] ) );
  DFF \Reg_Bank/registers_reg[12][29]  ( .D(\Reg_Bank/n3411 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][29] ) );
  DFF \Reg_Bank/registers_reg[12][30]  ( .D(\Reg_Bank/n3412 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][30] ) );
  DFF \Reg_Bank/registers_reg[12][31]  ( .D(\Reg_Bank/n3413 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][31] ) );
  DFF \Reg_Bank/registers_reg[13][0]  ( .D(\Reg_Bank/n3414 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][0] ) );
  DFF \Reg_Bank/registers_reg[13][1]  ( .D(\Reg_Bank/n3415 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][1] ) );
  DFF \Reg_Bank/registers_reg[13][2]  ( .D(\Reg_Bank/n3416 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][2] ) );
  DFF \Reg_Bank/registers_reg[13][3]  ( .D(\Reg_Bank/n3417 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][3] ) );
  DFF \Reg_Bank/registers_reg[13][4]  ( .D(\Reg_Bank/n3418 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][4] ) );
  DFF \Reg_Bank/registers_reg[13][5]  ( .D(\Reg_Bank/n3419 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][5] ) );
  DFF \Reg_Bank/registers_reg[13][6]  ( .D(\Reg_Bank/n3420 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][6] ) );
  DFF \Reg_Bank/registers_reg[13][7]  ( .D(\Reg_Bank/n3421 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][7] ) );
  DFF \Reg_Bank/registers_reg[13][8]  ( .D(\Reg_Bank/n3422 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][8] ) );
  DFF \Reg_Bank/registers_reg[13][9]  ( .D(\Reg_Bank/n3423 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][9] ) );
  DFF \Reg_Bank/registers_reg[13][10]  ( .D(\Reg_Bank/n3424 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][10] ) );
  DFF \Reg_Bank/registers_reg[13][11]  ( .D(\Reg_Bank/n3425 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][11] ) );
  DFF \Reg_Bank/registers_reg[13][12]  ( .D(\Reg_Bank/n3426 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][12] ) );
  DFF \Reg_Bank/registers_reg[13][13]  ( .D(\Reg_Bank/n3427 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][13] ) );
  DFF \Reg_Bank/registers_reg[13][14]  ( .D(\Reg_Bank/n3428 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][14] ) );
  DFF \Reg_Bank/registers_reg[13][15]  ( .D(\Reg_Bank/n3429 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][15] ) );
  DFF \Reg_Bank/registers_reg[13][16]  ( .D(\Reg_Bank/n3430 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][16] ) );
  DFF \Reg_Bank/registers_reg[13][17]  ( .D(\Reg_Bank/n3431 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][17] ) );
  DFF \Reg_Bank/registers_reg[13][18]  ( .D(\Reg_Bank/n3432 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][18] ) );
  DFF \Reg_Bank/registers_reg[13][19]  ( .D(\Reg_Bank/n3433 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][19] ) );
  DFF \Reg_Bank/registers_reg[13][20]  ( .D(\Reg_Bank/n3434 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][20] ) );
  DFF \Reg_Bank/registers_reg[13][21]  ( .D(\Reg_Bank/n3435 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][21] ) );
  DFF \Reg_Bank/registers_reg[13][22]  ( .D(\Reg_Bank/n3436 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][22] ) );
  DFF \Reg_Bank/registers_reg[13][23]  ( .D(\Reg_Bank/n3437 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][23] ) );
  DFF \Reg_Bank/registers_reg[13][24]  ( .D(\Reg_Bank/n3438 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][24] ) );
  DFF \Reg_Bank/registers_reg[13][25]  ( .D(\Reg_Bank/n3439 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][25] ) );
  DFF \Reg_Bank/registers_reg[13][26]  ( .D(\Reg_Bank/n3440 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][26] ) );
  DFF \Reg_Bank/registers_reg[13][27]  ( .D(\Reg_Bank/n3441 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][27] ) );
  DFF \Reg_Bank/registers_reg[13][28]  ( .D(\Reg_Bank/n3442 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][28] ) );
  DFF \Reg_Bank/registers_reg[13][29]  ( .D(\Reg_Bank/n3443 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][29] ) );
  DFF \Reg_Bank/registers_reg[13][30]  ( .D(\Reg_Bank/n3444 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][30] ) );
  DFF \Reg_Bank/registers_reg[13][31]  ( .D(\Reg_Bank/n3445 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][31] ) );
  DFF \Reg_Bank/registers_reg[14][0]  ( .D(\Reg_Bank/n3446 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][0] ) );
  DFF \Reg_Bank/registers_reg[14][1]  ( .D(\Reg_Bank/n3447 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][1] ) );
  DFF \Reg_Bank/registers_reg[14][2]  ( .D(\Reg_Bank/n3448 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][2] ) );
  DFF \Reg_Bank/registers_reg[14][3]  ( .D(\Reg_Bank/n3449 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][3] ) );
  DFF \Reg_Bank/registers_reg[14][4]  ( .D(\Reg_Bank/n3450 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][4] ) );
  DFF \Reg_Bank/registers_reg[14][5]  ( .D(\Reg_Bank/n3451 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][5] ) );
  DFF \Reg_Bank/registers_reg[14][6]  ( .D(\Reg_Bank/n3452 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][6] ) );
  DFF \Reg_Bank/registers_reg[14][7]  ( .D(\Reg_Bank/n3453 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][7] ) );
  DFF \Reg_Bank/registers_reg[14][8]  ( .D(\Reg_Bank/n3454 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][8] ) );
  DFF \Reg_Bank/registers_reg[14][9]  ( .D(\Reg_Bank/n3455 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][9] ) );
  DFF \Reg_Bank/registers_reg[14][10]  ( .D(\Reg_Bank/n3456 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][10] ) );
  DFF \Reg_Bank/registers_reg[14][11]  ( .D(\Reg_Bank/n3457 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][11] ) );
  DFF \Reg_Bank/registers_reg[14][12]  ( .D(\Reg_Bank/n3458 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][12] ) );
  DFF \Reg_Bank/registers_reg[14][13]  ( .D(\Reg_Bank/n3459 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][13] ) );
  DFF \Reg_Bank/registers_reg[14][14]  ( .D(\Reg_Bank/n3460 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][14] ) );
  DFF \Reg_Bank/registers_reg[14][15]  ( .D(\Reg_Bank/n3461 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][15] ) );
  DFF \Reg_Bank/registers_reg[14][16]  ( .D(\Reg_Bank/n3462 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][16] ) );
  DFF \Reg_Bank/registers_reg[14][17]  ( .D(\Reg_Bank/n3463 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][17] ) );
  DFF \Reg_Bank/registers_reg[14][18]  ( .D(\Reg_Bank/n3464 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][18] ) );
  DFF \Reg_Bank/registers_reg[14][19]  ( .D(\Reg_Bank/n3465 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][19] ) );
  DFF \Reg_Bank/registers_reg[14][20]  ( .D(\Reg_Bank/n3466 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][20] ) );
  DFF \Reg_Bank/registers_reg[14][21]  ( .D(\Reg_Bank/n3467 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][21] ) );
  DFF \Reg_Bank/registers_reg[14][22]  ( .D(\Reg_Bank/n3468 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][22] ) );
  DFF \Reg_Bank/registers_reg[14][23]  ( .D(\Reg_Bank/n3469 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][23] ) );
  DFF \Reg_Bank/registers_reg[14][24]  ( .D(\Reg_Bank/n3470 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][24] ) );
  DFF \Reg_Bank/registers_reg[14][25]  ( .D(\Reg_Bank/n3471 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][25] ) );
  DFF \Reg_Bank/registers_reg[14][26]  ( .D(\Reg_Bank/n3472 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][26] ) );
  DFF \Reg_Bank/registers_reg[14][27]  ( .D(\Reg_Bank/n3473 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][27] ) );
  DFF \Reg_Bank/registers_reg[14][28]  ( .D(\Reg_Bank/n3474 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][28] ) );
  DFF \Reg_Bank/registers_reg[14][29]  ( .D(\Reg_Bank/n3475 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][29] ) );
  DFF \Reg_Bank/registers_reg[14][30]  ( .D(\Reg_Bank/n3476 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][30] ) );
  DFF \Reg_Bank/registers_reg[14][31]  ( .D(\Reg_Bank/n3477 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][31] ) );
  DFF \Reg_Bank/registers_reg[15][0]  ( .D(\Reg_Bank/n3478 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][0] ) );
  DFF \Reg_Bank/registers_reg[15][1]  ( .D(\Reg_Bank/n3479 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][1] ) );
  DFF \Reg_Bank/registers_reg[15][2]  ( .D(\Reg_Bank/n3480 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][2] ) );
  DFF \Reg_Bank/registers_reg[15][3]  ( .D(\Reg_Bank/n3481 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][3] ) );
  DFF \Reg_Bank/registers_reg[15][4]  ( .D(\Reg_Bank/n3482 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][4] ) );
  DFF \Reg_Bank/registers_reg[15][5]  ( .D(\Reg_Bank/n3483 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][5] ) );
  DFF \Reg_Bank/registers_reg[15][6]  ( .D(\Reg_Bank/n3484 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][6] ) );
  DFF \Reg_Bank/registers_reg[15][7]  ( .D(\Reg_Bank/n3485 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][7] ) );
  DFF \Reg_Bank/registers_reg[15][8]  ( .D(\Reg_Bank/n3486 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][8] ) );
  DFF \Reg_Bank/registers_reg[15][9]  ( .D(\Reg_Bank/n3487 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][9] ) );
  DFF \Reg_Bank/registers_reg[15][10]  ( .D(\Reg_Bank/n3488 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][10] ) );
  DFF \Reg_Bank/registers_reg[15][11]  ( .D(\Reg_Bank/n3489 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][11] ) );
  DFF \Reg_Bank/registers_reg[15][12]  ( .D(\Reg_Bank/n3490 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][12] ) );
  DFF \Reg_Bank/registers_reg[15][13]  ( .D(\Reg_Bank/n3491 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][13] ) );
  DFF \Reg_Bank/registers_reg[15][14]  ( .D(\Reg_Bank/n3492 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][14] ) );
  DFF \Reg_Bank/registers_reg[15][15]  ( .D(\Reg_Bank/n3493 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][15] ) );
  DFF \Reg_Bank/registers_reg[15][16]  ( .D(\Reg_Bank/n3494 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][16] ) );
  DFF \Reg_Bank/registers_reg[15][17]  ( .D(\Reg_Bank/n3495 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][17] ) );
  DFF \Reg_Bank/registers_reg[15][18]  ( .D(\Reg_Bank/n3496 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][18] ) );
  DFF \Reg_Bank/registers_reg[15][19]  ( .D(\Reg_Bank/n3497 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][19] ) );
  DFF \Reg_Bank/registers_reg[15][20]  ( .D(\Reg_Bank/n3498 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][20] ) );
  DFF \Reg_Bank/registers_reg[15][21]  ( .D(\Reg_Bank/n3499 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][21] ) );
  DFF \Reg_Bank/registers_reg[15][22]  ( .D(\Reg_Bank/n3500 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][22] ) );
  DFF \Reg_Bank/registers_reg[15][23]  ( .D(\Reg_Bank/n3501 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][23] ) );
  DFF \Reg_Bank/registers_reg[15][24]  ( .D(\Reg_Bank/n3502 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][24] ) );
  DFF \Reg_Bank/registers_reg[15][25]  ( .D(\Reg_Bank/n3503 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][25] ) );
  DFF \Reg_Bank/registers_reg[15][26]  ( .D(\Reg_Bank/n3504 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][26] ) );
  DFF \Reg_Bank/registers_reg[15][27]  ( .D(\Reg_Bank/n3505 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][27] ) );
  DFF \Reg_Bank/registers_reg[15][28]  ( .D(\Reg_Bank/n3506 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][28] ) );
  DFF \Reg_Bank/registers_reg[15][29]  ( .D(\Reg_Bank/n3507 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][29] ) );
  DFF \Reg_Bank/registers_reg[15][30]  ( .D(\Reg_Bank/n3508 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][30] ) );
  DFF \Reg_Bank/registers_reg[15][31]  ( .D(\Reg_Bank/n3509 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][31] ) );
  DFF \Reg_Bank/registers_reg[16][0]  ( .D(\Reg_Bank/n3510 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][0] ) );
  DFF \Reg_Bank/registers_reg[16][1]  ( .D(\Reg_Bank/n3511 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][1] ) );
  DFF \Reg_Bank/registers_reg[16][2]  ( .D(\Reg_Bank/n3512 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][2] ) );
  DFF \Reg_Bank/registers_reg[16][3]  ( .D(\Reg_Bank/n3513 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][3] ) );
  DFF \Reg_Bank/registers_reg[16][4]  ( .D(\Reg_Bank/n3514 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][4] ) );
  DFF \Reg_Bank/registers_reg[16][5]  ( .D(\Reg_Bank/n3515 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][5] ) );
  DFF \Reg_Bank/registers_reg[16][6]  ( .D(\Reg_Bank/n3516 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][6] ) );
  DFF \Reg_Bank/registers_reg[16][7]  ( .D(\Reg_Bank/n3517 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][7] ) );
  DFF \Reg_Bank/registers_reg[16][8]  ( .D(\Reg_Bank/n3518 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][8] ) );
  DFF \Reg_Bank/registers_reg[16][9]  ( .D(\Reg_Bank/n3519 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][9] ) );
  DFF \Reg_Bank/registers_reg[16][10]  ( .D(\Reg_Bank/n3520 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][10] ) );
  DFF \Reg_Bank/registers_reg[16][11]  ( .D(\Reg_Bank/n3521 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][11] ) );
  DFF \Reg_Bank/registers_reg[16][12]  ( .D(\Reg_Bank/n3522 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][12] ) );
  DFF \Reg_Bank/registers_reg[16][13]  ( .D(\Reg_Bank/n3523 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][13] ) );
  DFF \Reg_Bank/registers_reg[16][14]  ( .D(\Reg_Bank/n3524 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][14] ) );
  DFF \Reg_Bank/registers_reg[16][15]  ( .D(\Reg_Bank/n3525 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][15] ) );
  DFF \Reg_Bank/registers_reg[16][16]  ( .D(\Reg_Bank/n3526 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][16] ) );
  DFF \Reg_Bank/registers_reg[16][17]  ( .D(\Reg_Bank/n3527 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][17] ) );
  DFF \Reg_Bank/registers_reg[16][18]  ( .D(\Reg_Bank/n3528 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][18] ) );
  DFF \Reg_Bank/registers_reg[16][19]  ( .D(\Reg_Bank/n3529 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][19] ) );
  DFF \Reg_Bank/registers_reg[16][20]  ( .D(\Reg_Bank/n3530 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][20] ) );
  DFF \Reg_Bank/registers_reg[16][21]  ( .D(\Reg_Bank/n3531 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][21] ) );
  DFF \Reg_Bank/registers_reg[16][22]  ( .D(\Reg_Bank/n3532 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][22] ) );
  DFF \Reg_Bank/registers_reg[16][23]  ( .D(\Reg_Bank/n3533 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][23] ) );
  DFF \Reg_Bank/registers_reg[16][24]  ( .D(\Reg_Bank/n3534 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][24] ) );
  DFF \Reg_Bank/registers_reg[16][25]  ( .D(\Reg_Bank/n3535 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][25] ) );
  DFF \Reg_Bank/registers_reg[16][26]  ( .D(\Reg_Bank/n3536 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][26] ) );
  DFF \Reg_Bank/registers_reg[16][27]  ( .D(\Reg_Bank/n3537 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][27] ) );
  DFF \Reg_Bank/registers_reg[16][28]  ( .D(\Reg_Bank/n3538 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][28] ) );
  DFF \Reg_Bank/registers_reg[16][29]  ( .D(\Reg_Bank/n3539 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][29] ) );
  DFF \Reg_Bank/registers_reg[16][30]  ( .D(\Reg_Bank/n3540 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][30] ) );
  DFF \Reg_Bank/registers_reg[16][31]  ( .D(\Reg_Bank/n3541 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][31] ) );
  DFF \Reg_Bank/registers_reg[17][0]  ( .D(\Reg_Bank/n3542 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][0] ) );
  DFF \Reg_Bank/registers_reg[17][1]  ( .D(\Reg_Bank/n3543 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][1] ) );
  DFF \Reg_Bank/registers_reg[17][2]  ( .D(\Reg_Bank/n3544 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][2] ) );
  DFF \Reg_Bank/registers_reg[17][3]  ( .D(\Reg_Bank/n3545 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][3] ) );
  DFF \Reg_Bank/registers_reg[17][4]  ( .D(\Reg_Bank/n3546 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][4] ) );
  DFF \Reg_Bank/registers_reg[17][5]  ( .D(\Reg_Bank/n3547 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][5] ) );
  DFF \Reg_Bank/registers_reg[17][6]  ( .D(\Reg_Bank/n3548 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][6] ) );
  DFF \Reg_Bank/registers_reg[17][7]  ( .D(\Reg_Bank/n3549 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][7] ) );
  DFF \Reg_Bank/registers_reg[17][8]  ( .D(\Reg_Bank/n3550 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][8] ) );
  DFF \Reg_Bank/registers_reg[17][9]  ( .D(\Reg_Bank/n3551 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][9] ) );
  DFF \Reg_Bank/registers_reg[17][10]  ( .D(\Reg_Bank/n3552 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][10] ) );
  DFF \Reg_Bank/registers_reg[17][11]  ( .D(\Reg_Bank/n3553 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][11] ) );
  DFF \Reg_Bank/registers_reg[17][12]  ( .D(\Reg_Bank/n3554 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][12] ) );
  DFF \Reg_Bank/registers_reg[17][13]  ( .D(\Reg_Bank/n3555 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][13] ) );
  DFF \Reg_Bank/registers_reg[17][14]  ( .D(\Reg_Bank/n3556 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][14] ) );
  DFF \Reg_Bank/registers_reg[17][15]  ( .D(\Reg_Bank/n3557 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][15] ) );
  DFF \Reg_Bank/registers_reg[17][16]  ( .D(\Reg_Bank/n3558 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][16] ) );
  DFF \Reg_Bank/registers_reg[17][17]  ( .D(\Reg_Bank/n3559 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][17] ) );
  DFF \Reg_Bank/registers_reg[17][18]  ( .D(\Reg_Bank/n3560 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][18] ) );
  DFF \Reg_Bank/registers_reg[17][19]  ( .D(\Reg_Bank/n3561 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][19] ) );
  DFF \Reg_Bank/registers_reg[17][20]  ( .D(\Reg_Bank/n3562 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][20] ) );
  DFF \Reg_Bank/registers_reg[17][21]  ( .D(\Reg_Bank/n3563 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][21] ) );
  DFF \Reg_Bank/registers_reg[17][22]  ( .D(\Reg_Bank/n3564 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][22] ) );
  DFF \Reg_Bank/registers_reg[17][23]  ( .D(\Reg_Bank/n3565 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][23] ) );
  DFF \Reg_Bank/registers_reg[17][24]  ( .D(\Reg_Bank/n3566 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][24] ) );
  DFF \Reg_Bank/registers_reg[17][25]  ( .D(\Reg_Bank/n3567 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][25] ) );
  DFF \Reg_Bank/registers_reg[17][26]  ( .D(\Reg_Bank/n3568 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][26] ) );
  DFF \Reg_Bank/registers_reg[17][27]  ( .D(\Reg_Bank/n3569 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][27] ) );
  DFF \Reg_Bank/registers_reg[17][28]  ( .D(\Reg_Bank/n3570 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][28] ) );
  DFF \Reg_Bank/registers_reg[17][29]  ( .D(\Reg_Bank/n3571 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][29] ) );
  DFF \Reg_Bank/registers_reg[17][30]  ( .D(\Reg_Bank/n3572 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][30] ) );
  DFF \Reg_Bank/registers_reg[17][31]  ( .D(\Reg_Bank/n3573 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][31] ) );
  DFF \Reg_Bank/registers_reg[18][0]  ( .D(\Reg_Bank/n3574 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][0] ) );
  DFF \Reg_Bank/registers_reg[18][1]  ( .D(\Reg_Bank/n3575 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][1] ) );
  DFF \Reg_Bank/registers_reg[18][2]  ( .D(\Reg_Bank/n3576 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][2] ) );
  DFF \Reg_Bank/registers_reg[18][3]  ( .D(\Reg_Bank/n3577 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][3] ) );
  DFF \Reg_Bank/registers_reg[18][4]  ( .D(\Reg_Bank/n3578 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][4] ) );
  DFF \Reg_Bank/registers_reg[18][5]  ( .D(\Reg_Bank/n3579 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][5] ) );
  DFF \Reg_Bank/registers_reg[18][6]  ( .D(\Reg_Bank/n3580 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][6] ) );
  DFF \Reg_Bank/registers_reg[18][7]  ( .D(\Reg_Bank/n3581 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][7] ) );
  DFF \Reg_Bank/registers_reg[18][8]  ( .D(\Reg_Bank/n3582 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][8] ) );
  DFF \Reg_Bank/registers_reg[18][9]  ( .D(\Reg_Bank/n3583 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][9] ) );
  DFF \Reg_Bank/registers_reg[18][10]  ( .D(\Reg_Bank/n3584 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][10] ) );
  DFF \Reg_Bank/registers_reg[18][11]  ( .D(\Reg_Bank/n3585 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][11] ) );
  DFF \Reg_Bank/registers_reg[18][12]  ( .D(\Reg_Bank/n3586 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][12] ) );
  DFF \Reg_Bank/registers_reg[18][13]  ( .D(\Reg_Bank/n3587 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][13] ) );
  DFF \Reg_Bank/registers_reg[18][14]  ( .D(\Reg_Bank/n3588 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][14] ) );
  DFF \Reg_Bank/registers_reg[18][15]  ( .D(\Reg_Bank/n3589 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][15] ) );
  DFF \Reg_Bank/registers_reg[18][16]  ( .D(\Reg_Bank/n3590 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][16] ) );
  DFF \Reg_Bank/registers_reg[18][17]  ( .D(\Reg_Bank/n3591 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][17] ) );
  DFF \Reg_Bank/registers_reg[18][18]  ( .D(\Reg_Bank/n3592 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][18] ) );
  DFF \Reg_Bank/registers_reg[18][19]  ( .D(\Reg_Bank/n3593 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][19] ) );
  DFF \Reg_Bank/registers_reg[18][20]  ( .D(\Reg_Bank/n3594 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][20] ) );
  DFF \Reg_Bank/registers_reg[18][21]  ( .D(\Reg_Bank/n3595 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][21] ) );
  DFF \Reg_Bank/registers_reg[18][22]  ( .D(\Reg_Bank/n3596 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][22] ) );
  DFF \Reg_Bank/registers_reg[18][23]  ( .D(\Reg_Bank/n3597 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][23] ) );
  DFF \Reg_Bank/registers_reg[18][24]  ( .D(\Reg_Bank/n3598 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][24] ) );
  DFF \Reg_Bank/registers_reg[18][25]  ( .D(\Reg_Bank/n3599 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][25] ) );
  DFF \Reg_Bank/registers_reg[18][26]  ( .D(\Reg_Bank/n3600 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][26] ) );
  DFF \Reg_Bank/registers_reg[18][27]  ( .D(\Reg_Bank/n3601 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][27] ) );
  DFF \Reg_Bank/registers_reg[18][28]  ( .D(\Reg_Bank/n3602 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][28] ) );
  DFF \Reg_Bank/registers_reg[18][29]  ( .D(\Reg_Bank/n3603 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][29] ) );
  DFF \Reg_Bank/registers_reg[18][30]  ( .D(\Reg_Bank/n3604 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][30] ) );
  DFF \Reg_Bank/registers_reg[18][31]  ( .D(\Reg_Bank/n3605 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][31] ) );
  DFF \Reg_Bank/registers_reg[19][0]  ( .D(\Reg_Bank/n3606 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][0] ) );
  DFF \Reg_Bank/registers_reg[19][1]  ( .D(\Reg_Bank/n3607 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][1] ) );
  DFF \Reg_Bank/registers_reg[19][2]  ( .D(\Reg_Bank/n3608 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][2] ) );
  DFF \Reg_Bank/registers_reg[19][3]  ( .D(\Reg_Bank/n3609 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][3] ) );
  DFF \Reg_Bank/registers_reg[19][4]  ( .D(\Reg_Bank/n3610 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][4] ) );
  DFF \Reg_Bank/registers_reg[19][5]  ( .D(\Reg_Bank/n3611 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][5] ) );
  DFF \Reg_Bank/registers_reg[19][6]  ( .D(\Reg_Bank/n3612 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][6] ) );
  DFF \Reg_Bank/registers_reg[19][7]  ( .D(\Reg_Bank/n3613 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][7] ) );
  DFF \Reg_Bank/registers_reg[19][8]  ( .D(\Reg_Bank/n3614 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][8] ) );
  DFF \Reg_Bank/registers_reg[19][9]  ( .D(\Reg_Bank/n3615 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][9] ) );
  DFF \Reg_Bank/registers_reg[19][10]  ( .D(\Reg_Bank/n3616 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][10] ) );
  DFF \Reg_Bank/registers_reg[19][11]  ( .D(\Reg_Bank/n3617 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][11] ) );
  DFF \Reg_Bank/registers_reg[19][12]  ( .D(\Reg_Bank/n3618 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][12] ) );
  DFF \Reg_Bank/registers_reg[19][13]  ( .D(\Reg_Bank/n3619 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][13] ) );
  DFF \Reg_Bank/registers_reg[19][14]  ( .D(\Reg_Bank/n3620 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][14] ) );
  DFF \Reg_Bank/registers_reg[19][15]  ( .D(\Reg_Bank/n3621 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][15] ) );
  DFF \Reg_Bank/registers_reg[19][16]  ( .D(\Reg_Bank/n3622 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][16] ) );
  DFF \Reg_Bank/registers_reg[19][17]  ( .D(\Reg_Bank/n3623 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][17] ) );
  DFF \Reg_Bank/registers_reg[19][18]  ( .D(\Reg_Bank/n3624 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][18] ) );
  DFF \Reg_Bank/registers_reg[19][19]  ( .D(\Reg_Bank/n3625 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][19] ) );
  DFF \Reg_Bank/registers_reg[19][20]  ( .D(\Reg_Bank/n3626 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][20] ) );
  DFF \Reg_Bank/registers_reg[19][21]  ( .D(\Reg_Bank/n3627 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][21] ) );
  DFF \Reg_Bank/registers_reg[19][22]  ( .D(\Reg_Bank/n3628 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][22] ) );
  DFF \Reg_Bank/registers_reg[19][23]  ( .D(\Reg_Bank/n3629 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][23] ) );
  DFF \Reg_Bank/registers_reg[19][24]  ( .D(\Reg_Bank/n3630 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][24] ) );
  DFF \Reg_Bank/registers_reg[19][25]  ( .D(\Reg_Bank/n3631 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][25] ) );
  DFF \Reg_Bank/registers_reg[19][26]  ( .D(\Reg_Bank/n3632 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][26] ) );
  DFF \Reg_Bank/registers_reg[19][27]  ( .D(\Reg_Bank/n3633 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][27] ) );
  DFF \Reg_Bank/registers_reg[19][28]  ( .D(\Reg_Bank/n3634 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][28] ) );
  DFF \Reg_Bank/registers_reg[19][29]  ( .D(\Reg_Bank/n3635 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][29] ) );
  DFF \Reg_Bank/registers_reg[19][30]  ( .D(\Reg_Bank/n3636 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][30] ) );
  DFF \Reg_Bank/registers_reg[19][31]  ( .D(\Reg_Bank/n3637 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][31] ) );
  DFF \Reg_Bank/registers_reg[20][0]  ( .D(\Reg_Bank/n3638 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][0] ) );
  DFF \Reg_Bank/registers_reg[20][1]  ( .D(\Reg_Bank/n3639 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][1] ) );
  DFF \Reg_Bank/registers_reg[20][2]  ( .D(\Reg_Bank/n3640 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][2] ) );
  DFF \Reg_Bank/registers_reg[20][3]  ( .D(\Reg_Bank/n3641 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][3] ) );
  DFF \Reg_Bank/registers_reg[20][4]  ( .D(\Reg_Bank/n3642 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][4] ) );
  DFF \Reg_Bank/registers_reg[20][5]  ( .D(\Reg_Bank/n3643 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][5] ) );
  DFF \Reg_Bank/registers_reg[20][6]  ( .D(\Reg_Bank/n3644 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][6] ) );
  DFF \Reg_Bank/registers_reg[20][7]  ( .D(\Reg_Bank/n3645 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][7] ) );
  DFF \Reg_Bank/registers_reg[20][8]  ( .D(\Reg_Bank/n3646 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][8] ) );
  DFF \Reg_Bank/registers_reg[20][9]  ( .D(\Reg_Bank/n3647 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][9] ) );
  DFF \Reg_Bank/registers_reg[20][10]  ( .D(\Reg_Bank/n3648 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][10] ) );
  DFF \Reg_Bank/registers_reg[20][11]  ( .D(\Reg_Bank/n3649 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][11] ) );
  DFF \Reg_Bank/registers_reg[20][12]  ( .D(\Reg_Bank/n3650 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][12] ) );
  DFF \Reg_Bank/registers_reg[20][13]  ( .D(\Reg_Bank/n3651 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][13] ) );
  DFF \Reg_Bank/registers_reg[20][14]  ( .D(\Reg_Bank/n3652 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][14] ) );
  DFF \Reg_Bank/registers_reg[20][15]  ( .D(\Reg_Bank/n3653 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][15] ) );
  DFF \Reg_Bank/registers_reg[20][16]  ( .D(\Reg_Bank/n3654 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][16] ) );
  DFF \Reg_Bank/registers_reg[20][17]  ( .D(\Reg_Bank/n3655 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][17] ) );
  DFF \Reg_Bank/registers_reg[20][18]  ( .D(\Reg_Bank/n3656 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][18] ) );
  DFF \Reg_Bank/registers_reg[20][19]  ( .D(\Reg_Bank/n3657 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][19] ) );
  DFF \Reg_Bank/registers_reg[20][20]  ( .D(\Reg_Bank/n3658 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][20] ) );
  DFF \Reg_Bank/registers_reg[20][21]  ( .D(\Reg_Bank/n3659 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][21] ) );
  DFF \Reg_Bank/registers_reg[20][22]  ( .D(\Reg_Bank/n3660 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][22] ) );
  DFF \Reg_Bank/registers_reg[20][23]  ( .D(\Reg_Bank/n3661 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][23] ) );
  DFF \Reg_Bank/registers_reg[20][24]  ( .D(\Reg_Bank/n3662 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][24] ) );
  DFF \Reg_Bank/registers_reg[20][25]  ( .D(\Reg_Bank/n3663 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][25] ) );
  DFF \Reg_Bank/registers_reg[20][26]  ( .D(\Reg_Bank/n3664 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][26] ) );
  DFF \Reg_Bank/registers_reg[20][27]  ( .D(\Reg_Bank/n3665 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][27] ) );
  DFF \Reg_Bank/registers_reg[20][28]  ( .D(\Reg_Bank/n3666 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][28] ) );
  DFF \Reg_Bank/registers_reg[20][29]  ( .D(\Reg_Bank/n3667 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][29] ) );
  DFF \Reg_Bank/registers_reg[20][30]  ( .D(\Reg_Bank/n3668 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][30] ) );
  DFF \Reg_Bank/registers_reg[20][31]  ( .D(\Reg_Bank/n3669 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][31] ) );
  DFF \Reg_Bank/registers_reg[21][0]  ( .D(\Reg_Bank/n3670 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][0] ) );
  DFF \Reg_Bank/registers_reg[21][1]  ( .D(\Reg_Bank/n3671 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][1] ) );
  DFF \Reg_Bank/registers_reg[21][2]  ( .D(\Reg_Bank/n3672 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][2] ) );
  DFF \Reg_Bank/registers_reg[21][3]  ( .D(\Reg_Bank/n3673 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][3] ) );
  DFF \Reg_Bank/registers_reg[21][4]  ( .D(\Reg_Bank/n3674 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][4] ) );
  DFF \Reg_Bank/registers_reg[21][5]  ( .D(\Reg_Bank/n3675 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][5] ) );
  DFF \Reg_Bank/registers_reg[21][6]  ( .D(\Reg_Bank/n3676 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][6] ) );
  DFF \Reg_Bank/registers_reg[21][7]  ( .D(\Reg_Bank/n3677 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][7] ) );
  DFF \Reg_Bank/registers_reg[21][8]  ( .D(\Reg_Bank/n3678 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][8] ) );
  DFF \Reg_Bank/registers_reg[21][9]  ( .D(\Reg_Bank/n3679 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][9] ) );
  DFF \Reg_Bank/registers_reg[21][10]  ( .D(\Reg_Bank/n3680 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][10] ) );
  DFF \Reg_Bank/registers_reg[21][11]  ( .D(\Reg_Bank/n3681 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][11] ) );
  DFF \Reg_Bank/registers_reg[21][12]  ( .D(\Reg_Bank/n3682 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][12] ) );
  DFF \Reg_Bank/registers_reg[21][13]  ( .D(\Reg_Bank/n3683 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][13] ) );
  DFF \Reg_Bank/registers_reg[21][14]  ( .D(\Reg_Bank/n3684 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][14] ) );
  DFF \Reg_Bank/registers_reg[21][15]  ( .D(\Reg_Bank/n3685 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][15] ) );
  DFF \Reg_Bank/registers_reg[21][16]  ( .D(\Reg_Bank/n3686 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][16] ) );
  DFF \Reg_Bank/registers_reg[21][17]  ( .D(\Reg_Bank/n3687 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][17] ) );
  DFF \Reg_Bank/registers_reg[21][18]  ( .D(\Reg_Bank/n3688 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][18] ) );
  DFF \Reg_Bank/registers_reg[21][19]  ( .D(\Reg_Bank/n3689 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][19] ) );
  DFF \Reg_Bank/registers_reg[21][20]  ( .D(\Reg_Bank/n3690 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][20] ) );
  DFF \Reg_Bank/registers_reg[21][21]  ( .D(\Reg_Bank/n3691 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][21] ) );
  DFF \Reg_Bank/registers_reg[21][22]  ( .D(\Reg_Bank/n3692 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][22] ) );
  DFF \Reg_Bank/registers_reg[21][23]  ( .D(\Reg_Bank/n3693 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][23] ) );
  DFF \Reg_Bank/registers_reg[21][24]  ( .D(\Reg_Bank/n3694 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][24] ) );
  DFF \Reg_Bank/registers_reg[21][25]  ( .D(\Reg_Bank/n3695 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][25] ) );
  DFF \Reg_Bank/registers_reg[21][26]  ( .D(\Reg_Bank/n3696 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][26] ) );
  DFF \Reg_Bank/registers_reg[21][27]  ( .D(\Reg_Bank/n3697 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][27] ) );
  DFF \Reg_Bank/registers_reg[21][28]  ( .D(\Reg_Bank/n3698 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][28] ) );
  DFF \Reg_Bank/registers_reg[21][29]  ( .D(\Reg_Bank/n3699 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][29] ) );
  DFF \Reg_Bank/registers_reg[21][30]  ( .D(\Reg_Bank/n3700 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][30] ) );
  DFF \Reg_Bank/registers_reg[21][31]  ( .D(\Reg_Bank/n3701 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][31] ) );
  DFF \Reg_Bank/registers_reg[22][0]  ( .D(\Reg_Bank/n3702 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][0] ) );
  DFF \Reg_Bank/registers_reg[22][1]  ( .D(\Reg_Bank/n3703 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][1] ) );
  DFF \Reg_Bank/registers_reg[22][2]  ( .D(\Reg_Bank/n3704 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][2] ) );
  DFF \Reg_Bank/registers_reg[22][3]  ( .D(\Reg_Bank/n3705 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][3] ) );
  DFF \Reg_Bank/registers_reg[22][4]  ( .D(\Reg_Bank/n3706 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][4] ) );
  DFF \Reg_Bank/registers_reg[22][5]  ( .D(\Reg_Bank/n3707 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][5] ) );
  DFF \Reg_Bank/registers_reg[22][6]  ( .D(\Reg_Bank/n3708 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][6] ) );
  DFF \Reg_Bank/registers_reg[22][7]  ( .D(\Reg_Bank/n3709 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][7] ) );
  DFF \Reg_Bank/registers_reg[22][8]  ( .D(\Reg_Bank/n3710 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][8] ) );
  DFF \Reg_Bank/registers_reg[22][9]  ( .D(\Reg_Bank/n3711 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][9] ) );
  DFF \Reg_Bank/registers_reg[22][10]  ( .D(\Reg_Bank/n3712 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][10] ) );
  DFF \Reg_Bank/registers_reg[22][11]  ( .D(\Reg_Bank/n3713 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][11] ) );
  DFF \Reg_Bank/registers_reg[22][12]  ( .D(\Reg_Bank/n3714 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][12] ) );
  DFF \Reg_Bank/registers_reg[22][13]  ( .D(\Reg_Bank/n3715 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][13] ) );
  DFF \Reg_Bank/registers_reg[22][14]  ( .D(\Reg_Bank/n3716 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][14] ) );
  DFF \Reg_Bank/registers_reg[22][15]  ( .D(\Reg_Bank/n3717 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][15] ) );
  DFF \Reg_Bank/registers_reg[22][16]  ( .D(\Reg_Bank/n3718 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][16] ) );
  DFF \Reg_Bank/registers_reg[22][17]  ( .D(\Reg_Bank/n3719 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][17] ) );
  DFF \Reg_Bank/registers_reg[22][18]  ( .D(\Reg_Bank/n3720 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][18] ) );
  DFF \Reg_Bank/registers_reg[22][19]  ( .D(\Reg_Bank/n3721 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][19] ) );
  DFF \Reg_Bank/registers_reg[22][20]  ( .D(\Reg_Bank/n3722 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][20] ) );
  DFF \Reg_Bank/registers_reg[22][21]  ( .D(\Reg_Bank/n3723 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][21] ) );
  DFF \Reg_Bank/registers_reg[22][22]  ( .D(\Reg_Bank/n3724 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][22] ) );
  DFF \Reg_Bank/registers_reg[22][23]  ( .D(\Reg_Bank/n3725 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][23] ) );
  DFF \Reg_Bank/registers_reg[22][24]  ( .D(\Reg_Bank/n3726 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][24] ) );
  DFF \Reg_Bank/registers_reg[22][25]  ( .D(\Reg_Bank/n3727 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][25] ) );
  DFF \Reg_Bank/registers_reg[22][26]  ( .D(\Reg_Bank/n3728 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][26] ) );
  DFF \Reg_Bank/registers_reg[22][27]  ( .D(\Reg_Bank/n3729 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][27] ) );
  DFF \Reg_Bank/registers_reg[22][28]  ( .D(\Reg_Bank/n3730 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][28] ) );
  DFF \Reg_Bank/registers_reg[22][29]  ( .D(\Reg_Bank/n3731 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][29] ) );
  DFF \Reg_Bank/registers_reg[22][30]  ( .D(\Reg_Bank/n3732 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][30] ) );
  DFF \Reg_Bank/registers_reg[22][31]  ( .D(\Reg_Bank/n3733 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][31] ) );
  DFF \Reg_Bank/registers_reg[23][0]  ( .D(\Reg_Bank/n3734 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][0] ) );
  DFF \Reg_Bank/registers_reg[23][1]  ( .D(\Reg_Bank/n3735 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][1] ) );
  DFF \Reg_Bank/registers_reg[23][2]  ( .D(\Reg_Bank/n3736 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][2] ) );
  DFF \Reg_Bank/registers_reg[23][3]  ( .D(\Reg_Bank/n3737 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][3] ) );
  DFF \Reg_Bank/registers_reg[23][4]  ( .D(\Reg_Bank/n3738 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][4] ) );
  DFF \Reg_Bank/registers_reg[23][5]  ( .D(\Reg_Bank/n3739 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][5] ) );
  DFF \Reg_Bank/registers_reg[23][6]  ( .D(\Reg_Bank/n3740 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][6] ) );
  DFF \Reg_Bank/registers_reg[23][7]  ( .D(\Reg_Bank/n3741 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][7] ) );
  DFF \Reg_Bank/registers_reg[23][8]  ( .D(\Reg_Bank/n3742 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][8] ) );
  DFF \Reg_Bank/registers_reg[23][9]  ( .D(\Reg_Bank/n3743 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][9] ) );
  DFF \Reg_Bank/registers_reg[23][10]  ( .D(\Reg_Bank/n3744 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][10] ) );
  DFF \Reg_Bank/registers_reg[23][11]  ( .D(\Reg_Bank/n3745 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][11] ) );
  DFF \Reg_Bank/registers_reg[23][12]  ( .D(\Reg_Bank/n3746 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][12] ) );
  DFF \Reg_Bank/registers_reg[23][13]  ( .D(\Reg_Bank/n3747 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][13] ) );
  DFF \Reg_Bank/registers_reg[23][14]  ( .D(\Reg_Bank/n3748 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][14] ) );
  DFF \Reg_Bank/registers_reg[23][15]  ( .D(\Reg_Bank/n3749 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][15] ) );
  DFF \Reg_Bank/registers_reg[23][16]  ( .D(\Reg_Bank/n3750 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][16] ) );
  DFF \Reg_Bank/registers_reg[23][17]  ( .D(\Reg_Bank/n3751 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][17] ) );
  DFF \Reg_Bank/registers_reg[23][18]  ( .D(\Reg_Bank/n3752 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][18] ) );
  DFF \Reg_Bank/registers_reg[23][19]  ( .D(\Reg_Bank/n3753 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][19] ) );
  DFF \Reg_Bank/registers_reg[23][20]  ( .D(\Reg_Bank/n3754 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][20] ) );
  DFF \Reg_Bank/registers_reg[23][21]  ( .D(\Reg_Bank/n3755 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][21] ) );
  DFF \Reg_Bank/registers_reg[23][22]  ( .D(\Reg_Bank/n3756 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][22] ) );
  DFF \Reg_Bank/registers_reg[23][23]  ( .D(\Reg_Bank/n3757 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][23] ) );
  DFF \Reg_Bank/registers_reg[23][24]  ( .D(\Reg_Bank/n3758 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][24] ) );
  DFF \Reg_Bank/registers_reg[23][25]  ( .D(\Reg_Bank/n3759 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][25] ) );
  DFF \Reg_Bank/registers_reg[23][26]  ( .D(\Reg_Bank/n3760 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][26] ) );
  DFF \Reg_Bank/registers_reg[23][27]  ( .D(\Reg_Bank/n3761 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][27] ) );
  DFF \Reg_Bank/registers_reg[23][28]  ( .D(\Reg_Bank/n3762 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][28] ) );
  DFF \Reg_Bank/registers_reg[23][29]  ( .D(\Reg_Bank/n3763 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][29] ) );
  DFF \Reg_Bank/registers_reg[23][30]  ( .D(\Reg_Bank/n3764 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][30] ) );
  DFF \Reg_Bank/registers_reg[23][31]  ( .D(\Reg_Bank/n3765 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][31] ) );
  DFF \Reg_Bank/registers_reg[24][0]  ( .D(\Reg_Bank/n3766 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][0] ) );
  DFF \Reg_Bank/registers_reg[24][1]  ( .D(\Reg_Bank/n3767 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][1] ) );
  DFF \Reg_Bank/registers_reg[24][2]  ( .D(\Reg_Bank/n3768 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][2] ) );
  DFF \Reg_Bank/registers_reg[24][3]  ( .D(\Reg_Bank/n3769 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][3] ) );
  DFF \Reg_Bank/registers_reg[24][4]  ( .D(\Reg_Bank/n3770 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][4] ) );
  DFF \Reg_Bank/registers_reg[24][5]  ( .D(\Reg_Bank/n3771 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][5] ) );
  DFF \Reg_Bank/registers_reg[24][6]  ( .D(\Reg_Bank/n3772 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][6] ) );
  DFF \Reg_Bank/registers_reg[24][7]  ( .D(\Reg_Bank/n3773 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][7] ) );
  DFF \Reg_Bank/registers_reg[24][8]  ( .D(\Reg_Bank/n3774 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][8] ) );
  DFF \Reg_Bank/registers_reg[24][9]  ( .D(\Reg_Bank/n3775 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][9] ) );
  DFF \Reg_Bank/registers_reg[24][10]  ( .D(\Reg_Bank/n3776 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][10] ) );
  DFF \Reg_Bank/registers_reg[24][11]  ( .D(\Reg_Bank/n3777 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][11] ) );
  DFF \Reg_Bank/registers_reg[24][12]  ( .D(\Reg_Bank/n3778 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][12] ) );
  DFF \Reg_Bank/registers_reg[24][13]  ( .D(\Reg_Bank/n3779 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][13] ) );
  DFF \Reg_Bank/registers_reg[24][14]  ( .D(\Reg_Bank/n3780 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][14] ) );
  DFF \Reg_Bank/registers_reg[24][15]  ( .D(\Reg_Bank/n3781 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][15] ) );
  DFF \Reg_Bank/registers_reg[24][16]  ( .D(\Reg_Bank/n3782 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][16] ) );
  DFF \Reg_Bank/registers_reg[24][17]  ( .D(\Reg_Bank/n3783 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][17] ) );
  DFF \Reg_Bank/registers_reg[24][18]  ( .D(\Reg_Bank/n3784 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][18] ) );
  DFF \Reg_Bank/registers_reg[24][19]  ( .D(\Reg_Bank/n3785 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][19] ) );
  DFF \Reg_Bank/registers_reg[24][20]  ( .D(\Reg_Bank/n3786 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][20] ) );
  DFF \Reg_Bank/registers_reg[24][21]  ( .D(\Reg_Bank/n3787 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][21] ) );
  DFF \Reg_Bank/registers_reg[24][22]  ( .D(\Reg_Bank/n3788 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][22] ) );
  DFF \Reg_Bank/registers_reg[24][23]  ( .D(\Reg_Bank/n3789 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][23] ) );
  DFF \Reg_Bank/registers_reg[24][24]  ( .D(\Reg_Bank/n3790 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][24] ) );
  DFF \Reg_Bank/registers_reg[24][25]  ( .D(\Reg_Bank/n3791 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][25] ) );
  DFF \Reg_Bank/registers_reg[24][26]  ( .D(\Reg_Bank/n3792 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][26] ) );
  DFF \Reg_Bank/registers_reg[24][27]  ( .D(\Reg_Bank/n3793 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][27] ) );
  DFF \Reg_Bank/registers_reg[24][28]  ( .D(\Reg_Bank/n3794 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][28] ) );
  DFF \Reg_Bank/registers_reg[24][29]  ( .D(\Reg_Bank/n3795 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][29] ) );
  DFF \Reg_Bank/registers_reg[24][30]  ( .D(\Reg_Bank/n3796 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][30] ) );
  DFF \Reg_Bank/registers_reg[24][31]  ( .D(\Reg_Bank/n3797 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][31] ) );
  DFF \Reg_Bank/registers_reg[25][0]  ( .D(\Reg_Bank/n3798 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][0] ) );
  DFF \Reg_Bank/registers_reg[25][1]  ( .D(\Reg_Bank/n3799 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][1] ) );
  DFF \Reg_Bank/registers_reg[25][2]  ( .D(\Reg_Bank/n3800 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][2] ) );
  DFF \Reg_Bank/registers_reg[25][3]  ( .D(\Reg_Bank/n3801 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][3] ) );
  DFF \Reg_Bank/registers_reg[25][4]  ( .D(\Reg_Bank/n3802 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][4] ) );
  DFF \Reg_Bank/registers_reg[25][5]  ( .D(\Reg_Bank/n3803 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][5] ) );
  DFF \Reg_Bank/registers_reg[25][6]  ( .D(\Reg_Bank/n3804 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][6] ) );
  DFF \Reg_Bank/registers_reg[25][7]  ( .D(\Reg_Bank/n3805 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][7] ) );
  DFF \Reg_Bank/registers_reg[25][8]  ( .D(\Reg_Bank/n3806 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][8] ) );
  DFF \Reg_Bank/registers_reg[25][9]  ( .D(\Reg_Bank/n3807 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][9] ) );
  DFF \Reg_Bank/registers_reg[25][10]  ( .D(\Reg_Bank/n3808 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][10] ) );
  DFF \Reg_Bank/registers_reg[25][11]  ( .D(\Reg_Bank/n3809 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][11] ) );
  DFF \Reg_Bank/registers_reg[25][12]  ( .D(\Reg_Bank/n3810 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][12] ) );
  DFF \Reg_Bank/registers_reg[25][13]  ( .D(\Reg_Bank/n3811 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][13] ) );
  DFF \Reg_Bank/registers_reg[25][14]  ( .D(\Reg_Bank/n3812 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][14] ) );
  DFF \Reg_Bank/registers_reg[25][15]  ( .D(\Reg_Bank/n3813 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][15] ) );
  DFF \Reg_Bank/registers_reg[25][16]  ( .D(\Reg_Bank/n3814 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][16] ) );
  DFF \Reg_Bank/registers_reg[25][17]  ( .D(\Reg_Bank/n3815 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][17] ) );
  DFF \Reg_Bank/registers_reg[25][18]  ( .D(\Reg_Bank/n3816 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][18] ) );
  DFF \Reg_Bank/registers_reg[25][19]  ( .D(\Reg_Bank/n3817 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][19] ) );
  DFF \Reg_Bank/registers_reg[25][20]  ( .D(\Reg_Bank/n3818 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][20] ) );
  DFF \Reg_Bank/registers_reg[25][21]  ( .D(\Reg_Bank/n3819 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][21] ) );
  DFF \Reg_Bank/registers_reg[25][22]  ( .D(\Reg_Bank/n3820 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][22] ) );
  DFF \Reg_Bank/registers_reg[25][23]  ( .D(\Reg_Bank/n3821 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][23] ) );
  DFF \Reg_Bank/registers_reg[25][24]  ( .D(\Reg_Bank/n3822 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][24] ) );
  DFF \Reg_Bank/registers_reg[25][25]  ( .D(\Reg_Bank/n3823 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][25] ) );
  DFF \Reg_Bank/registers_reg[25][26]  ( .D(\Reg_Bank/n3824 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][26] ) );
  DFF \Reg_Bank/registers_reg[25][27]  ( .D(\Reg_Bank/n3825 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][27] ) );
  DFF \Reg_Bank/registers_reg[25][28]  ( .D(\Reg_Bank/n3826 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][28] ) );
  DFF \Reg_Bank/registers_reg[25][29]  ( .D(\Reg_Bank/n3827 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][29] ) );
  DFF \Reg_Bank/registers_reg[25][30]  ( .D(\Reg_Bank/n3828 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][30] ) );
  DFF \Reg_Bank/registers_reg[25][31]  ( .D(\Reg_Bank/n3829 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][31] ) );
  DFF \Reg_Bank/registers_reg[26][0]  ( .D(\Reg_Bank/n3830 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][0] ) );
  DFF \Reg_Bank/registers_reg[26][1]  ( .D(\Reg_Bank/n3831 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][1] ) );
  DFF \Reg_Bank/registers_reg[26][2]  ( .D(\Reg_Bank/n3832 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][2] ) );
  DFF \Reg_Bank/registers_reg[26][3]  ( .D(\Reg_Bank/n3833 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][3] ) );
  DFF \Reg_Bank/registers_reg[26][4]  ( .D(\Reg_Bank/n3834 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][4] ) );
  DFF \Reg_Bank/registers_reg[26][5]  ( .D(\Reg_Bank/n3835 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][5] ) );
  DFF \Reg_Bank/registers_reg[26][6]  ( .D(\Reg_Bank/n3836 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][6] ) );
  DFF \Reg_Bank/registers_reg[26][7]  ( .D(\Reg_Bank/n3837 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][7] ) );
  DFF \Reg_Bank/registers_reg[26][8]  ( .D(\Reg_Bank/n3838 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][8] ) );
  DFF \Reg_Bank/registers_reg[26][9]  ( .D(\Reg_Bank/n3839 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][9] ) );
  DFF \Reg_Bank/registers_reg[26][10]  ( .D(\Reg_Bank/n3840 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][10] ) );
  DFF \Reg_Bank/registers_reg[26][11]  ( .D(\Reg_Bank/n3841 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][11] ) );
  DFF \Reg_Bank/registers_reg[26][12]  ( .D(\Reg_Bank/n3842 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][12] ) );
  DFF \Reg_Bank/registers_reg[26][13]  ( .D(\Reg_Bank/n3843 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][13] ) );
  DFF \Reg_Bank/registers_reg[26][14]  ( .D(\Reg_Bank/n3844 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][14] ) );
  DFF \Reg_Bank/registers_reg[26][15]  ( .D(\Reg_Bank/n3845 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][15] ) );
  DFF \Reg_Bank/registers_reg[26][16]  ( .D(\Reg_Bank/n3846 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][16] ) );
  DFF \Reg_Bank/registers_reg[26][17]  ( .D(\Reg_Bank/n3847 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][17] ) );
  DFF \Reg_Bank/registers_reg[26][18]  ( .D(\Reg_Bank/n3848 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][18] ) );
  DFF \Reg_Bank/registers_reg[26][19]  ( .D(\Reg_Bank/n3849 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][19] ) );
  DFF \Reg_Bank/registers_reg[26][20]  ( .D(\Reg_Bank/n3850 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][20] ) );
  DFF \Reg_Bank/registers_reg[26][21]  ( .D(\Reg_Bank/n3851 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][21] ) );
  DFF \Reg_Bank/registers_reg[26][22]  ( .D(\Reg_Bank/n3852 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][22] ) );
  DFF \Reg_Bank/registers_reg[26][23]  ( .D(\Reg_Bank/n3853 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][23] ) );
  DFF \Reg_Bank/registers_reg[26][24]  ( .D(\Reg_Bank/n3854 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][24] ) );
  DFF \Reg_Bank/registers_reg[26][25]  ( .D(\Reg_Bank/n3855 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][25] ) );
  DFF \Reg_Bank/registers_reg[26][26]  ( .D(\Reg_Bank/n3856 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][26] ) );
  DFF \Reg_Bank/registers_reg[26][27]  ( .D(\Reg_Bank/n3857 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][27] ) );
  DFF \Reg_Bank/registers_reg[26][28]  ( .D(\Reg_Bank/n3858 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][28] ) );
  DFF \Reg_Bank/registers_reg[26][29]  ( .D(\Reg_Bank/n3859 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][29] ) );
  DFF \Reg_Bank/registers_reg[26][30]  ( .D(\Reg_Bank/n3860 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][30] ) );
  DFF \Reg_Bank/registers_reg[26][31]  ( .D(\Reg_Bank/n3861 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][31] ) );
  DFF \Reg_Bank/registers_reg[27][0]  ( .D(\Reg_Bank/n3862 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][0] ) );
  DFF \Reg_Bank/registers_reg[27][1]  ( .D(\Reg_Bank/n3863 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][1] ) );
  DFF \Reg_Bank/registers_reg[27][2]  ( .D(\Reg_Bank/n3864 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][2] ) );
  DFF \Reg_Bank/registers_reg[27][3]  ( .D(\Reg_Bank/n3865 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][3] ) );
  DFF \Reg_Bank/registers_reg[27][4]  ( .D(\Reg_Bank/n3866 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][4] ) );
  DFF \Reg_Bank/registers_reg[27][5]  ( .D(\Reg_Bank/n3867 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][5] ) );
  DFF \Reg_Bank/registers_reg[27][6]  ( .D(\Reg_Bank/n3868 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][6] ) );
  DFF \Reg_Bank/registers_reg[27][7]  ( .D(\Reg_Bank/n3869 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][7] ) );
  DFF \Reg_Bank/registers_reg[27][8]  ( .D(\Reg_Bank/n3870 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][8] ) );
  DFF \Reg_Bank/registers_reg[27][9]  ( .D(\Reg_Bank/n3871 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][9] ) );
  DFF \Reg_Bank/registers_reg[27][10]  ( .D(\Reg_Bank/n3872 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][10] ) );
  DFF \Reg_Bank/registers_reg[27][11]  ( .D(\Reg_Bank/n3873 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][11] ) );
  DFF \Reg_Bank/registers_reg[27][12]  ( .D(\Reg_Bank/n3874 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][12] ) );
  DFF \Reg_Bank/registers_reg[27][13]  ( .D(\Reg_Bank/n3875 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][13] ) );
  DFF \Reg_Bank/registers_reg[27][14]  ( .D(\Reg_Bank/n3876 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][14] ) );
  DFF \Reg_Bank/registers_reg[27][15]  ( .D(\Reg_Bank/n3877 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][15] ) );
  DFF \Reg_Bank/registers_reg[27][16]  ( .D(\Reg_Bank/n3878 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][16] ) );
  DFF \Reg_Bank/registers_reg[27][17]  ( .D(\Reg_Bank/n3879 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][17] ) );
  DFF \Reg_Bank/registers_reg[27][18]  ( .D(\Reg_Bank/n3880 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][18] ) );
  DFF \Reg_Bank/registers_reg[27][19]  ( .D(\Reg_Bank/n3881 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][19] ) );
  DFF \Reg_Bank/registers_reg[27][20]  ( .D(\Reg_Bank/n3882 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][20] ) );
  DFF \Reg_Bank/registers_reg[27][21]  ( .D(\Reg_Bank/n3883 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][21] ) );
  DFF \Reg_Bank/registers_reg[27][22]  ( .D(\Reg_Bank/n3884 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][22] ) );
  DFF \Reg_Bank/registers_reg[27][23]  ( .D(\Reg_Bank/n3885 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][23] ) );
  DFF \Reg_Bank/registers_reg[27][24]  ( .D(\Reg_Bank/n3886 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][24] ) );
  DFF \Reg_Bank/registers_reg[27][25]  ( .D(\Reg_Bank/n3887 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][25] ) );
  DFF \Reg_Bank/registers_reg[27][26]  ( .D(\Reg_Bank/n3888 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][26] ) );
  DFF \Reg_Bank/registers_reg[27][27]  ( .D(\Reg_Bank/n3889 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][27] ) );
  DFF \Reg_Bank/registers_reg[27][28]  ( .D(\Reg_Bank/n3890 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][28] ) );
  DFF \Reg_Bank/registers_reg[27][29]  ( .D(\Reg_Bank/n3891 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][29] ) );
  DFF \Reg_Bank/registers_reg[27][30]  ( .D(\Reg_Bank/n3892 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][30] ) );
  DFF \Reg_Bank/registers_reg[27][31]  ( .D(\Reg_Bank/n3893 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][31] ) );
  DFF \Reg_Bank/registers_reg[28][0]  ( .D(\Reg_Bank/n3894 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][0] ) );
  DFF \Reg_Bank/registers_reg[28][1]  ( .D(\Reg_Bank/n3895 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][1] ) );
  DFF \Reg_Bank/registers_reg[28][2]  ( .D(\Reg_Bank/n3896 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][2] ) );
  DFF \Reg_Bank/registers_reg[28][3]  ( .D(\Reg_Bank/n3897 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][3] ) );
  DFF \Reg_Bank/registers_reg[28][4]  ( .D(\Reg_Bank/n3898 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][4] ) );
  DFF \Reg_Bank/registers_reg[28][5]  ( .D(\Reg_Bank/n3899 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][5] ) );
  DFF \Reg_Bank/registers_reg[28][6]  ( .D(\Reg_Bank/n3900 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][6] ) );
  DFF \Reg_Bank/registers_reg[28][7]  ( .D(\Reg_Bank/n3901 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][7] ) );
  DFF \Reg_Bank/registers_reg[28][8]  ( .D(\Reg_Bank/n3902 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][8] ) );
  DFF \Reg_Bank/registers_reg[28][9]  ( .D(\Reg_Bank/n3903 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][9] ) );
  DFF \Reg_Bank/registers_reg[28][10]  ( .D(\Reg_Bank/n3904 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][10] ) );
  DFF \Reg_Bank/registers_reg[28][11]  ( .D(\Reg_Bank/n3905 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][11] ) );
  DFF \Reg_Bank/registers_reg[28][12]  ( .D(\Reg_Bank/n3906 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][12] ) );
  DFF \Reg_Bank/registers_reg[28][13]  ( .D(\Reg_Bank/n3907 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][13] ) );
  DFF \Reg_Bank/registers_reg[28][14]  ( .D(\Reg_Bank/n3908 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][14] ) );
  DFF \Reg_Bank/registers_reg[28][15]  ( .D(\Reg_Bank/n3909 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][15] ) );
  DFF \Reg_Bank/registers_reg[28][16]  ( .D(\Reg_Bank/n3910 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][16] ) );
  DFF \Reg_Bank/registers_reg[28][17]  ( .D(\Reg_Bank/n3911 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][17] ) );
  DFF \Reg_Bank/registers_reg[28][18]  ( .D(\Reg_Bank/n3912 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][18] ) );
  DFF \Reg_Bank/registers_reg[28][19]  ( .D(\Reg_Bank/n3913 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][19] ) );
  DFF \Reg_Bank/registers_reg[28][20]  ( .D(\Reg_Bank/n3914 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][20] ) );
  DFF \Reg_Bank/registers_reg[28][21]  ( .D(\Reg_Bank/n3915 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][21] ) );
  DFF \Reg_Bank/registers_reg[28][22]  ( .D(\Reg_Bank/n3916 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][22] ) );
  DFF \Reg_Bank/registers_reg[28][23]  ( .D(\Reg_Bank/n3917 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][23] ) );
  DFF \Reg_Bank/registers_reg[28][24]  ( .D(\Reg_Bank/n3918 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][24] ) );
  DFF \Reg_Bank/registers_reg[28][25]  ( .D(\Reg_Bank/n3919 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][25] ) );
  DFF \Reg_Bank/registers_reg[28][26]  ( .D(\Reg_Bank/n3920 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][26] ) );
  DFF \Reg_Bank/registers_reg[28][27]  ( .D(\Reg_Bank/n3921 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][27] ) );
  DFF \Reg_Bank/registers_reg[28][28]  ( .D(\Reg_Bank/n3922 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][28] ) );
  DFF \Reg_Bank/registers_reg[28][29]  ( .D(\Reg_Bank/n3923 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][29] ) );
  DFF \Reg_Bank/registers_reg[28][30]  ( .D(\Reg_Bank/n3924 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][30] ) );
  DFF \Reg_Bank/registers_reg[28][31]  ( .D(\Reg_Bank/n3925 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][31] ) );
  DFF \Reg_Bank/registers_reg[29][0]  ( .D(\Reg_Bank/n3926 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][0] ) );
  DFF \Reg_Bank/registers_reg[29][1]  ( .D(\Reg_Bank/n3927 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][1] ) );
  DFF \Reg_Bank/registers_reg[29][2]  ( .D(\Reg_Bank/n3928 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][2] ) );
  DFF \Reg_Bank/registers_reg[29][3]  ( .D(\Reg_Bank/n3929 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][3] ) );
  DFF \Reg_Bank/registers_reg[29][4]  ( .D(\Reg_Bank/n3930 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][4] ) );
  DFF \Reg_Bank/registers_reg[29][5]  ( .D(\Reg_Bank/n3931 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][5] ) );
  DFF \Reg_Bank/registers_reg[29][6]  ( .D(\Reg_Bank/n3932 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][6] ) );
  DFF \Reg_Bank/registers_reg[29][7]  ( .D(\Reg_Bank/n3933 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][7] ) );
  DFF \Reg_Bank/registers_reg[29][8]  ( .D(\Reg_Bank/n3934 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][8] ) );
  DFF \Reg_Bank/registers_reg[29][9]  ( .D(\Reg_Bank/n3935 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][9] ) );
  DFF \Reg_Bank/registers_reg[29][10]  ( .D(\Reg_Bank/n3936 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][10] ) );
  DFF \Reg_Bank/registers_reg[29][11]  ( .D(\Reg_Bank/n3937 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][11] ) );
  DFF \Reg_Bank/registers_reg[29][12]  ( .D(\Reg_Bank/n3938 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][12] ) );
  DFF \Reg_Bank/registers_reg[29][13]  ( .D(\Reg_Bank/n3939 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][13] ) );
  DFF \Reg_Bank/registers_reg[29][14]  ( .D(\Reg_Bank/n3940 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][14] ) );
  DFF \Reg_Bank/registers_reg[29][15]  ( .D(\Reg_Bank/n3941 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][15] ) );
  DFF \Reg_Bank/registers_reg[29][16]  ( .D(\Reg_Bank/n3942 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][16] ) );
  DFF \Reg_Bank/registers_reg[29][17]  ( .D(\Reg_Bank/n3943 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][17] ) );
  DFF \Reg_Bank/registers_reg[29][18]  ( .D(\Reg_Bank/n3944 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][18] ) );
  DFF \Reg_Bank/registers_reg[29][19]  ( .D(\Reg_Bank/n3945 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][19] ) );
  DFF \Reg_Bank/registers_reg[29][20]  ( .D(\Reg_Bank/n3946 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][20] ) );
  DFF \Reg_Bank/registers_reg[29][21]  ( .D(\Reg_Bank/n3947 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][21] ) );
  DFF \Reg_Bank/registers_reg[29][22]  ( .D(\Reg_Bank/n3948 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][22] ) );
  DFF \Reg_Bank/registers_reg[29][23]  ( .D(\Reg_Bank/n3949 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][23] ) );
  DFF \Reg_Bank/registers_reg[29][24]  ( .D(\Reg_Bank/n3950 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][24] ) );
  DFF \Reg_Bank/registers_reg[29][25]  ( .D(\Reg_Bank/n3951 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][25] ) );
  DFF \Reg_Bank/registers_reg[29][26]  ( .D(\Reg_Bank/n3952 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][26] ) );
  DFF \Reg_Bank/registers_reg[29][27]  ( .D(\Reg_Bank/n3953 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][27] ) );
  DFF \Reg_Bank/registers_reg[29][28]  ( .D(\Reg_Bank/n3954 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][28] ) );
  DFF \Reg_Bank/registers_reg[29][29]  ( .D(\Reg_Bank/n3955 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][29] ) );
  DFF \Reg_Bank/registers_reg[29][30]  ( .D(\Reg_Bank/n3956 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][30] ) );
  DFF \Reg_Bank/registers_reg[29][31]  ( .D(\Reg_Bank/n3957 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][31] ) );
  DFF \Reg_Bank/registers_reg[30][0]  ( .D(\Reg_Bank/n3958 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][0] ) );
  DFF \Reg_Bank/registers_reg[30][1]  ( .D(\Reg_Bank/n3959 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][1] ) );
  DFF \Reg_Bank/registers_reg[30][2]  ( .D(\Reg_Bank/n3960 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][2] ) );
  DFF \Reg_Bank/registers_reg[30][3]  ( .D(\Reg_Bank/n3961 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][3] ) );
  DFF \Reg_Bank/registers_reg[30][4]  ( .D(\Reg_Bank/n3962 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][4] ) );
  DFF \Reg_Bank/registers_reg[30][5]  ( .D(\Reg_Bank/n3963 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][5] ) );
  DFF \Reg_Bank/registers_reg[30][6]  ( .D(\Reg_Bank/n3964 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][6] ) );
  DFF \Reg_Bank/registers_reg[30][7]  ( .D(\Reg_Bank/n3965 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][7] ) );
  DFF \Reg_Bank/registers_reg[30][8]  ( .D(\Reg_Bank/n3966 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][8] ) );
  DFF \Reg_Bank/registers_reg[30][9]  ( .D(\Reg_Bank/n3967 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][9] ) );
  DFF \Reg_Bank/registers_reg[30][10]  ( .D(\Reg_Bank/n3968 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][10] ) );
  DFF \Reg_Bank/registers_reg[30][11]  ( .D(\Reg_Bank/n3969 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][11] ) );
  DFF \Reg_Bank/registers_reg[30][12]  ( .D(\Reg_Bank/n3970 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][12] ) );
  DFF \Reg_Bank/registers_reg[30][13]  ( .D(\Reg_Bank/n3971 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][13] ) );
  DFF \Reg_Bank/registers_reg[30][14]  ( .D(\Reg_Bank/n3972 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][14] ) );
  DFF \Reg_Bank/registers_reg[30][15]  ( .D(\Reg_Bank/n3973 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][15] ) );
  DFF \Reg_Bank/registers_reg[30][16]  ( .D(\Reg_Bank/n3974 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][16] ) );
  DFF \Reg_Bank/registers_reg[30][17]  ( .D(\Reg_Bank/n3975 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][17] ) );
  DFF \Reg_Bank/registers_reg[30][18]  ( .D(\Reg_Bank/n3976 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][18] ) );
  DFF \Reg_Bank/registers_reg[30][19]  ( .D(\Reg_Bank/n3977 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][19] ) );
  DFF \Reg_Bank/registers_reg[30][20]  ( .D(\Reg_Bank/n3978 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][20] ) );
  DFF \Reg_Bank/registers_reg[30][21]  ( .D(\Reg_Bank/n3979 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][21] ) );
  DFF \Reg_Bank/registers_reg[30][22]  ( .D(\Reg_Bank/n3980 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][22] ) );
  DFF \Reg_Bank/registers_reg[30][23]  ( .D(\Reg_Bank/n3981 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][23] ) );
  DFF \Reg_Bank/registers_reg[30][24]  ( .D(\Reg_Bank/n3982 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][24] ) );
  DFF \Reg_Bank/registers_reg[30][25]  ( .D(\Reg_Bank/n3983 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][25] ) );
  DFF \Reg_Bank/registers_reg[30][26]  ( .D(\Reg_Bank/n3984 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][26] ) );
  DFF \Reg_Bank/registers_reg[30][27]  ( .D(\Reg_Bank/n3985 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][27] ) );
  DFF \Reg_Bank/registers_reg[30][28]  ( .D(\Reg_Bank/n3986 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][28] ) );
  DFF \Reg_Bank/registers_reg[30][29]  ( .D(\Reg_Bank/n3987 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][29] ) );
  DFF \Reg_Bank/registers_reg[30][30]  ( .D(\Reg_Bank/n3988 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][30] ) );
  DFF \Reg_Bank/registers_reg[30][31]  ( .D(\Reg_Bank/n3989 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][31] ) );
  DFF \Reg_Bank/registers_reg[31][0]  ( .D(\Reg_Bank/n3990 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][0] ) );
  DFF \Reg_Bank/registers_reg[31][1]  ( .D(\Reg_Bank/n3991 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][1] ) );
  DFF \Reg_Bank/registers_reg[31][2]  ( .D(\Reg_Bank/n3992 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][2] ) );
  DFF \Reg_Bank/registers_reg[31][3]  ( .D(\Reg_Bank/n3993 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][3] ) );
  DFF \Reg_Bank/registers_reg[31][4]  ( .D(\Reg_Bank/n3994 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][4] ) );
  DFF \Reg_Bank/registers_reg[31][5]  ( .D(\Reg_Bank/n3995 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][5] ) );
  DFF \Reg_Bank/registers_reg[31][6]  ( .D(\Reg_Bank/n3996 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][6] ) );
  DFF \Reg_Bank/registers_reg[31][7]  ( .D(\Reg_Bank/n3997 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][7] ) );
  DFF \Reg_Bank/registers_reg[31][8]  ( .D(\Reg_Bank/n3998 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][8] ) );
  DFF \Reg_Bank/registers_reg[31][9]  ( .D(\Reg_Bank/n3999 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][9] ) );
  DFF \Reg_Bank/registers_reg[31][10]  ( .D(\Reg_Bank/n4000 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][10] ) );
  DFF \Reg_Bank/registers_reg[31][11]  ( .D(\Reg_Bank/n4001 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][11] ) );
  DFF \Reg_Bank/registers_reg[31][12]  ( .D(\Reg_Bank/n4002 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][12] ) );
  DFF \Reg_Bank/registers_reg[31][13]  ( .D(\Reg_Bank/n4003 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][13] ) );
  DFF \Reg_Bank/registers_reg[31][14]  ( .D(\Reg_Bank/n4004 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][14] ) );
  DFF \Reg_Bank/registers_reg[31][15]  ( .D(\Reg_Bank/n4005 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][15] ) );
  DFF \Reg_Bank/registers_reg[31][16]  ( .D(\Reg_Bank/n4006 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][16] ) );
  DFF \Reg_Bank/registers_reg[31][17]  ( .D(\Reg_Bank/n4007 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][17] ) );
  DFF \Reg_Bank/registers_reg[31][18]  ( .D(\Reg_Bank/n4008 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][18] ) );
  DFF \Reg_Bank/registers_reg[31][19]  ( .D(\Reg_Bank/n4009 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][19] ) );
  DFF \Reg_Bank/registers_reg[31][20]  ( .D(\Reg_Bank/n4010 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][20] ) );
  DFF \Reg_Bank/registers_reg[31][21]  ( .D(\Reg_Bank/n4011 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][21] ) );
  DFF \Reg_Bank/registers_reg[31][22]  ( .D(\Reg_Bank/n4012 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][22] ) );
  DFF \Reg_Bank/registers_reg[31][23]  ( .D(\Reg_Bank/n4013 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][23] ) );
  DFF \Reg_Bank/registers_reg[31][24]  ( .D(\Reg_Bank/n4014 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][24] ) );
  DFF \Reg_Bank/registers_reg[31][25]  ( .D(\Reg_Bank/n4015 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][25] ) );
  DFF \Reg_Bank/registers_reg[31][26]  ( .D(\Reg_Bank/n4016 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][26] ) );
  DFF \Reg_Bank/registers_reg[31][27]  ( .D(\Reg_Bank/n4017 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][27] ) );
  DFF \Reg_Bank/registers_reg[31][28]  ( .D(\Reg_Bank/n4018 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][28] ) );
  DFF \Reg_Bank/registers_reg[31][29]  ( .D(\Reg_Bank/n4019 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][29] ) );
  DFF \Reg_Bank/registers_reg[31][30]  ( .D(\Reg_Bank/n4020 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][30] ) );
  DFF \Reg_Bank/registers_reg[31][31]  ( .D(\Reg_Bank/n4021 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][31] ) );
  MUX \Shifter/sll_27/M1_0_1  ( .A(b_bus[1]), .B(b_bus[0]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][1] ) );
  MUX \Shifter/sll_27/M1_0_2  ( .A(b_bus[2]), .B(b_bus[1]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][2] ) );
  MUX \Shifter/sll_27/M1_0_3  ( .A(b_bus[3]), .B(b_bus[2]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][3] ) );
  MUX \Shifter/sll_27/M1_0_4  ( .A(b_bus[4]), .B(b_bus[3]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][4] ) );
  MUX \Shifter/sll_27/M1_0_5  ( .A(b_bus[5]), .B(b_bus[4]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][5] ) );
  MUX \Shifter/sll_27/M1_0_6  ( .A(b_bus[6]), .B(b_bus[5]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][6] ) );
  MUX \Shifter/sll_27/M1_0_7  ( .A(b_bus[7]), .B(b_bus[6]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][7] ) );
  MUX \Shifter/sll_27/M1_0_8  ( .A(b_bus[8]), .B(b_bus[7]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][8] ) );
  MUX \Shifter/sll_27/M1_0_9  ( .A(b_bus[9]), .B(b_bus[8]), .S(a_bus[0]), .Z(
        \Shifter/sll_27/ML_int[1][9] ) );
  MUX \Shifter/sll_27/M1_0_10  ( .A(b_bus[10]), .B(b_bus[9]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][10] ) );
  MUX \Shifter/sll_27/M1_0_11  ( .A(b_bus[11]), .B(b_bus[10]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][11] ) );
  MUX \Shifter/sll_27/M1_0_12  ( .A(b_bus[12]), .B(b_bus[11]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][12] ) );
  MUX \Shifter/sll_27/M1_0_13  ( .A(b_bus[13]), .B(b_bus[12]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][13] ) );
  MUX \Shifter/sll_27/M1_0_14  ( .A(b_bus[14]), .B(b_bus[13]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][14] ) );
  MUX \Shifter/sll_27/M1_0_15  ( .A(b_bus[15]), .B(b_bus[14]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][15] ) );
  MUX \Shifter/sll_27/M1_0_16  ( .A(b_bus[16]), .B(b_bus[15]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][16] ) );
  MUX \Shifter/sll_27/M1_0_17  ( .A(b_bus[17]), .B(b_bus[16]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][17] ) );
  MUX \Shifter/sll_27/M1_0_18  ( .A(b_bus[18]), .B(b_bus[17]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][18] ) );
  MUX \Shifter/sll_27/M1_0_19  ( .A(b_bus[19]), .B(b_bus[18]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][19] ) );
  MUX \Shifter/sll_27/M1_0_20  ( .A(b_bus[20]), .B(b_bus[19]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][20] ) );
  MUX \Shifter/sll_27/M1_0_21  ( .A(b_bus[21]), .B(b_bus[20]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][21] ) );
  MUX \Shifter/sll_27/M1_0_22  ( .A(b_bus[22]), .B(b_bus[21]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][22] ) );
  MUX \Shifter/sll_27/M1_0_23  ( .A(b_bus[23]), .B(b_bus[22]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][23] ) );
  MUX \Shifter/sll_27/M1_0_24  ( .A(b_bus[24]), .B(b_bus[23]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][24] ) );
  MUX \Shifter/sll_27/M1_0_25  ( .A(b_bus[25]), .B(b_bus[24]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][25] ) );
  MUX \Shifter/sll_27/M1_0_26  ( .A(b_bus[26]), .B(b_bus[25]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][26] ) );
  MUX \Shifter/sll_27/M1_0_27  ( .A(b_bus[27]), .B(b_bus[26]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][27] ) );
  MUX \Shifter/sll_27/M1_0_28  ( .A(b_bus[28]), .B(b_bus[27]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][28] ) );
  MUX \Shifter/sll_27/M1_0_29  ( .A(b_bus[29]), .B(b_bus[28]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][29] ) );
  MUX \Shifter/sll_27/M1_0_30  ( .A(b_bus[30]), .B(b_bus[29]), .S(a_bus[0]), 
        .Z(\Shifter/sll_27/ML_int[1][30] ) );
  MUX \Shifter/sll_27/M1_0_31  ( .A(\Shifter/N75 ), .B(b_bus[30]), .S(a_bus[0]), .Z(\Shifter/sll_27/ML_int[1][31] ) );
  MUX \Shifter/sll_27/M1_1_2  ( .A(\Shifter/sll_27/ML_int[1][2] ), .B(
        \Shifter/sll_27/ML_int[1][0] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][2] ) );
  MUX \Shifter/sll_27/M1_1_3  ( .A(\Shifter/sll_27/ML_int[1][3] ), .B(
        \Shifter/sll_27/ML_int[1][1] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][3] ) );
  MUX \Shifter/sll_27/M1_1_4  ( .A(\Shifter/sll_27/ML_int[1][4] ), .B(
        \Shifter/sll_27/ML_int[1][2] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][4] ) );
  MUX \Shifter/sll_27/M1_1_5  ( .A(\Shifter/sll_27/ML_int[1][5] ), .B(
        \Shifter/sll_27/ML_int[1][3] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][5] ) );
  MUX \Shifter/sll_27/M1_1_6  ( .A(\Shifter/sll_27/ML_int[1][6] ), .B(
        \Shifter/sll_27/ML_int[1][4] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][6] ) );
  MUX \Shifter/sll_27/M1_1_7  ( .A(\Shifter/sll_27/ML_int[1][7] ), .B(
        \Shifter/sll_27/ML_int[1][5] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][7] ) );
  MUX \Shifter/sll_27/M1_1_8  ( .A(\Shifter/sll_27/ML_int[1][8] ), .B(
        \Shifter/sll_27/ML_int[1][6] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][8] ) );
  MUX \Shifter/sll_27/M1_1_9  ( .A(\Shifter/sll_27/ML_int[1][9] ), .B(
        \Shifter/sll_27/ML_int[1][7] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][9] ) );
  MUX \Shifter/sll_27/M1_1_10  ( .A(\Shifter/sll_27/ML_int[1][10] ), .B(
        \Shifter/sll_27/ML_int[1][8] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][10] ) );
  MUX \Shifter/sll_27/M1_1_11  ( .A(\Shifter/sll_27/ML_int[1][11] ), .B(
        \Shifter/sll_27/ML_int[1][9] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][11] ) );
  MUX \Shifter/sll_27/M1_1_12  ( .A(\Shifter/sll_27/ML_int[1][12] ), .B(
        \Shifter/sll_27/ML_int[1][10] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][12] ) );
  MUX \Shifter/sll_27/M1_1_13  ( .A(\Shifter/sll_27/ML_int[1][13] ), .B(
        \Shifter/sll_27/ML_int[1][11] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][13] ) );
  MUX \Shifter/sll_27/M1_1_14  ( .A(\Shifter/sll_27/ML_int[1][14] ), .B(
        \Shifter/sll_27/ML_int[1][12] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][14] ) );
  MUX \Shifter/sll_27/M1_1_15  ( .A(\Shifter/sll_27/ML_int[1][15] ), .B(
        \Shifter/sll_27/ML_int[1][13] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][15] ) );
  MUX \Shifter/sll_27/M1_1_16  ( .A(\Shifter/sll_27/ML_int[1][16] ), .B(
        \Shifter/sll_27/ML_int[1][14] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][16] ) );
  MUX \Shifter/sll_27/M1_1_17  ( .A(\Shifter/sll_27/ML_int[1][17] ), .B(
        \Shifter/sll_27/ML_int[1][15] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][17] ) );
  MUX \Shifter/sll_27/M1_1_18  ( .A(\Shifter/sll_27/ML_int[1][18] ), .B(
        \Shifter/sll_27/ML_int[1][16] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][18] ) );
  MUX \Shifter/sll_27/M1_1_19  ( .A(\Shifter/sll_27/ML_int[1][19] ), .B(
        \Shifter/sll_27/ML_int[1][17] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][19] ) );
  MUX \Shifter/sll_27/M1_1_20  ( .A(\Shifter/sll_27/ML_int[1][20] ), .B(
        \Shifter/sll_27/ML_int[1][18] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][20] ) );
  MUX \Shifter/sll_27/M1_1_21  ( .A(\Shifter/sll_27/ML_int[1][21] ), .B(
        \Shifter/sll_27/ML_int[1][19] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][21] ) );
  MUX \Shifter/sll_27/M1_1_22  ( .A(\Shifter/sll_27/ML_int[1][22] ), .B(
        \Shifter/sll_27/ML_int[1][20] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][22] ) );
  MUX \Shifter/sll_27/M1_1_23  ( .A(\Shifter/sll_27/ML_int[1][23] ), .B(
        \Shifter/sll_27/ML_int[1][21] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][23] ) );
  MUX \Shifter/sll_27/M1_1_24  ( .A(\Shifter/sll_27/ML_int[1][24] ), .B(
        \Shifter/sll_27/ML_int[1][22] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][24] ) );
  MUX \Shifter/sll_27/M1_1_25  ( .A(\Shifter/sll_27/ML_int[1][25] ), .B(
        \Shifter/sll_27/ML_int[1][23] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][25] ) );
  MUX \Shifter/sll_27/M1_1_26  ( .A(\Shifter/sll_27/ML_int[1][26] ), .B(
        \Shifter/sll_27/ML_int[1][24] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][26] ) );
  MUX \Shifter/sll_27/M1_1_27  ( .A(\Shifter/sll_27/ML_int[1][27] ), .B(
        \Shifter/sll_27/ML_int[1][25] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][27] ) );
  MUX \Shifter/sll_27/M1_1_28  ( .A(\Shifter/sll_27/ML_int[1][28] ), .B(
        \Shifter/sll_27/ML_int[1][26] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][28] ) );
  MUX \Shifter/sll_27/M1_1_29  ( .A(\Shifter/sll_27/ML_int[1][29] ), .B(
        \Shifter/sll_27/ML_int[1][27] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][29] ) );
  MUX \Shifter/sll_27/M1_1_30  ( .A(\Shifter/sll_27/ML_int[1][30] ), .B(
        \Shifter/sll_27/ML_int[1][28] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][30] ) );
  MUX \Shifter/sll_27/M1_1_31  ( .A(\Shifter/sll_27/ML_int[1][31] ), .B(
        \Shifter/sll_27/ML_int[1][29] ), .S(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][31] ) );
  MUX \Shifter/sll_27/M1_2_4  ( .A(\Shifter/sll_27/ML_int[2][4] ), .B(
        \Shifter/sll_27/ML_int[2][0] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][4] ) );
  MUX \Shifter/sll_27/M1_2_5  ( .A(\Shifter/sll_27/ML_int[2][5] ), .B(
        \Shifter/sll_27/ML_int[2][1] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][5] ) );
  MUX \Shifter/sll_27/M1_2_6  ( .A(\Shifter/sll_27/ML_int[2][6] ), .B(
        \Shifter/sll_27/ML_int[2][2] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][6] ) );
  MUX \Shifter/sll_27/M1_2_7  ( .A(\Shifter/sll_27/ML_int[2][7] ), .B(
        \Shifter/sll_27/ML_int[2][3] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][7] ) );
  MUX \Shifter/sll_27/M1_2_8  ( .A(\Shifter/sll_27/ML_int[2][8] ), .B(
        \Shifter/sll_27/ML_int[2][4] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][8] ) );
  MUX \Shifter/sll_27/M1_2_9  ( .A(\Shifter/sll_27/ML_int[2][9] ), .B(
        \Shifter/sll_27/ML_int[2][5] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][9] ) );
  MUX \Shifter/sll_27/M1_2_10  ( .A(\Shifter/sll_27/ML_int[2][10] ), .B(
        \Shifter/sll_27/ML_int[2][6] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][10] ) );
  MUX \Shifter/sll_27/M1_2_11  ( .A(\Shifter/sll_27/ML_int[2][11] ), .B(
        \Shifter/sll_27/ML_int[2][7] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][11] ) );
  MUX \Shifter/sll_27/M1_2_12  ( .A(\Shifter/sll_27/ML_int[2][12] ), .B(
        \Shifter/sll_27/ML_int[2][8] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][12] ) );
  MUX \Shifter/sll_27/M1_2_13  ( .A(\Shifter/sll_27/ML_int[2][13] ), .B(
        \Shifter/sll_27/ML_int[2][9] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][13] ) );
  MUX \Shifter/sll_27/M1_2_14  ( .A(\Shifter/sll_27/ML_int[2][14] ), .B(
        \Shifter/sll_27/ML_int[2][10] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][14] ) );
  MUX \Shifter/sll_27/M1_2_15  ( .A(\Shifter/sll_27/ML_int[2][15] ), .B(
        \Shifter/sll_27/ML_int[2][11] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][15] ) );
  MUX \Shifter/sll_27/M1_2_16  ( .A(\Shifter/sll_27/ML_int[2][16] ), .B(
        \Shifter/sll_27/ML_int[2][12] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][16] ) );
  MUX \Shifter/sll_27/M1_2_17  ( .A(\Shifter/sll_27/ML_int[2][17] ), .B(
        \Shifter/sll_27/ML_int[2][13] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][17] ) );
  MUX \Shifter/sll_27/M1_2_18  ( .A(\Shifter/sll_27/ML_int[2][18] ), .B(
        \Shifter/sll_27/ML_int[2][14] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][18] ) );
  MUX \Shifter/sll_27/M1_2_19  ( .A(\Shifter/sll_27/ML_int[2][19] ), .B(
        \Shifter/sll_27/ML_int[2][15] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][19] ) );
  MUX \Shifter/sll_27/M1_2_20  ( .A(\Shifter/sll_27/ML_int[2][20] ), .B(
        \Shifter/sll_27/ML_int[2][16] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][20] ) );
  MUX \Shifter/sll_27/M1_2_21  ( .A(\Shifter/sll_27/ML_int[2][21] ), .B(
        \Shifter/sll_27/ML_int[2][17] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][21] ) );
  MUX \Shifter/sll_27/M1_2_22  ( .A(\Shifter/sll_27/ML_int[2][22] ), .B(
        \Shifter/sll_27/ML_int[2][18] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][22] ) );
  MUX \Shifter/sll_27/M1_2_23  ( .A(\Shifter/sll_27/ML_int[2][23] ), .B(
        \Shifter/sll_27/ML_int[2][19] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][23] ) );
  MUX \Shifter/sll_27/M1_2_24  ( .A(\Shifter/sll_27/ML_int[2][24] ), .B(
        \Shifter/sll_27/ML_int[2][20] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][24] ) );
  MUX \Shifter/sll_27/M1_2_25  ( .A(\Shifter/sll_27/ML_int[2][25] ), .B(
        \Shifter/sll_27/ML_int[2][21] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][25] ) );
  MUX \Shifter/sll_27/M1_2_26  ( .A(\Shifter/sll_27/ML_int[2][26] ), .B(
        \Shifter/sll_27/ML_int[2][22] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][26] ) );
  MUX \Shifter/sll_27/M1_2_27  ( .A(\Shifter/sll_27/ML_int[2][27] ), .B(
        \Shifter/sll_27/ML_int[2][23] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][27] ) );
  MUX \Shifter/sll_27/M1_2_28  ( .A(\Shifter/sll_27/ML_int[2][28] ), .B(
        \Shifter/sll_27/ML_int[2][24] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][28] ) );
  MUX \Shifter/sll_27/M1_2_29  ( .A(\Shifter/sll_27/ML_int[2][29] ), .B(
        \Shifter/sll_27/ML_int[2][25] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][29] ) );
  MUX \Shifter/sll_27/M1_2_30  ( .A(\Shifter/sll_27/ML_int[2][30] ), .B(
        \Shifter/sll_27/ML_int[2][26] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][30] ) );
  MUX \Shifter/sll_27/M1_2_31  ( .A(\Shifter/sll_27/ML_int[2][31] ), .B(
        \Shifter/sll_27/ML_int[2][27] ), .S(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][31] ) );
  MUX \Shifter/sll_27/M1_3_8  ( .A(\Shifter/sll_27/ML_int[3][8] ), .B(
        \Shifter/sll_27/ML_int[3][0] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][8] ) );
  MUX \Shifter/sll_27/M1_3_9  ( .A(\Shifter/sll_27/ML_int[3][9] ), .B(
        \Shifter/sll_27/ML_int[3][1] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][9] ) );
  MUX \Shifter/sll_27/M1_3_10  ( .A(\Shifter/sll_27/ML_int[3][10] ), .B(
        \Shifter/sll_27/ML_int[3][2] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][10] ) );
  MUX \Shifter/sll_27/M1_3_11  ( .A(\Shifter/sll_27/ML_int[3][11] ), .B(
        \Shifter/sll_27/ML_int[3][3] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][11] ) );
  MUX \Shifter/sll_27/M1_3_12  ( .A(\Shifter/sll_27/ML_int[3][12] ), .B(
        \Shifter/sll_27/ML_int[3][4] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][12] ) );
  MUX \Shifter/sll_27/M1_3_13  ( .A(\Shifter/sll_27/ML_int[3][13] ), .B(
        \Shifter/sll_27/ML_int[3][5] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][13] ) );
  MUX \Shifter/sll_27/M1_3_14  ( .A(\Shifter/sll_27/ML_int[3][14] ), .B(
        \Shifter/sll_27/ML_int[3][6] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][14] ) );
  MUX \Shifter/sll_27/M1_3_15  ( .A(\Shifter/sll_27/ML_int[3][15] ), .B(
        \Shifter/sll_27/ML_int[3][7] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][15] ) );
  MUX \Shifter/sll_27/M1_3_16  ( .A(\Shifter/sll_27/ML_int[3][16] ), .B(
        \Shifter/sll_27/ML_int[3][8] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][16] ) );
  MUX \Shifter/sll_27/M1_3_17  ( .A(\Shifter/sll_27/ML_int[3][17] ), .B(
        \Shifter/sll_27/ML_int[3][9] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][17] ) );
  MUX \Shifter/sll_27/M1_3_18  ( .A(\Shifter/sll_27/ML_int[3][18] ), .B(
        \Shifter/sll_27/ML_int[3][10] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][18] ) );
  MUX \Shifter/sll_27/M1_3_19  ( .A(\Shifter/sll_27/ML_int[3][19] ), .B(
        \Shifter/sll_27/ML_int[3][11] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][19] ) );
  MUX \Shifter/sll_27/M1_3_20  ( .A(\Shifter/sll_27/ML_int[3][20] ), .B(
        \Shifter/sll_27/ML_int[3][12] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][20] ) );
  MUX \Shifter/sll_27/M1_3_21  ( .A(\Shifter/sll_27/ML_int[3][21] ), .B(
        \Shifter/sll_27/ML_int[3][13] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][21] ) );
  MUX \Shifter/sll_27/M1_3_22  ( .A(\Shifter/sll_27/ML_int[3][22] ), .B(
        \Shifter/sll_27/ML_int[3][14] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][22] ) );
  MUX \Shifter/sll_27/M1_3_23  ( .A(\Shifter/sll_27/ML_int[3][23] ), .B(
        \Shifter/sll_27/ML_int[3][15] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][23] ) );
  MUX \Shifter/sll_27/M1_3_24  ( .A(\Shifter/sll_27/ML_int[3][24] ), .B(
        \Shifter/sll_27/ML_int[3][16] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][24] ) );
  MUX \Shifter/sll_27/M1_3_25  ( .A(\Shifter/sll_27/ML_int[3][25] ), .B(
        \Shifter/sll_27/ML_int[3][17] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][25] ) );
  MUX \Shifter/sll_27/M1_3_26  ( .A(\Shifter/sll_27/ML_int[3][26] ), .B(
        \Shifter/sll_27/ML_int[3][18] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][26] ) );
  MUX \Shifter/sll_27/M1_3_27  ( .A(\Shifter/sll_27/ML_int[3][27] ), .B(
        \Shifter/sll_27/ML_int[3][19] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][27] ) );
  MUX \Shifter/sll_27/M1_3_28  ( .A(\Shifter/sll_27/ML_int[3][28] ), .B(
        \Shifter/sll_27/ML_int[3][20] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][28] ) );
  MUX \Shifter/sll_27/M1_3_29  ( .A(\Shifter/sll_27/ML_int[3][29] ), .B(
        \Shifter/sll_27/ML_int[3][21] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][29] ) );
  MUX \Shifter/sll_27/M1_3_30  ( .A(\Shifter/sll_27/ML_int[3][30] ), .B(
        \Shifter/sll_27/ML_int[3][22] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][30] ) );
  MUX \Shifter/sll_27/M1_3_31  ( .A(\Shifter/sll_27/ML_int[3][31] ), .B(
        \Shifter/sll_27/ML_int[3][23] ), .S(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][31] ) );
  MUX \Shifter/sll_27/M1_4_16  ( .A(\Shifter/sll_27/ML_int[4][16] ), .B(
        \Shifter/sll_27/ML_int[4][0] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][16] ) );
  MUX \Shifter/sll_27/M1_4_17  ( .A(\Shifter/sll_27/ML_int[4][17] ), .B(
        \Shifter/sll_27/ML_int[4][1] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][17] ) );
  MUX \Shifter/sll_27/M1_4_18  ( .A(\Shifter/sll_27/ML_int[4][18] ), .B(
        \Shifter/sll_27/ML_int[4][2] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][18] ) );
  MUX \Shifter/sll_27/M1_4_19  ( .A(\Shifter/sll_27/ML_int[4][19] ), .B(
        \Shifter/sll_27/ML_int[4][3] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][19] ) );
  MUX \Shifter/sll_27/M1_4_20  ( .A(\Shifter/sll_27/ML_int[4][20] ), .B(
        \Shifter/sll_27/ML_int[4][4] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][20] ) );
  MUX \Shifter/sll_27/M1_4_21  ( .A(\Shifter/sll_27/ML_int[4][21] ), .B(
        \Shifter/sll_27/ML_int[4][5] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][21] ) );
  MUX \Shifter/sll_27/M1_4_22  ( .A(\Shifter/sll_27/ML_int[4][22] ), .B(
        \Shifter/sll_27/ML_int[4][6] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][22] ) );
  MUX \Shifter/sll_27/M1_4_23  ( .A(\Shifter/sll_27/ML_int[4][23] ), .B(
        \Shifter/sll_27/ML_int[4][7] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][23] ) );
  MUX \Shifter/sll_27/M1_4_24  ( .A(\Shifter/sll_27/ML_int[4][24] ), .B(
        \Shifter/sll_27/ML_int[4][8] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][24] ) );
  MUX \Shifter/sll_27/M1_4_25  ( .A(\Shifter/sll_27/ML_int[4][25] ), .B(
        \Shifter/sll_27/ML_int[4][9] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][25] ) );
  MUX \Shifter/sll_27/M1_4_26  ( .A(\Shifter/sll_27/ML_int[4][26] ), .B(
        \Shifter/sll_27/ML_int[4][10] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][26] ) );
  MUX \Shifter/sll_27/M1_4_27  ( .A(\Shifter/sll_27/ML_int[4][27] ), .B(
        \Shifter/sll_27/ML_int[4][11] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][27] ) );
  MUX \Shifter/sll_27/M1_4_28  ( .A(\Shifter/sll_27/ML_int[4][28] ), .B(
        \Shifter/sll_27/ML_int[4][12] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][28] ) );
  MUX \Shifter/sll_27/M1_4_29  ( .A(\Shifter/sll_27/ML_int[4][29] ), .B(
        \Shifter/sll_27/ML_int[4][13] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][29] ) );
  MUX \Shifter/sll_27/M1_4_30  ( .A(\Shifter/sll_27/ML_int[4][30] ), .B(
        \Shifter/sll_27/ML_int[4][14] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][30] ) );
  MUX \Shifter/sll_27/M1_4_31  ( .A(\Shifter/sll_27/ML_int[4][31] ), .B(
        \Shifter/sll_27/ML_int[4][15] ), .S(a_bus[4]), .Z(
        \Shifter/sll_27/ML_int[5][31] ) );
  FA \ALU/r67/U1_0  ( .A(a_bus[0]), .B(\ALU/r67/B_AS[0] ), .CI(\ALU/U2/U1/Z_0 ), .CO(\ALU/r67/carry[1] ), .S(\ALU/N108 ) );
  FA \ALU/r67/U1_1  ( .A(a_bus[1]), .B(\ALU/r67/B_AS[1] ), .CI(
        \ALU/r67/carry[1] ), .CO(\ALU/r67/carry[2] ), .S(\ALU/N109 ) );
  FA \ALU/r67/U1_2  ( .A(a_bus[2]), .B(\ALU/r67/B_AS[2] ), .CI(
        \ALU/r67/carry[2] ), .CO(\ALU/r67/carry[3] ), .S(\ALU/N110 ) );
  FA \ALU/r67/U1_3  ( .A(a_bus[3]), .B(\ALU/r67/B_AS[3] ), .CI(
        \ALU/r67/carry[3] ), .CO(\ALU/r67/carry[4] ), .S(\ALU/N111 ) );
  FA \ALU/r67/U1_4  ( .A(a_bus[4]), .B(\ALU/r67/B_AS[4] ), .CI(
        \ALU/r67/carry[4] ), .CO(\ALU/r67/carry[5] ), .S(\ALU/N112 ) );
  FA \ALU/r67/U1_5  ( .A(n2485), .B(\ALU/r67/B_AS[5] ), .CI(\ALU/r67/carry[5] ), .CO(\ALU/r67/carry[6] ), .S(\ALU/N113 ) );
  FA \ALU/r67/U1_6  ( .A(n2484), .B(\ALU/r67/B_AS[6] ), .CI(\ALU/r67/carry[6] ), .CO(\ALU/r67/carry[7] ), .S(\ALU/N114 ) );
  FA \ALU/r67/U1_7  ( .A(n2483), .B(\ALU/r67/B_AS[7] ), .CI(\ALU/r67/carry[7] ), .CO(\ALU/r67/carry[8] ), .S(\ALU/N115 ) );
  FA \ALU/r67/U1_8  ( .A(n2482), .B(\ALU/r67/B_AS[8] ), .CI(\ALU/r67/carry[8] ), .CO(\ALU/r67/carry[9] ), .S(\ALU/N116 ) );
  FA \ALU/r67/U1_9  ( .A(n2481), .B(\ALU/r67/B_AS[9] ), .CI(\ALU/r67/carry[9] ), .CO(\ALU/r67/carry[10] ), .S(\ALU/N117 ) );
  FA \ALU/r67/U1_10  ( .A(n2507), .B(\ALU/r67/B_AS[10] ), .CI(
        \ALU/r67/carry[10] ), .CO(\ALU/r67/carry[11] ), .S(\ALU/N118 ) );
  FA \ALU/r67/U1_11  ( .A(n2506), .B(\ALU/r67/B_AS[11] ), .CI(
        \ALU/r67/carry[11] ), .CO(\ALU/r67/carry[12] ), .S(\ALU/N119 ) );
  FA \ALU/r67/U1_12  ( .A(n2505), .B(\ALU/r67/B_AS[12] ), .CI(
        \ALU/r67/carry[12] ), .CO(\ALU/r67/carry[13] ), .S(\ALU/N120 ) );
  FA \ALU/r67/U1_13  ( .A(n2504), .B(\ALU/r67/B_AS[13] ), .CI(
        \ALU/r67/carry[13] ), .CO(\ALU/r67/carry[14] ), .S(\ALU/N121 ) );
  FA \ALU/r67/U1_14  ( .A(n2503), .B(\ALU/r67/B_AS[14] ), .CI(
        \ALU/r67/carry[14] ), .CO(\ALU/r67/carry[15] ), .S(\ALU/N122 ) );
  FA \ALU/r67/U1_15  ( .A(n2502), .B(\ALU/r67/B_AS[15] ), .CI(
        \ALU/r67/carry[15] ), .CO(\ALU/r67/carry[16] ), .S(\ALU/N123 ) );
  FA \ALU/r67/U1_16  ( .A(n2501), .B(\ALU/r67/B_AS[16] ), .CI(
        \ALU/r67/carry[16] ), .CO(\ALU/r67/carry[17] ), .S(\ALU/N124 ) );
  FA \ALU/r67/U1_17  ( .A(n2500), .B(\ALU/r67/B_AS[17] ), .CI(
        \ALU/r67/carry[17] ), .CO(\ALU/r67/carry[18] ), .S(\ALU/N125 ) );
  FA \ALU/r67/U1_18  ( .A(n2499), .B(\ALU/r67/B_AS[18] ), .CI(
        \ALU/r67/carry[18] ), .CO(\ALU/r67/carry[19] ), .S(\ALU/N126 ) );
  FA \ALU/r67/U1_19  ( .A(n2498), .B(\ALU/r67/B_AS[19] ), .CI(
        \ALU/r67/carry[19] ), .CO(\ALU/r67/carry[20] ), .S(\ALU/N127 ) );
  FA \ALU/r67/U1_20  ( .A(n2497), .B(\ALU/r67/B_AS[20] ), .CI(
        \ALU/r67/carry[20] ), .CO(\ALU/r67/carry[21] ), .S(\ALU/N128 ) );
  FA \ALU/r67/U1_21  ( .A(n2496), .B(\ALU/r67/B_AS[21] ), .CI(
        \ALU/r67/carry[21] ), .CO(\ALU/r67/carry[22] ), .S(\ALU/N129 ) );
  FA \ALU/r67/U1_22  ( .A(n2495), .B(\ALU/r67/B_AS[22] ), .CI(
        \ALU/r67/carry[22] ), .CO(\ALU/r67/carry[23] ), .S(\ALU/N130 ) );
  FA \ALU/r67/U1_23  ( .A(n2494), .B(\ALU/r67/B_AS[23] ), .CI(
        \ALU/r67/carry[23] ), .CO(\ALU/r67/carry[24] ), .S(\ALU/N131 ) );
  FA \ALU/r67/U1_24  ( .A(n2493), .B(\ALU/r67/B_AS[24] ), .CI(
        \ALU/r67/carry[24] ), .CO(\ALU/r67/carry[25] ), .S(\ALU/N132 ) );
  FA \ALU/r67/U1_25  ( .A(n2492), .B(\ALU/r67/B_AS[25] ), .CI(
        \ALU/r67/carry[25] ), .CO(\ALU/r67/carry[26] ), .S(\ALU/N133 ) );
  FA \ALU/r67/U1_26  ( .A(n2491), .B(\ALU/r67/B_AS[26] ), .CI(
        \ALU/r67/carry[26] ), .CO(\ALU/r67/carry[27] ), .S(\ALU/N134 ) );
  FA \ALU/r67/U1_27  ( .A(n2490), .B(\ALU/r67/B_AS[27] ), .CI(
        \ALU/r67/carry[27] ), .CO(\ALU/r67/carry[28] ), .S(\ALU/N135 ) );
  FA \ALU/r67/U1_28  ( .A(n2489), .B(\ALU/r67/B_AS[28] ), .CI(
        \ALU/r67/carry[28] ), .CO(\ALU/r67/carry[29] ), .S(\ALU/N136 ) );
  FA \ALU/r67/U1_29  ( .A(n2488), .B(\ALU/r67/B_AS[29] ), .CI(
        \ALU/r67/carry[29] ), .CO(\ALU/r67/carry[30] ), .S(\ALU/N137 ) );
  FA \ALU/r67/U1_30  ( .A(n2487), .B(\ALU/r67/B_AS[30] ), .CI(
        \ALU/r67/carry[30] ), .CO(\ALU/r67/carry[31] ), .S(\ALU/N138 ) );
  FA \ALU/r67/U1_31  ( .A(n2486), .B(\ALU/r67/B_AS[31] ), .CI(
        \ALU/r67/carry[31] ), .S(\ALU/N139 ) );
  HA \PC_Next/add_30/U1_1_1  ( .A(pc_current[3]), .B(pc_current[2]), .CO(
        \PC_Next/add_30/carry[2] ), .S(pc_plus4[3]) );
  HA \PC_Next/add_30/U1_1_2  ( .A(pc_current[4]), .B(\PC_Next/add_30/carry[2] ), .CO(\PC_Next/add_30/carry[3] ), .S(pc_plus4[4]) );
  HA \PC_Next/add_30/U1_1_3  ( .A(pc_current[5]), .B(\PC_Next/add_30/carry[3] ), .CO(\PC_Next/add_30/carry[4] ), .S(pc_plus4[5]) );
  HA \PC_Next/add_30/U1_1_4  ( .A(pc_current[6]), .B(\PC_Next/add_30/carry[4] ), .CO(\PC_Next/add_30/carry[5] ), .S(pc_plus4[6]) );
  HA \PC_Next/add_30/U1_1_5  ( .A(pc_current[7]), .B(\PC_Next/add_30/carry[5] ), .CO(\PC_Next/add_30/carry[6] ), .S(pc_plus4[7]) );
  HA \PC_Next/add_30/U1_1_6  ( .A(pc_current[8]), .B(\PC_Next/add_30/carry[6] ), .CO(\PC_Next/add_30/carry[7] ), .S(pc_plus4[8]) );
  HA \PC_Next/add_30/U1_1_7  ( .A(pc_current[9]), .B(\PC_Next/add_30/carry[7] ), .CO(\PC_Next/add_30/carry[8] ), .S(pc_plus4[9]) );
  HA \PC_Next/add_30/U1_1_8  ( .A(pc_current[10]), .B(
        \PC_Next/add_30/carry[8] ), .CO(\PC_Next/add_30/carry[9] ), .S(
        pc_plus4[10]) );
  HA \PC_Next/add_30/U1_1_9  ( .A(pc_current[11]), .B(
        \PC_Next/add_30/carry[9] ), .CO(\PC_Next/add_30/carry[10] ), .S(
        pc_plus4[11]) );
  HA \PC_Next/add_30/U1_1_10  ( .A(pc_current[12]), .B(
        \PC_Next/add_30/carry[10] ), .CO(\PC_Next/add_30/carry[11] ), .S(
        pc_plus4[12]) );
  HA \PC_Next/add_30/U1_1_11  ( .A(pc_current[13]), .B(
        \PC_Next/add_30/carry[11] ), .CO(\PC_Next/add_30/carry[12] ), .S(
        pc_plus4[13]) );
  HA \PC_Next/add_30/U1_1_12  ( .A(pc_current[14]), .B(
        \PC_Next/add_30/carry[12] ), .CO(\PC_Next/add_30/carry[13] ), .S(
        pc_plus4[14]) );
  HA \PC_Next/add_30/U1_1_13  ( .A(pc_current[15]), .B(
        \PC_Next/add_30/carry[13] ), .CO(\PC_Next/add_30/carry[14] ), .S(
        pc_plus4[15]) );
  HA \PC_Next/add_30/U1_1_14  ( .A(pc_current[16]), .B(
        \PC_Next/add_30/carry[14] ), .CO(\PC_Next/add_30/carry[15] ), .S(
        pc_plus4[16]) );
  HA \PC_Next/add_30/U1_1_15  ( .A(pc_current[17]), .B(
        \PC_Next/add_30/carry[15] ), .CO(\PC_Next/add_30/carry[16] ), .S(
        pc_plus4[17]) );
  HA \PC_Next/add_30/U1_1_16  ( .A(pc_current[18]), .B(
        \PC_Next/add_30/carry[16] ), .CO(\PC_Next/add_30/carry[17] ), .S(
        pc_plus4[18]) );
  HA \PC_Next/add_30/U1_1_17  ( .A(pc_current[19]), .B(
        \PC_Next/add_30/carry[17] ), .CO(\PC_Next/add_30/carry[18] ), .S(
        pc_plus4[19]) );
  HA \PC_Next/add_30/U1_1_18  ( .A(pc_current[20]), .B(
        \PC_Next/add_30/carry[18] ), .CO(\PC_Next/add_30/carry[19] ), .S(
        pc_plus4[20]) );
  HA \PC_Next/add_30/U1_1_19  ( .A(pc_current[21]), .B(
        \PC_Next/add_30/carry[19] ), .CO(\PC_Next/add_30/carry[20] ), .S(
        pc_plus4[21]) );
  HA \PC_Next/add_30/U1_1_20  ( .A(pc_current[22]), .B(
        \PC_Next/add_30/carry[20] ), .CO(\PC_Next/add_30/carry[21] ), .S(
        pc_plus4[22]) );
  HA \PC_Next/add_30/U1_1_21  ( .A(pc_current[23]), .B(
        \PC_Next/add_30/carry[21] ), .CO(\PC_Next/add_30/carry[22] ), .S(
        pc_plus4[23]) );
  HA \PC_Next/add_30/U1_1_22  ( .A(pc_current[24]), .B(
        \PC_Next/add_30/carry[22] ), .CO(\PC_Next/add_30/carry[23] ), .S(
        pc_plus4[24]) );
  HA \PC_Next/add_30/U1_1_23  ( .A(pc_current[25]), .B(
        \PC_Next/add_30/carry[23] ), .CO(\PC_Next/add_30/carry[24] ), .S(
        pc_plus4[25]) );
  HA \PC_Next/add_30/U1_1_24  ( .A(pc_current[26]), .B(
        \PC_Next/add_30/carry[24] ), .CO(\PC_Next/add_30/carry[25] ), .S(
        pc_plus4[26]) );
  HA \PC_Next/add_30/U1_1_25  ( .A(pc_current[27]), .B(
        \PC_Next/add_30/carry[25] ), .CO(\PC_Next/add_30/carry[26] ), .S(
        pc_plus4[27]) );
  HA \PC_Next/add_30/U1_1_26  ( .A(pc_current[28]), .B(
        \PC_Next/add_30/carry[26] ), .CO(\PC_Next/add_30/carry[27] ), .S(
        pc_plus4[28]) );
  HA \PC_Next/add_30/U1_1_27  ( .A(pc_current[29]), .B(
        \PC_Next/add_30/carry[27] ), .CO(\PC_Next/add_30/carry[28] ), .S(
        pc_plus4[29]) );
  HA \PC_Next/add_30/U1_1_28  ( .A(pc_current[30]), .B(
        \PC_Next/add_30/carry[28] ), .CO(\PC_Next/add_30/carry[29] ), .S(
        pc_plus4[30]) );
  FA \PC_Next/add_41/U1_1  ( .A(pc_current[3]), .B(imm[1]), .CI(
        \PC_Next/add_41/carry[1] ), .CO(\PC_Next/add_41/carry[2] ), .S(
        \PC_Next/N17 ) );
  FA \PC_Next/add_41/U1_2  ( .A(pc_current[4]), .B(imm[2]), .CI(
        \PC_Next/add_41/carry[2] ), .CO(\PC_Next/add_41/carry[3] ), .S(
        \PC_Next/N18 ) );
  FA \PC_Next/add_41/U1_3  ( .A(pc_current[5]), .B(imm[3]), .CI(
        \PC_Next/add_41/carry[3] ), .CO(\PC_Next/add_41/carry[4] ), .S(
        \PC_Next/N19 ) );
  FA \PC_Next/add_41/U1_4  ( .A(pc_current[6]), .B(imm[4]), .CI(
        \PC_Next/add_41/carry[4] ), .CO(\PC_Next/add_41/carry[5] ), .S(
        \PC_Next/N20 ) );
  FA \PC_Next/add_41/U1_5  ( .A(pc_current[7]), .B(imm[5]), .CI(
        \PC_Next/add_41/carry[5] ), .CO(\PC_Next/add_41/carry[6] ), .S(
        \PC_Next/N21 ) );
  FA \PC_Next/add_41/U1_6  ( .A(pc_current[8]), .B(imm[6]), .CI(
        \PC_Next/add_41/carry[6] ), .CO(\PC_Next/add_41/carry[7] ), .S(
        \PC_Next/N22 ) );
  FA \PC_Next/add_41/U1_7  ( .A(pc_current[9]), .B(imm[7]), .CI(
        \PC_Next/add_41/carry[7] ), .CO(\PC_Next/add_41/carry[8] ), .S(
        \PC_Next/N23 ) );
  FA \PC_Next/add_41/U1_8  ( .A(pc_current[10]), .B(imm[8]), .CI(
        \PC_Next/add_41/carry[8] ), .CO(\PC_Next/add_41/carry[9] ), .S(
        \PC_Next/N24 ) );
  FA \PC_Next/add_41/U1_9  ( .A(pc_current[11]), .B(imm[9]), .CI(
        \PC_Next/add_41/carry[9] ), .CO(\PC_Next/add_41/carry[10] ), .S(
        \PC_Next/N25 ) );
  FA \PC_Next/add_41/U1_10  ( .A(pc_current[12]), .B(imm[10]), .CI(
        \PC_Next/add_41/carry[10] ), .CO(\PC_Next/add_41/carry[11] ), .S(
        \PC_Next/N26 ) );
  FA \PC_Next/add_41/U1_11  ( .A(pc_current[13]), .B(imm[11]), .CI(
        \PC_Next/add_41/carry[11] ), .CO(\PC_Next/add_41/carry[12] ), .S(
        \PC_Next/N27 ) );
  FA \PC_Next/add_41/U1_12  ( .A(pc_current[14]), .B(imm[12]), .CI(
        \PC_Next/add_41/carry[12] ), .CO(\PC_Next/add_41/carry[13] ), .S(
        \PC_Next/N28 ) );
  FA \PC_Next/add_41/U1_13  ( .A(pc_current[15]), .B(imm[13]), .CI(
        \PC_Next/add_41/carry[13] ), .CO(\PC_Next/add_41/carry[14] ), .S(
        \PC_Next/N29 ) );
  FA \PC_Next/add_41/U1_14  ( .A(pc_current[16]), .B(imm[14]), .CI(
        \PC_Next/add_41/carry[14] ), .CO(\PC_Next/add_41/carry[15] ), .S(
        \PC_Next/N30 ) );
  FA \PC_Next/add_41/U1_15  ( .A(pc_current[17]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[15] ), .CO(\PC_Next/add_41/carry[16] ), .S(
        \PC_Next/N31 ) );
  FA \PC_Next/add_41/U1_16  ( .A(pc_current[18]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[16] ), .CO(\PC_Next/add_41/carry[17] ), .S(
        \PC_Next/N32 ) );
  FA \PC_Next/add_41/U1_17  ( .A(pc_current[19]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[17] ), .CO(\PC_Next/add_41/carry[18] ), .S(
        \PC_Next/N33 ) );
  FA \PC_Next/add_41/U1_18  ( .A(pc_current[20]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[18] ), .CO(\PC_Next/add_41/carry[19] ), .S(
        \PC_Next/N34 ) );
  FA \PC_Next/add_41/U1_19  ( .A(pc_current[21]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[19] ), .CO(\PC_Next/add_41/carry[20] ), .S(
        \PC_Next/N35 ) );
  FA \PC_Next/add_41/U1_20  ( .A(pc_current[22]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[20] ), .CO(\PC_Next/add_41/carry[21] ), .S(
        \PC_Next/N36 ) );
  FA \PC_Next/add_41/U1_21  ( .A(pc_current[23]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[21] ), .CO(\PC_Next/add_41/carry[22] ), .S(
        \PC_Next/N37 ) );
  FA \PC_Next/add_41/U1_22  ( .A(pc_current[24]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[22] ), .CO(\PC_Next/add_41/carry[23] ), .S(
        \PC_Next/N38 ) );
  FA \PC_Next/add_41/U1_23  ( .A(pc_current[25]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[23] ), .CO(\PC_Next/add_41/carry[24] ), .S(
        \PC_Next/N39 ) );
  FA \PC_Next/add_41/U1_24  ( .A(pc_current[26]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[24] ), .CO(\PC_Next/add_41/carry[25] ), .S(
        \PC_Next/N40 ) );
  FA \PC_Next/add_41/U1_25  ( .A(pc_current[27]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[25] ), .CO(\PC_Next/add_41/carry[26] ), .S(
        \PC_Next/N41 ) );
  FA \PC_Next/add_41/U1_26  ( .A(pc_current[28]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[26] ), .CO(\PC_Next/add_41/carry[27] ), .S(
        \PC_Next/N42 ) );
  FA \PC_Next/add_41/U1_27  ( .A(pc_current[29]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[27] ), .CO(\PC_Next/add_41/carry[28] ), .S(
        \PC_Next/N43 ) );
  FA \PC_Next/add_41/U1_28  ( .A(pc_current[30]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[28] ), .CO(\PC_Next/add_41/carry[29] ), .S(
        \PC_Next/N44 ) );
  FA \PC_Next/add_41/U1_29  ( .A(pc_current[31]), .B(imm[15]), .CI(
        \PC_Next/add_41/carry[29] ), .S(\PC_Next/N45 ) );
  AND U34 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][31] ), .Z(
        \Reg_Bank/n5938 ) );
  AND U35 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][31] ), .Z(
        \Reg_Bank/n4978 ) );
  AND U36 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][30] ), .Z(
        \Reg_Bank/n5908 ) );
  AND U37 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][30] ), .Z(
        \Reg_Bank/n4948 ) );
  AND U38 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][29] ), .Z(
        \Reg_Bank/n5878 ) );
  AND U39 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][29] ), .Z(
        \Reg_Bank/n4918 ) );
  AND U40 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][28] ), .Z(
        \Reg_Bank/n5848 ) );
  AND U41 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][28] ), .Z(
        \Reg_Bank/n4888 ) );
  AND U42 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][27] ), .Z(
        \Reg_Bank/n5818 ) );
  AND U43 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][27] ), .Z(
        \Reg_Bank/n4858 ) );
  AND U44 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][26] ), .Z(
        \Reg_Bank/n5788 ) );
  AND U45 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][26] ), .Z(
        \Reg_Bank/n4828 ) );
  AND U46 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][25] ), .Z(
        \Reg_Bank/n5758 ) );
  AND U47 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][25] ), .Z(
        \Reg_Bank/n4798 ) );
  AND U48 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][24] ), .Z(
        \Reg_Bank/n5728 ) );
  AND U49 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][24] ), .Z(
        \Reg_Bank/n4768 ) );
  AND U50 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][23] ), .Z(
        \Reg_Bank/n5698 ) );
  AND U51 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][23] ), .Z(
        \Reg_Bank/n4738 ) );
  AND U52 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][22] ), .Z(
        \Reg_Bank/n5668 ) );
  AND U53 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][22] ), .Z(
        \Reg_Bank/n4708 ) );
  AND U54 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][21] ), .Z(
        \Reg_Bank/n5638 ) );
  AND U55 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][21] ), .Z(
        \Reg_Bank/n4678 ) );
  AND U56 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][20] ), .Z(
        \Reg_Bank/n5608 ) );
  AND U57 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][20] ), .Z(
        \Reg_Bank/n4648 ) );
  AND U58 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][19] ), .Z(
        \Reg_Bank/n5578 ) );
  AND U59 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][19] ), .Z(
        \Reg_Bank/n4618 ) );
  AND U60 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][18] ), .Z(
        \Reg_Bank/n5548 ) );
  AND U61 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][18] ), .Z(
        \Reg_Bank/n4588 ) );
  AND U62 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][17] ), .Z(
        \Reg_Bank/n5518 ) );
  AND U63 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][17] ), .Z(
        \Reg_Bank/n4558 ) );
  AND U64 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][16] ), .Z(
        \Reg_Bank/n5488 ) );
  AND U65 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][16] ), .Z(
        \Reg_Bank/n4528 ) );
  AND U66 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][15] ), .Z(
        \Reg_Bank/n5458 ) );
  AND U67 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][15] ), .Z(
        \Reg_Bank/n4498 ) );
  AND U68 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][14] ), .Z(
        \Reg_Bank/n5428 ) );
  AND U69 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][14] ), .Z(
        \Reg_Bank/n4468 ) );
  AND U70 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][13] ), .Z(
        \Reg_Bank/n5398 ) );
  AND U71 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][13] ), .Z(
        \Reg_Bank/n4438 ) );
  AND U72 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][12] ), .Z(
        \Reg_Bank/n5368 ) );
  AND U73 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][12] ), .Z(
        \Reg_Bank/n4408 ) );
  AND U74 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][11] ), .Z(
        \Reg_Bank/n5338 ) );
  AND U75 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][11] ), .Z(
        \Reg_Bank/n4378 ) );
  AND U76 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][10] ), .Z(
        \Reg_Bank/n5308 ) );
  AND U77 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][10] ), .Z(
        \Reg_Bank/n4348 ) );
  AND U78 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][9] ), .Z(
        \Reg_Bank/n5278 ) );
  AND U79 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][9] ), .Z(
        \Reg_Bank/n4318 ) );
  AND U80 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][8] ), .Z(
        \Reg_Bank/n5248 ) );
  AND U81 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][8] ), .Z(
        \Reg_Bank/n4288 ) );
  AND U82 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][7] ), .Z(
        \Reg_Bank/n5218 ) );
  AND U83 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][7] ), .Z(
        \Reg_Bank/n4258 ) );
  AND U84 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][6] ), .Z(
        \Reg_Bank/n5188 ) );
  AND U85 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][6] ), .Z(
        \Reg_Bank/n4228 ) );
  AND U86 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][5] ), .Z(
        \Reg_Bank/n5158 ) );
  AND U87 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][5] ), .Z(
        \Reg_Bank/n4198 ) );
  AND U88 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][4] ), .Z(
        \Reg_Bank/n5128 ) );
  AND U89 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][4] ), .Z(
        \Reg_Bank/n4168 ) );
  AND U90 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][3] ), .Z(
        \Reg_Bank/n5098 ) );
  AND U91 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][3] ), .Z(
        \Reg_Bank/n4138 ) );
  AND U92 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][2] ), .Z(
        \Reg_Bank/n5068 ) );
  AND U93 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][2] ), .Z(
        \Reg_Bank/n4108 ) );
  AND U94 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][1] ), .Z(
        \Reg_Bank/n5038 ) );
  AND U95 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][1] ), .Z(
        \Reg_Bank/n4078 ) );
  AND U96 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][0] ), .Z(
        \Reg_Bank/n5008 ) );
  AND U97 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][0] ), .Z(
        \Reg_Bank/n4048 ) );
  AND U98 ( .A(imm[0]), .B(pc_current[2]), .Z(\PC_Next/add_41/carry[1] ) );
  XOR U99 ( .A(imm[0]), .B(pc_current[2]), .Z(\PC_Next/N16 ) );
  NAND U100 ( .A(n1), .B(n2), .Z(rt_index[4]) );
  NAND U101 ( .A(n3), .B(opcode[20]), .Z(n2) );
  AND U102 ( .A(n4), .B(n5), .Z(n1) );
  NAND U103 ( .A(n6), .B(n7), .Z(n5) );
  NAND U104 ( .A(n8), .B(n9), .Z(n6) );
  NAND U105 ( .A(n10), .B(n11), .Z(n9) );
  NAND U106 ( .A(n12), .B(n13), .Z(n11) );
  NAND U107 ( .A(imm[1]), .B(opcode[20]), .Z(n13) );
  NAND U108 ( .A(n14), .B(opcode[20]), .Z(n12) );
  AND U109 ( .A(n15), .B(n16), .Z(n8) );
  NAND U110 ( .A(n17), .B(n18), .Z(n16) );
  NAND U111 ( .A(n19), .B(n20), .Z(n18) );
  NANDN U112 ( .A(n21), .B(opcode[20]), .Z(n20) );
  NAND U113 ( .A(opcode[19]), .B(opcode[20]), .Z(n19) );
  NAND U114 ( .A(n22), .B(opcode[20]), .Z(n15) );
  NAND U115 ( .A(n23), .B(n24), .Z(n4) );
  NAND U116 ( .A(n25), .B(n26), .Z(n23) );
  NAND U117 ( .A(n27), .B(opcode[20]), .Z(n26) );
  NAND U118 ( .A(n28), .B(opcode[20]), .Z(n25) );
  NAND U119 ( .A(n29), .B(n30), .Z(rt_index[3]) );
  NAND U120 ( .A(opcode[19]), .B(n3), .Z(n30) );
  AND U121 ( .A(n31), .B(n32), .Z(n29) );
  NAND U122 ( .A(n33), .B(n7), .Z(n32) );
  NAND U123 ( .A(n34), .B(n35), .Z(n33) );
  NAND U124 ( .A(n10), .B(n36), .Z(n35) );
  NAND U125 ( .A(n37), .B(n38), .Z(n36) );
  NAND U126 ( .A(imm[1]), .B(opcode[19]), .Z(n38) );
  NAND U127 ( .A(opcode[19]), .B(n14), .Z(n37) );
  AND U128 ( .A(n39), .B(n40), .Z(n34) );
  NAND U129 ( .A(n17), .B(opcode[19]), .Z(n40) );
  NAND U130 ( .A(opcode[19]), .B(n22), .Z(n39) );
  NAND U131 ( .A(n41), .B(n24), .Z(n31) );
  NAND U132 ( .A(n42), .B(n43), .Z(n41) );
  NAND U133 ( .A(opcode[19]), .B(n27), .Z(n43) );
  NAND U134 ( .A(opcode[19]), .B(n28), .Z(n42) );
  NAND U135 ( .A(n44), .B(n45), .Z(rt_index[2]) );
  NAND U136 ( .A(n3), .B(opcode[18]), .Z(n45) );
  AND U137 ( .A(n46), .B(n47), .Z(n44) );
  NAND U138 ( .A(n48), .B(n7), .Z(n47) );
  NAND U139 ( .A(n49), .B(n50), .Z(n48) );
  NAND U140 ( .A(n10), .B(n51), .Z(n50) );
  NAND U141 ( .A(n52), .B(n53), .Z(n51) );
  NAND U142 ( .A(imm[1]), .B(opcode[18]), .Z(n53) );
  NAND U143 ( .A(n14), .B(opcode[18]), .Z(n52) );
  AND U144 ( .A(n54), .B(n55), .Z(n49) );
  NAND U145 ( .A(n17), .B(opcode[18]), .Z(n55) );
  NAND U146 ( .A(n22), .B(opcode[18]), .Z(n54) );
  NAND U147 ( .A(n56), .B(n24), .Z(n46) );
  NAND U148 ( .A(n57), .B(n58), .Z(n56) );
  NAND U149 ( .A(n27), .B(opcode[18]), .Z(n58) );
  NAND U150 ( .A(n28), .B(opcode[18]), .Z(n57) );
  NAND U151 ( .A(n59), .B(n60), .Z(rt_index[1]) );
  NAND U152 ( .A(n3), .B(opcode[17]), .Z(n60) );
  AND U153 ( .A(n61), .B(n62), .Z(n59) );
  NAND U154 ( .A(n63), .B(n7), .Z(n62) );
  NAND U155 ( .A(n64), .B(n65), .Z(n63) );
  NAND U156 ( .A(n10), .B(n66), .Z(n65) );
  NAND U157 ( .A(n67), .B(n68), .Z(n66) );
  NAND U158 ( .A(imm[1]), .B(opcode[17]), .Z(n68) );
  NAND U159 ( .A(n14), .B(opcode[17]), .Z(n67) );
  AND U160 ( .A(n69), .B(n70), .Z(n64) );
  NAND U161 ( .A(n17), .B(opcode[17]), .Z(n70) );
  NAND U162 ( .A(n22), .B(opcode[17]), .Z(n69) );
  NAND U163 ( .A(n71), .B(n24), .Z(n61) );
  NAND U164 ( .A(n72), .B(n73), .Z(n71) );
  NAND U165 ( .A(n27), .B(opcode[17]), .Z(n73) );
  NAND U166 ( .A(n28), .B(opcode[17]), .Z(n72) );
  NAND U167 ( .A(n74), .B(n75), .Z(rt_index[0]) );
  NAND U168 ( .A(n3), .B(opcode[16]), .Z(n75) );
  AND U169 ( .A(n76), .B(n77), .Z(n74) );
  NAND U170 ( .A(n78), .B(n7), .Z(n77) );
  NAND U171 ( .A(n79), .B(n80), .Z(n78) );
  NAND U172 ( .A(n10), .B(n81), .Z(n80) );
  NAND U173 ( .A(n82), .B(n83), .Z(n81) );
  NAND U174 ( .A(imm[1]), .B(opcode[16]), .Z(n83) );
  NAND U175 ( .A(n14), .B(opcode[16]), .Z(n82) );
  AND U176 ( .A(n84), .B(n85), .Z(n79) );
  NAND U177 ( .A(n17), .B(n86), .Z(n85) );
  NAND U178 ( .A(n87), .B(n88), .Z(n86) );
  NANDN U179 ( .A(n21), .B(opcode[16]), .Z(n88) );
  NAND U180 ( .A(opcode[19]), .B(opcode[16]), .Z(n87) );
  NAND U181 ( .A(opcode[16]), .B(n22), .Z(n84) );
  NANDN U182 ( .A(n89), .B(n90), .Z(n22) );
  NAND U183 ( .A(n91), .B(n24), .Z(n76) );
  NAND U184 ( .A(n92), .B(n93), .Z(n91) );
  NAND U185 ( .A(n27), .B(opcode[16]), .Z(n93) );
  NAND U186 ( .A(opcode[16]), .B(n28), .Z(n92) );
  NAND U187 ( .A(n94), .B(n95), .Z(rs_index[4]) );
  AND U188 ( .A(n96), .B(n97), .Z(n94) );
  IV U189 ( .A(opcode[25]), .Z(n97) );
  NAND U190 ( .A(n98), .B(n99), .Z(n96) );
  MUX U191 ( .A(opcode[20]), .B(imm[15]), .S(n100), .Z(n99) );
  NAND U192 ( .A(n101), .B(n102), .Z(rs_index[3]) );
  NAND U193 ( .A(n98), .B(n103), .Z(n102) );
  MUX U194 ( .A(opcode[19]), .B(imm[14]), .S(n100), .Z(n103) );
  ANDN U195 ( .B(n95), .A(opcode[24]), .Z(n101) );
  NAND U196 ( .A(n104), .B(n105), .Z(rs_index[2]) );
  NAND U197 ( .A(n106), .B(n7), .Z(n105) );
  NAND U198 ( .A(n100), .B(n107), .Z(n106) );
  NAND U199 ( .A(n108), .B(n109), .Z(n107) );
  AND U200 ( .A(n110), .B(n10), .Z(n109) );
  AND U201 ( .A(n111), .B(n112), .Z(n104) );
  NAND U202 ( .A(n113), .B(n24), .Z(n112) );
  NAND U203 ( .A(n114), .B(n115), .Z(n113) );
  NAND U204 ( .A(n10), .B(n116), .Z(n115) );
  NAND U205 ( .A(n117), .B(n118), .Z(n116) );
  NAND U206 ( .A(n119), .B(n120), .Z(n118) );
  MUX U207 ( .A(opcode[18]), .B(imm[13]), .S(n100), .Z(n119) );
  NAND U208 ( .A(opcode[23]), .B(n27), .Z(n117) );
  NANDN U209 ( .A(n121), .B(n122), .Z(n27) );
  NAND U210 ( .A(opcode[23]), .B(n28), .Z(n114) );
  NAND U211 ( .A(n123), .B(n124), .Z(n28) );
  AND U212 ( .A(n125), .B(n126), .Z(n124) );
  AND U213 ( .A(n127), .B(n128), .Z(n126) );
  AND U214 ( .A(n90), .B(n129), .Z(n123) );
  AND U215 ( .A(n130), .B(n131), .Z(n129) );
  NAND U216 ( .A(opcode[23]), .B(n3), .Z(n111) );
  NANDN U217 ( .A(opcode[29]), .B(n132), .Z(n3) );
  NAND U218 ( .A(n133), .B(n134), .Z(rs_index[1]) );
  NAND U219 ( .A(n98), .B(n135), .Z(n134) );
  MUX U220 ( .A(opcode[17]), .B(imm[12]), .S(n100), .Z(n135) );
  AND U221 ( .A(n95), .B(n136), .Z(n133) );
  IV U222 ( .A(opcode[22]), .Z(n136) );
  NAND U223 ( .A(n137), .B(n138), .Z(rs_index[0]) );
  NAND U224 ( .A(n98), .B(n139), .Z(n138) );
  MUX U225 ( .A(opcode[16]), .B(imm[11]), .S(n100), .Z(n139) );
  ANDN U226 ( .B(n95), .A(opcode[21]), .Z(n137) );
  NAND U227 ( .A(n140), .B(n141), .Z(n95) );
  AND U228 ( .A(n7), .B(n10), .Z(n141) );
  AND U229 ( .A(n110), .B(n108), .Z(n140) );
  MUX U230 ( .A(n142), .B(\Reg_Bank/registers[31][31] ), .S(n143), .Z(
        \Reg_Bank/n4021 ) );
  MUX U231 ( .A(n144), .B(\Reg_Bank/registers[31][30] ), .S(n143), .Z(
        \Reg_Bank/n4020 ) );
  MUX U232 ( .A(n145), .B(\Reg_Bank/registers[31][29] ), .S(n143), .Z(
        \Reg_Bank/n4019 ) );
  MUX U233 ( .A(n146), .B(\Reg_Bank/registers[31][28] ), .S(n143), .Z(
        \Reg_Bank/n4018 ) );
  MUX U234 ( .A(n147), .B(\Reg_Bank/registers[31][27] ), .S(n143), .Z(
        \Reg_Bank/n4017 ) );
  MUX U235 ( .A(n148), .B(\Reg_Bank/registers[31][26] ), .S(n143), .Z(
        \Reg_Bank/n4016 ) );
  MUX U236 ( .A(n149), .B(\Reg_Bank/registers[31][25] ), .S(n143), .Z(
        \Reg_Bank/n4015 ) );
  MUX U237 ( .A(n150), .B(\Reg_Bank/registers[31][24] ), .S(n143), .Z(
        \Reg_Bank/n4014 ) );
  MUX U238 ( .A(n151), .B(\Reg_Bank/registers[31][23] ), .S(n143), .Z(
        \Reg_Bank/n4013 ) );
  MUX U239 ( .A(n152), .B(\Reg_Bank/registers[31][22] ), .S(n143), .Z(
        \Reg_Bank/n4012 ) );
  MUX U240 ( .A(n153), .B(\Reg_Bank/registers[31][21] ), .S(n143), .Z(
        \Reg_Bank/n4011 ) );
  MUX U241 ( .A(n154), .B(\Reg_Bank/registers[31][20] ), .S(n143), .Z(
        \Reg_Bank/n4010 ) );
  MUX U242 ( .A(n155), .B(\Reg_Bank/registers[31][19] ), .S(n143), .Z(
        \Reg_Bank/n4009 ) );
  MUX U243 ( .A(n156), .B(\Reg_Bank/registers[31][18] ), .S(n143), .Z(
        \Reg_Bank/n4008 ) );
  MUX U244 ( .A(n157), .B(\Reg_Bank/registers[31][17] ), .S(n143), .Z(
        \Reg_Bank/n4007 ) );
  MUX U245 ( .A(n158), .B(\Reg_Bank/registers[31][16] ), .S(n143), .Z(
        \Reg_Bank/n4006 ) );
  MUX U246 ( .A(n159), .B(\Reg_Bank/registers[31][15] ), .S(n143), .Z(
        \Reg_Bank/n4005 ) );
  MUX U247 ( .A(n160), .B(\Reg_Bank/registers[31][14] ), .S(n143), .Z(
        \Reg_Bank/n4004 ) );
  MUX U248 ( .A(n161), .B(\Reg_Bank/registers[31][13] ), .S(n143), .Z(
        \Reg_Bank/n4003 ) );
  MUX U249 ( .A(n162), .B(\Reg_Bank/registers[31][12] ), .S(n143), .Z(
        \Reg_Bank/n4002 ) );
  MUX U250 ( .A(n163), .B(\Reg_Bank/registers[31][11] ), .S(n143), .Z(
        \Reg_Bank/n4001 ) );
  MUX U251 ( .A(n164), .B(\Reg_Bank/registers[31][10] ), .S(n143), .Z(
        \Reg_Bank/n4000 ) );
  MUX U252 ( .A(n165), .B(\Reg_Bank/registers[31][9] ), .S(n143), .Z(
        \Reg_Bank/n3999 ) );
  MUX U253 ( .A(n166), .B(\Reg_Bank/registers[31][8] ), .S(n143), .Z(
        \Reg_Bank/n3998 ) );
  MUX U254 ( .A(n167), .B(\Reg_Bank/registers[31][7] ), .S(n143), .Z(
        \Reg_Bank/n3997 ) );
  MUX U255 ( .A(n168), .B(\Reg_Bank/registers[31][6] ), .S(n143), .Z(
        \Reg_Bank/n3996 ) );
  MUX U256 ( .A(n169), .B(\Reg_Bank/registers[31][5] ), .S(n143), .Z(
        \Reg_Bank/n3995 ) );
  MUX U257 ( .A(n170), .B(\Reg_Bank/registers[31][4] ), .S(n143), .Z(
        \Reg_Bank/n3994 ) );
  MUX U258 ( .A(n171), .B(\Reg_Bank/registers[31][3] ), .S(n143), .Z(
        \Reg_Bank/n3993 ) );
  MUX U259 ( .A(n172), .B(\Reg_Bank/registers[31][2] ), .S(n143), .Z(
        \Reg_Bank/n3992 ) );
  IV U260 ( .A(n173), .Z(n143) );
  MUX U261 ( .A(\Reg_Bank/registers[31][1] ), .B(n174), .S(n173), .Z(
        \Reg_Bank/n3991 ) );
  MUX U262 ( .A(\Reg_Bank/registers[31][0] ), .B(n175), .S(n173), .Z(
        \Reg_Bank/n3990 ) );
  ANDN U263 ( .B(n176), .A(n177), .Z(n173) );
  MUX U264 ( .A(n142), .B(\Reg_Bank/registers[30][31] ), .S(n178), .Z(
        \Reg_Bank/n3989 ) );
  MUX U265 ( .A(n144), .B(\Reg_Bank/registers[30][30] ), .S(n178), .Z(
        \Reg_Bank/n3988 ) );
  MUX U266 ( .A(n145), .B(\Reg_Bank/registers[30][29] ), .S(n178), .Z(
        \Reg_Bank/n3987 ) );
  MUX U267 ( .A(n146), .B(\Reg_Bank/registers[30][28] ), .S(n178), .Z(
        \Reg_Bank/n3986 ) );
  MUX U268 ( .A(n147), .B(\Reg_Bank/registers[30][27] ), .S(n178), .Z(
        \Reg_Bank/n3985 ) );
  MUX U269 ( .A(n148), .B(\Reg_Bank/registers[30][26] ), .S(n178), .Z(
        \Reg_Bank/n3984 ) );
  MUX U270 ( .A(n149), .B(\Reg_Bank/registers[30][25] ), .S(n178), .Z(
        \Reg_Bank/n3983 ) );
  MUX U271 ( .A(n150), .B(\Reg_Bank/registers[30][24] ), .S(n178), .Z(
        \Reg_Bank/n3982 ) );
  MUX U272 ( .A(n151), .B(\Reg_Bank/registers[30][23] ), .S(n178), .Z(
        \Reg_Bank/n3981 ) );
  MUX U273 ( .A(n152), .B(\Reg_Bank/registers[30][22] ), .S(n178), .Z(
        \Reg_Bank/n3980 ) );
  MUX U274 ( .A(n153), .B(\Reg_Bank/registers[30][21] ), .S(n178), .Z(
        \Reg_Bank/n3979 ) );
  MUX U275 ( .A(n154), .B(\Reg_Bank/registers[30][20] ), .S(n178), .Z(
        \Reg_Bank/n3978 ) );
  MUX U276 ( .A(n155), .B(\Reg_Bank/registers[30][19] ), .S(n178), .Z(
        \Reg_Bank/n3977 ) );
  MUX U277 ( .A(n156), .B(\Reg_Bank/registers[30][18] ), .S(n178), .Z(
        \Reg_Bank/n3976 ) );
  MUX U278 ( .A(n157), .B(\Reg_Bank/registers[30][17] ), .S(n178), .Z(
        \Reg_Bank/n3975 ) );
  MUX U279 ( .A(n158), .B(\Reg_Bank/registers[30][16] ), .S(n178), .Z(
        \Reg_Bank/n3974 ) );
  MUX U280 ( .A(n159), .B(\Reg_Bank/registers[30][15] ), .S(n178), .Z(
        \Reg_Bank/n3973 ) );
  MUX U281 ( .A(n160), .B(\Reg_Bank/registers[30][14] ), .S(n178), .Z(
        \Reg_Bank/n3972 ) );
  MUX U282 ( .A(n161), .B(\Reg_Bank/registers[30][13] ), .S(n178), .Z(
        \Reg_Bank/n3971 ) );
  MUX U283 ( .A(n162), .B(\Reg_Bank/registers[30][12] ), .S(n178), .Z(
        \Reg_Bank/n3970 ) );
  MUX U284 ( .A(n163), .B(\Reg_Bank/registers[30][11] ), .S(n178), .Z(
        \Reg_Bank/n3969 ) );
  MUX U285 ( .A(n164), .B(\Reg_Bank/registers[30][10] ), .S(n178), .Z(
        \Reg_Bank/n3968 ) );
  MUX U286 ( .A(n165), .B(\Reg_Bank/registers[30][9] ), .S(n178), .Z(
        \Reg_Bank/n3967 ) );
  MUX U287 ( .A(n166), .B(\Reg_Bank/registers[30][8] ), .S(n178), .Z(
        \Reg_Bank/n3966 ) );
  MUX U288 ( .A(n167), .B(\Reg_Bank/registers[30][7] ), .S(n178), .Z(
        \Reg_Bank/n3965 ) );
  MUX U289 ( .A(n168), .B(\Reg_Bank/registers[30][6] ), .S(n178), .Z(
        \Reg_Bank/n3964 ) );
  MUX U290 ( .A(n169), .B(\Reg_Bank/registers[30][5] ), .S(n178), .Z(
        \Reg_Bank/n3963 ) );
  MUX U291 ( .A(n170), .B(\Reg_Bank/registers[30][4] ), .S(n178), .Z(
        \Reg_Bank/n3962 ) );
  MUX U292 ( .A(n171), .B(\Reg_Bank/registers[30][3] ), .S(n178), .Z(
        \Reg_Bank/n3961 ) );
  MUX U293 ( .A(n172), .B(\Reg_Bank/registers[30][2] ), .S(n178), .Z(
        \Reg_Bank/n3960 ) );
  IV U294 ( .A(n179), .Z(n178) );
  MUX U295 ( .A(\Reg_Bank/registers[30][1] ), .B(n174), .S(n179), .Z(
        \Reg_Bank/n3959 ) );
  MUX U296 ( .A(\Reg_Bank/registers[30][0] ), .B(n175), .S(n179), .Z(
        \Reg_Bank/n3958 ) );
  AND U297 ( .A(n176), .B(n180), .Z(n179) );
  MUX U298 ( .A(n142), .B(\Reg_Bank/registers[29][31] ), .S(n181), .Z(
        \Reg_Bank/n3957 ) );
  MUX U299 ( .A(n144), .B(\Reg_Bank/registers[29][30] ), .S(n181), .Z(
        \Reg_Bank/n3956 ) );
  MUX U300 ( .A(n145), .B(\Reg_Bank/registers[29][29] ), .S(n181), .Z(
        \Reg_Bank/n3955 ) );
  MUX U301 ( .A(n146), .B(\Reg_Bank/registers[29][28] ), .S(n181), .Z(
        \Reg_Bank/n3954 ) );
  MUX U302 ( .A(n147), .B(\Reg_Bank/registers[29][27] ), .S(n181), .Z(
        \Reg_Bank/n3953 ) );
  MUX U303 ( .A(n148), .B(\Reg_Bank/registers[29][26] ), .S(n181), .Z(
        \Reg_Bank/n3952 ) );
  MUX U304 ( .A(n149), .B(\Reg_Bank/registers[29][25] ), .S(n181), .Z(
        \Reg_Bank/n3951 ) );
  MUX U305 ( .A(n150), .B(\Reg_Bank/registers[29][24] ), .S(n181), .Z(
        \Reg_Bank/n3950 ) );
  MUX U306 ( .A(n151), .B(\Reg_Bank/registers[29][23] ), .S(n181), .Z(
        \Reg_Bank/n3949 ) );
  MUX U307 ( .A(n152), .B(\Reg_Bank/registers[29][22] ), .S(n181), .Z(
        \Reg_Bank/n3948 ) );
  MUX U308 ( .A(n153), .B(\Reg_Bank/registers[29][21] ), .S(n181), .Z(
        \Reg_Bank/n3947 ) );
  MUX U309 ( .A(n154), .B(\Reg_Bank/registers[29][20] ), .S(n181), .Z(
        \Reg_Bank/n3946 ) );
  MUX U310 ( .A(n155), .B(\Reg_Bank/registers[29][19] ), .S(n181), .Z(
        \Reg_Bank/n3945 ) );
  MUX U311 ( .A(n156), .B(\Reg_Bank/registers[29][18] ), .S(n181), .Z(
        \Reg_Bank/n3944 ) );
  MUX U312 ( .A(n157), .B(\Reg_Bank/registers[29][17] ), .S(n181), .Z(
        \Reg_Bank/n3943 ) );
  MUX U313 ( .A(n158), .B(\Reg_Bank/registers[29][16] ), .S(n181), .Z(
        \Reg_Bank/n3942 ) );
  MUX U314 ( .A(n159), .B(\Reg_Bank/registers[29][15] ), .S(n181), .Z(
        \Reg_Bank/n3941 ) );
  MUX U315 ( .A(n160), .B(\Reg_Bank/registers[29][14] ), .S(n181), .Z(
        \Reg_Bank/n3940 ) );
  MUX U316 ( .A(n161), .B(\Reg_Bank/registers[29][13] ), .S(n181), .Z(
        \Reg_Bank/n3939 ) );
  MUX U317 ( .A(n162), .B(\Reg_Bank/registers[29][12] ), .S(n181), .Z(
        \Reg_Bank/n3938 ) );
  MUX U318 ( .A(n163), .B(\Reg_Bank/registers[29][11] ), .S(n181), .Z(
        \Reg_Bank/n3937 ) );
  MUX U319 ( .A(n164), .B(\Reg_Bank/registers[29][10] ), .S(n181), .Z(
        \Reg_Bank/n3936 ) );
  MUX U320 ( .A(n165), .B(\Reg_Bank/registers[29][9] ), .S(n181), .Z(
        \Reg_Bank/n3935 ) );
  MUX U321 ( .A(n166), .B(\Reg_Bank/registers[29][8] ), .S(n181), .Z(
        \Reg_Bank/n3934 ) );
  MUX U322 ( .A(n167), .B(\Reg_Bank/registers[29][7] ), .S(n181), .Z(
        \Reg_Bank/n3933 ) );
  MUX U323 ( .A(n168), .B(\Reg_Bank/registers[29][6] ), .S(n181), .Z(
        \Reg_Bank/n3932 ) );
  MUX U324 ( .A(n169), .B(\Reg_Bank/registers[29][5] ), .S(n181), .Z(
        \Reg_Bank/n3931 ) );
  MUX U325 ( .A(n170), .B(\Reg_Bank/registers[29][4] ), .S(n181), .Z(
        \Reg_Bank/n3930 ) );
  MUX U326 ( .A(n171), .B(\Reg_Bank/registers[29][3] ), .S(n181), .Z(
        \Reg_Bank/n3929 ) );
  MUX U327 ( .A(n172), .B(\Reg_Bank/registers[29][2] ), .S(n181), .Z(
        \Reg_Bank/n3928 ) );
  IV U328 ( .A(n182), .Z(n181) );
  MUX U329 ( .A(\Reg_Bank/registers[29][1] ), .B(n174), .S(n182), .Z(
        \Reg_Bank/n3927 ) );
  MUX U330 ( .A(\Reg_Bank/registers[29][0] ), .B(n175), .S(n182), .Z(
        \Reg_Bank/n3926 ) );
  AND U331 ( .A(n176), .B(n183), .Z(n182) );
  MUX U332 ( .A(n142), .B(\Reg_Bank/registers[28][31] ), .S(n184), .Z(
        \Reg_Bank/n3925 ) );
  MUX U333 ( .A(n144), .B(\Reg_Bank/registers[28][30] ), .S(n184), .Z(
        \Reg_Bank/n3924 ) );
  MUX U334 ( .A(n145), .B(\Reg_Bank/registers[28][29] ), .S(n184), .Z(
        \Reg_Bank/n3923 ) );
  MUX U335 ( .A(n146), .B(\Reg_Bank/registers[28][28] ), .S(n184), .Z(
        \Reg_Bank/n3922 ) );
  MUX U336 ( .A(n147), .B(\Reg_Bank/registers[28][27] ), .S(n184), .Z(
        \Reg_Bank/n3921 ) );
  MUX U337 ( .A(n148), .B(\Reg_Bank/registers[28][26] ), .S(n184), .Z(
        \Reg_Bank/n3920 ) );
  MUX U338 ( .A(n149), .B(\Reg_Bank/registers[28][25] ), .S(n184), .Z(
        \Reg_Bank/n3919 ) );
  MUX U339 ( .A(n150), .B(\Reg_Bank/registers[28][24] ), .S(n184), .Z(
        \Reg_Bank/n3918 ) );
  MUX U340 ( .A(n151), .B(\Reg_Bank/registers[28][23] ), .S(n184), .Z(
        \Reg_Bank/n3917 ) );
  MUX U341 ( .A(n152), .B(\Reg_Bank/registers[28][22] ), .S(n184), .Z(
        \Reg_Bank/n3916 ) );
  MUX U342 ( .A(n153), .B(\Reg_Bank/registers[28][21] ), .S(n184), .Z(
        \Reg_Bank/n3915 ) );
  MUX U343 ( .A(n154), .B(\Reg_Bank/registers[28][20] ), .S(n184), .Z(
        \Reg_Bank/n3914 ) );
  MUX U344 ( .A(n155), .B(\Reg_Bank/registers[28][19] ), .S(n184), .Z(
        \Reg_Bank/n3913 ) );
  MUX U345 ( .A(n156), .B(\Reg_Bank/registers[28][18] ), .S(n184), .Z(
        \Reg_Bank/n3912 ) );
  MUX U346 ( .A(n157), .B(\Reg_Bank/registers[28][17] ), .S(n184), .Z(
        \Reg_Bank/n3911 ) );
  MUX U347 ( .A(n158), .B(\Reg_Bank/registers[28][16] ), .S(n184), .Z(
        \Reg_Bank/n3910 ) );
  MUX U348 ( .A(n159), .B(\Reg_Bank/registers[28][15] ), .S(n184), .Z(
        \Reg_Bank/n3909 ) );
  MUX U349 ( .A(n160), .B(\Reg_Bank/registers[28][14] ), .S(n184), .Z(
        \Reg_Bank/n3908 ) );
  MUX U350 ( .A(n161), .B(\Reg_Bank/registers[28][13] ), .S(n184), .Z(
        \Reg_Bank/n3907 ) );
  MUX U351 ( .A(n162), .B(\Reg_Bank/registers[28][12] ), .S(n184), .Z(
        \Reg_Bank/n3906 ) );
  MUX U352 ( .A(n163), .B(\Reg_Bank/registers[28][11] ), .S(n184), .Z(
        \Reg_Bank/n3905 ) );
  MUX U353 ( .A(n164), .B(\Reg_Bank/registers[28][10] ), .S(n184), .Z(
        \Reg_Bank/n3904 ) );
  MUX U354 ( .A(n165), .B(\Reg_Bank/registers[28][9] ), .S(n184), .Z(
        \Reg_Bank/n3903 ) );
  MUX U355 ( .A(n166), .B(\Reg_Bank/registers[28][8] ), .S(n184), .Z(
        \Reg_Bank/n3902 ) );
  MUX U356 ( .A(n167), .B(\Reg_Bank/registers[28][7] ), .S(n184), .Z(
        \Reg_Bank/n3901 ) );
  MUX U357 ( .A(n168), .B(\Reg_Bank/registers[28][6] ), .S(n184), .Z(
        \Reg_Bank/n3900 ) );
  MUX U358 ( .A(n169), .B(\Reg_Bank/registers[28][5] ), .S(n184), .Z(
        \Reg_Bank/n3899 ) );
  MUX U359 ( .A(n170), .B(\Reg_Bank/registers[28][4] ), .S(n184), .Z(
        \Reg_Bank/n3898 ) );
  MUX U360 ( .A(n171), .B(\Reg_Bank/registers[28][3] ), .S(n184), .Z(
        \Reg_Bank/n3897 ) );
  MUX U361 ( .A(n172), .B(\Reg_Bank/registers[28][2] ), .S(n184), .Z(
        \Reg_Bank/n3896 ) );
  IV U362 ( .A(n185), .Z(n184) );
  MUX U363 ( .A(\Reg_Bank/registers[28][1] ), .B(n174), .S(n185), .Z(
        \Reg_Bank/n3895 ) );
  MUX U364 ( .A(\Reg_Bank/registers[28][0] ), .B(n175), .S(n185), .Z(
        \Reg_Bank/n3894 ) );
  AND U365 ( .A(n176), .B(n186), .Z(n185) );
  MUX U366 ( .A(\Reg_Bank/registers[27][31] ), .B(n142), .S(n187), .Z(
        \Reg_Bank/n3893 ) );
  MUX U367 ( .A(\Reg_Bank/registers[27][30] ), .B(n144), .S(n187), .Z(
        \Reg_Bank/n3892 ) );
  MUX U368 ( .A(\Reg_Bank/registers[27][29] ), .B(n145), .S(n187), .Z(
        \Reg_Bank/n3891 ) );
  MUX U369 ( .A(\Reg_Bank/registers[27][28] ), .B(n146), .S(n187), .Z(
        \Reg_Bank/n3890 ) );
  MUX U370 ( .A(\Reg_Bank/registers[27][27] ), .B(n147), .S(n187), .Z(
        \Reg_Bank/n3889 ) );
  MUX U371 ( .A(\Reg_Bank/registers[27][26] ), .B(n148), .S(n187), .Z(
        \Reg_Bank/n3888 ) );
  MUX U372 ( .A(\Reg_Bank/registers[27][25] ), .B(n149), .S(n187), .Z(
        \Reg_Bank/n3887 ) );
  MUX U373 ( .A(\Reg_Bank/registers[27][24] ), .B(n150), .S(n187), .Z(
        \Reg_Bank/n3886 ) );
  MUX U374 ( .A(\Reg_Bank/registers[27][23] ), .B(n151), .S(n187), .Z(
        \Reg_Bank/n3885 ) );
  MUX U375 ( .A(\Reg_Bank/registers[27][22] ), .B(n152), .S(n187), .Z(
        \Reg_Bank/n3884 ) );
  MUX U376 ( .A(\Reg_Bank/registers[27][21] ), .B(n153), .S(n187), .Z(
        \Reg_Bank/n3883 ) );
  MUX U377 ( .A(\Reg_Bank/registers[27][20] ), .B(n154), .S(n187), .Z(
        \Reg_Bank/n3882 ) );
  MUX U378 ( .A(\Reg_Bank/registers[27][19] ), .B(n155), .S(n187), .Z(
        \Reg_Bank/n3881 ) );
  MUX U379 ( .A(\Reg_Bank/registers[27][18] ), .B(n156), .S(n187), .Z(
        \Reg_Bank/n3880 ) );
  MUX U380 ( .A(\Reg_Bank/registers[27][17] ), .B(n157), .S(n187), .Z(
        \Reg_Bank/n3879 ) );
  MUX U381 ( .A(\Reg_Bank/registers[27][16] ), .B(n158), .S(n187), .Z(
        \Reg_Bank/n3878 ) );
  MUX U382 ( .A(\Reg_Bank/registers[27][15] ), .B(n159), .S(n187), .Z(
        \Reg_Bank/n3877 ) );
  MUX U383 ( .A(\Reg_Bank/registers[27][14] ), .B(n160), .S(n187), .Z(
        \Reg_Bank/n3876 ) );
  MUX U384 ( .A(\Reg_Bank/registers[27][13] ), .B(n161), .S(n187), .Z(
        \Reg_Bank/n3875 ) );
  MUX U385 ( .A(\Reg_Bank/registers[27][12] ), .B(n162), .S(n187), .Z(
        \Reg_Bank/n3874 ) );
  MUX U386 ( .A(\Reg_Bank/registers[27][11] ), .B(n163), .S(n187), .Z(
        \Reg_Bank/n3873 ) );
  MUX U387 ( .A(\Reg_Bank/registers[27][10] ), .B(n164), .S(n187), .Z(
        \Reg_Bank/n3872 ) );
  MUX U388 ( .A(\Reg_Bank/registers[27][9] ), .B(n165), .S(n187), .Z(
        \Reg_Bank/n3871 ) );
  MUX U389 ( .A(\Reg_Bank/registers[27][8] ), .B(n166), .S(n187), .Z(
        \Reg_Bank/n3870 ) );
  MUX U390 ( .A(\Reg_Bank/registers[27][7] ), .B(n167), .S(n187), .Z(
        \Reg_Bank/n3869 ) );
  MUX U391 ( .A(\Reg_Bank/registers[27][6] ), .B(n168), .S(n187), .Z(
        \Reg_Bank/n3868 ) );
  MUX U392 ( .A(\Reg_Bank/registers[27][5] ), .B(n169), .S(n187), .Z(
        \Reg_Bank/n3867 ) );
  MUX U393 ( .A(\Reg_Bank/registers[27][4] ), .B(n170), .S(n187), .Z(
        \Reg_Bank/n3866 ) );
  MUX U394 ( .A(\Reg_Bank/registers[27][3] ), .B(n171), .S(n187), .Z(
        \Reg_Bank/n3865 ) );
  MUX U395 ( .A(\Reg_Bank/registers[27][2] ), .B(n172), .S(n187), .Z(
        \Reg_Bank/n3864 ) );
  MUX U396 ( .A(\Reg_Bank/registers[27][1] ), .B(n174), .S(n187), .Z(
        \Reg_Bank/n3863 ) );
  MUX U397 ( .A(\Reg_Bank/registers[27][0] ), .B(n175), .S(n187), .Z(
        \Reg_Bank/n3862 ) );
  AND U398 ( .A(n176), .B(n188), .Z(n187) );
  MUX U399 ( .A(\Reg_Bank/registers[26][31] ), .B(n142), .S(n189), .Z(
        \Reg_Bank/n3861 ) );
  MUX U400 ( .A(\Reg_Bank/registers[26][30] ), .B(n144), .S(n189), .Z(
        \Reg_Bank/n3860 ) );
  MUX U401 ( .A(\Reg_Bank/registers[26][29] ), .B(n145), .S(n189), .Z(
        \Reg_Bank/n3859 ) );
  MUX U402 ( .A(\Reg_Bank/registers[26][28] ), .B(n146), .S(n189), .Z(
        \Reg_Bank/n3858 ) );
  MUX U403 ( .A(\Reg_Bank/registers[26][27] ), .B(n147), .S(n189), .Z(
        \Reg_Bank/n3857 ) );
  MUX U404 ( .A(\Reg_Bank/registers[26][26] ), .B(n148), .S(n189), .Z(
        \Reg_Bank/n3856 ) );
  MUX U405 ( .A(\Reg_Bank/registers[26][25] ), .B(n149), .S(n189), .Z(
        \Reg_Bank/n3855 ) );
  MUX U406 ( .A(\Reg_Bank/registers[26][24] ), .B(n150), .S(n189), .Z(
        \Reg_Bank/n3854 ) );
  MUX U407 ( .A(\Reg_Bank/registers[26][23] ), .B(n151), .S(n189), .Z(
        \Reg_Bank/n3853 ) );
  MUX U408 ( .A(\Reg_Bank/registers[26][22] ), .B(n152), .S(n189), .Z(
        \Reg_Bank/n3852 ) );
  MUX U409 ( .A(\Reg_Bank/registers[26][21] ), .B(n153), .S(n189), .Z(
        \Reg_Bank/n3851 ) );
  MUX U410 ( .A(\Reg_Bank/registers[26][20] ), .B(n154), .S(n189), .Z(
        \Reg_Bank/n3850 ) );
  MUX U411 ( .A(\Reg_Bank/registers[26][19] ), .B(n155), .S(n189), .Z(
        \Reg_Bank/n3849 ) );
  MUX U412 ( .A(\Reg_Bank/registers[26][18] ), .B(n156), .S(n189), .Z(
        \Reg_Bank/n3848 ) );
  MUX U413 ( .A(\Reg_Bank/registers[26][17] ), .B(n157), .S(n189), .Z(
        \Reg_Bank/n3847 ) );
  MUX U414 ( .A(\Reg_Bank/registers[26][16] ), .B(n158), .S(n189), .Z(
        \Reg_Bank/n3846 ) );
  MUX U415 ( .A(\Reg_Bank/registers[26][15] ), .B(n159), .S(n189), .Z(
        \Reg_Bank/n3845 ) );
  MUX U416 ( .A(\Reg_Bank/registers[26][14] ), .B(n160), .S(n189), .Z(
        \Reg_Bank/n3844 ) );
  MUX U417 ( .A(\Reg_Bank/registers[26][13] ), .B(n161), .S(n189), .Z(
        \Reg_Bank/n3843 ) );
  MUX U418 ( .A(\Reg_Bank/registers[26][12] ), .B(n162), .S(n189), .Z(
        \Reg_Bank/n3842 ) );
  MUX U419 ( .A(\Reg_Bank/registers[26][11] ), .B(n163), .S(n189), .Z(
        \Reg_Bank/n3841 ) );
  MUX U420 ( .A(\Reg_Bank/registers[26][10] ), .B(n164), .S(n189), .Z(
        \Reg_Bank/n3840 ) );
  MUX U421 ( .A(\Reg_Bank/registers[26][9] ), .B(n165), .S(n189), .Z(
        \Reg_Bank/n3839 ) );
  MUX U422 ( .A(\Reg_Bank/registers[26][8] ), .B(n166), .S(n189), .Z(
        \Reg_Bank/n3838 ) );
  MUX U423 ( .A(\Reg_Bank/registers[26][7] ), .B(n167), .S(n189), .Z(
        \Reg_Bank/n3837 ) );
  MUX U424 ( .A(\Reg_Bank/registers[26][6] ), .B(n168), .S(n189), .Z(
        \Reg_Bank/n3836 ) );
  MUX U425 ( .A(\Reg_Bank/registers[26][5] ), .B(n169), .S(n189), .Z(
        \Reg_Bank/n3835 ) );
  MUX U426 ( .A(\Reg_Bank/registers[26][4] ), .B(n170), .S(n189), .Z(
        \Reg_Bank/n3834 ) );
  MUX U427 ( .A(\Reg_Bank/registers[26][3] ), .B(n171), .S(n189), .Z(
        \Reg_Bank/n3833 ) );
  MUX U428 ( .A(\Reg_Bank/registers[26][2] ), .B(n172), .S(n189), .Z(
        \Reg_Bank/n3832 ) );
  MUX U429 ( .A(\Reg_Bank/registers[26][1] ), .B(n174), .S(n189), .Z(
        \Reg_Bank/n3831 ) );
  MUX U430 ( .A(\Reg_Bank/registers[26][0] ), .B(n175), .S(n189), .Z(
        \Reg_Bank/n3830 ) );
  AND U431 ( .A(n176), .B(n190), .Z(n189) );
  MUX U432 ( .A(\Reg_Bank/registers[25][31] ), .B(n142), .S(n191), .Z(
        \Reg_Bank/n3829 ) );
  MUX U433 ( .A(\Reg_Bank/registers[25][30] ), .B(n144), .S(n191), .Z(
        \Reg_Bank/n3828 ) );
  MUX U434 ( .A(\Reg_Bank/registers[25][29] ), .B(n145), .S(n191), .Z(
        \Reg_Bank/n3827 ) );
  MUX U435 ( .A(\Reg_Bank/registers[25][28] ), .B(n146), .S(n191), .Z(
        \Reg_Bank/n3826 ) );
  MUX U436 ( .A(\Reg_Bank/registers[25][27] ), .B(n147), .S(n191), .Z(
        \Reg_Bank/n3825 ) );
  MUX U437 ( .A(\Reg_Bank/registers[25][26] ), .B(n148), .S(n191), .Z(
        \Reg_Bank/n3824 ) );
  MUX U438 ( .A(\Reg_Bank/registers[25][25] ), .B(n149), .S(n191), .Z(
        \Reg_Bank/n3823 ) );
  MUX U439 ( .A(\Reg_Bank/registers[25][24] ), .B(n150), .S(n191), .Z(
        \Reg_Bank/n3822 ) );
  MUX U440 ( .A(\Reg_Bank/registers[25][23] ), .B(n151), .S(n191), .Z(
        \Reg_Bank/n3821 ) );
  MUX U441 ( .A(\Reg_Bank/registers[25][22] ), .B(n152), .S(n191), .Z(
        \Reg_Bank/n3820 ) );
  MUX U442 ( .A(\Reg_Bank/registers[25][21] ), .B(n153), .S(n191), .Z(
        \Reg_Bank/n3819 ) );
  MUX U443 ( .A(\Reg_Bank/registers[25][20] ), .B(n154), .S(n191), .Z(
        \Reg_Bank/n3818 ) );
  MUX U444 ( .A(\Reg_Bank/registers[25][19] ), .B(n155), .S(n191), .Z(
        \Reg_Bank/n3817 ) );
  MUX U445 ( .A(\Reg_Bank/registers[25][18] ), .B(n156), .S(n191), .Z(
        \Reg_Bank/n3816 ) );
  MUX U446 ( .A(\Reg_Bank/registers[25][17] ), .B(n157), .S(n191), .Z(
        \Reg_Bank/n3815 ) );
  MUX U447 ( .A(\Reg_Bank/registers[25][16] ), .B(n158), .S(n191), .Z(
        \Reg_Bank/n3814 ) );
  MUX U448 ( .A(\Reg_Bank/registers[25][15] ), .B(n159), .S(n191), .Z(
        \Reg_Bank/n3813 ) );
  MUX U449 ( .A(\Reg_Bank/registers[25][14] ), .B(n160), .S(n191), .Z(
        \Reg_Bank/n3812 ) );
  MUX U450 ( .A(\Reg_Bank/registers[25][13] ), .B(n161), .S(n191), .Z(
        \Reg_Bank/n3811 ) );
  MUX U451 ( .A(\Reg_Bank/registers[25][12] ), .B(n162), .S(n191), .Z(
        \Reg_Bank/n3810 ) );
  MUX U452 ( .A(\Reg_Bank/registers[25][11] ), .B(n163), .S(n191), .Z(
        \Reg_Bank/n3809 ) );
  MUX U453 ( .A(\Reg_Bank/registers[25][10] ), .B(n164), .S(n191), .Z(
        \Reg_Bank/n3808 ) );
  MUX U454 ( .A(\Reg_Bank/registers[25][9] ), .B(n165), .S(n191), .Z(
        \Reg_Bank/n3807 ) );
  MUX U455 ( .A(\Reg_Bank/registers[25][8] ), .B(n166), .S(n191), .Z(
        \Reg_Bank/n3806 ) );
  MUX U456 ( .A(\Reg_Bank/registers[25][7] ), .B(n167), .S(n191), .Z(
        \Reg_Bank/n3805 ) );
  MUX U457 ( .A(\Reg_Bank/registers[25][6] ), .B(n168), .S(n191), .Z(
        \Reg_Bank/n3804 ) );
  MUX U458 ( .A(\Reg_Bank/registers[25][5] ), .B(n169), .S(n191), .Z(
        \Reg_Bank/n3803 ) );
  MUX U459 ( .A(\Reg_Bank/registers[25][4] ), .B(n170), .S(n191), .Z(
        \Reg_Bank/n3802 ) );
  MUX U460 ( .A(\Reg_Bank/registers[25][3] ), .B(n171), .S(n191), .Z(
        \Reg_Bank/n3801 ) );
  MUX U461 ( .A(\Reg_Bank/registers[25][2] ), .B(n172), .S(n191), .Z(
        \Reg_Bank/n3800 ) );
  MUX U462 ( .A(\Reg_Bank/registers[25][1] ), .B(n174), .S(n191), .Z(
        \Reg_Bank/n3799 ) );
  MUX U463 ( .A(\Reg_Bank/registers[25][0] ), .B(n175), .S(n191), .Z(
        \Reg_Bank/n3798 ) );
  AND U464 ( .A(n176), .B(n192), .Z(n191) );
  MUX U465 ( .A(\Reg_Bank/registers[24][31] ), .B(n142), .S(n193), .Z(
        \Reg_Bank/n3797 ) );
  MUX U466 ( .A(\Reg_Bank/registers[24][30] ), .B(n144), .S(n193), .Z(
        \Reg_Bank/n3796 ) );
  MUX U467 ( .A(\Reg_Bank/registers[24][29] ), .B(n145), .S(n193), .Z(
        \Reg_Bank/n3795 ) );
  MUX U468 ( .A(\Reg_Bank/registers[24][28] ), .B(n146), .S(n193), .Z(
        \Reg_Bank/n3794 ) );
  MUX U469 ( .A(\Reg_Bank/registers[24][27] ), .B(n147), .S(n193), .Z(
        \Reg_Bank/n3793 ) );
  MUX U470 ( .A(\Reg_Bank/registers[24][26] ), .B(n148), .S(n193), .Z(
        \Reg_Bank/n3792 ) );
  MUX U471 ( .A(\Reg_Bank/registers[24][25] ), .B(n149), .S(n193), .Z(
        \Reg_Bank/n3791 ) );
  MUX U472 ( .A(\Reg_Bank/registers[24][24] ), .B(n150), .S(n193), .Z(
        \Reg_Bank/n3790 ) );
  MUX U473 ( .A(\Reg_Bank/registers[24][23] ), .B(n151), .S(n193), .Z(
        \Reg_Bank/n3789 ) );
  MUX U474 ( .A(\Reg_Bank/registers[24][22] ), .B(n152), .S(n193), .Z(
        \Reg_Bank/n3788 ) );
  MUX U475 ( .A(\Reg_Bank/registers[24][21] ), .B(n153), .S(n193), .Z(
        \Reg_Bank/n3787 ) );
  MUX U476 ( .A(\Reg_Bank/registers[24][20] ), .B(n154), .S(n193), .Z(
        \Reg_Bank/n3786 ) );
  MUX U477 ( .A(\Reg_Bank/registers[24][19] ), .B(n155), .S(n193), .Z(
        \Reg_Bank/n3785 ) );
  MUX U478 ( .A(\Reg_Bank/registers[24][18] ), .B(n156), .S(n193), .Z(
        \Reg_Bank/n3784 ) );
  MUX U479 ( .A(\Reg_Bank/registers[24][17] ), .B(n157), .S(n193), .Z(
        \Reg_Bank/n3783 ) );
  MUX U480 ( .A(\Reg_Bank/registers[24][16] ), .B(n158), .S(n193), .Z(
        \Reg_Bank/n3782 ) );
  MUX U481 ( .A(\Reg_Bank/registers[24][15] ), .B(n159), .S(n193), .Z(
        \Reg_Bank/n3781 ) );
  MUX U482 ( .A(\Reg_Bank/registers[24][14] ), .B(n160), .S(n193), .Z(
        \Reg_Bank/n3780 ) );
  MUX U483 ( .A(\Reg_Bank/registers[24][13] ), .B(n161), .S(n193), .Z(
        \Reg_Bank/n3779 ) );
  MUX U484 ( .A(\Reg_Bank/registers[24][12] ), .B(n162), .S(n193), .Z(
        \Reg_Bank/n3778 ) );
  MUX U485 ( .A(\Reg_Bank/registers[24][11] ), .B(n163), .S(n193), .Z(
        \Reg_Bank/n3777 ) );
  MUX U486 ( .A(\Reg_Bank/registers[24][10] ), .B(n164), .S(n193), .Z(
        \Reg_Bank/n3776 ) );
  MUX U487 ( .A(\Reg_Bank/registers[24][9] ), .B(n165), .S(n193), .Z(
        \Reg_Bank/n3775 ) );
  MUX U488 ( .A(\Reg_Bank/registers[24][8] ), .B(n166), .S(n193), .Z(
        \Reg_Bank/n3774 ) );
  MUX U489 ( .A(\Reg_Bank/registers[24][7] ), .B(n167), .S(n193), .Z(
        \Reg_Bank/n3773 ) );
  MUX U490 ( .A(\Reg_Bank/registers[24][6] ), .B(n168), .S(n193), .Z(
        \Reg_Bank/n3772 ) );
  MUX U491 ( .A(\Reg_Bank/registers[24][5] ), .B(n169), .S(n193), .Z(
        \Reg_Bank/n3771 ) );
  MUX U492 ( .A(\Reg_Bank/registers[24][4] ), .B(n170), .S(n193), .Z(
        \Reg_Bank/n3770 ) );
  MUX U493 ( .A(\Reg_Bank/registers[24][3] ), .B(n171), .S(n193), .Z(
        \Reg_Bank/n3769 ) );
  MUX U494 ( .A(\Reg_Bank/registers[24][2] ), .B(n172), .S(n193), .Z(
        \Reg_Bank/n3768 ) );
  MUX U495 ( .A(\Reg_Bank/registers[24][1] ), .B(n174), .S(n193), .Z(
        \Reg_Bank/n3767 ) );
  MUX U496 ( .A(\Reg_Bank/registers[24][0] ), .B(n175), .S(n193), .Z(
        \Reg_Bank/n3766 ) );
  AND U497 ( .A(n176), .B(n194), .Z(n193) );
  ANDN U498 ( .B(n195), .A(n196), .Z(n176) );
  MUX U499 ( .A(\Reg_Bank/registers[23][31] ), .B(n142), .S(n197), .Z(
        \Reg_Bank/n3765 ) );
  MUX U500 ( .A(\Reg_Bank/registers[23][30] ), .B(n144), .S(n197), .Z(
        \Reg_Bank/n3764 ) );
  MUX U501 ( .A(\Reg_Bank/registers[23][29] ), .B(n145), .S(n197), .Z(
        \Reg_Bank/n3763 ) );
  MUX U502 ( .A(\Reg_Bank/registers[23][28] ), .B(n146), .S(n197), .Z(
        \Reg_Bank/n3762 ) );
  MUX U503 ( .A(\Reg_Bank/registers[23][27] ), .B(n147), .S(n197), .Z(
        \Reg_Bank/n3761 ) );
  MUX U504 ( .A(\Reg_Bank/registers[23][26] ), .B(n148), .S(n197), .Z(
        \Reg_Bank/n3760 ) );
  MUX U505 ( .A(\Reg_Bank/registers[23][25] ), .B(n149), .S(n197), .Z(
        \Reg_Bank/n3759 ) );
  MUX U506 ( .A(\Reg_Bank/registers[23][24] ), .B(n150), .S(n197), .Z(
        \Reg_Bank/n3758 ) );
  MUX U507 ( .A(\Reg_Bank/registers[23][23] ), .B(n151), .S(n197), .Z(
        \Reg_Bank/n3757 ) );
  MUX U508 ( .A(\Reg_Bank/registers[23][22] ), .B(n152), .S(n197), .Z(
        \Reg_Bank/n3756 ) );
  MUX U509 ( .A(\Reg_Bank/registers[23][21] ), .B(n153), .S(n197), .Z(
        \Reg_Bank/n3755 ) );
  MUX U510 ( .A(\Reg_Bank/registers[23][20] ), .B(n154), .S(n197), .Z(
        \Reg_Bank/n3754 ) );
  MUX U511 ( .A(\Reg_Bank/registers[23][19] ), .B(n155), .S(n197), .Z(
        \Reg_Bank/n3753 ) );
  MUX U512 ( .A(\Reg_Bank/registers[23][18] ), .B(n156), .S(n197), .Z(
        \Reg_Bank/n3752 ) );
  MUX U513 ( .A(\Reg_Bank/registers[23][17] ), .B(n157), .S(n197), .Z(
        \Reg_Bank/n3751 ) );
  MUX U514 ( .A(\Reg_Bank/registers[23][16] ), .B(n158), .S(n197), .Z(
        \Reg_Bank/n3750 ) );
  MUX U515 ( .A(\Reg_Bank/registers[23][15] ), .B(n159), .S(n197), .Z(
        \Reg_Bank/n3749 ) );
  MUX U516 ( .A(\Reg_Bank/registers[23][14] ), .B(n160), .S(n197), .Z(
        \Reg_Bank/n3748 ) );
  MUX U517 ( .A(\Reg_Bank/registers[23][13] ), .B(n161), .S(n197), .Z(
        \Reg_Bank/n3747 ) );
  MUX U518 ( .A(\Reg_Bank/registers[23][12] ), .B(n162), .S(n197), .Z(
        \Reg_Bank/n3746 ) );
  MUX U519 ( .A(\Reg_Bank/registers[23][11] ), .B(n163), .S(n197), .Z(
        \Reg_Bank/n3745 ) );
  MUX U520 ( .A(\Reg_Bank/registers[23][10] ), .B(n164), .S(n197), .Z(
        \Reg_Bank/n3744 ) );
  MUX U521 ( .A(\Reg_Bank/registers[23][9] ), .B(n165), .S(n197), .Z(
        \Reg_Bank/n3743 ) );
  MUX U522 ( .A(\Reg_Bank/registers[23][8] ), .B(n166), .S(n197), .Z(
        \Reg_Bank/n3742 ) );
  MUX U523 ( .A(\Reg_Bank/registers[23][7] ), .B(n167), .S(n197), .Z(
        \Reg_Bank/n3741 ) );
  MUX U524 ( .A(\Reg_Bank/registers[23][6] ), .B(n168), .S(n197), .Z(
        \Reg_Bank/n3740 ) );
  MUX U525 ( .A(\Reg_Bank/registers[23][5] ), .B(n169), .S(n197), .Z(
        \Reg_Bank/n3739 ) );
  MUX U526 ( .A(\Reg_Bank/registers[23][4] ), .B(n170), .S(n197), .Z(
        \Reg_Bank/n3738 ) );
  MUX U527 ( .A(\Reg_Bank/registers[23][3] ), .B(n171), .S(n197), .Z(
        \Reg_Bank/n3737 ) );
  MUX U528 ( .A(\Reg_Bank/registers[23][2] ), .B(n172), .S(n197), .Z(
        \Reg_Bank/n3736 ) );
  MUX U529 ( .A(\Reg_Bank/registers[23][1] ), .B(n174), .S(n197), .Z(
        \Reg_Bank/n3735 ) );
  MUX U530 ( .A(\Reg_Bank/registers[23][0] ), .B(n175), .S(n197), .Z(
        \Reg_Bank/n3734 ) );
  ANDN U531 ( .B(n198), .A(n177), .Z(n197) );
  MUX U532 ( .A(\Reg_Bank/registers[22][31] ), .B(n142), .S(n199), .Z(
        \Reg_Bank/n3733 ) );
  MUX U533 ( .A(\Reg_Bank/registers[22][30] ), .B(n144), .S(n199), .Z(
        \Reg_Bank/n3732 ) );
  MUX U534 ( .A(\Reg_Bank/registers[22][29] ), .B(n145), .S(n199), .Z(
        \Reg_Bank/n3731 ) );
  MUX U535 ( .A(\Reg_Bank/registers[22][28] ), .B(n146), .S(n199), .Z(
        \Reg_Bank/n3730 ) );
  MUX U536 ( .A(\Reg_Bank/registers[22][27] ), .B(n147), .S(n199), .Z(
        \Reg_Bank/n3729 ) );
  MUX U537 ( .A(\Reg_Bank/registers[22][26] ), .B(n148), .S(n199), .Z(
        \Reg_Bank/n3728 ) );
  MUX U538 ( .A(\Reg_Bank/registers[22][25] ), .B(n149), .S(n199), .Z(
        \Reg_Bank/n3727 ) );
  MUX U539 ( .A(\Reg_Bank/registers[22][24] ), .B(n150), .S(n199), .Z(
        \Reg_Bank/n3726 ) );
  MUX U540 ( .A(\Reg_Bank/registers[22][23] ), .B(n151), .S(n199), .Z(
        \Reg_Bank/n3725 ) );
  MUX U541 ( .A(\Reg_Bank/registers[22][22] ), .B(n152), .S(n199), .Z(
        \Reg_Bank/n3724 ) );
  MUX U542 ( .A(\Reg_Bank/registers[22][21] ), .B(n153), .S(n199), .Z(
        \Reg_Bank/n3723 ) );
  MUX U543 ( .A(\Reg_Bank/registers[22][20] ), .B(n154), .S(n199), .Z(
        \Reg_Bank/n3722 ) );
  MUX U544 ( .A(\Reg_Bank/registers[22][19] ), .B(n155), .S(n199), .Z(
        \Reg_Bank/n3721 ) );
  MUX U545 ( .A(\Reg_Bank/registers[22][18] ), .B(n156), .S(n199), .Z(
        \Reg_Bank/n3720 ) );
  MUX U546 ( .A(\Reg_Bank/registers[22][17] ), .B(n157), .S(n199), .Z(
        \Reg_Bank/n3719 ) );
  MUX U547 ( .A(\Reg_Bank/registers[22][16] ), .B(n158), .S(n199), .Z(
        \Reg_Bank/n3718 ) );
  MUX U548 ( .A(\Reg_Bank/registers[22][15] ), .B(n159), .S(n199), .Z(
        \Reg_Bank/n3717 ) );
  MUX U549 ( .A(\Reg_Bank/registers[22][14] ), .B(n160), .S(n199), .Z(
        \Reg_Bank/n3716 ) );
  MUX U550 ( .A(\Reg_Bank/registers[22][13] ), .B(n161), .S(n199), .Z(
        \Reg_Bank/n3715 ) );
  MUX U551 ( .A(\Reg_Bank/registers[22][12] ), .B(n162), .S(n199), .Z(
        \Reg_Bank/n3714 ) );
  MUX U552 ( .A(\Reg_Bank/registers[22][11] ), .B(n163), .S(n199), .Z(
        \Reg_Bank/n3713 ) );
  MUX U553 ( .A(\Reg_Bank/registers[22][10] ), .B(n164), .S(n199), .Z(
        \Reg_Bank/n3712 ) );
  MUX U554 ( .A(\Reg_Bank/registers[22][9] ), .B(n165), .S(n199), .Z(
        \Reg_Bank/n3711 ) );
  MUX U555 ( .A(\Reg_Bank/registers[22][8] ), .B(n166), .S(n199), .Z(
        \Reg_Bank/n3710 ) );
  MUX U556 ( .A(\Reg_Bank/registers[22][7] ), .B(n167), .S(n199), .Z(
        \Reg_Bank/n3709 ) );
  MUX U557 ( .A(\Reg_Bank/registers[22][6] ), .B(n168), .S(n199), .Z(
        \Reg_Bank/n3708 ) );
  MUX U558 ( .A(\Reg_Bank/registers[22][5] ), .B(n169), .S(n199), .Z(
        \Reg_Bank/n3707 ) );
  MUX U559 ( .A(\Reg_Bank/registers[22][4] ), .B(n170), .S(n199), .Z(
        \Reg_Bank/n3706 ) );
  MUX U560 ( .A(\Reg_Bank/registers[22][3] ), .B(n171), .S(n199), .Z(
        \Reg_Bank/n3705 ) );
  MUX U561 ( .A(\Reg_Bank/registers[22][2] ), .B(n172), .S(n199), .Z(
        \Reg_Bank/n3704 ) );
  MUX U562 ( .A(\Reg_Bank/registers[22][1] ), .B(n174), .S(n199), .Z(
        \Reg_Bank/n3703 ) );
  MUX U563 ( .A(\Reg_Bank/registers[22][0] ), .B(n175), .S(n199), .Z(
        \Reg_Bank/n3702 ) );
  AND U564 ( .A(n180), .B(n198), .Z(n199) );
  MUX U565 ( .A(\Reg_Bank/registers[21][31] ), .B(n142), .S(n200), .Z(
        \Reg_Bank/n3701 ) );
  MUX U566 ( .A(\Reg_Bank/registers[21][30] ), .B(n144), .S(n200), .Z(
        \Reg_Bank/n3700 ) );
  MUX U567 ( .A(\Reg_Bank/registers[21][29] ), .B(n145), .S(n200), .Z(
        \Reg_Bank/n3699 ) );
  MUX U568 ( .A(\Reg_Bank/registers[21][28] ), .B(n146), .S(n200), .Z(
        \Reg_Bank/n3698 ) );
  MUX U569 ( .A(\Reg_Bank/registers[21][27] ), .B(n147), .S(n200), .Z(
        \Reg_Bank/n3697 ) );
  MUX U570 ( .A(\Reg_Bank/registers[21][26] ), .B(n148), .S(n200), .Z(
        \Reg_Bank/n3696 ) );
  MUX U571 ( .A(\Reg_Bank/registers[21][25] ), .B(n149), .S(n200), .Z(
        \Reg_Bank/n3695 ) );
  MUX U572 ( .A(\Reg_Bank/registers[21][24] ), .B(n150), .S(n200), .Z(
        \Reg_Bank/n3694 ) );
  MUX U573 ( .A(\Reg_Bank/registers[21][23] ), .B(n151), .S(n200), .Z(
        \Reg_Bank/n3693 ) );
  MUX U574 ( .A(\Reg_Bank/registers[21][22] ), .B(n152), .S(n200), .Z(
        \Reg_Bank/n3692 ) );
  MUX U575 ( .A(\Reg_Bank/registers[21][21] ), .B(n153), .S(n200), .Z(
        \Reg_Bank/n3691 ) );
  MUX U576 ( .A(\Reg_Bank/registers[21][20] ), .B(n154), .S(n200), .Z(
        \Reg_Bank/n3690 ) );
  MUX U577 ( .A(\Reg_Bank/registers[21][19] ), .B(n155), .S(n200), .Z(
        \Reg_Bank/n3689 ) );
  MUX U578 ( .A(\Reg_Bank/registers[21][18] ), .B(n156), .S(n200), .Z(
        \Reg_Bank/n3688 ) );
  MUX U579 ( .A(\Reg_Bank/registers[21][17] ), .B(n157), .S(n200), .Z(
        \Reg_Bank/n3687 ) );
  MUX U580 ( .A(\Reg_Bank/registers[21][16] ), .B(n158), .S(n200), .Z(
        \Reg_Bank/n3686 ) );
  MUX U581 ( .A(\Reg_Bank/registers[21][15] ), .B(n159), .S(n200), .Z(
        \Reg_Bank/n3685 ) );
  MUX U582 ( .A(\Reg_Bank/registers[21][14] ), .B(n160), .S(n200), .Z(
        \Reg_Bank/n3684 ) );
  MUX U583 ( .A(\Reg_Bank/registers[21][13] ), .B(n161), .S(n200), .Z(
        \Reg_Bank/n3683 ) );
  MUX U584 ( .A(\Reg_Bank/registers[21][12] ), .B(n162), .S(n200), .Z(
        \Reg_Bank/n3682 ) );
  MUX U585 ( .A(\Reg_Bank/registers[21][11] ), .B(n163), .S(n200), .Z(
        \Reg_Bank/n3681 ) );
  MUX U586 ( .A(\Reg_Bank/registers[21][10] ), .B(n164), .S(n200), .Z(
        \Reg_Bank/n3680 ) );
  MUX U587 ( .A(\Reg_Bank/registers[21][9] ), .B(n165), .S(n200), .Z(
        \Reg_Bank/n3679 ) );
  MUX U588 ( .A(\Reg_Bank/registers[21][8] ), .B(n166), .S(n200), .Z(
        \Reg_Bank/n3678 ) );
  MUX U589 ( .A(\Reg_Bank/registers[21][7] ), .B(n167), .S(n200), .Z(
        \Reg_Bank/n3677 ) );
  MUX U590 ( .A(\Reg_Bank/registers[21][6] ), .B(n168), .S(n200), .Z(
        \Reg_Bank/n3676 ) );
  MUX U591 ( .A(\Reg_Bank/registers[21][5] ), .B(n169), .S(n200), .Z(
        \Reg_Bank/n3675 ) );
  MUX U592 ( .A(\Reg_Bank/registers[21][4] ), .B(n170), .S(n200), .Z(
        \Reg_Bank/n3674 ) );
  MUX U593 ( .A(\Reg_Bank/registers[21][3] ), .B(n171), .S(n200), .Z(
        \Reg_Bank/n3673 ) );
  MUX U594 ( .A(\Reg_Bank/registers[21][2] ), .B(n172), .S(n200), .Z(
        \Reg_Bank/n3672 ) );
  MUX U595 ( .A(\Reg_Bank/registers[21][1] ), .B(n174), .S(n200), .Z(
        \Reg_Bank/n3671 ) );
  MUX U596 ( .A(\Reg_Bank/registers[21][0] ), .B(n175), .S(n200), .Z(
        \Reg_Bank/n3670 ) );
  AND U597 ( .A(n183), .B(n198), .Z(n200) );
  MUX U598 ( .A(\Reg_Bank/registers[20][31] ), .B(n142), .S(n201), .Z(
        \Reg_Bank/n3669 ) );
  MUX U599 ( .A(\Reg_Bank/registers[20][30] ), .B(n144), .S(n201), .Z(
        \Reg_Bank/n3668 ) );
  MUX U600 ( .A(\Reg_Bank/registers[20][29] ), .B(n145), .S(n201), .Z(
        \Reg_Bank/n3667 ) );
  MUX U601 ( .A(\Reg_Bank/registers[20][28] ), .B(n146), .S(n201), .Z(
        \Reg_Bank/n3666 ) );
  MUX U602 ( .A(\Reg_Bank/registers[20][27] ), .B(n147), .S(n201), .Z(
        \Reg_Bank/n3665 ) );
  MUX U603 ( .A(\Reg_Bank/registers[20][26] ), .B(n148), .S(n201), .Z(
        \Reg_Bank/n3664 ) );
  MUX U604 ( .A(\Reg_Bank/registers[20][25] ), .B(n149), .S(n201), .Z(
        \Reg_Bank/n3663 ) );
  MUX U605 ( .A(\Reg_Bank/registers[20][24] ), .B(n150), .S(n201), .Z(
        \Reg_Bank/n3662 ) );
  MUX U606 ( .A(\Reg_Bank/registers[20][23] ), .B(n151), .S(n201), .Z(
        \Reg_Bank/n3661 ) );
  MUX U607 ( .A(\Reg_Bank/registers[20][22] ), .B(n152), .S(n201), .Z(
        \Reg_Bank/n3660 ) );
  MUX U608 ( .A(\Reg_Bank/registers[20][21] ), .B(n153), .S(n201), .Z(
        \Reg_Bank/n3659 ) );
  MUX U609 ( .A(\Reg_Bank/registers[20][20] ), .B(n154), .S(n201), .Z(
        \Reg_Bank/n3658 ) );
  MUX U610 ( .A(\Reg_Bank/registers[20][19] ), .B(n155), .S(n201), .Z(
        \Reg_Bank/n3657 ) );
  MUX U611 ( .A(\Reg_Bank/registers[20][18] ), .B(n156), .S(n201), .Z(
        \Reg_Bank/n3656 ) );
  MUX U612 ( .A(\Reg_Bank/registers[20][17] ), .B(n157), .S(n201), .Z(
        \Reg_Bank/n3655 ) );
  MUX U613 ( .A(\Reg_Bank/registers[20][16] ), .B(n158), .S(n201), .Z(
        \Reg_Bank/n3654 ) );
  MUX U614 ( .A(\Reg_Bank/registers[20][15] ), .B(n159), .S(n201), .Z(
        \Reg_Bank/n3653 ) );
  MUX U615 ( .A(\Reg_Bank/registers[20][14] ), .B(n160), .S(n201), .Z(
        \Reg_Bank/n3652 ) );
  MUX U616 ( .A(\Reg_Bank/registers[20][13] ), .B(n161), .S(n201), .Z(
        \Reg_Bank/n3651 ) );
  MUX U617 ( .A(\Reg_Bank/registers[20][12] ), .B(n162), .S(n201), .Z(
        \Reg_Bank/n3650 ) );
  MUX U618 ( .A(\Reg_Bank/registers[20][11] ), .B(n163), .S(n201), .Z(
        \Reg_Bank/n3649 ) );
  MUX U619 ( .A(\Reg_Bank/registers[20][10] ), .B(n164), .S(n201), .Z(
        \Reg_Bank/n3648 ) );
  MUX U620 ( .A(\Reg_Bank/registers[20][9] ), .B(n165), .S(n201), .Z(
        \Reg_Bank/n3647 ) );
  MUX U621 ( .A(\Reg_Bank/registers[20][8] ), .B(n166), .S(n201), .Z(
        \Reg_Bank/n3646 ) );
  MUX U622 ( .A(\Reg_Bank/registers[20][7] ), .B(n167), .S(n201), .Z(
        \Reg_Bank/n3645 ) );
  MUX U623 ( .A(\Reg_Bank/registers[20][6] ), .B(n168), .S(n201), .Z(
        \Reg_Bank/n3644 ) );
  MUX U624 ( .A(\Reg_Bank/registers[20][5] ), .B(n169), .S(n201), .Z(
        \Reg_Bank/n3643 ) );
  MUX U625 ( .A(\Reg_Bank/registers[20][4] ), .B(n170), .S(n201), .Z(
        \Reg_Bank/n3642 ) );
  MUX U626 ( .A(\Reg_Bank/registers[20][3] ), .B(n171), .S(n201), .Z(
        \Reg_Bank/n3641 ) );
  MUX U627 ( .A(\Reg_Bank/registers[20][2] ), .B(n172), .S(n201), .Z(
        \Reg_Bank/n3640 ) );
  MUX U628 ( .A(\Reg_Bank/registers[20][1] ), .B(n174), .S(n201), .Z(
        \Reg_Bank/n3639 ) );
  MUX U629 ( .A(\Reg_Bank/registers[20][0] ), .B(n175), .S(n201), .Z(
        \Reg_Bank/n3638 ) );
  AND U630 ( .A(n186), .B(n198), .Z(n201) );
  MUX U631 ( .A(\Reg_Bank/registers[19][31] ), .B(n142), .S(n202), .Z(
        \Reg_Bank/n3637 ) );
  MUX U632 ( .A(\Reg_Bank/registers[19][30] ), .B(n144), .S(n202), .Z(
        \Reg_Bank/n3636 ) );
  MUX U633 ( .A(\Reg_Bank/registers[19][29] ), .B(n145), .S(n202), .Z(
        \Reg_Bank/n3635 ) );
  MUX U634 ( .A(\Reg_Bank/registers[19][28] ), .B(n146), .S(n202), .Z(
        \Reg_Bank/n3634 ) );
  MUX U635 ( .A(\Reg_Bank/registers[19][27] ), .B(n147), .S(n202), .Z(
        \Reg_Bank/n3633 ) );
  MUX U636 ( .A(\Reg_Bank/registers[19][26] ), .B(n148), .S(n202), .Z(
        \Reg_Bank/n3632 ) );
  MUX U637 ( .A(\Reg_Bank/registers[19][25] ), .B(n149), .S(n202), .Z(
        \Reg_Bank/n3631 ) );
  MUX U638 ( .A(\Reg_Bank/registers[19][24] ), .B(n150), .S(n202), .Z(
        \Reg_Bank/n3630 ) );
  MUX U639 ( .A(\Reg_Bank/registers[19][23] ), .B(n151), .S(n202), .Z(
        \Reg_Bank/n3629 ) );
  MUX U640 ( .A(\Reg_Bank/registers[19][22] ), .B(n152), .S(n202), .Z(
        \Reg_Bank/n3628 ) );
  MUX U641 ( .A(\Reg_Bank/registers[19][21] ), .B(n153), .S(n202), .Z(
        \Reg_Bank/n3627 ) );
  MUX U642 ( .A(\Reg_Bank/registers[19][20] ), .B(n154), .S(n202), .Z(
        \Reg_Bank/n3626 ) );
  MUX U643 ( .A(\Reg_Bank/registers[19][19] ), .B(n155), .S(n202), .Z(
        \Reg_Bank/n3625 ) );
  MUX U644 ( .A(\Reg_Bank/registers[19][18] ), .B(n156), .S(n202), .Z(
        \Reg_Bank/n3624 ) );
  MUX U645 ( .A(\Reg_Bank/registers[19][17] ), .B(n157), .S(n202), .Z(
        \Reg_Bank/n3623 ) );
  MUX U646 ( .A(\Reg_Bank/registers[19][16] ), .B(n158), .S(n202), .Z(
        \Reg_Bank/n3622 ) );
  MUX U647 ( .A(\Reg_Bank/registers[19][15] ), .B(n159), .S(n202), .Z(
        \Reg_Bank/n3621 ) );
  MUX U648 ( .A(\Reg_Bank/registers[19][14] ), .B(n160), .S(n202), .Z(
        \Reg_Bank/n3620 ) );
  MUX U649 ( .A(\Reg_Bank/registers[19][13] ), .B(n161), .S(n202), .Z(
        \Reg_Bank/n3619 ) );
  MUX U650 ( .A(\Reg_Bank/registers[19][12] ), .B(n162), .S(n202), .Z(
        \Reg_Bank/n3618 ) );
  MUX U651 ( .A(\Reg_Bank/registers[19][11] ), .B(n163), .S(n202), .Z(
        \Reg_Bank/n3617 ) );
  MUX U652 ( .A(\Reg_Bank/registers[19][10] ), .B(n164), .S(n202), .Z(
        \Reg_Bank/n3616 ) );
  MUX U653 ( .A(\Reg_Bank/registers[19][9] ), .B(n165), .S(n202), .Z(
        \Reg_Bank/n3615 ) );
  MUX U654 ( .A(\Reg_Bank/registers[19][8] ), .B(n166), .S(n202), .Z(
        \Reg_Bank/n3614 ) );
  MUX U655 ( .A(\Reg_Bank/registers[19][7] ), .B(n167), .S(n202), .Z(
        \Reg_Bank/n3613 ) );
  MUX U656 ( .A(\Reg_Bank/registers[19][6] ), .B(n168), .S(n202), .Z(
        \Reg_Bank/n3612 ) );
  MUX U657 ( .A(\Reg_Bank/registers[19][5] ), .B(n169), .S(n202), .Z(
        \Reg_Bank/n3611 ) );
  MUX U658 ( .A(\Reg_Bank/registers[19][4] ), .B(n170), .S(n202), .Z(
        \Reg_Bank/n3610 ) );
  MUX U659 ( .A(\Reg_Bank/registers[19][3] ), .B(n171), .S(n202), .Z(
        \Reg_Bank/n3609 ) );
  MUX U660 ( .A(\Reg_Bank/registers[19][2] ), .B(n172), .S(n202), .Z(
        \Reg_Bank/n3608 ) );
  MUX U661 ( .A(\Reg_Bank/registers[19][1] ), .B(n174), .S(n202), .Z(
        \Reg_Bank/n3607 ) );
  MUX U662 ( .A(\Reg_Bank/registers[19][0] ), .B(n175), .S(n202), .Z(
        \Reg_Bank/n3606 ) );
  AND U663 ( .A(n198), .B(n188), .Z(n202) );
  MUX U664 ( .A(\Reg_Bank/registers[18][31] ), .B(n142), .S(n203), .Z(
        \Reg_Bank/n3605 ) );
  MUX U665 ( .A(\Reg_Bank/registers[18][30] ), .B(n144), .S(n203), .Z(
        \Reg_Bank/n3604 ) );
  MUX U666 ( .A(\Reg_Bank/registers[18][29] ), .B(n145), .S(n203), .Z(
        \Reg_Bank/n3603 ) );
  MUX U667 ( .A(\Reg_Bank/registers[18][28] ), .B(n146), .S(n203), .Z(
        \Reg_Bank/n3602 ) );
  MUX U668 ( .A(\Reg_Bank/registers[18][27] ), .B(n147), .S(n203), .Z(
        \Reg_Bank/n3601 ) );
  MUX U669 ( .A(\Reg_Bank/registers[18][26] ), .B(n148), .S(n203), .Z(
        \Reg_Bank/n3600 ) );
  MUX U670 ( .A(\Reg_Bank/registers[18][25] ), .B(n149), .S(n203), .Z(
        \Reg_Bank/n3599 ) );
  MUX U671 ( .A(\Reg_Bank/registers[18][24] ), .B(n150), .S(n203), .Z(
        \Reg_Bank/n3598 ) );
  MUX U672 ( .A(\Reg_Bank/registers[18][23] ), .B(n151), .S(n203), .Z(
        \Reg_Bank/n3597 ) );
  MUX U673 ( .A(\Reg_Bank/registers[18][22] ), .B(n152), .S(n203), .Z(
        \Reg_Bank/n3596 ) );
  MUX U674 ( .A(\Reg_Bank/registers[18][21] ), .B(n153), .S(n203), .Z(
        \Reg_Bank/n3595 ) );
  MUX U675 ( .A(\Reg_Bank/registers[18][20] ), .B(n154), .S(n203), .Z(
        \Reg_Bank/n3594 ) );
  MUX U676 ( .A(\Reg_Bank/registers[18][19] ), .B(n155), .S(n203), .Z(
        \Reg_Bank/n3593 ) );
  MUX U677 ( .A(\Reg_Bank/registers[18][18] ), .B(n156), .S(n203), .Z(
        \Reg_Bank/n3592 ) );
  MUX U678 ( .A(\Reg_Bank/registers[18][17] ), .B(n157), .S(n203), .Z(
        \Reg_Bank/n3591 ) );
  MUX U679 ( .A(\Reg_Bank/registers[18][16] ), .B(n158), .S(n203), .Z(
        \Reg_Bank/n3590 ) );
  MUX U680 ( .A(\Reg_Bank/registers[18][15] ), .B(n159), .S(n203), .Z(
        \Reg_Bank/n3589 ) );
  MUX U681 ( .A(\Reg_Bank/registers[18][14] ), .B(n160), .S(n203), .Z(
        \Reg_Bank/n3588 ) );
  MUX U682 ( .A(\Reg_Bank/registers[18][13] ), .B(n161), .S(n203), .Z(
        \Reg_Bank/n3587 ) );
  MUX U683 ( .A(\Reg_Bank/registers[18][12] ), .B(n162), .S(n203), .Z(
        \Reg_Bank/n3586 ) );
  MUX U684 ( .A(\Reg_Bank/registers[18][11] ), .B(n163), .S(n203), .Z(
        \Reg_Bank/n3585 ) );
  MUX U685 ( .A(\Reg_Bank/registers[18][10] ), .B(n164), .S(n203), .Z(
        \Reg_Bank/n3584 ) );
  MUX U686 ( .A(\Reg_Bank/registers[18][9] ), .B(n165), .S(n203), .Z(
        \Reg_Bank/n3583 ) );
  MUX U687 ( .A(\Reg_Bank/registers[18][8] ), .B(n166), .S(n203), .Z(
        \Reg_Bank/n3582 ) );
  MUX U688 ( .A(\Reg_Bank/registers[18][7] ), .B(n167), .S(n203), .Z(
        \Reg_Bank/n3581 ) );
  MUX U689 ( .A(\Reg_Bank/registers[18][6] ), .B(n168), .S(n203), .Z(
        \Reg_Bank/n3580 ) );
  MUX U690 ( .A(\Reg_Bank/registers[18][5] ), .B(n169), .S(n203), .Z(
        \Reg_Bank/n3579 ) );
  MUX U691 ( .A(\Reg_Bank/registers[18][4] ), .B(n170), .S(n203), .Z(
        \Reg_Bank/n3578 ) );
  MUX U692 ( .A(\Reg_Bank/registers[18][3] ), .B(n171), .S(n203), .Z(
        \Reg_Bank/n3577 ) );
  MUX U693 ( .A(\Reg_Bank/registers[18][2] ), .B(n172), .S(n203), .Z(
        \Reg_Bank/n3576 ) );
  MUX U694 ( .A(\Reg_Bank/registers[18][1] ), .B(n174), .S(n203), .Z(
        \Reg_Bank/n3575 ) );
  MUX U695 ( .A(\Reg_Bank/registers[18][0] ), .B(n175), .S(n203), .Z(
        \Reg_Bank/n3574 ) );
  AND U696 ( .A(n198), .B(n190), .Z(n203) );
  MUX U697 ( .A(\Reg_Bank/registers[17][31] ), .B(n142), .S(n204), .Z(
        \Reg_Bank/n3573 ) );
  MUX U698 ( .A(\Reg_Bank/registers[17][30] ), .B(n144), .S(n204), .Z(
        \Reg_Bank/n3572 ) );
  MUX U699 ( .A(\Reg_Bank/registers[17][29] ), .B(n145), .S(n204), .Z(
        \Reg_Bank/n3571 ) );
  MUX U700 ( .A(\Reg_Bank/registers[17][28] ), .B(n146), .S(n204), .Z(
        \Reg_Bank/n3570 ) );
  MUX U701 ( .A(\Reg_Bank/registers[17][27] ), .B(n147), .S(n204), .Z(
        \Reg_Bank/n3569 ) );
  MUX U702 ( .A(\Reg_Bank/registers[17][26] ), .B(n148), .S(n204), .Z(
        \Reg_Bank/n3568 ) );
  MUX U703 ( .A(\Reg_Bank/registers[17][25] ), .B(n149), .S(n204), .Z(
        \Reg_Bank/n3567 ) );
  MUX U704 ( .A(\Reg_Bank/registers[17][24] ), .B(n150), .S(n204), .Z(
        \Reg_Bank/n3566 ) );
  MUX U705 ( .A(\Reg_Bank/registers[17][23] ), .B(n151), .S(n204), .Z(
        \Reg_Bank/n3565 ) );
  MUX U706 ( .A(\Reg_Bank/registers[17][22] ), .B(n152), .S(n204), .Z(
        \Reg_Bank/n3564 ) );
  MUX U707 ( .A(\Reg_Bank/registers[17][21] ), .B(n153), .S(n204), .Z(
        \Reg_Bank/n3563 ) );
  MUX U708 ( .A(\Reg_Bank/registers[17][20] ), .B(n154), .S(n204), .Z(
        \Reg_Bank/n3562 ) );
  MUX U709 ( .A(\Reg_Bank/registers[17][19] ), .B(n155), .S(n204), .Z(
        \Reg_Bank/n3561 ) );
  MUX U710 ( .A(\Reg_Bank/registers[17][18] ), .B(n156), .S(n204), .Z(
        \Reg_Bank/n3560 ) );
  MUX U711 ( .A(\Reg_Bank/registers[17][17] ), .B(n157), .S(n204), .Z(
        \Reg_Bank/n3559 ) );
  MUX U712 ( .A(\Reg_Bank/registers[17][16] ), .B(n158), .S(n204), .Z(
        \Reg_Bank/n3558 ) );
  MUX U713 ( .A(\Reg_Bank/registers[17][15] ), .B(n159), .S(n204), .Z(
        \Reg_Bank/n3557 ) );
  MUX U714 ( .A(\Reg_Bank/registers[17][14] ), .B(n160), .S(n204), .Z(
        \Reg_Bank/n3556 ) );
  MUX U715 ( .A(\Reg_Bank/registers[17][13] ), .B(n161), .S(n204), .Z(
        \Reg_Bank/n3555 ) );
  MUX U716 ( .A(\Reg_Bank/registers[17][12] ), .B(n162), .S(n204), .Z(
        \Reg_Bank/n3554 ) );
  MUX U717 ( .A(\Reg_Bank/registers[17][11] ), .B(n163), .S(n204), .Z(
        \Reg_Bank/n3553 ) );
  MUX U718 ( .A(\Reg_Bank/registers[17][10] ), .B(n164), .S(n204), .Z(
        \Reg_Bank/n3552 ) );
  MUX U719 ( .A(\Reg_Bank/registers[17][9] ), .B(n165), .S(n204), .Z(
        \Reg_Bank/n3551 ) );
  MUX U720 ( .A(\Reg_Bank/registers[17][8] ), .B(n166), .S(n204), .Z(
        \Reg_Bank/n3550 ) );
  MUX U721 ( .A(\Reg_Bank/registers[17][7] ), .B(n167), .S(n204), .Z(
        \Reg_Bank/n3549 ) );
  MUX U722 ( .A(\Reg_Bank/registers[17][6] ), .B(n168), .S(n204), .Z(
        \Reg_Bank/n3548 ) );
  MUX U723 ( .A(\Reg_Bank/registers[17][5] ), .B(n169), .S(n204), .Z(
        \Reg_Bank/n3547 ) );
  MUX U724 ( .A(\Reg_Bank/registers[17][4] ), .B(n170), .S(n204), .Z(
        \Reg_Bank/n3546 ) );
  MUX U725 ( .A(\Reg_Bank/registers[17][3] ), .B(n171), .S(n204), .Z(
        \Reg_Bank/n3545 ) );
  MUX U726 ( .A(\Reg_Bank/registers[17][2] ), .B(n172), .S(n204), .Z(
        \Reg_Bank/n3544 ) );
  MUX U727 ( .A(\Reg_Bank/registers[17][1] ), .B(n174), .S(n204), .Z(
        \Reg_Bank/n3543 ) );
  MUX U728 ( .A(\Reg_Bank/registers[17][0] ), .B(n175), .S(n204), .Z(
        \Reg_Bank/n3542 ) );
  AND U729 ( .A(n198), .B(n192), .Z(n204) );
  MUX U730 ( .A(\Reg_Bank/registers[16][31] ), .B(n142), .S(n205), .Z(
        \Reg_Bank/n3541 ) );
  MUX U731 ( .A(\Reg_Bank/registers[16][30] ), .B(n144), .S(n205), .Z(
        \Reg_Bank/n3540 ) );
  MUX U732 ( .A(\Reg_Bank/registers[16][29] ), .B(n145), .S(n205), .Z(
        \Reg_Bank/n3539 ) );
  MUX U733 ( .A(\Reg_Bank/registers[16][28] ), .B(n146), .S(n205), .Z(
        \Reg_Bank/n3538 ) );
  MUX U734 ( .A(\Reg_Bank/registers[16][27] ), .B(n147), .S(n205), .Z(
        \Reg_Bank/n3537 ) );
  MUX U735 ( .A(\Reg_Bank/registers[16][26] ), .B(n148), .S(n205), .Z(
        \Reg_Bank/n3536 ) );
  MUX U736 ( .A(\Reg_Bank/registers[16][25] ), .B(n149), .S(n205), .Z(
        \Reg_Bank/n3535 ) );
  MUX U737 ( .A(\Reg_Bank/registers[16][24] ), .B(n150), .S(n205), .Z(
        \Reg_Bank/n3534 ) );
  MUX U738 ( .A(\Reg_Bank/registers[16][23] ), .B(n151), .S(n205), .Z(
        \Reg_Bank/n3533 ) );
  MUX U739 ( .A(\Reg_Bank/registers[16][22] ), .B(n152), .S(n205), .Z(
        \Reg_Bank/n3532 ) );
  MUX U740 ( .A(\Reg_Bank/registers[16][21] ), .B(n153), .S(n205), .Z(
        \Reg_Bank/n3531 ) );
  MUX U741 ( .A(\Reg_Bank/registers[16][20] ), .B(n154), .S(n205), .Z(
        \Reg_Bank/n3530 ) );
  MUX U742 ( .A(\Reg_Bank/registers[16][19] ), .B(n155), .S(n205), .Z(
        \Reg_Bank/n3529 ) );
  MUX U743 ( .A(\Reg_Bank/registers[16][18] ), .B(n156), .S(n205), .Z(
        \Reg_Bank/n3528 ) );
  MUX U744 ( .A(\Reg_Bank/registers[16][17] ), .B(n157), .S(n205), .Z(
        \Reg_Bank/n3527 ) );
  MUX U745 ( .A(\Reg_Bank/registers[16][16] ), .B(n158), .S(n205), .Z(
        \Reg_Bank/n3526 ) );
  MUX U746 ( .A(\Reg_Bank/registers[16][15] ), .B(n159), .S(n205), .Z(
        \Reg_Bank/n3525 ) );
  MUX U747 ( .A(\Reg_Bank/registers[16][14] ), .B(n160), .S(n205), .Z(
        \Reg_Bank/n3524 ) );
  MUX U748 ( .A(\Reg_Bank/registers[16][13] ), .B(n161), .S(n205), .Z(
        \Reg_Bank/n3523 ) );
  MUX U749 ( .A(\Reg_Bank/registers[16][12] ), .B(n162), .S(n205), .Z(
        \Reg_Bank/n3522 ) );
  MUX U750 ( .A(\Reg_Bank/registers[16][11] ), .B(n163), .S(n205), .Z(
        \Reg_Bank/n3521 ) );
  MUX U751 ( .A(\Reg_Bank/registers[16][10] ), .B(n164), .S(n205), .Z(
        \Reg_Bank/n3520 ) );
  MUX U752 ( .A(\Reg_Bank/registers[16][9] ), .B(n165), .S(n205), .Z(
        \Reg_Bank/n3519 ) );
  MUX U753 ( .A(\Reg_Bank/registers[16][8] ), .B(n166), .S(n205), .Z(
        \Reg_Bank/n3518 ) );
  MUX U754 ( .A(\Reg_Bank/registers[16][7] ), .B(n167), .S(n205), .Z(
        \Reg_Bank/n3517 ) );
  MUX U755 ( .A(\Reg_Bank/registers[16][6] ), .B(n168), .S(n205), .Z(
        \Reg_Bank/n3516 ) );
  MUX U756 ( .A(\Reg_Bank/registers[16][5] ), .B(n169), .S(n205), .Z(
        \Reg_Bank/n3515 ) );
  MUX U757 ( .A(\Reg_Bank/registers[16][4] ), .B(n170), .S(n205), .Z(
        \Reg_Bank/n3514 ) );
  MUX U758 ( .A(\Reg_Bank/registers[16][3] ), .B(n171), .S(n205), .Z(
        \Reg_Bank/n3513 ) );
  MUX U759 ( .A(\Reg_Bank/registers[16][2] ), .B(n172), .S(n205), .Z(
        \Reg_Bank/n3512 ) );
  MUX U760 ( .A(\Reg_Bank/registers[16][1] ), .B(n174), .S(n205), .Z(
        \Reg_Bank/n3511 ) );
  MUX U761 ( .A(\Reg_Bank/registers[16][0] ), .B(n175), .S(n205), .Z(
        \Reg_Bank/n3510 ) );
  AND U762 ( .A(n198), .B(n194), .Z(n205) );
  IV U763 ( .A(n206), .Z(n194) );
  AND U764 ( .A(n195), .B(n196), .Z(n198) );
  IV U765 ( .A(n207), .Z(n196) );
  MUX U766 ( .A(n142), .B(\Reg_Bank/registers[15][31] ), .S(n208), .Z(
        \Reg_Bank/n3509 ) );
  MUX U767 ( .A(n144), .B(\Reg_Bank/registers[15][30] ), .S(n208), .Z(
        \Reg_Bank/n3508 ) );
  MUX U768 ( .A(n145), .B(\Reg_Bank/registers[15][29] ), .S(n208), .Z(
        \Reg_Bank/n3507 ) );
  MUX U769 ( .A(n146), .B(\Reg_Bank/registers[15][28] ), .S(n208), .Z(
        \Reg_Bank/n3506 ) );
  MUX U770 ( .A(n147), .B(\Reg_Bank/registers[15][27] ), .S(n208), .Z(
        \Reg_Bank/n3505 ) );
  MUX U771 ( .A(n148), .B(\Reg_Bank/registers[15][26] ), .S(n208), .Z(
        \Reg_Bank/n3504 ) );
  MUX U772 ( .A(n149), .B(\Reg_Bank/registers[15][25] ), .S(n208), .Z(
        \Reg_Bank/n3503 ) );
  MUX U773 ( .A(n150), .B(\Reg_Bank/registers[15][24] ), .S(n208), .Z(
        \Reg_Bank/n3502 ) );
  MUX U774 ( .A(n151), .B(\Reg_Bank/registers[15][23] ), .S(n208), .Z(
        \Reg_Bank/n3501 ) );
  MUX U775 ( .A(n152), .B(\Reg_Bank/registers[15][22] ), .S(n208), .Z(
        \Reg_Bank/n3500 ) );
  MUX U776 ( .A(n153), .B(\Reg_Bank/registers[15][21] ), .S(n208), .Z(
        \Reg_Bank/n3499 ) );
  MUX U777 ( .A(n154), .B(\Reg_Bank/registers[15][20] ), .S(n208), .Z(
        \Reg_Bank/n3498 ) );
  MUX U778 ( .A(n155), .B(\Reg_Bank/registers[15][19] ), .S(n208), .Z(
        \Reg_Bank/n3497 ) );
  MUX U779 ( .A(n156), .B(\Reg_Bank/registers[15][18] ), .S(n208), .Z(
        \Reg_Bank/n3496 ) );
  MUX U780 ( .A(n157), .B(\Reg_Bank/registers[15][17] ), .S(n208), .Z(
        \Reg_Bank/n3495 ) );
  MUX U781 ( .A(n158), .B(\Reg_Bank/registers[15][16] ), .S(n208), .Z(
        \Reg_Bank/n3494 ) );
  MUX U782 ( .A(n159), .B(\Reg_Bank/registers[15][15] ), .S(n208), .Z(
        \Reg_Bank/n3493 ) );
  MUX U783 ( .A(n160), .B(\Reg_Bank/registers[15][14] ), .S(n208), .Z(
        \Reg_Bank/n3492 ) );
  MUX U784 ( .A(n161), .B(\Reg_Bank/registers[15][13] ), .S(n208), .Z(
        \Reg_Bank/n3491 ) );
  MUX U785 ( .A(n162), .B(\Reg_Bank/registers[15][12] ), .S(n208), .Z(
        \Reg_Bank/n3490 ) );
  MUX U786 ( .A(n163), .B(\Reg_Bank/registers[15][11] ), .S(n208), .Z(
        \Reg_Bank/n3489 ) );
  MUX U787 ( .A(n164), .B(\Reg_Bank/registers[15][10] ), .S(n208), .Z(
        \Reg_Bank/n3488 ) );
  MUX U788 ( .A(n165), .B(\Reg_Bank/registers[15][9] ), .S(n208), .Z(
        \Reg_Bank/n3487 ) );
  MUX U789 ( .A(n166), .B(\Reg_Bank/registers[15][8] ), .S(n208), .Z(
        \Reg_Bank/n3486 ) );
  MUX U790 ( .A(n167), .B(\Reg_Bank/registers[15][7] ), .S(n208), .Z(
        \Reg_Bank/n3485 ) );
  MUX U791 ( .A(n168), .B(\Reg_Bank/registers[15][6] ), .S(n208), .Z(
        \Reg_Bank/n3484 ) );
  MUX U792 ( .A(n169), .B(\Reg_Bank/registers[15][5] ), .S(n208), .Z(
        \Reg_Bank/n3483 ) );
  MUX U793 ( .A(n170), .B(\Reg_Bank/registers[15][4] ), .S(n208), .Z(
        \Reg_Bank/n3482 ) );
  MUX U794 ( .A(n171), .B(\Reg_Bank/registers[15][3] ), .S(n208), .Z(
        \Reg_Bank/n3481 ) );
  MUX U795 ( .A(n172), .B(\Reg_Bank/registers[15][2] ), .S(n208), .Z(
        \Reg_Bank/n3480 ) );
  IV U796 ( .A(n209), .Z(n208) );
  MUX U797 ( .A(\Reg_Bank/registers[15][1] ), .B(n174), .S(n209), .Z(
        \Reg_Bank/n3479 ) );
  MUX U798 ( .A(\Reg_Bank/registers[15][0] ), .B(n175), .S(n209), .Z(
        \Reg_Bank/n3478 ) );
  NOR U799 ( .A(n177), .B(n210), .Z(n209) );
  MUX U800 ( .A(\Reg_Bank/registers[14][31] ), .B(n142), .S(n211), .Z(
        \Reg_Bank/n3477 ) );
  MUX U801 ( .A(\Reg_Bank/registers[14][30] ), .B(n144), .S(n211), .Z(
        \Reg_Bank/n3476 ) );
  MUX U802 ( .A(\Reg_Bank/registers[14][29] ), .B(n145), .S(n211), .Z(
        \Reg_Bank/n3475 ) );
  MUX U803 ( .A(\Reg_Bank/registers[14][28] ), .B(n146), .S(n211), .Z(
        \Reg_Bank/n3474 ) );
  MUX U804 ( .A(\Reg_Bank/registers[14][27] ), .B(n147), .S(n211), .Z(
        \Reg_Bank/n3473 ) );
  MUX U805 ( .A(\Reg_Bank/registers[14][26] ), .B(n148), .S(n211), .Z(
        \Reg_Bank/n3472 ) );
  MUX U806 ( .A(\Reg_Bank/registers[14][25] ), .B(n149), .S(n211), .Z(
        \Reg_Bank/n3471 ) );
  MUX U807 ( .A(\Reg_Bank/registers[14][24] ), .B(n150), .S(n211), .Z(
        \Reg_Bank/n3470 ) );
  MUX U808 ( .A(\Reg_Bank/registers[14][23] ), .B(n151), .S(n211), .Z(
        \Reg_Bank/n3469 ) );
  MUX U809 ( .A(\Reg_Bank/registers[14][22] ), .B(n152), .S(n211), .Z(
        \Reg_Bank/n3468 ) );
  MUX U810 ( .A(\Reg_Bank/registers[14][21] ), .B(n153), .S(n211), .Z(
        \Reg_Bank/n3467 ) );
  MUX U811 ( .A(\Reg_Bank/registers[14][20] ), .B(n154), .S(n211), .Z(
        \Reg_Bank/n3466 ) );
  MUX U812 ( .A(\Reg_Bank/registers[14][19] ), .B(n155), .S(n211), .Z(
        \Reg_Bank/n3465 ) );
  MUX U813 ( .A(\Reg_Bank/registers[14][18] ), .B(n156), .S(n211), .Z(
        \Reg_Bank/n3464 ) );
  MUX U814 ( .A(\Reg_Bank/registers[14][17] ), .B(n157), .S(n211), .Z(
        \Reg_Bank/n3463 ) );
  MUX U815 ( .A(\Reg_Bank/registers[14][16] ), .B(n158), .S(n211), .Z(
        \Reg_Bank/n3462 ) );
  MUX U816 ( .A(\Reg_Bank/registers[14][15] ), .B(n159), .S(n211), .Z(
        \Reg_Bank/n3461 ) );
  MUX U817 ( .A(\Reg_Bank/registers[14][14] ), .B(n160), .S(n211), .Z(
        \Reg_Bank/n3460 ) );
  MUX U818 ( .A(\Reg_Bank/registers[14][13] ), .B(n161), .S(n211), .Z(
        \Reg_Bank/n3459 ) );
  MUX U819 ( .A(\Reg_Bank/registers[14][12] ), .B(n162), .S(n211), .Z(
        \Reg_Bank/n3458 ) );
  MUX U820 ( .A(\Reg_Bank/registers[14][11] ), .B(n163), .S(n211), .Z(
        \Reg_Bank/n3457 ) );
  MUX U821 ( .A(\Reg_Bank/registers[14][10] ), .B(n164), .S(n211), .Z(
        \Reg_Bank/n3456 ) );
  MUX U822 ( .A(\Reg_Bank/registers[14][9] ), .B(n165), .S(n211), .Z(
        \Reg_Bank/n3455 ) );
  MUX U823 ( .A(\Reg_Bank/registers[14][8] ), .B(n166), .S(n211), .Z(
        \Reg_Bank/n3454 ) );
  MUX U824 ( .A(\Reg_Bank/registers[14][7] ), .B(n167), .S(n211), .Z(
        \Reg_Bank/n3453 ) );
  MUX U825 ( .A(\Reg_Bank/registers[14][6] ), .B(n168), .S(n211), .Z(
        \Reg_Bank/n3452 ) );
  MUX U826 ( .A(\Reg_Bank/registers[14][5] ), .B(n169), .S(n211), .Z(
        \Reg_Bank/n3451 ) );
  MUX U827 ( .A(\Reg_Bank/registers[14][4] ), .B(n170), .S(n211), .Z(
        \Reg_Bank/n3450 ) );
  MUX U828 ( .A(\Reg_Bank/registers[14][3] ), .B(n171), .S(n211), .Z(
        \Reg_Bank/n3449 ) );
  MUX U829 ( .A(\Reg_Bank/registers[14][2] ), .B(n172), .S(n211), .Z(
        \Reg_Bank/n3448 ) );
  MUX U830 ( .A(\Reg_Bank/registers[14][1] ), .B(n174), .S(n211), .Z(
        \Reg_Bank/n3447 ) );
  MUX U831 ( .A(\Reg_Bank/registers[14][0] ), .B(n175), .S(n211), .Z(
        \Reg_Bank/n3446 ) );
  ANDN U832 ( .B(n180), .A(n210), .Z(n211) );
  MUX U833 ( .A(\Reg_Bank/registers[13][31] ), .B(n142), .S(n212), .Z(
        \Reg_Bank/n3445 ) );
  MUX U834 ( .A(\Reg_Bank/registers[13][30] ), .B(n144), .S(n212), .Z(
        \Reg_Bank/n3444 ) );
  MUX U835 ( .A(\Reg_Bank/registers[13][29] ), .B(n145), .S(n212), .Z(
        \Reg_Bank/n3443 ) );
  MUX U836 ( .A(\Reg_Bank/registers[13][28] ), .B(n146), .S(n212), .Z(
        \Reg_Bank/n3442 ) );
  MUX U837 ( .A(\Reg_Bank/registers[13][27] ), .B(n147), .S(n212), .Z(
        \Reg_Bank/n3441 ) );
  MUX U838 ( .A(\Reg_Bank/registers[13][26] ), .B(n148), .S(n212), .Z(
        \Reg_Bank/n3440 ) );
  MUX U839 ( .A(\Reg_Bank/registers[13][25] ), .B(n149), .S(n212), .Z(
        \Reg_Bank/n3439 ) );
  MUX U840 ( .A(\Reg_Bank/registers[13][24] ), .B(n150), .S(n212), .Z(
        \Reg_Bank/n3438 ) );
  MUX U841 ( .A(\Reg_Bank/registers[13][23] ), .B(n151), .S(n212), .Z(
        \Reg_Bank/n3437 ) );
  MUX U842 ( .A(\Reg_Bank/registers[13][22] ), .B(n152), .S(n212), .Z(
        \Reg_Bank/n3436 ) );
  MUX U843 ( .A(\Reg_Bank/registers[13][21] ), .B(n153), .S(n212), .Z(
        \Reg_Bank/n3435 ) );
  MUX U844 ( .A(\Reg_Bank/registers[13][20] ), .B(n154), .S(n212), .Z(
        \Reg_Bank/n3434 ) );
  MUX U845 ( .A(\Reg_Bank/registers[13][19] ), .B(n155), .S(n212), .Z(
        \Reg_Bank/n3433 ) );
  MUX U846 ( .A(\Reg_Bank/registers[13][18] ), .B(n156), .S(n212), .Z(
        \Reg_Bank/n3432 ) );
  MUX U847 ( .A(\Reg_Bank/registers[13][17] ), .B(n157), .S(n212), .Z(
        \Reg_Bank/n3431 ) );
  MUX U848 ( .A(\Reg_Bank/registers[13][16] ), .B(n158), .S(n212), .Z(
        \Reg_Bank/n3430 ) );
  MUX U849 ( .A(\Reg_Bank/registers[13][15] ), .B(n159), .S(n212), .Z(
        \Reg_Bank/n3429 ) );
  MUX U850 ( .A(\Reg_Bank/registers[13][14] ), .B(n160), .S(n212), .Z(
        \Reg_Bank/n3428 ) );
  MUX U851 ( .A(\Reg_Bank/registers[13][13] ), .B(n161), .S(n212), .Z(
        \Reg_Bank/n3427 ) );
  MUX U852 ( .A(\Reg_Bank/registers[13][12] ), .B(n162), .S(n212), .Z(
        \Reg_Bank/n3426 ) );
  MUX U853 ( .A(\Reg_Bank/registers[13][11] ), .B(n163), .S(n212), .Z(
        \Reg_Bank/n3425 ) );
  MUX U854 ( .A(\Reg_Bank/registers[13][10] ), .B(n164), .S(n212), .Z(
        \Reg_Bank/n3424 ) );
  MUX U855 ( .A(\Reg_Bank/registers[13][9] ), .B(n165), .S(n212), .Z(
        \Reg_Bank/n3423 ) );
  MUX U856 ( .A(\Reg_Bank/registers[13][8] ), .B(n166), .S(n212), .Z(
        \Reg_Bank/n3422 ) );
  MUX U857 ( .A(\Reg_Bank/registers[13][7] ), .B(n167), .S(n212), .Z(
        \Reg_Bank/n3421 ) );
  MUX U858 ( .A(\Reg_Bank/registers[13][6] ), .B(n168), .S(n212), .Z(
        \Reg_Bank/n3420 ) );
  MUX U859 ( .A(\Reg_Bank/registers[13][5] ), .B(n169), .S(n212), .Z(
        \Reg_Bank/n3419 ) );
  MUX U860 ( .A(\Reg_Bank/registers[13][4] ), .B(n170), .S(n212), .Z(
        \Reg_Bank/n3418 ) );
  MUX U861 ( .A(\Reg_Bank/registers[13][3] ), .B(n171), .S(n212), .Z(
        \Reg_Bank/n3417 ) );
  MUX U862 ( .A(\Reg_Bank/registers[13][2] ), .B(n172), .S(n212), .Z(
        \Reg_Bank/n3416 ) );
  MUX U863 ( .A(\Reg_Bank/registers[13][1] ), .B(n174), .S(n212), .Z(
        \Reg_Bank/n3415 ) );
  MUX U864 ( .A(\Reg_Bank/registers[13][0] ), .B(n175), .S(n212), .Z(
        \Reg_Bank/n3414 ) );
  ANDN U865 ( .B(n183), .A(n210), .Z(n212) );
  MUX U866 ( .A(\Reg_Bank/registers[12][31] ), .B(n142), .S(n213), .Z(
        \Reg_Bank/n3413 ) );
  MUX U867 ( .A(\Reg_Bank/registers[12][30] ), .B(n144), .S(n213), .Z(
        \Reg_Bank/n3412 ) );
  MUX U868 ( .A(\Reg_Bank/registers[12][29] ), .B(n145), .S(n213), .Z(
        \Reg_Bank/n3411 ) );
  MUX U869 ( .A(\Reg_Bank/registers[12][28] ), .B(n146), .S(n213), .Z(
        \Reg_Bank/n3410 ) );
  MUX U870 ( .A(\Reg_Bank/registers[12][27] ), .B(n147), .S(n213), .Z(
        \Reg_Bank/n3409 ) );
  MUX U871 ( .A(\Reg_Bank/registers[12][26] ), .B(n148), .S(n213), .Z(
        \Reg_Bank/n3408 ) );
  MUX U872 ( .A(\Reg_Bank/registers[12][25] ), .B(n149), .S(n213), .Z(
        \Reg_Bank/n3407 ) );
  MUX U873 ( .A(\Reg_Bank/registers[12][24] ), .B(n150), .S(n213), .Z(
        \Reg_Bank/n3406 ) );
  MUX U874 ( .A(\Reg_Bank/registers[12][23] ), .B(n151), .S(n213), .Z(
        \Reg_Bank/n3405 ) );
  MUX U875 ( .A(\Reg_Bank/registers[12][22] ), .B(n152), .S(n213), .Z(
        \Reg_Bank/n3404 ) );
  MUX U876 ( .A(\Reg_Bank/registers[12][21] ), .B(n153), .S(n213), .Z(
        \Reg_Bank/n3403 ) );
  MUX U877 ( .A(\Reg_Bank/registers[12][20] ), .B(n154), .S(n213), .Z(
        \Reg_Bank/n3402 ) );
  MUX U878 ( .A(\Reg_Bank/registers[12][19] ), .B(n155), .S(n213), .Z(
        \Reg_Bank/n3401 ) );
  MUX U879 ( .A(\Reg_Bank/registers[12][18] ), .B(n156), .S(n213), .Z(
        \Reg_Bank/n3400 ) );
  MUX U880 ( .A(\Reg_Bank/registers[12][17] ), .B(n157), .S(n213), .Z(
        \Reg_Bank/n3399 ) );
  MUX U881 ( .A(\Reg_Bank/registers[12][16] ), .B(n158), .S(n213), .Z(
        \Reg_Bank/n3398 ) );
  MUX U882 ( .A(\Reg_Bank/registers[12][15] ), .B(n159), .S(n213), .Z(
        \Reg_Bank/n3397 ) );
  MUX U883 ( .A(\Reg_Bank/registers[12][14] ), .B(n160), .S(n213), .Z(
        \Reg_Bank/n3396 ) );
  MUX U884 ( .A(\Reg_Bank/registers[12][13] ), .B(n161), .S(n213), .Z(
        \Reg_Bank/n3395 ) );
  MUX U885 ( .A(\Reg_Bank/registers[12][12] ), .B(n162), .S(n213), .Z(
        \Reg_Bank/n3394 ) );
  MUX U886 ( .A(\Reg_Bank/registers[12][11] ), .B(n163), .S(n213), .Z(
        \Reg_Bank/n3393 ) );
  MUX U887 ( .A(\Reg_Bank/registers[12][10] ), .B(n164), .S(n213), .Z(
        \Reg_Bank/n3392 ) );
  MUX U888 ( .A(\Reg_Bank/registers[12][9] ), .B(n165), .S(n213), .Z(
        \Reg_Bank/n3391 ) );
  MUX U889 ( .A(\Reg_Bank/registers[12][8] ), .B(n166), .S(n213), .Z(
        \Reg_Bank/n3390 ) );
  MUX U890 ( .A(\Reg_Bank/registers[12][7] ), .B(n167), .S(n213), .Z(
        \Reg_Bank/n3389 ) );
  MUX U891 ( .A(\Reg_Bank/registers[12][6] ), .B(n168), .S(n213), .Z(
        \Reg_Bank/n3388 ) );
  MUX U892 ( .A(\Reg_Bank/registers[12][5] ), .B(n169), .S(n213), .Z(
        \Reg_Bank/n3387 ) );
  MUX U893 ( .A(\Reg_Bank/registers[12][4] ), .B(n170), .S(n213), .Z(
        \Reg_Bank/n3386 ) );
  MUX U894 ( .A(\Reg_Bank/registers[12][3] ), .B(n171), .S(n213), .Z(
        \Reg_Bank/n3385 ) );
  MUX U895 ( .A(\Reg_Bank/registers[12][2] ), .B(n172), .S(n213), .Z(
        \Reg_Bank/n3384 ) );
  MUX U896 ( .A(\Reg_Bank/registers[12][1] ), .B(n174), .S(n213), .Z(
        \Reg_Bank/n3383 ) );
  MUX U897 ( .A(\Reg_Bank/registers[12][0] ), .B(n175), .S(n213), .Z(
        \Reg_Bank/n3382 ) );
  ANDN U898 ( .B(n186), .A(n210), .Z(n213) );
  MUX U899 ( .A(\Reg_Bank/registers[11][31] ), .B(n142), .S(n214), .Z(
        \Reg_Bank/n3381 ) );
  MUX U900 ( .A(\Reg_Bank/registers[11][30] ), .B(n144), .S(n214), .Z(
        \Reg_Bank/n3380 ) );
  MUX U901 ( .A(\Reg_Bank/registers[11][29] ), .B(n145), .S(n214), .Z(
        \Reg_Bank/n3379 ) );
  MUX U902 ( .A(\Reg_Bank/registers[11][28] ), .B(n146), .S(n214), .Z(
        \Reg_Bank/n3378 ) );
  MUX U903 ( .A(\Reg_Bank/registers[11][27] ), .B(n147), .S(n214), .Z(
        \Reg_Bank/n3377 ) );
  MUX U904 ( .A(\Reg_Bank/registers[11][26] ), .B(n148), .S(n214), .Z(
        \Reg_Bank/n3376 ) );
  MUX U905 ( .A(\Reg_Bank/registers[11][25] ), .B(n149), .S(n214), .Z(
        \Reg_Bank/n3375 ) );
  MUX U906 ( .A(\Reg_Bank/registers[11][24] ), .B(n150), .S(n214), .Z(
        \Reg_Bank/n3374 ) );
  MUX U907 ( .A(\Reg_Bank/registers[11][23] ), .B(n151), .S(n214), .Z(
        \Reg_Bank/n3373 ) );
  MUX U908 ( .A(\Reg_Bank/registers[11][22] ), .B(n152), .S(n214), .Z(
        \Reg_Bank/n3372 ) );
  MUX U909 ( .A(\Reg_Bank/registers[11][21] ), .B(n153), .S(n214), .Z(
        \Reg_Bank/n3371 ) );
  MUX U910 ( .A(\Reg_Bank/registers[11][20] ), .B(n154), .S(n214), .Z(
        \Reg_Bank/n3370 ) );
  MUX U911 ( .A(\Reg_Bank/registers[11][19] ), .B(n155), .S(n214), .Z(
        \Reg_Bank/n3369 ) );
  MUX U912 ( .A(\Reg_Bank/registers[11][18] ), .B(n156), .S(n214), .Z(
        \Reg_Bank/n3368 ) );
  MUX U913 ( .A(\Reg_Bank/registers[11][17] ), .B(n157), .S(n214), .Z(
        \Reg_Bank/n3367 ) );
  MUX U914 ( .A(\Reg_Bank/registers[11][16] ), .B(n158), .S(n214), .Z(
        \Reg_Bank/n3366 ) );
  MUX U915 ( .A(\Reg_Bank/registers[11][15] ), .B(n159), .S(n214), .Z(
        \Reg_Bank/n3365 ) );
  MUX U916 ( .A(\Reg_Bank/registers[11][14] ), .B(n160), .S(n214), .Z(
        \Reg_Bank/n3364 ) );
  MUX U917 ( .A(\Reg_Bank/registers[11][13] ), .B(n161), .S(n214), .Z(
        \Reg_Bank/n3363 ) );
  MUX U918 ( .A(\Reg_Bank/registers[11][12] ), .B(n162), .S(n214), .Z(
        \Reg_Bank/n3362 ) );
  MUX U919 ( .A(\Reg_Bank/registers[11][11] ), .B(n163), .S(n214), .Z(
        \Reg_Bank/n3361 ) );
  MUX U920 ( .A(\Reg_Bank/registers[11][10] ), .B(n164), .S(n214), .Z(
        \Reg_Bank/n3360 ) );
  MUX U921 ( .A(\Reg_Bank/registers[11][9] ), .B(n165), .S(n214), .Z(
        \Reg_Bank/n3359 ) );
  MUX U922 ( .A(\Reg_Bank/registers[11][8] ), .B(n166), .S(n214), .Z(
        \Reg_Bank/n3358 ) );
  MUX U923 ( .A(\Reg_Bank/registers[11][7] ), .B(n167), .S(n214), .Z(
        \Reg_Bank/n3357 ) );
  MUX U924 ( .A(\Reg_Bank/registers[11][6] ), .B(n168), .S(n214), .Z(
        \Reg_Bank/n3356 ) );
  MUX U925 ( .A(\Reg_Bank/registers[11][5] ), .B(n169), .S(n214), .Z(
        \Reg_Bank/n3355 ) );
  MUX U926 ( .A(\Reg_Bank/registers[11][4] ), .B(n170), .S(n214), .Z(
        \Reg_Bank/n3354 ) );
  MUX U927 ( .A(\Reg_Bank/registers[11][3] ), .B(n171), .S(n214), .Z(
        \Reg_Bank/n3353 ) );
  MUX U928 ( .A(\Reg_Bank/registers[11][2] ), .B(n172), .S(n214), .Z(
        \Reg_Bank/n3352 ) );
  MUX U929 ( .A(\Reg_Bank/registers[11][1] ), .B(n174), .S(n214), .Z(
        \Reg_Bank/n3351 ) );
  MUX U930 ( .A(\Reg_Bank/registers[11][0] ), .B(n175), .S(n214), .Z(
        \Reg_Bank/n3350 ) );
  NOR U931 ( .A(n215), .B(n210), .Z(n214) );
  MUX U932 ( .A(\Reg_Bank/registers[10][31] ), .B(n142), .S(n216), .Z(
        \Reg_Bank/n3349 ) );
  MUX U933 ( .A(\Reg_Bank/registers[10][30] ), .B(n144), .S(n216), .Z(
        \Reg_Bank/n3348 ) );
  MUX U934 ( .A(\Reg_Bank/registers[10][29] ), .B(n145), .S(n216), .Z(
        \Reg_Bank/n3347 ) );
  MUX U935 ( .A(\Reg_Bank/registers[10][28] ), .B(n146), .S(n216), .Z(
        \Reg_Bank/n3346 ) );
  MUX U936 ( .A(\Reg_Bank/registers[10][27] ), .B(n147), .S(n216), .Z(
        \Reg_Bank/n3345 ) );
  MUX U937 ( .A(\Reg_Bank/registers[10][26] ), .B(n148), .S(n216), .Z(
        \Reg_Bank/n3344 ) );
  MUX U938 ( .A(\Reg_Bank/registers[10][25] ), .B(n149), .S(n216), .Z(
        \Reg_Bank/n3343 ) );
  MUX U939 ( .A(\Reg_Bank/registers[10][24] ), .B(n150), .S(n216), .Z(
        \Reg_Bank/n3342 ) );
  MUX U940 ( .A(\Reg_Bank/registers[10][23] ), .B(n151), .S(n216), .Z(
        \Reg_Bank/n3341 ) );
  MUX U941 ( .A(\Reg_Bank/registers[10][22] ), .B(n152), .S(n216), .Z(
        \Reg_Bank/n3340 ) );
  MUX U942 ( .A(\Reg_Bank/registers[10][21] ), .B(n153), .S(n216), .Z(
        \Reg_Bank/n3339 ) );
  MUX U943 ( .A(\Reg_Bank/registers[10][20] ), .B(n154), .S(n216), .Z(
        \Reg_Bank/n3338 ) );
  MUX U944 ( .A(\Reg_Bank/registers[10][19] ), .B(n155), .S(n216), .Z(
        \Reg_Bank/n3337 ) );
  MUX U945 ( .A(\Reg_Bank/registers[10][18] ), .B(n156), .S(n216), .Z(
        \Reg_Bank/n3336 ) );
  MUX U946 ( .A(\Reg_Bank/registers[10][17] ), .B(n157), .S(n216), .Z(
        \Reg_Bank/n3335 ) );
  MUX U947 ( .A(\Reg_Bank/registers[10][16] ), .B(n158), .S(n216), .Z(
        \Reg_Bank/n3334 ) );
  MUX U948 ( .A(\Reg_Bank/registers[10][15] ), .B(n159), .S(n216), .Z(
        \Reg_Bank/n3333 ) );
  MUX U949 ( .A(\Reg_Bank/registers[10][14] ), .B(n160), .S(n216), .Z(
        \Reg_Bank/n3332 ) );
  MUX U950 ( .A(\Reg_Bank/registers[10][13] ), .B(n161), .S(n216), .Z(
        \Reg_Bank/n3331 ) );
  MUX U951 ( .A(\Reg_Bank/registers[10][12] ), .B(n162), .S(n216), .Z(
        \Reg_Bank/n3330 ) );
  MUX U952 ( .A(\Reg_Bank/registers[10][11] ), .B(n163), .S(n216), .Z(
        \Reg_Bank/n3329 ) );
  MUX U953 ( .A(\Reg_Bank/registers[10][10] ), .B(n164), .S(n216), .Z(
        \Reg_Bank/n3328 ) );
  MUX U954 ( .A(\Reg_Bank/registers[10][9] ), .B(n165), .S(n216), .Z(
        \Reg_Bank/n3327 ) );
  MUX U955 ( .A(\Reg_Bank/registers[10][8] ), .B(n166), .S(n216), .Z(
        \Reg_Bank/n3326 ) );
  MUX U956 ( .A(\Reg_Bank/registers[10][7] ), .B(n167), .S(n216), .Z(
        \Reg_Bank/n3325 ) );
  MUX U957 ( .A(\Reg_Bank/registers[10][6] ), .B(n168), .S(n216), .Z(
        \Reg_Bank/n3324 ) );
  MUX U958 ( .A(\Reg_Bank/registers[10][5] ), .B(n169), .S(n216), .Z(
        \Reg_Bank/n3323 ) );
  MUX U959 ( .A(\Reg_Bank/registers[10][4] ), .B(n170), .S(n216), .Z(
        \Reg_Bank/n3322 ) );
  MUX U960 ( .A(\Reg_Bank/registers[10][3] ), .B(n171), .S(n216), .Z(
        \Reg_Bank/n3321 ) );
  MUX U961 ( .A(\Reg_Bank/registers[10][2] ), .B(n172), .S(n216), .Z(
        \Reg_Bank/n3320 ) );
  MUX U962 ( .A(\Reg_Bank/registers[10][1] ), .B(n174), .S(n216), .Z(
        \Reg_Bank/n3319 ) );
  MUX U963 ( .A(\Reg_Bank/registers[10][0] ), .B(n175), .S(n216), .Z(
        \Reg_Bank/n3318 ) );
  NOR U964 ( .A(n217), .B(n210), .Z(n216) );
  MUX U965 ( .A(\Reg_Bank/registers[9][31] ), .B(n142), .S(n218), .Z(
        \Reg_Bank/n3317 ) );
  MUX U966 ( .A(\Reg_Bank/registers[9][30] ), .B(n144), .S(n218), .Z(
        \Reg_Bank/n3316 ) );
  MUX U967 ( .A(\Reg_Bank/registers[9][29] ), .B(n145), .S(n218), .Z(
        \Reg_Bank/n3315 ) );
  MUX U968 ( .A(\Reg_Bank/registers[9][28] ), .B(n146), .S(n218), .Z(
        \Reg_Bank/n3314 ) );
  MUX U969 ( .A(\Reg_Bank/registers[9][27] ), .B(n147), .S(n218), .Z(
        \Reg_Bank/n3313 ) );
  MUX U970 ( .A(\Reg_Bank/registers[9][26] ), .B(n148), .S(n218), .Z(
        \Reg_Bank/n3312 ) );
  MUX U971 ( .A(\Reg_Bank/registers[9][25] ), .B(n149), .S(n218), .Z(
        \Reg_Bank/n3311 ) );
  MUX U972 ( .A(\Reg_Bank/registers[9][24] ), .B(n150), .S(n218), .Z(
        \Reg_Bank/n3310 ) );
  MUX U973 ( .A(\Reg_Bank/registers[9][23] ), .B(n151), .S(n218), .Z(
        \Reg_Bank/n3309 ) );
  MUX U974 ( .A(\Reg_Bank/registers[9][22] ), .B(n152), .S(n218), .Z(
        \Reg_Bank/n3308 ) );
  MUX U975 ( .A(\Reg_Bank/registers[9][21] ), .B(n153), .S(n218), .Z(
        \Reg_Bank/n3307 ) );
  MUX U976 ( .A(\Reg_Bank/registers[9][20] ), .B(n154), .S(n218), .Z(
        \Reg_Bank/n3306 ) );
  MUX U977 ( .A(\Reg_Bank/registers[9][19] ), .B(n155), .S(n218), .Z(
        \Reg_Bank/n3305 ) );
  MUX U978 ( .A(\Reg_Bank/registers[9][18] ), .B(n156), .S(n218), .Z(
        \Reg_Bank/n3304 ) );
  MUX U979 ( .A(\Reg_Bank/registers[9][17] ), .B(n157), .S(n218), .Z(
        \Reg_Bank/n3303 ) );
  MUX U980 ( .A(\Reg_Bank/registers[9][16] ), .B(n158), .S(n218), .Z(
        \Reg_Bank/n3302 ) );
  MUX U981 ( .A(\Reg_Bank/registers[9][15] ), .B(n159), .S(n218), .Z(
        \Reg_Bank/n3301 ) );
  MUX U982 ( .A(\Reg_Bank/registers[9][14] ), .B(n160), .S(n218), .Z(
        \Reg_Bank/n3300 ) );
  MUX U983 ( .A(\Reg_Bank/registers[9][13] ), .B(n161), .S(n218), .Z(
        \Reg_Bank/n3299 ) );
  MUX U984 ( .A(\Reg_Bank/registers[9][12] ), .B(n162), .S(n218), .Z(
        \Reg_Bank/n3298 ) );
  MUX U985 ( .A(\Reg_Bank/registers[9][11] ), .B(n163), .S(n218), .Z(
        \Reg_Bank/n3297 ) );
  MUX U986 ( .A(\Reg_Bank/registers[9][10] ), .B(n164), .S(n218), .Z(
        \Reg_Bank/n3296 ) );
  MUX U987 ( .A(\Reg_Bank/registers[9][9] ), .B(n165), .S(n218), .Z(
        \Reg_Bank/n3295 ) );
  MUX U988 ( .A(\Reg_Bank/registers[9][8] ), .B(n166), .S(n218), .Z(
        \Reg_Bank/n3294 ) );
  MUX U989 ( .A(\Reg_Bank/registers[9][7] ), .B(n167), .S(n218), .Z(
        \Reg_Bank/n3293 ) );
  MUX U990 ( .A(\Reg_Bank/registers[9][6] ), .B(n168), .S(n218), .Z(
        \Reg_Bank/n3292 ) );
  MUX U991 ( .A(\Reg_Bank/registers[9][5] ), .B(n169), .S(n218), .Z(
        \Reg_Bank/n3291 ) );
  MUX U992 ( .A(\Reg_Bank/registers[9][4] ), .B(n170), .S(n218), .Z(
        \Reg_Bank/n3290 ) );
  MUX U993 ( .A(\Reg_Bank/registers[9][3] ), .B(n171), .S(n218), .Z(
        \Reg_Bank/n3289 ) );
  MUX U994 ( .A(\Reg_Bank/registers[9][2] ), .B(n172), .S(n218), .Z(
        \Reg_Bank/n3288 ) );
  MUX U995 ( .A(\Reg_Bank/registers[9][1] ), .B(n174), .S(n218), .Z(
        \Reg_Bank/n3287 ) );
  MUX U996 ( .A(\Reg_Bank/registers[9][0] ), .B(n175), .S(n218), .Z(
        \Reg_Bank/n3286 ) );
  NOR U997 ( .A(n219), .B(n210), .Z(n218) );
  MUX U998 ( .A(\Reg_Bank/registers[8][31] ), .B(n142), .S(n220), .Z(
        \Reg_Bank/n3285 ) );
  MUX U999 ( .A(\Reg_Bank/registers[8][30] ), .B(n144), .S(n220), .Z(
        \Reg_Bank/n3284 ) );
  MUX U1000 ( .A(\Reg_Bank/registers[8][29] ), .B(n145), .S(n220), .Z(
        \Reg_Bank/n3283 ) );
  MUX U1001 ( .A(\Reg_Bank/registers[8][28] ), .B(n146), .S(n220), .Z(
        \Reg_Bank/n3282 ) );
  MUX U1002 ( .A(\Reg_Bank/registers[8][27] ), .B(n147), .S(n220), .Z(
        \Reg_Bank/n3281 ) );
  MUX U1003 ( .A(\Reg_Bank/registers[8][26] ), .B(n148), .S(n220), .Z(
        \Reg_Bank/n3280 ) );
  MUX U1004 ( .A(\Reg_Bank/registers[8][25] ), .B(n149), .S(n220), .Z(
        \Reg_Bank/n3279 ) );
  MUX U1005 ( .A(\Reg_Bank/registers[8][24] ), .B(n150), .S(n220), .Z(
        \Reg_Bank/n3278 ) );
  MUX U1006 ( .A(\Reg_Bank/registers[8][23] ), .B(n151), .S(n220), .Z(
        \Reg_Bank/n3277 ) );
  MUX U1007 ( .A(\Reg_Bank/registers[8][22] ), .B(n152), .S(n220), .Z(
        \Reg_Bank/n3276 ) );
  MUX U1008 ( .A(\Reg_Bank/registers[8][21] ), .B(n153), .S(n220), .Z(
        \Reg_Bank/n3275 ) );
  MUX U1009 ( .A(\Reg_Bank/registers[8][20] ), .B(n154), .S(n220), .Z(
        \Reg_Bank/n3274 ) );
  MUX U1010 ( .A(\Reg_Bank/registers[8][19] ), .B(n155), .S(n220), .Z(
        \Reg_Bank/n3273 ) );
  MUX U1011 ( .A(\Reg_Bank/registers[8][18] ), .B(n156), .S(n220), .Z(
        \Reg_Bank/n3272 ) );
  MUX U1012 ( .A(\Reg_Bank/registers[8][17] ), .B(n157), .S(n220), .Z(
        \Reg_Bank/n3271 ) );
  MUX U1013 ( .A(\Reg_Bank/registers[8][16] ), .B(n158), .S(n220), .Z(
        \Reg_Bank/n3270 ) );
  MUX U1014 ( .A(\Reg_Bank/registers[8][15] ), .B(n159), .S(n220), .Z(
        \Reg_Bank/n3269 ) );
  MUX U1015 ( .A(\Reg_Bank/registers[8][14] ), .B(n160), .S(n220), .Z(
        \Reg_Bank/n3268 ) );
  MUX U1016 ( .A(\Reg_Bank/registers[8][13] ), .B(n161), .S(n220), .Z(
        \Reg_Bank/n3267 ) );
  MUX U1017 ( .A(\Reg_Bank/registers[8][12] ), .B(n162), .S(n220), .Z(
        \Reg_Bank/n3266 ) );
  MUX U1018 ( .A(\Reg_Bank/registers[8][11] ), .B(n163), .S(n220), .Z(
        \Reg_Bank/n3265 ) );
  MUX U1019 ( .A(\Reg_Bank/registers[8][10] ), .B(n164), .S(n220), .Z(
        \Reg_Bank/n3264 ) );
  MUX U1020 ( .A(\Reg_Bank/registers[8][9] ), .B(n165), .S(n220), .Z(
        \Reg_Bank/n3263 ) );
  MUX U1021 ( .A(\Reg_Bank/registers[8][8] ), .B(n166), .S(n220), .Z(
        \Reg_Bank/n3262 ) );
  MUX U1022 ( .A(\Reg_Bank/registers[8][7] ), .B(n167), .S(n220), .Z(
        \Reg_Bank/n3261 ) );
  MUX U1023 ( .A(\Reg_Bank/registers[8][6] ), .B(n168), .S(n220), .Z(
        \Reg_Bank/n3260 ) );
  MUX U1024 ( .A(\Reg_Bank/registers[8][5] ), .B(n169), .S(n220), .Z(
        \Reg_Bank/n3259 ) );
  MUX U1025 ( .A(\Reg_Bank/registers[8][4] ), .B(n170), .S(n220), .Z(
        \Reg_Bank/n3258 ) );
  MUX U1026 ( .A(\Reg_Bank/registers[8][3] ), .B(n171), .S(n220), .Z(
        \Reg_Bank/n3257 ) );
  MUX U1027 ( .A(\Reg_Bank/registers[8][2] ), .B(n172), .S(n220), .Z(
        \Reg_Bank/n3256 ) );
  MUX U1028 ( .A(\Reg_Bank/registers[8][1] ), .B(n174), .S(n220), .Z(
        \Reg_Bank/n3255 ) );
  MUX U1029 ( .A(\Reg_Bank/registers[8][0] ), .B(n175), .S(n220), .Z(
        \Reg_Bank/n3254 ) );
  NOR U1030 ( .A(n206), .B(n210), .Z(n220) );
  NANDN U1031 ( .A(n195), .B(n207), .Z(n210) );
  NANDN U1032 ( .A(n221), .B(n222), .Z(n206) );
  MUX U1033 ( .A(\Reg_Bank/registers[7][31] ), .B(n142), .S(n223), .Z(
        \Reg_Bank/n3253 ) );
  MUX U1034 ( .A(\Reg_Bank/registers[7][30] ), .B(n144), .S(n223), .Z(
        \Reg_Bank/n3252 ) );
  MUX U1035 ( .A(\Reg_Bank/registers[7][29] ), .B(n145), .S(n223), .Z(
        \Reg_Bank/n3251 ) );
  MUX U1036 ( .A(\Reg_Bank/registers[7][28] ), .B(n146), .S(n223), .Z(
        \Reg_Bank/n3250 ) );
  MUX U1037 ( .A(\Reg_Bank/registers[7][27] ), .B(n147), .S(n223), .Z(
        \Reg_Bank/n3249 ) );
  MUX U1038 ( .A(\Reg_Bank/registers[7][26] ), .B(n148), .S(n223), .Z(
        \Reg_Bank/n3248 ) );
  MUX U1039 ( .A(\Reg_Bank/registers[7][25] ), .B(n149), .S(n223), .Z(
        \Reg_Bank/n3247 ) );
  MUX U1040 ( .A(\Reg_Bank/registers[7][24] ), .B(n150), .S(n223), .Z(
        \Reg_Bank/n3246 ) );
  MUX U1041 ( .A(\Reg_Bank/registers[7][23] ), .B(n151), .S(n223), .Z(
        \Reg_Bank/n3245 ) );
  MUX U1042 ( .A(\Reg_Bank/registers[7][22] ), .B(n152), .S(n223), .Z(
        \Reg_Bank/n3244 ) );
  MUX U1043 ( .A(\Reg_Bank/registers[7][21] ), .B(n153), .S(n223), .Z(
        \Reg_Bank/n3243 ) );
  MUX U1044 ( .A(\Reg_Bank/registers[7][20] ), .B(n154), .S(n223), .Z(
        \Reg_Bank/n3242 ) );
  MUX U1045 ( .A(\Reg_Bank/registers[7][19] ), .B(n155), .S(n223), .Z(
        \Reg_Bank/n3241 ) );
  MUX U1046 ( .A(\Reg_Bank/registers[7][18] ), .B(n156), .S(n223), .Z(
        \Reg_Bank/n3240 ) );
  MUX U1047 ( .A(\Reg_Bank/registers[7][17] ), .B(n157), .S(n223), .Z(
        \Reg_Bank/n3239 ) );
  MUX U1048 ( .A(\Reg_Bank/registers[7][16] ), .B(n158), .S(n223), .Z(
        \Reg_Bank/n3238 ) );
  MUX U1049 ( .A(\Reg_Bank/registers[7][15] ), .B(n159), .S(n223), .Z(
        \Reg_Bank/n3237 ) );
  MUX U1050 ( .A(\Reg_Bank/registers[7][14] ), .B(n160), .S(n223), .Z(
        \Reg_Bank/n3236 ) );
  MUX U1051 ( .A(\Reg_Bank/registers[7][13] ), .B(n161), .S(n223), .Z(
        \Reg_Bank/n3235 ) );
  MUX U1052 ( .A(\Reg_Bank/registers[7][12] ), .B(n162), .S(n223), .Z(
        \Reg_Bank/n3234 ) );
  MUX U1053 ( .A(\Reg_Bank/registers[7][11] ), .B(n163), .S(n223), .Z(
        \Reg_Bank/n3233 ) );
  MUX U1054 ( .A(\Reg_Bank/registers[7][10] ), .B(n164), .S(n223), .Z(
        \Reg_Bank/n3232 ) );
  MUX U1055 ( .A(\Reg_Bank/registers[7][9] ), .B(n165), .S(n223), .Z(
        \Reg_Bank/n3231 ) );
  MUX U1056 ( .A(\Reg_Bank/registers[7][8] ), .B(n166), .S(n223), .Z(
        \Reg_Bank/n3230 ) );
  MUX U1057 ( .A(\Reg_Bank/registers[7][7] ), .B(n167), .S(n223), .Z(
        \Reg_Bank/n3229 ) );
  MUX U1058 ( .A(\Reg_Bank/registers[7][6] ), .B(n168), .S(n223), .Z(
        \Reg_Bank/n3228 ) );
  MUX U1059 ( .A(\Reg_Bank/registers[7][5] ), .B(n169), .S(n223), .Z(
        \Reg_Bank/n3227 ) );
  MUX U1060 ( .A(\Reg_Bank/registers[7][4] ), .B(n170), .S(n223), .Z(
        \Reg_Bank/n3226 ) );
  MUX U1061 ( .A(\Reg_Bank/registers[7][3] ), .B(n171), .S(n223), .Z(
        \Reg_Bank/n3225 ) );
  MUX U1062 ( .A(\Reg_Bank/registers[7][2] ), .B(n172), .S(n223), .Z(
        \Reg_Bank/n3224 ) );
  MUX U1063 ( .A(\Reg_Bank/registers[7][1] ), .B(n174), .S(n223), .Z(
        \Reg_Bank/n3223 ) );
  MUX U1064 ( .A(\Reg_Bank/registers[7][0] ), .B(n175), .S(n223), .Z(
        \Reg_Bank/n3222 ) );
  ANDN U1065 ( .B(n224), .A(n177), .Z(n223) );
  NAND U1066 ( .A(n221), .B(n225), .Z(n177) );
  MUX U1067 ( .A(\Reg_Bank/registers[6][31] ), .B(n142), .S(n226), .Z(
        \Reg_Bank/n3221 ) );
  MUX U1068 ( .A(\Reg_Bank/registers[6][30] ), .B(n144), .S(n226), .Z(
        \Reg_Bank/n3220 ) );
  MUX U1069 ( .A(\Reg_Bank/registers[6][29] ), .B(n145), .S(n226), .Z(
        \Reg_Bank/n3219 ) );
  MUX U1070 ( .A(\Reg_Bank/registers[6][28] ), .B(n146), .S(n226), .Z(
        \Reg_Bank/n3218 ) );
  MUX U1071 ( .A(\Reg_Bank/registers[6][27] ), .B(n147), .S(n226), .Z(
        \Reg_Bank/n3217 ) );
  MUX U1072 ( .A(\Reg_Bank/registers[6][26] ), .B(n148), .S(n226), .Z(
        \Reg_Bank/n3216 ) );
  MUX U1073 ( .A(\Reg_Bank/registers[6][25] ), .B(n149), .S(n226), .Z(
        \Reg_Bank/n3215 ) );
  MUX U1074 ( .A(\Reg_Bank/registers[6][24] ), .B(n150), .S(n226), .Z(
        \Reg_Bank/n3214 ) );
  MUX U1075 ( .A(\Reg_Bank/registers[6][23] ), .B(n151), .S(n226), .Z(
        \Reg_Bank/n3213 ) );
  MUX U1076 ( .A(\Reg_Bank/registers[6][22] ), .B(n152), .S(n226), .Z(
        \Reg_Bank/n3212 ) );
  MUX U1077 ( .A(\Reg_Bank/registers[6][21] ), .B(n153), .S(n226), .Z(
        \Reg_Bank/n3211 ) );
  MUX U1078 ( .A(\Reg_Bank/registers[6][20] ), .B(n154), .S(n226), .Z(
        \Reg_Bank/n3210 ) );
  MUX U1079 ( .A(\Reg_Bank/registers[6][19] ), .B(n155), .S(n226), .Z(
        \Reg_Bank/n3209 ) );
  MUX U1080 ( .A(\Reg_Bank/registers[6][18] ), .B(n156), .S(n226), .Z(
        \Reg_Bank/n3208 ) );
  MUX U1081 ( .A(\Reg_Bank/registers[6][17] ), .B(n157), .S(n226), .Z(
        \Reg_Bank/n3207 ) );
  MUX U1082 ( .A(\Reg_Bank/registers[6][16] ), .B(n158), .S(n226), .Z(
        \Reg_Bank/n3206 ) );
  MUX U1083 ( .A(\Reg_Bank/registers[6][15] ), .B(n159), .S(n226), .Z(
        \Reg_Bank/n3205 ) );
  MUX U1084 ( .A(\Reg_Bank/registers[6][14] ), .B(n160), .S(n226), .Z(
        \Reg_Bank/n3204 ) );
  MUX U1085 ( .A(\Reg_Bank/registers[6][13] ), .B(n161), .S(n226), .Z(
        \Reg_Bank/n3203 ) );
  MUX U1086 ( .A(\Reg_Bank/registers[6][12] ), .B(n162), .S(n226), .Z(
        \Reg_Bank/n3202 ) );
  MUX U1087 ( .A(\Reg_Bank/registers[6][11] ), .B(n163), .S(n226), .Z(
        \Reg_Bank/n3201 ) );
  MUX U1088 ( .A(\Reg_Bank/registers[6][10] ), .B(n164), .S(n226), .Z(
        \Reg_Bank/n3200 ) );
  MUX U1089 ( .A(\Reg_Bank/registers[6][9] ), .B(n165), .S(n226), .Z(
        \Reg_Bank/n3199 ) );
  MUX U1090 ( .A(\Reg_Bank/registers[6][8] ), .B(n166), .S(n226), .Z(
        \Reg_Bank/n3198 ) );
  MUX U1091 ( .A(\Reg_Bank/registers[6][7] ), .B(n167), .S(n226), .Z(
        \Reg_Bank/n3197 ) );
  MUX U1092 ( .A(\Reg_Bank/registers[6][6] ), .B(n168), .S(n226), .Z(
        \Reg_Bank/n3196 ) );
  MUX U1093 ( .A(\Reg_Bank/registers[6][5] ), .B(n169), .S(n226), .Z(
        \Reg_Bank/n3195 ) );
  MUX U1094 ( .A(\Reg_Bank/registers[6][4] ), .B(n170), .S(n226), .Z(
        \Reg_Bank/n3194 ) );
  MUX U1095 ( .A(\Reg_Bank/registers[6][3] ), .B(n171), .S(n226), .Z(
        \Reg_Bank/n3193 ) );
  MUX U1096 ( .A(\Reg_Bank/registers[6][2] ), .B(n172), .S(n226), .Z(
        \Reg_Bank/n3192 ) );
  MUX U1097 ( .A(\Reg_Bank/registers[6][1] ), .B(n174), .S(n226), .Z(
        \Reg_Bank/n3191 ) );
  MUX U1098 ( .A(\Reg_Bank/registers[6][0] ), .B(n175), .S(n226), .Z(
        \Reg_Bank/n3190 ) );
  AND U1099 ( .A(n180), .B(n224), .Z(n226) );
  AND U1100 ( .A(n221), .B(n227), .Z(n180) );
  MUX U1101 ( .A(\Reg_Bank/registers[5][31] ), .B(n142), .S(n228), .Z(
        \Reg_Bank/n3189 ) );
  MUX U1102 ( .A(\Reg_Bank/registers[5][30] ), .B(n144), .S(n228), .Z(
        \Reg_Bank/n3188 ) );
  MUX U1103 ( .A(\Reg_Bank/registers[5][29] ), .B(n145), .S(n228), .Z(
        \Reg_Bank/n3187 ) );
  MUX U1104 ( .A(\Reg_Bank/registers[5][28] ), .B(n146), .S(n228), .Z(
        \Reg_Bank/n3186 ) );
  MUX U1105 ( .A(\Reg_Bank/registers[5][27] ), .B(n147), .S(n228), .Z(
        \Reg_Bank/n3185 ) );
  MUX U1106 ( .A(\Reg_Bank/registers[5][26] ), .B(n148), .S(n228), .Z(
        \Reg_Bank/n3184 ) );
  MUX U1107 ( .A(\Reg_Bank/registers[5][25] ), .B(n149), .S(n228), .Z(
        \Reg_Bank/n3183 ) );
  MUX U1108 ( .A(\Reg_Bank/registers[5][24] ), .B(n150), .S(n228), .Z(
        \Reg_Bank/n3182 ) );
  MUX U1109 ( .A(\Reg_Bank/registers[5][23] ), .B(n151), .S(n228), .Z(
        \Reg_Bank/n3181 ) );
  MUX U1110 ( .A(\Reg_Bank/registers[5][22] ), .B(n152), .S(n228), .Z(
        \Reg_Bank/n3180 ) );
  MUX U1111 ( .A(\Reg_Bank/registers[5][21] ), .B(n153), .S(n228), .Z(
        \Reg_Bank/n3179 ) );
  MUX U1112 ( .A(\Reg_Bank/registers[5][20] ), .B(n154), .S(n228), .Z(
        \Reg_Bank/n3178 ) );
  MUX U1113 ( .A(\Reg_Bank/registers[5][19] ), .B(n155), .S(n228), .Z(
        \Reg_Bank/n3177 ) );
  MUX U1114 ( .A(\Reg_Bank/registers[5][18] ), .B(n156), .S(n228), .Z(
        \Reg_Bank/n3176 ) );
  MUX U1115 ( .A(\Reg_Bank/registers[5][17] ), .B(n157), .S(n228), .Z(
        \Reg_Bank/n3175 ) );
  MUX U1116 ( .A(\Reg_Bank/registers[5][16] ), .B(n158), .S(n228), .Z(
        \Reg_Bank/n3174 ) );
  MUX U1117 ( .A(\Reg_Bank/registers[5][15] ), .B(n159), .S(n228), .Z(
        \Reg_Bank/n3173 ) );
  MUX U1118 ( .A(\Reg_Bank/registers[5][14] ), .B(n160), .S(n228), .Z(
        \Reg_Bank/n3172 ) );
  MUX U1119 ( .A(\Reg_Bank/registers[5][13] ), .B(n161), .S(n228), .Z(
        \Reg_Bank/n3171 ) );
  MUX U1120 ( .A(\Reg_Bank/registers[5][12] ), .B(n162), .S(n228), .Z(
        \Reg_Bank/n3170 ) );
  MUX U1121 ( .A(\Reg_Bank/registers[5][11] ), .B(n163), .S(n228), .Z(
        \Reg_Bank/n3169 ) );
  MUX U1122 ( .A(\Reg_Bank/registers[5][10] ), .B(n164), .S(n228), .Z(
        \Reg_Bank/n3168 ) );
  MUX U1123 ( .A(\Reg_Bank/registers[5][9] ), .B(n165), .S(n228), .Z(
        \Reg_Bank/n3167 ) );
  MUX U1124 ( .A(\Reg_Bank/registers[5][8] ), .B(n166), .S(n228), .Z(
        \Reg_Bank/n3166 ) );
  MUX U1125 ( .A(\Reg_Bank/registers[5][7] ), .B(n167), .S(n228), .Z(
        \Reg_Bank/n3165 ) );
  MUX U1126 ( .A(\Reg_Bank/registers[5][6] ), .B(n168), .S(n228), .Z(
        \Reg_Bank/n3164 ) );
  MUX U1127 ( .A(\Reg_Bank/registers[5][5] ), .B(n169), .S(n228), .Z(
        \Reg_Bank/n3163 ) );
  MUX U1128 ( .A(\Reg_Bank/registers[5][4] ), .B(n170), .S(n228), .Z(
        \Reg_Bank/n3162 ) );
  MUX U1129 ( .A(\Reg_Bank/registers[5][3] ), .B(n171), .S(n228), .Z(
        \Reg_Bank/n3161 ) );
  MUX U1130 ( .A(\Reg_Bank/registers[5][2] ), .B(n172), .S(n228), .Z(
        \Reg_Bank/n3160 ) );
  MUX U1131 ( .A(\Reg_Bank/registers[5][1] ), .B(n174), .S(n228), .Z(
        \Reg_Bank/n3159 ) );
  MUX U1132 ( .A(\Reg_Bank/registers[5][0] ), .B(n175), .S(n228), .Z(
        \Reg_Bank/n3158 ) );
  AND U1133 ( .A(n183), .B(n224), .Z(n228) );
  AND U1134 ( .A(n221), .B(n229), .Z(n183) );
  MUX U1135 ( .A(\Reg_Bank/registers[4][31] ), .B(n142), .S(n230), .Z(
        \Reg_Bank/n3157 ) );
  MUX U1136 ( .A(\Reg_Bank/registers[4][30] ), .B(n144), .S(n230), .Z(
        \Reg_Bank/n3156 ) );
  MUX U1137 ( .A(\Reg_Bank/registers[4][29] ), .B(n145), .S(n230), .Z(
        \Reg_Bank/n3155 ) );
  MUX U1138 ( .A(\Reg_Bank/registers[4][28] ), .B(n146), .S(n230), .Z(
        \Reg_Bank/n3154 ) );
  MUX U1139 ( .A(\Reg_Bank/registers[4][27] ), .B(n147), .S(n230), .Z(
        \Reg_Bank/n3153 ) );
  MUX U1140 ( .A(\Reg_Bank/registers[4][26] ), .B(n148), .S(n230), .Z(
        \Reg_Bank/n3152 ) );
  MUX U1141 ( .A(\Reg_Bank/registers[4][25] ), .B(n149), .S(n230), .Z(
        \Reg_Bank/n3151 ) );
  MUX U1142 ( .A(\Reg_Bank/registers[4][24] ), .B(n150), .S(n230), .Z(
        \Reg_Bank/n3150 ) );
  MUX U1143 ( .A(\Reg_Bank/registers[4][23] ), .B(n151), .S(n230), .Z(
        \Reg_Bank/n3149 ) );
  MUX U1144 ( .A(\Reg_Bank/registers[4][22] ), .B(n152), .S(n230), .Z(
        \Reg_Bank/n3148 ) );
  MUX U1145 ( .A(\Reg_Bank/registers[4][21] ), .B(n153), .S(n230), .Z(
        \Reg_Bank/n3147 ) );
  MUX U1146 ( .A(\Reg_Bank/registers[4][20] ), .B(n154), .S(n230), .Z(
        \Reg_Bank/n3146 ) );
  MUX U1147 ( .A(\Reg_Bank/registers[4][19] ), .B(n155), .S(n230), .Z(
        \Reg_Bank/n3145 ) );
  MUX U1148 ( .A(\Reg_Bank/registers[4][18] ), .B(n156), .S(n230), .Z(
        \Reg_Bank/n3144 ) );
  MUX U1149 ( .A(\Reg_Bank/registers[4][17] ), .B(n157), .S(n230), .Z(
        \Reg_Bank/n3143 ) );
  MUX U1150 ( .A(\Reg_Bank/registers[4][16] ), .B(n158), .S(n230), .Z(
        \Reg_Bank/n3142 ) );
  MUX U1151 ( .A(\Reg_Bank/registers[4][15] ), .B(n159), .S(n230), .Z(
        \Reg_Bank/n3141 ) );
  MUX U1152 ( .A(\Reg_Bank/registers[4][14] ), .B(n160), .S(n230), .Z(
        \Reg_Bank/n3140 ) );
  MUX U1153 ( .A(\Reg_Bank/registers[4][13] ), .B(n161), .S(n230), .Z(
        \Reg_Bank/n3139 ) );
  MUX U1154 ( .A(\Reg_Bank/registers[4][12] ), .B(n162), .S(n230), .Z(
        \Reg_Bank/n3138 ) );
  MUX U1155 ( .A(\Reg_Bank/registers[4][11] ), .B(n163), .S(n230), .Z(
        \Reg_Bank/n3137 ) );
  MUX U1156 ( .A(\Reg_Bank/registers[4][10] ), .B(n164), .S(n230), .Z(
        \Reg_Bank/n3136 ) );
  MUX U1157 ( .A(\Reg_Bank/registers[4][9] ), .B(n165), .S(n230), .Z(
        \Reg_Bank/n3135 ) );
  MUX U1158 ( .A(\Reg_Bank/registers[4][8] ), .B(n166), .S(n230), .Z(
        \Reg_Bank/n3134 ) );
  MUX U1159 ( .A(\Reg_Bank/registers[4][7] ), .B(n167), .S(n230), .Z(
        \Reg_Bank/n3133 ) );
  MUX U1160 ( .A(\Reg_Bank/registers[4][6] ), .B(n168), .S(n230), .Z(
        \Reg_Bank/n3132 ) );
  MUX U1161 ( .A(\Reg_Bank/registers[4][5] ), .B(n169), .S(n230), .Z(
        \Reg_Bank/n3131 ) );
  MUX U1162 ( .A(\Reg_Bank/registers[4][4] ), .B(n170), .S(n230), .Z(
        \Reg_Bank/n3130 ) );
  MUX U1163 ( .A(\Reg_Bank/registers[4][3] ), .B(n171), .S(n230), .Z(
        \Reg_Bank/n3129 ) );
  MUX U1164 ( .A(\Reg_Bank/registers[4][2] ), .B(n172), .S(n230), .Z(
        \Reg_Bank/n3128 ) );
  MUX U1165 ( .A(\Reg_Bank/registers[4][1] ), .B(n174), .S(n230), .Z(
        \Reg_Bank/n3127 ) );
  MUX U1166 ( .A(\Reg_Bank/registers[4][0] ), .B(n175), .S(n230), .Z(
        \Reg_Bank/n3126 ) );
  AND U1167 ( .A(n186), .B(n224), .Z(n230) );
  AND U1168 ( .A(n221), .B(n222), .Z(n186) );
  NOR U1169 ( .A(n231), .B(n232), .Z(n222) );
  MUX U1170 ( .A(\Reg_Bank/registers[3][31] ), .B(n142), .S(n233), .Z(
        \Reg_Bank/n3125 ) );
  MUX U1171 ( .A(\Reg_Bank/registers[3][30] ), .B(n144), .S(n233), .Z(
        \Reg_Bank/n3124 ) );
  MUX U1172 ( .A(\Reg_Bank/registers[3][29] ), .B(n145), .S(n233), .Z(
        \Reg_Bank/n3123 ) );
  MUX U1173 ( .A(\Reg_Bank/registers[3][28] ), .B(n146), .S(n233), .Z(
        \Reg_Bank/n3122 ) );
  MUX U1174 ( .A(\Reg_Bank/registers[3][27] ), .B(n147), .S(n233), .Z(
        \Reg_Bank/n3121 ) );
  MUX U1175 ( .A(\Reg_Bank/registers[3][26] ), .B(n148), .S(n233), .Z(
        \Reg_Bank/n3120 ) );
  MUX U1176 ( .A(\Reg_Bank/registers[3][25] ), .B(n149), .S(n233), .Z(
        \Reg_Bank/n3119 ) );
  MUX U1177 ( .A(\Reg_Bank/registers[3][24] ), .B(n150), .S(n233), .Z(
        \Reg_Bank/n3118 ) );
  MUX U1178 ( .A(\Reg_Bank/registers[3][23] ), .B(n151), .S(n233), .Z(
        \Reg_Bank/n3117 ) );
  MUX U1179 ( .A(\Reg_Bank/registers[3][22] ), .B(n152), .S(n233), .Z(
        \Reg_Bank/n3116 ) );
  MUX U1180 ( .A(\Reg_Bank/registers[3][21] ), .B(n153), .S(n233), .Z(
        \Reg_Bank/n3115 ) );
  MUX U1181 ( .A(\Reg_Bank/registers[3][20] ), .B(n154), .S(n233), .Z(
        \Reg_Bank/n3114 ) );
  MUX U1182 ( .A(\Reg_Bank/registers[3][19] ), .B(n155), .S(n233), .Z(
        \Reg_Bank/n3113 ) );
  MUX U1183 ( .A(\Reg_Bank/registers[3][18] ), .B(n156), .S(n233), .Z(
        \Reg_Bank/n3112 ) );
  MUX U1184 ( .A(\Reg_Bank/registers[3][17] ), .B(n157), .S(n233), .Z(
        \Reg_Bank/n3111 ) );
  MUX U1185 ( .A(\Reg_Bank/registers[3][16] ), .B(n158), .S(n233), .Z(
        \Reg_Bank/n3110 ) );
  MUX U1186 ( .A(\Reg_Bank/registers[3][15] ), .B(n159), .S(n233), .Z(
        \Reg_Bank/n3109 ) );
  MUX U1187 ( .A(\Reg_Bank/registers[3][14] ), .B(n160), .S(n233), .Z(
        \Reg_Bank/n3108 ) );
  MUX U1188 ( .A(\Reg_Bank/registers[3][13] ), .B(n161), .S(n233), .Z(
        \Reg_Bank/n3107 ) );
  MUX U1189 ( .A(\Reg_Bank/registers[3][12] ), .B(n162), .S(n233), .Z(
        \Reg_Bank/n3106 ) );
  MUX U1190 ( .A(\Reg_Bank/registers[3][11] ), .B(n163), .S(n233), .Z(
        \Reg_Bank/n3105 ) );
  MUX U1191 ( .A(\Reg_Bank/registers[3][10] ), .B(n164), .S(n233), .Z(
        \Reg_Bank/n3104 ) );
  MUX U1192 ( .A(\Reg_Bank/registers[3][9] ), .B(n165), .S(n233), .Z(
        \Reg_Bank/n3103 ) );
  MUX U1193 ( .A(\Reg_Bank/registers[3][8] ), .B(n166), .S(n233), .Z(
        \Reg_Bank/n3102 ) );
  MUX U1194 ( .A(\Reg_Bank/registers[3][7] ), .B(n167), .S(n233), .Z(
        \Reg_Bank/n3101 ) );
  MUX U1195 ( .A(\Reg_Bank/registers[3][6] ), .B(n168), .S(n233), .Z(
        \Reg_Bank/n3100 ) );
  MUX U1196 ( .A(\Reg_Bank/registers[3][5] ), .B(n169), .S(n233), .Z(
        \Reg_Bank/n3099 ) );
  MUX U1197 ( .A(\Reg_Bank/registers[3][4] ), .B(n170), .S(n233), .Z(
        \Reg_Bank/n3098 ) );
  MUX U1198 ( .A(\Reg_Bank/registers[3][3] ), .B(n171), .S(n233), .Z(
        \Reg_Bank/n3097 ) );
  MUX U1199 ( .A(\Reg_Bank/registers[3][2] ), .B(n172), .S(n233), .Z(
        \Reg_Bank/n3096 ) );
  MUX U1200 ( .A(\Reg_Bank/registers[3][1] ), .B(n174), .S(n233), .Z(
        \Reg_Bank/n3095 ) );
  MUX U1201 ( .A(\Reg_Bank/registers[3][0] ), .B(n175), .S(n233), .Z(
        \Reg_Bank/n3094 ) );
  AND U1202 ( .A(n224), .B(n188), .Z(n233) );
  IV U1203 ( .A(n215), .Z(n188) );
  NANDN U1204 ( .A(n221), .B(n225), .Z(n215) );
  AND U1205 ( .A(n232), .B(n231), .Z(n225) );
  MUX U1206 ( .A(\Reg_Bank/registers[2][31] ), .B(n142), .S(n234), .Z(
        \Reg_Bank/n3093 ) );
  MUX U1207 ( .A(\Reg_Bank/registers[2][30] ), .B(n144), .S(n234), .Z(
        \Reg_Bank/n3092 ) );
  MUX U1208 ( .A(\Reg_Bank/registers[2][29] ), .B(n145), .S(n234), .Z(
        \Reg_Bank/n3091 ) );
  MUX U1209 ( .A(\Reg_Bank/registers[2][28] ), .B(n146), .S(n234), .Z(
        \Reg_Bank/n3090 ) );
  MUX U1210 ( .A(\Reg_Bank/registers[2][27] ), .B(n147), .S(n234), .Z(
        \Reg_Bank/n3089 ) );
  MUX U1211 ( .A(\Reg_Bank/registers[2][26] ), .B(n148), .S(n234), .Z(
        \Reg_Bank/n3088 ) );
  MUX U1212 ( .A(\Reg_Bank/registers[2][25] ), .B(n149), .S(n234), .Z(
        \Reg_Bank/n3087 ) );
  MUX U1213 ( .A(\Reg_Bank/registers[2][24] ), .B(n150), .S(n234), .Z(
        \Reg_Bank/n3086 ) );
  MUX U1214 ( .A(\Reg_Bank/registers[2][23] ), .B(n151), .S(n234), .Z(
        \Reg_Bank/n3085 ) );
  MUX U1215 ( .A(\Reg_Bank/registers[2][22] ), .B(n152), .S(n234), .Z(
        \Reg_Bank/n3084 ) );
  MUX U1216 ( .A(\Reg_Bank/registers[2][21] ), .B(n153), .S(n234), .Z(
        \Reg_Bank/n3083 ) );
  MUX U1217 ( .A(\Reg_Bank/registers[2][20] ), .B(n154), .S(n234), .Z(
        \Reg_Bank/n3082 ) );
  MUX U1218 ( .A(\Reg_Bank/registers[2][19] ), .B(n155), .S(n234), .Z(
        \Reg_Bank/n3081 ) );
  MUX U1219 ( .A(\Reg_Bank/registers[2][18] ), .B(n156), .S(n234), .Z(
        \Reg_Bank/n3080 ) );
  MUX U1220 ( .A(\Reg_Bank/registers[2][17] ), .B(n157), .S(n234), .Z(
        \Reg_Bank/n3079 ) );
  MUX U1221 ( .A(\Reg_Bank/registers[2][16] ), .B(n158), .S(n234), .Z(
        \Reg_Bank/n3078 ) );
  MUX U1222 ( .A(\Reg_Bank/registers[2][15] ), .B(n159), .S(n234), .Z(
        \Reg_Bank/n3077 ) );
  MUX U1223 ( .A(\Reg_Bank/registers[2][14] ), .B(n160), .S(n234), .Z(
        \Reg_Bank/n3076 ) );
  MUX U1224 ( .A(\Reg_Bank/registers[2][13] ), .B(n161), .S(n234), .Z(
        \Reg_Bank/n3075 ) );
  MUX U1225 ( .A(\Reg_Bank/registers[2][12] ), .B(n162), .S(n234), .Z(
        \Reg_Bank/n3074 ) );
  MUX U1226 ( .A(\Reg_Bank/registers[2][11] ), .B(n163), .S(n234), .Z(
        \Reg_Bank/n3073 ) );
  MUX U1227 ( .A(\Reg_Bank/registers[2][10] ), .B(n164), .S(n234), .Z(
        \Reg_Bank/n3072 ) );
  MUX U1228 ( .A(\Reg_Bank/registers[2][9] ), .B(n165), .S(n234), .Z(
        \Reg_Bank/n3071 ) );
  MUX U1229 ( .A(\Reg_Bank/registers[2][8] ), .B(n166), .S(n234), .Z(
        \Reg_Bank/n3070 ) );
  MUX U1230 ( .A(\Reg_Bank/registers[2][7] ), .B(n167), .S(n234), .Z(
        \Reg_Bank/n3069 ) );
  MUX U1231 ( .A(\Reg_Bank/registers[2][6] ), .B(n168), .S(n234), .Z(
        \Reg_Bank/n3068 ) );
  MUX U1232 ( .A(\Reg_Bank/registers[2][5] ), .B(n169), .S(n234), .Z(
        \Reg_Bank/n3067 ) );
  MUX U1233 ( .A(\Reg_Bank/registers[2][4] ), .B(n170), .S(n234), .Z(
        \Reg_Bank/n3066 ) );
  MUX U1234 ( .A(\Reg_Bank/registers[2][3] ), .B(n171), .S(n234), .Z(
        \Reg_Bank/n3065 ) );
  MUX U1235 ( .A(\Reg_Bank/registers[2][2] ), .B(n172), .S(n234), .Z(
        \Reg_Bank/n3064 ) );
  MUX U1236 ( .A(\Reg_Bank/registers[2][1] ), .B(n174), .S(n234), .Z(
        \Reg_Bank/n3063 ) );
  MUX U1237 ( .A(\Reg_Bank/registers[2][0] ), .B(n175), .S(n234), .Z(
        \Reg_Bank/n3062 ) );
  AND U1238 ( .A(n224), .B(n190), .Z(n234) );
  IV U1239 ( .A(n217), .Z(n190) );
  NANDN U1240 ( .A(n221), .B(n227), .Z(n217) );
  AND U1241 ( .A(n232), .B(n235), .Z(n227) );
  MUX U1242 ( .A(\Reg_Bank/registers[1][31] ), .B(n142), .S(n236), .Z(
        \Reg_Bank/n3061 ) );
  NAND U1243 ( .A(n237), .B(n238), .Z(n142) );
  AND U1244 ( .A(n239), .B(n240), .Z(n238) );
  NAND U1245 ( .A(n241), .B(c_memory[31]), .Z(n240) );
  NAND U1246 ( .A(n242), .B(n243), .Z(n239) );
  AND U1247 ( .A(n244), .B(n245), .Z(n237) );
  NANDN U1248 ( .A(n246), .B(n247), .Z(n245) );
  NANDN U1249 ( .A(n248), .B(imm[15]), .Z(n244) );
  MUX U1250 ( .A(\Reg_Bank/registers[1][30] ), .B(n144), .S(n236), .Z(
        \Reg_Bank/n3060 ) );
  NAND U1251 ( .A(n249), .B(n250), .Z(n144) );
  AND U1252 ( .A(n251), .B(n252), .Z(n250) );
  NAND U1253 ( .A(n241), .B(c_memory[30]), .Z(n252) );
  NAND U1254 ( .A(n242), .B(n253), .Z(n251) );
  AND U1255 ( .A(n254), .B(n255), .Z(n249) );
  NANDN U1256 ( .A(n246), .B(pc_plus4[30]), .Z(n255) );
  NANDN U1257 ( .A(n248), .B(imm[14]), .Z(n254) );
  MUX U1258 ( .A(\Reg_Bank/registers[1][29] ), .B(n145), .S(n236), .Z(
        \Reg_Bank/n3059 ) );
  NAND U1259 ( .A(n256), .B(n257), .Z(n145) );
  AND U1260 ( .A(n258), .B(n259), .Z(n257) );
  NAND U1261 ( .A(n241), .B(c_memory[29]), .Z(n259) );
  NAND U1262 ( .A(n242), .B(n260), .Z(n258) );
  AND U1263 ( .A(n261), .B(n262), .Z(n256) );
  NANDN U1264 ( .A(n246), .B(pc_plus4[29]), .Z(n262) );
  NANDN U1265 ( .A(n248), .B(imm[13]), .Z(n261) );
  MUX U1266 ( .A(\Reg_Bank/registers[1][28] ), .B(n146), .S(n236), .Z(
        \Reg_Bank/n3058 ) );
  NAND U1267 ( .A(n263), .B(n264), .Z(n146) );
  AND U1268 ( .A(n265), .B(n266), .Z(n264) );
  NAND U1269 ( .A(n241), .B(c_memory[28]), .Z(n266) );
  NAND U1270 ( .A(n242), .B(n267), .Z(n265) );
  AND U1271 ( .A(n268), .B(n269), .Z(n263) );
  NANDN U1272 ( .A(n246), .B(pc_plus4[28]), .Z(n269) );
  NANDN U1273 ( .A(n248), .B(imm[12]), .Z(n268) );
  MUX U1274 ( .A(\Reg_Bank/registers[1][27] ), .B(n147), .S(n236), .Z(
        \Reg_Bank/n3057 ) );
  NAND U1275 ( .A(n270), .B(n271), .Z(n147) );
  AND U1276 ( .A(n272), .B(n273), .Z(n271) );
  NAND U1277 ( .A(n241), .B(c_memory[27]), .Z(n273) );
  NAND U1278 ( .A(n242), .B(n274), .Z(n272) );
  AND U1279 ( .A(n275), .B(n276), .Z(n270) );
  NANDN U1280 ( .A(n246), .B(pc_plus4[27]), .Z(n276) );
  NANDN U1281 ( .A(n248), .B(imm[11]), .Z(n275) );
  MUX U1282 ( .A(\Reg_Bank/registers[1][26] ), .B(n148), .S(n236), .Z(
        \Reg_Bank/n3056 ) );
  NAND U1283 ( .A(n277), .B(n278), .Z(n148) );
  AND U1284 ( .A(n279), .B(n280), .Z(n278) );
  NAND U1285 ( .A(n241), .B(c_memory[26]), .Z(n280) );
  NAND U1286 ( .A(n242), .B(n281), .Z(n279) );
  AND U1287 ( .A(n282), .B(n283), .Z(n277) );
  NANDN U1288 ( .A(n246), .B(pc_plus4[26]), .Z(n283) );
  NANDN U1289 ( .A(n248), .B(imm[10]), .Z(n282) );
  MUX U1290 ( .A(\Reg_Bank/registers[1][25] ), .B(n149), .S(n236), .Z(
        \Reg_Bank/n3055 ) );
  NAND U1291 ( .A(n284), .B(n285), .Z(n149) );
  AND U1292 ( .A(n286), .B(n287), .Z(n285) );
  NAND U1293 ( .A(n241), .B(c_memory[25]), .Z(n287) );
  NAND U1294 ( .A(n242), .B(n288), .Z(n286) );
  AND U1295 ( .A(n289), .B(n290), .Z(n284) );
  NANDN U1296 ( .A(n246), .B(pc_plus4[25]), .Z(n290) );
  NANDN U1297 ( .A(n248), .B(imm[9]), .Z(n289) );
  MUX U1298 ( .A(\Reg_Bank/registers[1][24] ), .B(n150), .S(n236), .Z(
        \Reg_Bank/n3054 ) );
  NAND U1299 ( .A(n291), .B(n292), .Z(n150) );
  AND U1300 ( .A(n293), .B(n294), .Z(n292) );
  NAND U1301 ( .A(n241), .B(c_memory[24]), .Z(n294) );
  NAND U1302 ( .A(n242), .B(n295), .Z(n293) );
  AND U1303 ( .A(n296), .B(n297), .Z(n291) );
  NANDN U1304 ( .A(n246), .B(pc_plus4[24]), .Z(n297) );
  NANDN U1305 ( .A(n248), .B(imm[8]), .Z(n296) );
  MUX U1306 ( .A(\Reg_Bank/registers[1][23] ), .B(n151), .S(n236), .Z(
        \Reg_Bank/n3053 ) );
  NAND U1307 ( .A(n298), .B(n299), .Z(n151) );
  AND U1308 ( .A(n300), .B(n301), .Z(n299) );
  NAND U1309 ( .A(n241), .B(c_memory[23]), .Z(n301) );
  NAND U1310 ( .A(n242), .B(n302), .Z(n300) );
  AND U1311 ( .A(n303), .B(n304), .Z(n298) );
  NANDN U1312 ( .A(n246), .B(pc_plus4[23]), .Z(n304) );
  NANDN U1313 ( .A(n248), .B(imm[7]), .Z(n303) );
  MUX U1314 ( .A(\Reg_Bank/registers[1][22] ), .B(n152), .S(n236), .Z(
        \Reg_Bank/n3052 ) );
  NAND U1315 ( .A(n305), .B(n306), .Z(n152) );
  AND U1316 ( .A(n307), .B(n308), .Z(n306) );
  NAND U1317 ( .A(n241), .B(c_memory[22]), .Z(n308) );
  NAND U1318 ( .A(n242), .B(n309), .Z(n307) );
  AND U1319 ( .A(n310), .B(n311), .Z(n305) );
  NANDN U1320 ( .A(n246), .B(pc_plus4[22]), .Z(n311) );
  NANDN U1321 ( .A(n248), .B(imm[6]), .Z(n310) );
  MUX U1322 ( .A(\Reg_Bank/registers[1][21] ), .B(n153), .S(n236), .Z(
        \Reg_Bank/n3051 ) );
  NAND U1323 ( .A(n312), .B(n313), .Z(n153) );
  AND U1324 ( .A(n314), .B(n315), .Z(n313) );
  NAND U1325 ( .A(n241), .B(c_memory[21]), .Z(n315) );
  NAND U1326 ( .A(n242), .B(n316), .Z(n314) );
  AND U1327 ( .A(n317), .B(n318), .Z(n312) );
  NANDN U1328 ( .A(n246), .B(pc_plus4[21]), .Z(n318) );
  NANDN U1329 ( .A(n248), .B(imm[5]), .Z(n317) );
  MUX U1330 ( .A(\Reg_Bank/registers[1][20] ), .B(n154), .S(n236), .Z(
        \Reg_Bank/n3050 ) );
  NAND U1331 ( .A(n319), .B(n320), .Z(n154) );
  AND U1332 ( .A(n321), .B(n322), .Z(n320) );
  NAND U1333 ( .A(n241), .B(c_memory[20]), .Z(n322) );
  NAND U1334 ( .A(n242), .B(n323), .Z(n321) );
  AND U1335 ( .A(n324), .B(n325), .Z(n319) );
  NANDN U1336 ( .A(n246), .B(pc_plus4[20]), .Z(n325) );
  NANDN U1337 ( .A(n248), .B(imm[4]), .Z(n324) );
  MUX U1338 ( .A(\Reg_Bank/registers[1][19] ), .B(n155), .S(n236), .Z(
        \Reg_Bank/n3049 ) );
  NAND U1339 ( .A(n326), .B(n327), .Z(n155) );
  AND U1340 ( .A(n328), .B(n329), .Z(n327) );
  NAND U1341 ( .A(n241), .B(c_memory[19]), .Z(n329) );
  NAND U1342 ( .A(n242), .B(n330), .Z(n328) );
  AND U1343 ( .A(n331), .B(n332), .Z(n326) );
  NANDN U1344 ( .A(n246), .B(pc_plus4[19]), .Z(n332) );
  NANDN U1345 ( .A(n248), .B(imm[3]), .Z(n331) );
  MUX U1346 ( .A(\Reg_Bank/registers[1][18] ), .B(n156), .S(n236), .Z(
        \Reg_Bank/n3048 ) );
  NAND U1347 ( .A(n333), .B(n334), .Z(n156) );
  AND U1348 ( .A(n335), .B(n336), .Z(n334) );
  NAND U1349 ( .A(n241), .B(c_memory[18]), .Z(n336) );
  NAND U1350 ( .A(n242), .B(n337), .Z(n335) );
  AND U1351 ( .A(n338), .B(n339), .Z(n333) );
  NANDN U1352 ( .A(n246), .B(pc_plus4[18]), .Z(n339) );
  NANDN U1353 ( .A(n248), .B(imm[2]), .Z(n338) );
  MUX U1354 ( .A(\Reg_Bank/registers[1][17] ), .B(n157), .S(n236), .Z(
        \Reg_Bank/n3047 ) );
  NAND U1355 ( .A(n340), .B(n341), .Z(n157) );
  AND U1356 ( .A(n342), .B(n343), .Z(n341) );
  NAND U1357 ( .A(n241), .B(c_memory[17]), .Z(n343) );
  NAND U1358 ( .A(n242), .B(n344), .Z(n342) );
  AND U1359 ( .A(n345), .B(n346), .Z(n340) );
  NANDN U1360 ( .A(n246), .B(pc_plus4[17]), .Z(n346) );
  NANDN U1361 ( .A(n248), .B(imm[1]), .Z(n345) );
  MUX U1362 ( .A(\Reg_Bank/registers[1][16] ), .B(n158), .S(n236), .Z(
        \Reg_Bank/n3046 ) );
  NAND U1363 ( .A(n347), .B(n348), .Z(n158) );
  AND U1364 ( .A(n349), .B(n350), .Z(n348) );
  NAND U1365 ( .A(n241), .B(c_memory[16]), .Z(n350) );
  NAND U1366 ( .A(n242), .B(n351), .Z(n349) );
  AND U1367 ( .A(n352), .B(n353), .Z(n347) );
  NANDN U1368 ( .A(n246), .B(pc_plus4[16]), .Z(n353) );
  NANDN U1369 ( .A(n248), .B(imm[0]), .Z(n352) );
  NAND U1370 ( .A(n242), .B(n354), .Z(n248) );
  MUX U1371 ( .A(\Reg_Bank/registers[1][15] ), .B(n159), .S(n236), .Z(
        \Reg_Bank/n3045 ) );
  NAND U1372 ( .A(n355), .B(n356), .Z(n159) );
  NANDN U1373 ( .A(n246), .B(pc_plus4[15]), .Z(n356) );
  AND U1374 ( .A(n357), .B(n358), .Z(n355) );
  NAND U1375 ( .A(n242), .B(n359), .Z(n358) );
  NAND U1376 ( .A(n241), .B(c_memory[15]), .Z(n357) );
  MUX U1377 ( .A(\Reg_Bank/registers[1][14] ), .B(n160), .S(n236), .Z(
        \Reg_Bank/n3044 ) );
  NAND U1378 ( .A(n360), .B(n361), .Z(n160) );
  NANDN U1379 ( .A(n246), .B(pc_plus4[14]), .Z(n361) );
  AND U1380 ( .A(n362), .B(n363), .Z(n360) );
  NAND U1381 ( .A(n242), .B(n364), .Z(n363) );
  NAND U1382 ( .A(n241), .B(c_memory[14]), .Z(n362) );
  MUX U1383 ( .A(\Reg_Bank/registers[1][13] ), .B(n161), .S(n236), .Z(
        \Reg_Bank/n3043 ) );
  NAND U1384 ( .A(n365), .B(n366), .Z(n161) );
  NANDN U1385 ( .A(n246), .B(pc_plus4[13]), .Z(n366) );
  AND U1386 ( .A(n367), .B(n368), .Z(n365) );
  NAND U1387 ( .A(n242), .B(n369), .Z(n368) );
  NAND U1388 ( .A(n241), .B(c_memory[13]), .Z(n367) );
  MUX U1389 ( .A(\Reg_Bank/registers[1][12] ), .B(n162), .S(n236), .Z(
        \Reg_Bank/n3042 ) );
  NAND U1390 ( .A(n370), .B(n371), .Z(n162) );
  NANDN U1391 ( .A(n246), .B(pc_plus4[12]), .Z(n371) );
  AND U1392 ( .A(n372), .B(n373), .Z(n370) );
  NAND U1393 ( .A(n242), .B(n374), .Z(n373) );
  NAND U1394 ( .A(n241), .B(c_memory[12]), .Z(n372) );
  MUX U1395 ( .A(\Reg_Bank/registers[1][11] ), .B(n163), .S(n236), .Z(
        \Reg_Bank/n3041 ) );
  NAND U1396 ( .A(n375), .B(n376), .Z(n163) );
  NANDN U1397 ( .A(n246), .B(pc_plus4[11]), .Z(n376) );
  AND U1398 ( .A(n377), .B(n378), .Z(n375) );
  NAND U1399 ( .A(n242), .B(n379), .Z(n378) );
  NAND U1400 ( .A(n241), .B(c_memory[11]), .Z(n377) );
  MUX U1401 ( .A(\Reg_Bank/registers[1][10] ), .B(n164), .S(n236), .Z(
        \Reg_Bank/n3040 ) );
  NAND U1402 ( .A(n380), .B(n381), .Z(n164) );
  NANDN U1403 ( .A(n246), .B(pc_plus4[10]), .Z(n381) );
  AND U1404 ( .A(n382), .B(n383), .Z(n380) );
  NAND U1405 ( .A(n242), .B(n384), .Z(n383) );
  NAND U1406 ( .A(n241), .B(c_memory[10]), .Z(n382) );
  MUX U1407 ( .A(\Reg_Bank/registers[1][9] ), .B(n165), .S(n236), .Z(
        \Reg_Bank/n3039 ) );
  NAND U1408 ( .A(n385), .B(n386), .Z(n165) );
  NANDN U1409 ( .A(n246), .B(pc_plus4[9]), .Z(n386) );
  AND U1410 ( .A(n387), .B(n388), .Z(n385) );
  NAND U1411 ( .A(n242), .B(n389), .Z(n388) );
  NAND U1412 ( .A(n241), .B(c_memory[9]), .Z(n387) );
  MUX U1413 ( .A(\Reg_Bank/registers[1][8] ), .B(n166), .S(n236), .Z(
        \Reg_Bank/n3038 ) );
  NAND U1414 ( .A(n390), .B(n391), .Z(n166) );
  NANDN U1415 ( .A(n246), .B(pc_plus4[8]), .Z(n391) );
  AND U1416 ( .A(n392), .B(n393), .Z(n390) );
  NAND U1417 ( .A(n242), .B(n394), .Z(n393) );
  NAND U1418 ( .A(n241), .B(c_memory[8]), .Z(n392) );
  MUX U1419 ( .A(\Reg_Bank/registers[1][7] ), .B(n167), .S(n236), .Z(
        \Reg_Bank/n3037 ) );
  NAND U1420 ( .A(n395), .B(n396), .Z(n167) );
  NANDN U1421 ( .A(n246), .B(pc_plus4[7]), .Z(n396) );
  AND U1422 ( .A(n397), .B(n398), .Z(n395) );
  NAND U1423 ( .A(n242), .B(N24), .Z(n398) );
  NAND U1424 ( .A(n241), .B(c_memory[7]), .Z(n397) );
  MUX U1425 ( .A(\Reg_Bank/registers[1][6] ), .B(n168), .S(n236), .Z(
        \Reg_Bank/n3036 ) );
  NAND U1426 ( .A(n399), .B(n400), .Z(n168) );
  NANDN U1427 ( .A(n246), .B(pc_plus4[6]), .Z(n400) );
  AND U1428 ( .A(n401), .B(n402), .Z(n399) );
  NAND U1429 ( .A(n242), .B(N25), .Z(n402) );
  NAND U1430 ( .A(n241), .B(c_memory[6]), .Z(n401) );
  MUX U1431 ( .A(\Reg_Bank/registers[1][5] ), .B(n169), .S(n236), .Z(
        \Reg_Bank/n3035 ) );
  NAND U1432 ( .A(n403), .B(n404), .Z(n169) );
  NANDN U1433 ( .A(n246), .B(pc_plus4[5]), .Z(n404) );
  AND U1434 ( .A(n405), .B(n406), .Z(n403) );
  NAND U1435 ( .A(n242), .B(N26), .Z(n406) );
  NAND U1436 ( .A(n241), .B(c_memory[5]), .Z(n405) );
  MUX U1437 ( .A(\Reg_Bank/registers[1][4] ), .B(n170), .S(n236), .Z(
        \Reg_Bank/n3034 ) );
  NAND U1438 ( .A(n407), .B(n408), .Z(n170) );
  NANDN U1439 ( .A(n246), .B(pc_plus4[4]), .Z(n408) );
  AND U1440 ( .A(n409), .B(n410), .Z(n407) );
  NAND U1441 ( .A(n242), .B(N27), .Z(n410) );
  NAND U1442 ( .A(n241), .B(c_memory[4]), .Z(n409) );
  MUX U1443 ( .A(\Reg_Bank/registers[1][3] ), .B(n171), .S(n236), .Z(
        \Reg_Bank/n3033 ) );
  NAND U1444 ( .A(n411), .B(n412), .Z(n171) );
  NANDN U1445 ( .A(n246), .B(pc_plus4[3]), .Z(n412) );
  AND U1446 ( .A(n413), .B(n414), .Z(n411) );
  NAND U1447 ( .A(n242), .B(N28), .Z(n414) );
  NAND U1448 ( .A(n241), .B(c_memory[3]), .Z(n413) );
  MUX U1449 ( .A(\Reg_Bank/registers[1][2] ), .B(n172), .S(n236), .Z(
        \Reg_Bank/n3032 ) );
  NAND U1450 ( .A(n415), .B(n416), .Z(n172) );
  OR U1451 ( .A(n246), .B(pc_current[2]), .Z(n416) );
  NAND U1452 ( .A(n417), .B(n354), .Z(n246) );
  NAND U1453 ( .A(n418), .B(n127), .Z(n354) );
  NAND U1454 ( .A(n419), .B(n7), .Z(n418) );
  NAND U1455 ( .A(n420), .B(n421), .Z(n419) );
  IV U1456 ( .A(n108), .Z(n420) );
  AND U1457 ( .A(n422), .B(n423), .Z(n415) );
  NAND U1458 ( .A(n242), .B(N29), .Z(n423) );
  NAND U1459 ( .A(n241), .B(c_memory[2]), .Z(n422) );
  MUX U1460 ( .A(\Reg_Bank/registers[1][1] ), .B(n174), .S(n236), .Z(
        \Reg_Bank/n3031 ) );
  NAND U1461 ( .A(n424), .B(n425), .Z(n174) );
  NAND U1462 ( .A(n241), .B(c_memory[1]), .Z(n425) );
  NANDN U1463 ( .A(n426), .B(n242), .Z(n424) );
  MUX U1464 ( .A(\Reg_Bank/registers[1][0] ), .B(n175), .S(n236), .Z(
        \Reg_Bank/n3030 ) );
  AND U1465 ( .A(n224), .B(n192), .Z(n236) );
  IV U1466 ( .A(n219), .Z(n192) );
  NANDN U1467 ( .A(n221), .B(n229), .Z(n219) );
  NOR U1468 ( .A(n235), .B(n232), .Z(n229) );
  NAND U1469 ( .A(n427), .B(n428), .Z(n232) );
  AND U1470 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U1471 ( .A(n431), .B(opcode[17]), .Z(n430) );
  NAND U1472 ( .A(n432), .B(n7), .Z(n429) );
  NAND U1473 ( .A(n421), .B(n433), .Z(n432) );
  NAND U1474 ( .A(n10), .B(n434), .Z(n433) );
  NAND U1475 ( .A(n435), .B(n436), .Z(n434) );
  AND U1476 ( .A(n437), .B(n438), .Z(n436) );
  NAND U1477 ( .A(n439), .B(n440), .Z(n438) );
  AND U1478 ( .A(n441), .B(imm[12]), .Z(n439) );
  AND U1479 ( .A(n442), .B(n443), .Z(n437) );
  NANDN U1480 ( .A(n444), .B(imm[12]), .Z(n443) );
  NANDN U1481 ( .A(n445), .B(imm[12]), .Z(n442) );
  AND U1482 ( .A(n446), .B(n447), .Z(n435) );
  NAND U1483 ( .A(n448), .B(n449), .Z(n447) );
  AND U1484 ( .A(n450), .B(imm[12]), .Z(n449) );
  NAND U1485 ( .A(n108), .B(n451), .Z(n446) );
  NANDN U1486 ( .A(n110), .B(n452), .Z(n451) );
  NANDN U1487 ( .A(n453), .B(imm[12]), .Z(n452) );
  AND U1488 ( .A(n454), .B(n455), .Z(n427) );
  NAND U1489 ( .A(n98), .B(n456), .Z(n455) );
  MUX U1490 ( .A(imm[12]), .B(opcode[17]), .S(n100), .Z(n456) );
  NAND U1491 ( .A(n457), .B(n241), .Z(n454) );
  AND U1492 ( .A(n458), .B(opcode[17]), .Z(n457) );
  IV U1493 ( .A(n231), .Z(n235) );
  NAND U1494 ( .A(n459), .B(n460), .Z(n231) );
  AND U1495 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U1496 ( .A(n431), .B(opcode[16]), .Z(n462) );
  NAND U1497 ( .A(n463), .B(n7), .Z(n461) );
  NAND U1498 ( .A(n464), .B(n465), .Z(n463) );
  AND U1499 ( .A(n466), .B(n130), .Z(n464) );
  NAND U1500 ( .A(n10), .B(n467), .Z(n466) );
  NAND U1501 ( .A(n468), .B(n469), .Z(n467) );
  AND U1502 ( .A(n470), .B(n471), .Z(n469) );
  NAND U1503 ( .A(n472), .B(n440), .Z(n471) );
  AND U1504 ( .A(n441), .B(imm[11]), .Z(n472) );
  AND U1505 ( .A(n473), .B(n474), .Z(n470) );
  NANDN U1506 ( .A(n444), .B(imm[11]), .Z(n474) );
  NANDN U1507 ( .A(n445), .B(imm[11]), .Z(n473) );
  AND U1508 ( .A(n475), .B(n476), .Z(n468) );
  NAND U1509 ( .A(n448), .B(n477), .Z(n476) );
  AND U1510 ( .A(n450), .B(imm[11]), .Z(n477) );
  NANDN U1511 ( .A(n453), .B(n478), .Z(n475) );
  AND U1512 ( .A(imm[11]), .B(n108), .Z(n478) );
  AND U1513 ( .A(n479), .B(n480), .Z(n459) );
  NAND U1514 ( .A(n98), .B(n481), .Z(n480) );
  MUX U1515 ( .A(imm[11]), .B(opcode[16]), .S(n100), .Z(n481) );
  NAND U1516 ( .A(n482), .B(n241), .Z(n479) );
  AND U1517 ( .A(n458), .B(opcode[16]), .Z(n482) );
  NAND U1518 ( .A(n483), .B(n484), .Z(n221) );
  AND U1519 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U1520 ( .A(n431), .B(opcode[18]), .Z(n486) );
  NAND U1521 ( .A(n487), .B(n7), .Z(n485) );
  NAND U1522 ( .A(n421), .B(n488), .Z(n487) );
  NAND U1523 ( .A(n10), .B(n489), .Z(n488) );
  NAND U1524 ( .A(n490), .B(n491), .Z(n489) );
  AND U1525 ( .A(n492), .B(n493), .Z(n491) );
  NAND U1526 ( .A(n494), .B(n440), .Z(n493) );
  AND U1527 ( .A(imm[13]), .B(n441), .Z(n494) );
  AND U1528 ( .A(n495), .B(n496), .Z(n492) );
  NANDN U1529 ( .A(n444), .B(imm[13]), .Z(n496) );
  NANDN U1530 ( .A(n445), .B(imm[13]), .Z(n495) );
  AND U1531 ( .A(n497), .B(n498), .Z(n490) );
  NAND U1532 ( .A(n448), .B(n499), .Z(n498) );
  AND U1533 ( .A(imm[13]), .B(n450), .Z(n499) );
  NAND U1534 ( .A(n108), .B(n500), .Z(n497) );
  NANDN U1535 ( .A(n110), .B(n501), .Z(n500) );
  NANDN U1536 ( .A(n453), .B(imm[13]), .Z(n501) );
  AND U1537 ( .A(n502), .B(n503), .Z(n483) );
  NAND U1538 ( .A(n98), .B(n504), .Z(n503) );
  MUX U1539 ( .A(imm[13]), .B(opcode[18]), .S(n100), .Z(n504) );
  NAND U1540 ( .A(n505), .B(n241), .Z(n502) );
  AND U1541 ( .A(n458), .B(opcode[18]), .Z(n505) );
  NOR U1542 ( .A(n207), .B(n195), .Z(n224) );
  NAND U1543 ( .A(n506), .B(n507), .Z(n195) );
  AND U1544 ( .A(n508), .B(n509), .Z(n507) );
  NANDN U1545 ( .A(n431), .B(opcode[20]), .Z(n509) );
  NAND U1546 ( .A(n510), .B(n7), .Z(n508) );
  NAND U1547 ( .A(n421), .B(n511), .Z(n510) );
  NAND U1548 ( .A(n10), .B(n512), .Z(n511) );
  NAND U1549 ( .A(n513), .B(n514), .Z(n512) );
  AND U1550 ( .A(n515), .B(n516), .Z(n514) );
  NAND U1551 ( .A(n517), .B(n440), .Z(n516) );
  AND U1552 ( .A(n441), .B(imm[15]), .Z(n517) );
  AND U1553 ( .A(n518), .B(n519), .Z(n515) );
  NANDN U1554 ( .A(n444), .B(imm[15]), .Z(n519) );
  NANDN U1555 ( .A(n445), .B(imm[15]), .Z(n518) );
  AND U1556 ( .A(n520), .B(n521), .Z(n513) );
  NAND U1557 ( .A(n448), .B(n522), .Z(n521) );
  AND U1558 ( .A(n450), .B(imm[15]), .Z(n522) );
  NANDN U1559 ( .A(n453), .B(n523), .Z(n520) );
  AND U1560 ( .A(imm[15]), .B(n108), .Z(n523) );
  AND U1561 ( .A(n524), .B(n525), .Z(n506) );
  NAND U1562 ( .A(n98), .B(n526), .Z(n525) );
  MUX U1563 ( .A(imm[15]), .B(opcode[20]), .S(n100), .Z(n526) );
  NAND U1564 ( .A(n527), .B(n241), .Z(n524) );
  AND U1565 ( .A(n458), .B(opcode[20]), .Z(n527) );
  NAND U1566 ( .A(n528), .B(n529), .Z(n207) );
  AND U1567 ( .A(n530), .B(n531), .Z(n529) );
  NANDN U1568 ( .A(n431), .B(opcode[19]), .Z(n531) );
  NAND U1569 ( .A(n532), .B(n7), .Z(n530) );
  NAND U1570 ( .A(n421), .B(n533), .Z(n532) );
  NAND U1571 ( .A(n10), .B(n534), .Z(n533) );
  NAND U1572 ( .A(n535), .B(n536), .Z(n534) );
  AND U1573 ( .A(n537), .B(n538), .Z(n536) );
  NAND U1574 ( .A(n539), .B(n440), .Z(n538) );
  NOR U1575 ( .A(imm[3]), .B(imm[5]), .Z(n440) );
  AND U1576 ( .A(n441), .B(imm[14]), .Z(n539) );
  NANDN U1577 ( .A(n540), .B(n541), .Z(n441) );
  NANDN U1578 ( .A(n542), .B(n543), .Z(n541) );
  AND U1579 ( .A(n544), .B(n545), .Z(n537) );
  NANDN U1580 ( .A(n444), .B(imm[14]), .Z(n545) );
  NANDN U1581 ( .A(n445), .B(imm[14]), .Z(n544) );
  NAND U1582 ( .A(n546), .B(n547), .Z(n445) );
  NANDN U1583 ( .A(n548), .B(n549), .Z(n546) );
  AND U1584 ( .A(n550), .B(n551), .Z(n535) );
  NAND U1585 ( .A(n448), .B(n552), .Z(n551) );
  AND U1586 ( .A(n450), .B(imm[14]), .Z(n552) );
  OR U1587 ( .A(n553), .B(n540), .Z(n450) );
  NAND U1588 ( .A(n108), .B(n554), .Z(n550) );
  NANDN U1589 ( .A(n110), .B(n555), .Z(n554) );
  NANDN U1590 ( .A(n453), .B(imm[14]), .Z(n555) );
  NANDN U1591 ( .A(n542), .B(imm[0]), .Z(n453) );
  AND U1592 ( .A(n465), .B(n130), .Z(n421) );
  NAND U1593 ( .A(n556), .B(n557), .Z(n465) );
  AND U1594 ( .A(n21), .B(opcode[20]), .Z(n556) );
  AND U1595 ( .A(n558), .B(n559), .Z(n528) );
  NAND U1596 ( .A(n98), .B(n560), .Z(n559) );
  MUX U1597 ( .A(imm[14]), .B(opcode[19]), .S(n100), .Z(n560) );
  IV U1598 ( .A(opcode[23]), .Z(n100) );
  ANDN U1599 ( .B(n10), .A(n561), .Z(n98) );
  NAND U1600 ( .A(n24), .B(n120), .Z(n561) );
  ANDN U1601 ( .B(n122), .A(n121), .Z(n120) );
  NAND U1602 ( .A(n562), .B(n241), .Z(n558) );
  AND U1603 ( .A(n458), .B(opcode[19]), .Z(n562) );
  NAND U1604 ( .A(n563), .B(n564), .Z(n175) );
  NAND U1605 ( .A(n241), .B(c_memory[0]), .Z(n564) );
  NAND U1606 ( .A(n242), .B(n565), .Z(n563) );
  IV U1607 ( .A(n417), .Z(n242) );
  AND U1608 ( .A(n566), .B(n567), .Z(n417) );
  NAND U1609 ( .A(n568), .B(n7), .Z(n566) );
  AND U1610 ( .A(n14), .B(n10), .Z(n568) );
  NANDN U1611 ( .A(n569), .B(n570), .Z(n14) );
  AND U1612 ( .A(n571), .B(n572), .Z(n570) );
  NAND U1613 ( .A(n573), .B(n574), .Z(\PC_Next/pc_future[9] ) );
  AND U1614 ( .A(n575), .B(n576), .Z(n574) );
  NANDN U1615 ( .A(n577), .B(pc_plus4[9]), .Z(n576) );
  NANDN U1616 ( .A(n578), .B(imm[7]), .Z(n575) );
  AND U1617 ( .A(n579), .B(n580), .Z(n573) );
  NAND U1618 ( .A(n581), .B(n582), .Z(n580) );
  MUX U1619 ( .A(pc_plus4[9]), .B(\PC_Next/N23 ), .S(n583), .Z(n581) );
  NAND U1620 ( .A(n584), .B(n389), .Z(n579) );
  NAND U1621 ( .A(n585), .B(n586), .Z(\PC_Next/pc_future[8] ) );
  AND U1622 ( .A(n587), .B(n588), .Z(n586) );
  NANDN U1623 ( .A(n577), .B(pc_plus4[8]), .Z(n588) );
  NANDN U1624 ( .A(n578), .B(imm[6]), .Z(n587) );
  AND U1625 ( .A(n589), .B(n590), .Z(n585) );
  NAND U1626 ( .A(n591), .B(n582), .Z(n590) );
  MUX U1627 ( .A(pc_plus4[8]), .B(\PC_Next/N22 ), .S(n583), .Z(n591) );
  NAND U1628 ( .A(n394), .B(n584), .Z(n589) );
  NAND U1629 ( .A(n592), .B(n593), .Z(\PC_Next/pc_future[7] ) );
  AND U1630 ( .A(n594), .B(n595), .Z(n593) );
  NANDN U1631 ( .A(n577), .B(pc_plus4[7]), .Z(n595) );
  NANDN U1632 ( .A(n578), .B(imm[5]), .Z(n594) );
  AND U1633 ( .A(n596), .B(n597), .Z(n592) );
  NAND U1634 ( .A(n598), .B(n582), .Z(n597) );
  MUX U1635 ( .A(pc_plus4[7]), .B(\PC_Next/N21 ), .S(n583), .Z(n598) );
  NAND U1636 ( .A(N24), .B(n584), .Z(n596) );
  NAND U1637 ( .A(n599), .B(n600), .Z(\PC_Next/pc_future[6] ) );
  AND U1638 ( .A(n601), .B(n602), .Z(n600) );
  NANDN U1639 ( .A(n577), .B(pc_plus4[6]), .Z(n602) );
  NANDN U1640 ( .A(n578), .B(imm[4]), .Z(n601) );
  AND U1641 ( .A(n603), .B(n604), .Z(n599) );
  NAND U1642 ( .A(n605), .B(n582), .Z(n604) );
  MUX U1643 ( .A(pc_plus4[6]), .B(\PC_Next/N20 ), .S(n583), .Z(n605) );
  NAND U1644 ( .A(N25), .B(n584), .Z(n603) );
  NAND U1645 ( .A(n606), .B(n607), .Z(\PC_Next/pc_future[5] ) );
  AND U1646 ( .A(n608), .B(n609), .Z(n607) );
  NANDN U1647 ( .A(n577), .B(pc_plus4[5]), .Z(n609) );
  NANDN U1648 ( .A(n578), .B(imm[3]), .Z(n608) );
  AND U1649 ( .A(n610), .B(n611), .Z(n606) );
  NAND U1650 ( .A(n612), .B(n582), .Z(n611) );
  MUX U1651 ( .A(pc_plus4[5]), .B(\PC_Next/N19 ), .S(n583), .Z(n612) );
  NAND U1652 ( .A(N26), .B(n584), .Z(n610) );
  NAND U1653 ( .A(n613), .B(n614), .Z(\PC_Next/pc_future[4] ) );
  AND U1654 ( .A(n615), .B(n616), .Z(n614) );
  NANDN U1655 ( .A(n577), .B(pc_plus4[4]), .Z(n616) );
  NANDN U1656 ( .A(n578), .B(imm[2]), .Z(n615) );
  AND U1657 ( .A(n617), .B(n618), .Z(n613) );
  NAND U1658 ( .A(n619), .B(n582), .Z(n618) );
  MUX U1659 ( .A(pc_plus4[4]), .B(\PC_Next/N18 ), .S(n583), .Z(n619) );
  NAND U1660 ( .A(N27), .B(n584), .Z(n617) );
  NAND U1661 ( .A(n620), .B(n621), .Z(\PC_Next/pc_future[3] ) );
  AND U1662 ( .A(n622), .B(n623), .Z(n621) );
  NANDN U1663 ( .A(n577), .B(pc_plus4[3]), .Z(n623) );
  NANDN U1664 ( .A(n578), .B(imm[1]), .Z(n622) );
  AND U1665 ( .A(n624), .B(n625), .Z(n620) );
  NAND U1666 ( .A(n626), .B(n582), .Z(n625) );
  MUX U1667 ( .A(pc_plus4[3]), .B(\PC_Next/N17 ), .S(n583), .Z(n626) );
  NAND U1668 ( .A(N28), .B(n584), .Z(n624) );
  NAND U1669 ( .A(n627), .B(n628), .Z(\PC_Next/pc_future[2] ) );
  AND U1670 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U1671 ( .A(n577), .B(n631), .Z(n630) );
  NANDN U1672 ( .A(n578), .B(imm[0]), .Z(n629) );
  AND U1673 ( .A(n632), .B(n633), .Z(n627) );
  NAND U1674 ( .A(n634), .B(n582), .Z(n633) );
  MUX U1675 ( .A(n631), .B(\PC_Next/N16 ), .S(n583), .Z(n634) );
  IV U1676 ( .A(pc_current[2]), .Z(n631) );
  NAND U1677 ( .A(N29), .B(n584), .Z(n632) );
  NAND U1678 ( .A(n635), .B(n636), .Z(\PC_Next/pc_future[27] ) );
  AND U1679 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U1680 ( .A(n577), .B(pc_plus4[27]), .Z(n638) );
  NANDN U1681 ( .A(n578), .B(opcode[25]), .Z(n637) );
  AND U1682 ( .A(n639), .B(n640), .Z(n635) );
  NAND U1683 ( .A(n641), .B(n582), .Z(n640) );
  MUX U1684 ( .A(pc_plus4[27]), .B(\PC_Next/N41 ), .S(n583), .Z(n641) );
  NAND U1685 ( .A(n274), .B(n584), .Z(n639) );
  NAND U1686 ( .A(n642), .B(n643), .Z(\PC_Next/pc_future[26] ) );
  AND U1687 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U1688 ( .A(n577), .B(pc_plus4[26]), .Z(n645) );
  NANDN U1689 ( .A(n578), .B(opcode[24]), .Z(n644) );
  AND U1690 ( .A(n646), .B(n647), .Z(n642) );
  NAND U1691 ( .A(n648), .B(n582), .Z(n647) );
  MUX U1692 ( .A(pc_plus4[26]), .B(\PC_Next/N40 ), .S(n583), .Z(n648) );
  NAND U1693 ( .A(n281), .B(n584), .Z(n646) );
  NAND U1694 ( .A(n649), .B(n650), .Z(\PC_Next/pc_future[25] ) );
  AND U1695 ( .A(n651), .B(n652), .Z(n650) );
  NANDN U1696 ( .A(n577), .B(pc_plus4[25]), .Z(n652) );
  NANDN U1697 ( .A(n578), .B(opcode[23]), .Z(n651) );
  AND U1698 ( .A(n653), .B(n654), .Z(n649) );
  NAND U1699 ( .A(n655), .B(n582), .Z(n654) );
  MUX U1700 ( .A(pc_plus4[25]), .B(\PC_Next/N39 ), .S(n583), .Z(n655) );
  NAND U1701 ( .A(n288), .B(n584), .Z(n653) );
  NAND U1702 ( .A(n656), .B(n657), .Z(\PC_Next/pc_future[24] ) );
  AND U1703 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U1704 ( .A(n577), .B(pc_plus4[24]), .Z(n659) );
  NANDN U1705 ( .A(n578), .B(opcode[22]), .Z(n658) );
  AND U1706 ( .A(n660), .B(n661), .Z(n656) );
  NAND U1707 ( .A(n662), .B(n582), .Z(n661) );
  MUX U1708 ( .A(pc_plus4[24]), .B(\PC_Next/N38 ), .S(n583), .Z(n662) );
  NAND U1709 ( .A(n295), .B(n584), .Z(n660) );
  NAND U1710 ( .A(n663), .B(n664), .Z(\PC_Next/pc_future[23] ) );
  AND U1711 ( .A(n665), .B(n666), .Z(n664) );
  NANDN U1712 ( .A(n577), .B(pc_plus4[23]), .Z(n666) );
  NANDN U1713 ( .A(n578), .B(opcode[21]), .Z(n665) );
  AND U1714 ( .A(n667), .B(n668), .Z(n663) );
  NAND U1715 ( .A(n669), .B(n582), .Z(n668) );
  MUX U1716 ( .A(pc_plus4[23]), .B(\PC_Next/N37 ), .S(n583), .Z(n669) );
  NAND U1717 ( .A(n302), .B(n584), .Z(n667) );
  NAND U1718 ( .A(n670), .B(n671), .Z(\PC_Next/pc_future[22] ) );
  AND U1719 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U1720 ( .A(n577), .B(pc_plus4[22]), .Z(n673) );
  NANDN U1721 ( .A(n578), .B(opcode[20]), .Z(n672) );
  AND U1722 ( .A(n674), .B(n675), .Z(n670) );
  NAND U1723 ( .A(n676), .B(n582), .Z(n675) );
  MUX U1724 ( .A(pc_plus4[22]), .B(\PC_Next/N36 ), .S(n583), .Z(n676) );
  NAND U1725 ( .A(n309), .B(n584), .Z(n674) );
  NAND U1726 ( .A(n677), .B(n678), .Z(\PC_Next/pc_future[21] ) );
  AND U1727 ( .A(n679), .B(n680), .Z(n678) );
  NANDN U1728 ( .A(n577), .B(pc_plus4[21]), .Z(n680) );
  NANDN U1729 ( .A(n578), .B(opcode[19]), .Z(n679) );
  AND U1730 ( .A(n681), .B(n682), .Z(n677) );
  NAND U1731 ( .A(n683), .B(n582), .Z(n682) );
  MUX U1732 ( .A(pc_plus4[21]), .B(\PC_Next/N35 ), .S(n583), .Z(n683) );
  NAND U1733 ( .A(n316), .B(n584), .Z(n681) );
  NAND U1734 ( .A(n684), .B(n685), .Z(\PC_Next/pc_future[20] ) );
  AND U1735 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U1736 ( .A(n577), .B(pc_plus4[20]), .Z(n687) );
  NANDN U1737 ( .A(n578), .B(opcode[18]), .Z(n686) );
  AND U1738 ( .A(n688), .B(n689), .Z(n684) );
  NAND U1739 ( .A(n690), .B(n582), .Z(n689) );
  MUX U1740 ( .A(pc_plus4[20]), .B(\PC_Next/N34 ), .S(n583), .Z(n690) );
  NAND U1741 ( .A(n323), .B(n584), .Z(n688) );
  NAND U1742 ( .A(n691), .B(n692), .Z(\PC_Next/pc_future[19] ) );
  AND U1743 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U1744 ( .A(n577), .B(pc_plus4[19]), .Z(n694) );
  NANDN U1745 ( .A(n578), .B(opcode[17]), .Z(n693) );
  AND U1746 ( .A(n695), .B(n696), .Z(n691) );
  NAND U1747 ( .A(n697), .B(n582), .Z(n696) );
  MUX U1748 ( .A(pc_plus4[19]), .B(\PC_Next/N33 ), .S(n583), .Z(n697) );
  NAND U1749 ( .A(n330), .B(n584), .Z(n695) );
  NAND U1750 ( .A(n698), .B(n699), .Z(\PC_Next/pc_future[18] ) );
  AND U1751 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U1752 ( .A(n577), .B(pc_plus4[18]), .Z(n701) );
  NANDN U1753 ( .A(n578), .B(opcode[16]), .Z(n700) );
  AND U1754 ( .A(n702), .B(n703), .Z(n698) );
  NAND U1755 ( .A(n704), .B(n582), .Z(n703) );
  MUX U1756 ( .A(pc_plus4[18]), .B(\PC_Next/N32 ), .S(n583), .Z(n704) );
  NAND U1757 ( .A(n337), .B(n584), .Z(n702) );
  NAND U1758 ( .A(n705), .B(n706), .Z(\PC_Next/pc_future[17] ) );
  AND U1759 ( .A(n707), .B(n708), .Z(n706) );
  NANDN U1760 ( .A(n577), .B(pc_plus4[17]), .Z(n708) );
  NANDN U1761 ( .A(n578), .B(imm[15]), .Z(n707) );
  AND U1762 ( .A(n709), .B(n710), .Z(n705) );
  NAND U1763 ( .A(n711), .B(n582), .Z(n710) );
  MUX U1764 ( .A(pc_plus4[17]), .B(\PC_Next/N31 ), .S(n583), .Z(n711) );
  NAND U1765 ( .A(n344), .B(n584), .Z(n709) );
  NAND U1766 ( .A(n712), .B(n713), .Z(\PC_Next/pc_future[16] ) );
  AND U1767 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U1768 ( .A(n577), .B(pc_plus4[16]), .Z(n715) );
  NANDN U1769 ( .A(n578), .B(imm[14]), .Z(n714) );
  AND U1770 ( .A(n716), .B(n717), .Z(n712) );
  NAND U1771 ( .A(n718), .B(n582), .Z(n717) );
  MUX U1772 ( .A(pc_plus4[16]), .B(\PC_Next/N30 ), .S(n583), .Z(n718) );
  NAND U1773 ( .A(n351), .B(n584), .Z(n716) );
  NAND U1774 ( .A(n719), .B(n720), .Z(\PC_Next/pc_future[15] ) );
  AND U1775 ( .A(n721), .B(n722), .Z(n720) );
  NANDN U1776 ( .A(n577), .B(pc_plus4[15]), .Z(n722) );
  NANDN U1777 ( .A(n578), .B(imm[13]), .Z(n721) );
  AND U1778 ( .A(n723), .B(n724), .Z(n719) );
  NAND U1779 ( .A(n725), .B(n582), .Z(n724) );
  MUX U1780 ( .A(pc_plus4[15]), .B(\PC_Next/N29 ), .S(n583), .Z(n725) );
  NAND U1781 ( .A(n359), .B(n584), .Z(n723) );
  NAND U1782 ( .A(n726), .B(n727), .Z(\PC_Next/pc_future[14] ) );
  AND U1783 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U1784 ( .A(n577), .B(pc_plus4[14]), .Z(n729) );
  NANDN U1785 ( .A(n578), .B(imm[12]), .Z(n728) );
  AND U1786 ( .A(n730), .B(n731), .Z(n726) );
  NAND U1787 ( .A(n732), .B(n582), .Z(n731) );
  MUX U1788 ( .A(pc_plus4[14]), .B(\PC_Next/N28 ), .S(n583), .Z(n732) );
  NAND U1789 ( .A(n364), .B(n584), .Z(n730) );
  NAND U1790 ( .A(n733), .B(n734), .Z(\PC_Next/pc_future[13] ) );
  AND U1791 ( .A(n735), .B(n736), .Z(n734) );
  NANDN U1792 ( .A(n577), .B(pc_plus4[13]), .Z(n736) );
  NANDN U1793 ( .A(n578), .B(imm[11]), .Z(n735) );
  AND U1794 ( .A(n737), .B(n738), .Z(n733) );
  NAND U1795 ( .A(n739), .B(n582), .Z(n738) );
  MUX U1796 ( .A(pc_plus4[13]), .B(\PC_Next/N27 ), .S(n583), .Z(n739) );
  NAND U1797 ( .A(n369), .B(n584), .Z(n737) );
  NAND U1798 ( .A(n740), .B(n741), .Z(\PC_Next/pc_future[12] ) );
  AND U1799 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U1800 ( .A(n577), .B(pc_plus4[12]), .Z(n743) );
  NANDN U1801 ( .A(n578), .B(imm[10]), .Z(n742) );
  AND U1802 ( .A(n744), .B(n745), .Z(n740) );
  NAND U1803 ( .A(n746), .B(n582), .Z(n745) );
  MUX U1804 ( .A(pc_plus4[12]), .B(\PC_Next/N26 ), .S(n583), .Z(n746) );
  NAND U1805 ( .A(n374), .B(n584), .Z(n744) );
  NAND U1806 ( .A(n747), .B(n748), .Z(\PC_Next/pc_future[11] ) );
  AND U1807 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U1808 ( .A(n577), .B(pc_plus4[11]), .Z(n750) );
  NANDN U1809 ( .A(n578), .B(imm[9]), .Z(n749) );
  AND U1810 ( .A(n751), .B(n752), .Z(n747) );
  NAND U1811 ( .A(n753), .B(n582), .Z(n752) );
  MUX U1812 ( .A(pc_plus4[11]), .B(\PC_Next/N25 ), .S(n583), .Z(n753) );
  NAND U1813 ( .A(n379), .B(n584), .Z(n751) );
  NAND U1814 ( .A(n754), .B(n755), .Z(\PC_Next/pc_future[10] ) );
  AND U1815 ( .A(n756), .B(n757), .Z(n755) );
  NANDN U1816 ( .A(n577), .B(pc_plus4[10]), .Z(n757) );
  NANDN U1817 ( .A(n578), .B(imm[8]), .Z(n756) );
  AND U1818 ( .A(n758), .B(n759), .Z(n754) );
  NAND U1819 ( .A(n760), .B(n582), .Z(n759) );
  MUX U1820 ( .A(pc_plus4[10]), .B(\PC_Next/N24 ), .S(n583), .Z(n760) );
  NAND U1821 ( .A(n384), .B(n584), .Z(n758) );
  NAND U1822 ( .A(n761), .B(n762), .Z(\PC_Next/n311 ) );
  AND U1823 ( .A(n763), .B(n764), .Z(n762) );
  NANDN U1824 ( .A(n578), .B(pc_current[28]), .Z(n764) );
  NANDN U1825 ( .A(n577), .B(pc_plus4[28]), .Z(n763) );
  AND U1826 ( .A(n765), .B(n766), .Z(n761) );
  NAND U1827 ( .A(n767), .B(n582), .Z(n766) );
  MUX U1828 ( .A(pc_plus4[28]), .B(\PC_Next/N42 ), .S(n583), .Z(n767) );
  IV U1829 ( .A(n768), .Z(n583) );
  NAND U1830 ( .A(n267), .B(n584), .Z(n765) );
  NAND U1831 ( .A(n769), .B(n770), .Z(\PC_Next/n310 ) );
  AND U1832 ( .A(n771), .B(n772), .Z(n770) );
  NANDN U1833 ( .A(n578), .B(pc_current[29]), .Z(n772) );
  NANDN U1834 ( .A(n577), .B(pc_plus4[29]), .Z(n771) );
  AND U1835 ( .A(n773), .B(n774), .Z(n769) );
  NAND U1836 ( .A(n775), .B(n582), .Z(n774) );
  MUX U1837 ( .A(\PC_Next/N43 ), .B(pc_plus4[29]), .S(n768), .Z(n775) );
  NAND U1838 ( .A(n260), .B(n584), .Z(n773) );
  NAND U1839 ( .A(n776), .B(n777), .Z(\PC_Next/n309 ) );
  AND U1840 ( .A(n778), .B(n779), .Z(n777) );
  NANDN U1841 ( .A(n578), .B(pc_current[30]), .Z(n779) );
  NANDN U1842 ( .A(n577), .B(pc_plus4[30]), .Z(n778) );
  AND U1843 ( .A(n780), .B(n781), .Z(n776) );
  NAND U1844 ( .A(n782), .B(n582), .Z(n781) );
  MUX U1845 ( .A(\PC_Next/N44 ), .B(pc_plus4[30]), .S(n768), .Z(n782) );
  NAND U1846 ( .A(n253), .B(n584), .Z(n780) );
  NAND U1847 ( .A(n783), .B(n784), .Z(\PC_Next/n308 ) );
  AND U1848 ( .A(n785), .B(n786), .Z(n784) );
  NANDN U1849 ( .A(n578), .B(pc_current[31]), .Z(n786) );
  NAND U1850 ( .A(n584), .B(n787), .Z(n578) );
  NANDN U1851 ( .A(n577), .B(n247), .Z(n785) );
  NANDN U1852 ( .A(n584), .B(n787), .Z(n577) );
  AND U1853 ( .A(n788), .B(n789), .Z(n783) );
  NAND U1854 ( .A(n790), .B(n582), .Z(n789) );
  NOR U1855 ( .A(n584), .B(n787), .Z(n582) );
  NAND U1856 ( .A(n791), .B(n7), .Z(n787) );
  NAND U1857 ( .A(n792), .B(n793), .Z(n791) );
  ANDN U1858 ( .B(n794), .A(n795), .Z(n792) );
  MUX U1859 ( .A(\PC_Next/N45 ), .B(n247), .S(n768), .Z(n790) );
  AND U1860 ( .A(n796), .B(n797), .Z(n768) );
  AND U1861 ( .A(n798), .B(n799), .Z(n797) );
  NANDN U1862 ( .A(n800), .B(n243), .Z(n799) );
  MUX U1863 ( .A(n801), .B(n802), .S(n803), .Z(n798) );
  NAND U1864 ( .A(n804), .B(n805), .Z(n801) );
  AND U1865 ( .A(n806), .B(n807), .Z(n796) );
  MUX U1866 ( .A(n808), .B(n802), .S(n804), .Z(n807) );
  NANDN U1867 ( .A(n809), .B(n810), .Z(n802) );
  NAND U1868 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U1869 ( .A(n800), .B(n813), .Z(n808) );
  NANDN U1870 ( .A(n811), .B(n812), .Z(n800) );
  MUX U1871 ( .A(n814), .B(n815), .S(n804), .Z(n806) );
  ANDN U1872 ( .B(n816), .A(n817), .Z(n804) );
  ANDN U1873 ( .B(n127), .A(n818), .Z(n816) );
  NANDN U1874 ( .A(n812), .B(n811), .Z(n815) );
  NAND U1875 ( .A(n803), .B(n805), .Z(n814) );
  NOR U1876 ( .A(n812), .B(n811), .Z(n805) );
  NAND U1877 ( .A(n819), .B(n820), .Z(n811) );
  AND U1878 ( .A(n127), .B(n821), .Z(n820) );
  AND U1879 ( .A(n567), .B(n822), .Z(n819) );
  NAND U1880 ( .A(n17), .B(opcode[16]), .Z(n822) );
  NOR U1881 ( .A(opcode[29]), .B(n24), .Z(n567) );
  ANDN U1882 ( .B(n823), .A(n824), .Z(n812) );
  ANDN U1883 ( .B(n825), .A(n818), .Z(n823) );
  IV U1884 ( .A(n813), .Z(n803) );
  AND U1885 ( .A(n826), .B(n827), .Z(n813) );
  AND U1886 ( .A(n828), .B(n829), .Z(n827) );
  AND U1887 ( .A(n830), .B(n831), .Z(n829) );
  AND U1888 ( .A(n832), .B(n833), .Z(n831) );
  AND U1889 ( .A(n834), .B(n835), .Z(n833) );
  AND U1890 ( .A(n836), .B(n837), .Z(n832) );
  IV U1891 ( .A(N27), .Z(n836) );
  AND U1892 ( .A(n838), .B(n839), .Z(n830) );
  AND U1893 ( .A(n840), .B(n841), .Z(n839) );
  IV U1894 ( .A(N24), .Z(n841) );
  ANDN U1895 ( .B(n426), .A(n565), .Z(n838) );
  NAND U1896 ( .A(n842), .B(n843), .Z(n565) );
  AND U1897 ( .A(n844), .B(n845), .Z(n843) );
  AND U1898 ( .A(n846), .B(n847), .Z(n845) );
  NAND U1899 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][0] ), .Z(n847) );
  ANDN U1900 ( .B(\Shifter/sll_27/ML_int[3][0] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][0] ) );
  ANDN U1901 ( .B(\Shifter/sll_27/ML_int[2][0] ), .A(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][0] ) );
  ANDN U1902 ( .B(\Shifter/sll_27/ML_int[1][0] ), .A(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][0] ) );
  ANDN U1903 ( .B(b_bus[0]), .A(a_bus[0]), .Z(\Shifter/sll_27/ML_int[1][0] )
         );
  AND U1904 ( .A(n849), .B(n850), .Z(n846) );
  NAND U1905 ( .A(n851), .B(n852), .Z(n850) );
  NAND U1906 ( .A(n853), .B(n854), .Z(n851) );
  AND U1907 ( .A(n855), .B(n856), .Z(n854) );
  AND U1908 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U1909 ( .A(n859), .B(a_bus[4]), .Z(n858) );
  AND U1910 ( .A(n860), .B(n861), .Z(n853) );
  NAND U1911 ( .A(n862), .B(n863), .Z(n861) );
  NAND U1912 ( .A(n864), .B(n865), .Z(n849) );
  NAND U1913 ( .A(n866), .B(n867), .Z(n864) );
  AND U1914 ( .A(n868), .B(n856), .Z(n867) );
  NAND U1915 ( .A(n869), .B(n870), .Z(n856) );
  AND U1916 ( .A(n857), .B(n871), .Z(n868) );
  NANDN U1917 ( .A(n872), .B(a_bus[4]), .Z(n871) );
  NAND U1918 ( .A(n873), .B(n874), .Z(n857) );
  AND U1919 ( .A(n860), .B(n875), .Z(n866) );
  NAND U1920 ( .A(n862), .B(n876), .Z(n875) );
  NAND U1921 ( .A(n877), .B(n878), .Z(n862) );
  AND U1922 ( .A(n879), .B(n880), .Z(n878) );
  NANDN U1923 ( .A(n881), .B(b_bus[0]), .Z(n880) );
  NANDN U1924 ( .A(n882), .B(b_bus[1]), .Z(n879) );
  AND U1925 ( .A(n883), .B(n884), .Z(n877) );
  NANDN U1926 ( .A(n885), .B(b_bus[3]), .Z(n884) );
  NANDN U1927 ( .A(n886), .B(b_bus[2]), .Z(n883) );
  NAND U1928 ( .A(n887), .B(n888), .Z(n860) );
  AND U1929 ( .A(n889), .B(n890), .Z(n844) );
  NANDN U1930 ( .A(n891), .B(\ALU/N108 ), .Z(n890) );
  NAND U1931 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N108 ), .Z(n889) );
  AND U1932 ( .A(n892), .B(n893), .Z(n842) );
  AND U1933 ( .A(n894), .B(n895), .Z(n893) );
  NAND U1934 ( .A(n896), .B(n897), .Z(n895) );
  AND U1935 ( .A(b_bus[0]), .B(a_bus[0]), .Z(n896) );
  AND U1936 ( .A(n898), .B(n899), .Z(n894) );
  NAND U1937 ( .A(n900), .B(n901), .Z(n899) );
  AND U1938 ( .A(n902), .B(n903), .Z(n900) );
  NAND U1939 ( .A(n904), .B(n902), .Z(n898) );
  MUX U1940 ( .A(n905), .B(n906), .S(n907), .Z(n902) );
  MUX U1941 ( .A(n904), .B(n908), .S(n909), .Z(n906) );
  MUX U1942 ( .A(n910), .B(n908), .S(n2486), .Z(n905) );
  FA U1943 ( .A(b_bus[30]), .B(n911), .CI(n912), .CO(n908) );
  NAND U1944 ( .A(n913), .B(reg_source[30]), .Z(n912) );
  IV U1945 ( .A(n914), .Z(n911) );
  FA U1946 ( .A(n915), .B(n916), .CI(n917), .CO(n914) );
  AND U1947 ( .A(n918), .B(n919), .Z(n917) );
  FA U1948 ( .A(n920), .B(n921), .CI(n2489), .CO(n916) );
  FA U1949 ( .A(n922), .B(n923), .CI(n924), .CO(n921) );
  AND U1950 ( .A(n918), .B(n925), .Z(n924) );
  FA U1951 ( .A(n926), .B(n927), .CI(n2491), .CO(n923) );
  FA U1952 ( .A(n928), .B(n929), .CI(n930), .CO(n927) );
  AND U1953 ( .A(n918), .B(n931), .Z(n930) );
  FA U1954 ( .A(n932), .B(n933), .CI(n2493), .CO(n929) );
  FA U1955 ( .A(n934), .B(n935), .CI(n936), .CO(n933) );
  AND U1956 ( .A(n918), .B(n937), .Z(n936) );
  FA U1957 ( .A(n938), .B(n939), .CI(n2495), .CO(n935) );
  FA U1958 ( .A(n940), .B(n941), .CI(n942), .CO(n939) );
  AND U1959 ( .A(n918), .B(n943), .Z(n942) );
  FA U1960 ( .A(n944), .B(n945), .CI(n2497), .CO(n941) );
  FA U1961 ( .A(n946), .B(n947), .CI(n948), .CO(n945) );
  AND U1962 ( .A(n918), .B(n949), .Z(n948) );
  FA U1963 ( .A(n950), .B(n951), .CI(n2499), .CO(n947) );
  FA U1964 ( .A(n952), .B(n953), .CI(n954), .CO(n951) );
  FA U1965 ( .A(n955), .B(n956), .CI(n2501), .CO(n953) );
  FA U1966 ( .A(n957), .B(n958), .CI(n959), .CO(n956) );
  FA U1967 ( .A(n960), .B(n961), .CI(n2503), .CO(n958) );
  FA U1968 ( .A(n962), .B(n963), .CI(n964), .CO(n961) );
  FA U1969 ( .A(n965), .B(n966), .CI(n2505), .CO(n963) );
  FA U1970 ( .A(n967), .B(n968), .CI(n969), .CO(n966) );
  AND U1971 ( .A(n970), .B(n971), .Z(n968) );
  NAND U1972 ( .A(n972), .B(n973), .Z(n971) );
  NAND U1973 ( .A(n974), .B(n2481), .Z(n973) );
  AND U1974 ( .A(n975), .B(n976), .Z(n972) );
  NAND U1975 ( .A(n977), .B(n2507), .Z(n976) );
  NAND U1976 ( .A(n978), .B(n979), .Z(n975) );
  FA U1977 ( .A(n980), .B(n981), .CI(n982), .CO(n979) );
  AND U1978 ( .A(reg_source[8]), .B(n913), .Z(n982) );
  FA U1979 ( .A(n2483), .B(n983), .CI(n984), .CO(n981) );
  FA U1980 ( .A(n985), .B(n986), .CI(n987), .CO(n983) );
  AND U1981 ( .A(reg_source[6]), .B(n913), .Z(n987) );
  FA U1982 ( .A(n2485), .B(n988), .CI(n989), .CO(n986) );
  FA U1983 ( .A(n990), .B(n991), .CI(n992), .CO(n988) );
  MUX U1984 ( .A(imm[10]), .B(reg_source[4]), .S(n913), .Z(n992) );
  FA U1985 ( .A(a_bus[3]), .B(n993), .CI(n994), .CO(n991) );
  FA U1986 ( .A(n995), .B(n996), .CI(n997), .CO(n993) );
  MUX U1987 ( .A(imm[8]), .B(reg_source[2]), .S(n913), .Z(n997) );
  NAND U1988 ( .A(n998), .B(n999), .Z(n996) );
  NANDN U1989 ( .A(n1000), .B(a_bus[1]), .Z(n999) );
  NAND U1990 ( .A(n1001), .B(n1002), .Z(n998) );
  NAND U1991 ( .A(n1003), .B(n1000), .Z(n1002) );
  ANDN U1992 ( .B(n1004), .A(n1005), .Z(n1000) );
  NAND U1993 ( .A(b_bus[9]), .B(n1006), .Z(n978) );
  NAND U1994 ( .A(b_bus[10]), .B(n1007), .Z(n970) );
  AND U1995 ( .A(reg_source[11]), .B(n913), .Z(n967) );
  AND U1996 ( .A(reg_source[13]), .B(n913), .Z(n962) );
  AND U1997 ( .A(reg_source[15]), .B(n913), .Z(n957) );
  AND U1998 ( .A(n1008), .B(n918), .Z(n955) );
  AND U1999 ( .A(reg_source[17]), .B(n913), .Z(n952) );
  AND U2000 ( .A(n1009), .B(n918), .Z(n950) );
  AND U2001 ( .A(reg_source[19]), .B(n913), .Z(n946) );
  AND U2002 ( .A(n1010), .B(n918), .Z(n944) );
  AND U2003 ( .A(reg_source[21]), .B(n913), .Z(n940) );
  AND U2004 ( .A(n1011), .B(n918), .Z(n938) );
  AND U2005 ( .A(reg_source[23]), .B(n913), .Z(n934) );
  AND U2006 ( .A(n1012), .B(n918), .Z(n932) );
  AND U2007 ( .A(reg_source[25]), .B(n913), .Z(n928) );
  AND U2008 ( .A(n1013), .B(n918), .Z(n926) );
  AND U2009 ( .A(reg_source[27]), .B(n913), .Z(n922) );
  AND U2010 ( .A(n1014), .B(n918), .Z(n920) );
  AND U2011 ( .A(reg_source[29]), .B(n913), .Z(n915) );
  IV U2012 ( .A(n1015), .Z(n913) );
  IV U2013 ( .A(n904), .Z(n910) );
  AND U2014 ( .A(n1016), .B(n1017), .Z(n904) );
  ANDN U2015 ( .B(n1018), .A(n1019), .Z(n1016) );
  AND U2016 ( .A(n1020), .B(n1021), .Z(n892) );
  MUX U2017 ( .A(n1022), .B(n1023), .S(n1024), .Z(n1021) );
  AND U2018 ( .A(n1005), .B(n1004), .Z(n1024) );
  NAND U2019 ( .A(n1025), .B(n1026), .Z(n1020) );
  XOR U2020 ( .A(a_bus[0]), .B(b_bus[0]), .Z(n1025) );
  AND U2021 ( .A(n1027), .B(n1028), .Z(n426) );
  AND U2022 ( .A(n1029), .B(n1030), .Z(n1028) );
  AND U2023 ( .A(n1031), .B(n1032), .Z(n1030) );
  NAND U2024 ( .A(n1033), .B(n852), .Z(n1032) );
  NAND U2025 ( .A(n1034), .B(n1035), .Z(n1033) );
  AND U2026 ( .A(n1036), .B(n1037), .Z(n1035) );
  AND U2027 ( .A(n1038), .B(n1039), .Z(n1036) );
  NANDN U2028 ( .A(n1040), .B(a_bus[4]), .Z(n1039) );
  AND U2029 ( .A(n1041), .B(n1042), .Z(n1034) );
  NAND U2030 ( .A(n1043), .B(n863), .Z(n1042) );
  NAND U2031 ( .A(n1044), .B(n865), .Z(n1031) );
  NAND U2032 ( .A(n1045), .B(n1046), .Z(n1044) );
  AND U2033 ( .A(n1047), .B(n1037), .Z(n1046) );
  NAND U2034 ( .A(n870), .B(n1048), .Z(n1037) );
  AND U2035 ( .A(n1038), .B(n1049), .Z(n1047) );
  NANDN U2036 ( .A(n1050), .B(a_bus[4]), .Z(n1049) );
  NANDN U2037 ( .A(n1051), .B(n874), .Z(n1038) );
  AND U2038 ( .A(n1041), .B(n1052), .Z(n1045) );
  NAND U2039 ( .A(n1043), .B(n876), .Z(n1052) );
  NAND U2040 ( .A(n1053), .B(n1054), .Z(n1043) );
  AND U2041 ( .A(n1055), .B(n1056), .Z(n1054) );
  NANDN U2042 ( .A(n881), .B(b_bus[1]), .Z(n1056) );
  NANDN U2043 ( .A(n882), .B(b_bus[2]), .Z(n1055) );
  AND U2044 ( .A(n1057), .B(n1058), .Z(n1053) );
  NANDN U2045 ( .A(n885), .B(b_bus[4]), .Z(n1058) );
  NANDN U2046 ( .A(n886), .B(b_bus[3]), .Z(n1057) );
  NAND U2047 ( .A(n888), .B(n1059), .Z(n1041) );
  AND U2048 ( .A(n1060), .B(n1061), .Z(n1029) );
  NAND U2049 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][1] ), .Z(n1061) );
  ANDN U2050 ( .B(\Shifter/sll_27/ML_int[3][1] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][1] ) );
  ANDN U2051 ( .B(\Shifter/sll_27/ML_int[2][1] ), .A(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][1] ) );
  ANDN U2052 ( .B(\Shifter/sll_27/ML_int[1][1] ), .A(a_bus[1]), .Z(
        \Shifter/sll_27/ML_int[2][1] ) );
  NAND U2053 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N109 ), .Z(n1060) );
  AND U2054 ( .A(n1062), .B(n1063), .Z(n1027) );
  AND U2055 ( .A(n1064), .B(n1065), .Z(n1063) );
  NANDN U2056 ( .A(n891), .B(\ALU/N109 ), .Z(n1065) );
  NAND U2057 ( .A(n1066), .B(n1026), .Z(n1064) );
  XOR U2058 ( .A(a_bus[1]), .B(b_bus[1]), .Z(n1066) );
  AND U2059 ( .A(n1067), .B(n1068), .Z(n1062) );
  NAND U2060 ( .A(n1069), .B(n897), .Z(n1068) );
  AND U2061 ( .A(b_bus[1]), .B(a_bus[1]), .Z(n1069) );
  MUX U2062 ( .A(n1022), .B(n1023), .S(n1070), .Z(n1067) );
  AND U2063 ( .A(n1001), .B(n1003), .Z(n1070) );
  AND U2064 ( .A(n1071), .B(n1072), .Z(n828) );
  AND U2065 ( .A(n1073), .B(n1074), .Z(n1072) );
  NOR U2066 ( .A(n394), .B(n389), .Z(n1074) );
  NAND U2067 ( .A(n1075), .B(n1076), .Z(n389) );
  AND U2068 ( .A(n1077), .B(n1078), .Z(n1076) );
  AND U2069 ( .A(n1079), .B(n1080), .Z(n1078) );
  NAND U2070 ( .A(n1081), .B(n852), .Z(n1080) );
  NAND U2071 ( .A(n1082), .B(n1083), .Z(n1081) );
  AND U2072 ( .A(n1084), .B(n1085), .Z(n1083) );
  AND U2073 ( .A(n1086), .B(n1087), .Z(n1084) );
  NANDN U2074 ( .A(n1088), .B(a_bus[4]), .Z(n1087) );
  NAND U2075 ( .A(n1048), .B(n863), .Z(n1086) );
  NAND U2076 ( .A(n1089), .B(n865), .Z(n1079) );
  NAND U2077 ( .A(n1082), .B(n1090), .Z(n1089) );
  AND U2078 ( .A(n1091), .B(n1085), .Z(n1090) );
  NAND U2079 ( .A(n888), .B(n1092), .Z(n1085) );
  AND U2080 ( .A(n1093), .B(n1094), .Z(n1091) );
  NANDN U2081 ( .A(n1095), .B(a_bus[4]), .Z(n1094) );
  NAND U2082 ( .A(n1048), .B(n876), .Z(n1093) );
  AND U2083 ( .A(n1096), .B(n1097), .Z(n1082) );
  NAND U2084 ( .A(n870), .B(n1098), .Z(n1097) );
  NAND U2085 ( .A(n1059), .B(n874), .Z(n1096) );
  AND U2086 ( .A(n1099), .B(n1100), .Z(n1077) );
  NAND U2087 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][9] ), .Z(n1100) );
  NAND U2088 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N117 ), .Z(n1099) );
  AND U2089 ( .A(n1101), .B(n1102), .Z(n1075) );
  AND U2090 ( .A(n1103), .B(n1104), .Z(n1102) );
  NANDN U2091 ( .A(n891), .B(\ALU/N117 ), .Z(n1104) );
  NAND U2092 ( .A(n1105), .B(n1026), .Z(n1103) );
  XOR U2093 ( .A(n974), .B(n1006), .Z(n1105) );
  AND U2094 ( .A(n1106), .B(n1107), .Z(n1101) );
  NAND U2095 ( .A(n2481), .B(n1108), .Z(n1107) );
  AND U2096 ( .A(n897), .B(b_bus[9]), .Z(n1108) );
  MUX U2097 ( .A(n1022), .B(n1023), .S(n1109), .Z(n1106) );
  AND U2098 ( .A(n974), .B(n1006), .Z(n1109) );
  IV U2099 ( .A(n2481), .Z(n1006) );
  ANDN U2100 ( .B(reg_source[9]), .A(n1015), .Z(n2481) );
  NAND U2101 ( .A(n1110), .B(n1111), .Z(n394) );
  AND U2102 ( .A(n1112), .B(n1113), .Z(n1111) );
  AND U2103 ( .A(n1114), .B(n1115), .Z(n1113) );
  NAND U2104 ( .A(n1116), .B(n852), .Z(n1115) );
  NAND U2105 ( .A(n1117), .B(n1118), .Z(n1116) );
  AND U2106 ( .A(n1119), .B(n1120), .Z(n1118) );
  AND U2107 ( .A(n1121), .B(n1122), .Z(n1119) );
  NANDN U2108 ( .A(n1123), .B(a_bus[4]), .Z(n1122) );
  NAND U2109 ( .A(n869), .B(n863), .Z(n1121) );
  NAND U2110 ( .A(n1124), .B(n865), .Z(n1114) );
  NAND U2111 ( .A(n1117), .B(n1125), .Z(n1124) );
  AND U2112 ( .A(n1126), .B(n1120), .Z(n1125) );
  NAND U2113 ( .A(n888), .B(n1127), .Z(n1120) );
  AND U2114 ( .A(n1128), .B(n1129), .Z(n1126) );
  NANDN U2115 ( .A(n1130), .B(a_bus[4]), .Z(n1129) );
  NAND U2116 ( .A(n869), .B(n876), .Z(n1128) );
  AND U2117 ( .A(n1131), .B(n1132), .Z(n1117) );
  NAND U2118 ( .A(n870), .B(n1133), .Z(n1132) );
  NAND U2119 ( .A(n887), .B(n874), .Z(n1131) );
  AND U2120 ( .A(n1134), .B(n1135), .Z(n1112) );
  NAND U2121 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][8] ), .Z(n1135) );
  NAND U2122 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N116 ), .Z(n1134) );
  AND U2123 ( .A(n1136), .B(n1137), .Z(n1110) );
  AND U2124 ( .A(n1138), .B(n1139), .Z(n1137) );
  NANDN U2125 ( .A(n891), .B(\ALU/N116 ), .Z(n1139) );
  NAND U2126 ( .A(n1140), .B(n1026), .Z(n1138) );
  XNOR U2127 ( .A(n980), .B(n2482), .Z(n1140) );
  AND U2128 ( .A(n1141), .B(n1142), .Z(n1136) );
  NAND U2129 ( .A(n1143), .B(n2482), .Z(n1142) );
  AND U2130 ( .A(n897), .B(b_bus[8]), .Z(n1143) );
  MUX U2131 ( .A(n1022), .B(n1023), .S(n1144), .Z(n1141) );
  NOR U2132 ( .A(b_bus[8]), .B(n2482), .Z(n1144) );
  ANDN U2133 ( .B(reg_source[8]), .A(n1015), .Z(n2482) );
  AND U2134 ( .A(n1145), .B(n1146), .Z(n1073) );
  IV U2135 ( .A(n379), .Z(n1146) );
  NAND U2136 ( .A(n1147), .B(n1148), .Z(n379) );
  AND U2137 ( .A(n1149), .B(n1150), .Z(n1148) );
  AND U2138 ( .A(n1151), .B(n1152), .Z(n1150) );
  NAND U2139 ( .A(n1153), .B(n852), .Z(n1152) );
  NAND U2140 ( .A(n1154), .B(n1155), .Z(n1153) );
  AND U2141 ( .A(n1156), .B(n1157), .Z(n1155) );
  AND U2142 ( .A(n1158), .B(n1159), .Z(n1156) );
  NAND U2143 ( .A(a_bus[4]), .B(n1160), .Z(n1159) );
  NAND U2144 ( .A(n1161), .B(n863), .Z(n1158) );
  AND U2145 ( .A(n1162), .B(n1163), .Z(n1154) );
  NAND U2146 ( .A(n1164), .B(n865), .Z(n1151) );
  NAND U2147 ( .A(n1165), .B(n1166), .Z(n1164) );
  AND U2148 ( .A(n1167), .B(n1163), .Z(n1166) );
  NAND U2149 ( .A(n870), .B(n1168), .Z(n1163) );
  AND U2150 ( .A(n1162), .B(n1169), .Z(n1167) );
  NAND U2151 ( .A(n1161), .B(n876), .Z(n1169) );
  NAND U2152 ( .A(n1170), .B(n874), .Z(n1162) );
  AND U2153 ( .A(n1157), .B(n1171), .Z(n1165) );
  NAND U2154 ( .A(n1172), .B(n1173), .Z(n1171) );
  AND U2155 ( .A(a_bus[4]), .B(n1174), .Z(n1173) );
  NAND U2156 ( .A(n888), .B(n1175), .Z(n1157) );
  AND U2157 ( .A(n1176), .B(n1177), .Z(n1149) );
  NAND U2158 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][11] ), .Z(n1177) );
  NAND U2159 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N119 ), .Z(n1176) );
  AND U2160 ( .A(n1178), .B(n1179), .Z(n1147) );
  AND U2161 ( .A(n1180), .B(n1181), .Z(n1179) );
  NANDN U2162 ( .A(n891), .B(\ALU/N119 ), .Z(n1181) );
  NAND U2163 ( .A(n1182), .B(n1026), .Z(n1180) );
  XNOR U2164 ( .A(n969), .B(n2506), .Z(n1182) );
  AND U2165 ( .A(n1183), .B(n1184), .Z(n1178) );
  NAND U2166 ( .A(n1185), .B(n2506), .Z(n1184) );
  AND U2167 ( .A(n897), .B(b_bus[11]), .Z(n1185) );
  MUX U2168 ( .A(n1022), .B(n1023), .S(n1186), .Z(n1183) );
  NOR U2169 ( .A(b_bus[11]), .B(n2506), .Z(n1186) );
  ANDN U2170 ( .B(reg_source[11]), .A(n1015), .Z(n2506) );
  IV U2171 ( .A(n384), .Z(n1145) );
  NAND U2172 ( .A(n1187), .B(n1188), .Z(n384) );
  AND U2173 ( .A(n1189), .B(n1190), .Z(n1188) );
  AND U2174 ( .A(n1191), .B(n1192), .Z(n1190) );
  NAND U2175 ( .A(n1193), .B(n852), .Z(n1192) );
  NAND U2176 ( .A(n1194), .B(n1195), .Z(n1193) );
  AND U2177 ( .A(n1196), .B(n1197), .Z(n1195) );
  AND U2178 ( .A(n1198), .B(n1199), .Z(n1196) );
  NANDN U2179 ( .A(n1200), .B(a_bus[4]), .Z(n1199) );
  NAND U2180 ( .A(n1201), .B(n863), .Z(n1198) );
  NAND U2181 ( .A(n1202), .B(n865), .Z(n1191) );
  NAND U2182 ( .A(n1194), .B(n1203), .Z(n1202) );
  AND U2183 ( .A(n1204), .B(n1197), .Z(n1203) );
  NAND U2184 ( .A(n888), .B(n1205), .Z(n1197) );
  AND U2185 ( .A(n1206), .B(n1207), .Z(n1204) );
  NANDN U2186 ( .A(n1208), .B(a_bus[4]), .Z(n1207) );
  NAND U2187 ( .A(n1201), .B(n876), .Z(n1206) );
  AND U2188 ( .A(n1209), .B(n1210), .Z(n1194) );
  NAND U2189 ( .A(n870), .B(n1211), .Z(n1210) );
  NAND U2190 ( .A(n1212), .B(n874), .Z(n1209) );
  AND U2191 ( .A(n1213), .B(n1214), .Z(n1189) );
  NAND U2192 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][10] ), .Z(n1214) );
  NAND U2193 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N118 ), .Z(n1213) );
  AND U2194 ( .A(n1215), .B(n1216), .Z(n1187) );
  AND U2195 ( .A(n1217), .B(n1218), .Z(n1216) );
  NANDN U2196 ( .A(n891), .B(\ALU/N118 ), .Z(n1218) );
  NAND U2197 ( .A(n1219), .B(n1026), .Z(n1217) );
  XOR U2198 ( .A(n977), .B(n1007), .Z(n1219) );
  AND U2199 ( .A(n1220), .B(n1221), .Z(n1215) );
  NAND U2200 ( .A(n2507), .B(n1222), .Z(n1221) );
  AND U2201 ( .A(n897), .B(b_bus[10]), .Z(n1222) );
  MUX U2202 ( .A(n1022), .B(n1023), .S(n1223), .Z(n1220) );
  AND U2203 ( .A(n977), .B(n1007), .Z(n1223) );
  IV U2204 ( .A(n2507), .Z(n1007) );
  ANDN U2205 ( .B(reg_source[10]), .A(n1015), .Z(n2507) );
  AND U2206 ( .A(n1224), .B(n1225), .Z(n1071) );
  AND U2207 ( .A(n1226), .B(n1227), .Z(n1225) );
  IV U2208 ( .A(n369), .Z(n1227) );
  NAND U2209 ( .A(n1228), .B(n1229), .Z(n369) );
  AND U2210 ( .A(n1230), .B(n1231), .Z(n1229) );
  AND U2211 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U2212 ( .A(n1234), .B(n852), .Z(n1233) );
  NAND U2213 ( .A(n1235), .B(n1236), .Z(n1234) );
  AND U2214 ( .A(n1237), .B(n1238), .Z(n1236) );
  AND U2215 ( .A(n1239), .B(n1240), .Z(n1237) );
  NANDN U2216 ( .A(n1241), .B(a_bus[4]), .Z(n1240) );
  NAND U2217 ( .A(n1059), .B(n863), .Z(n1239) );
  AND U2218 ( .A(n1242), .B(n1243), .Z(n1235) );
  NAND U2219 ( .A(n1244), .B(n865), .Z(n1232) );
  NAND U2220 ( .A(n1245), .B(n1246), .Z(n1244) );
  AND U2221 ( .A(n1247), .B(n1243), .Z(n1246) );
  NAND U2222 ( .A(n870), .B(n1092), .Z(n1243) );
  AND U2223 ( .A(n1242), .B(n1248), .Z(n1247) );
  NAND U2224 ( .A(n1059), .B(n876), .Z(n1248) );
  NAND U2225 ( .A(n1098), .B(n874), .Z(n1242) );
  AND U2226 ( .A(n1238), .B(n1249), .Z(n1245) );
  NAND U2227 ( .A(n1250), .B(n1251), .Z(n1249) );
  NAND U2228 ( .A(n888), .B(n1252), .Z(n1238) );
  AND U2229 ( .A(n1253), .B(n1254), .Z(n1230) );
  NAND U2230 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][13] ), .Z(n1254) );
  NAND U2231 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N121 ), .Z(n1253) );
  AND U2232 ( .A(n1255), .B(n1256), .Z(n1228) );
  AND U2233 ( .A(n1257), .B(n1258), .Z(n1256) );
  NANDN U2234 ( .A(n891), .B(\ALU/N121 ), .Z(n1258) );
  NAND U2235 ( .A(n1259), .B(n1026), .Z(n1257) );
  XNOR U2236 ( .A(n964), .B(n2504), .Z(n1259) );
  AND U2237 ( .A(n1260), .B(n1261), .Z(n1255) );
  NAND U2238 ( .A(n1262), .B(n2504), .Z(n1261) );
  AND U2239 ( .A(n897), .B(b_bus[13]), .Z(n1262) );
  MUX U2240 ( .A(n1022), .B(n1023), .S(n1263), .Z(n1260) );
  NOR U2241 ( .A(b_bus[13]), .B(n2504), .Z(n1263) );
  ANDN U2242 ( .B(reg_source[13]), .A(n1015), .Z(n2504) );
  IV U2243 ( .A(n374), .Z(n1226) );
  NAND U2244 ( .A(n1264), .B(n1265), .Z(n374) );
  AND U2245 ( .A(n1266), .B(n1267), .Z(n1265) );
  AND U2246 ( .A(n1268), .B(n1269), .Z(n1267) );
  NAND U2247 ( .A(n1270), .B(n852), .Z(n1269) );
  NAND U2248 ( .A(n1271), .B(n1272), .Z(n1270) );
  AND U2249 ( .A(n1273), .B(n1274), .Z(n1272) );
  AND U2250 ( .A(n1275), .B(n1276), .Z(n1273) );
  NANDN U2251 ( .A(n1277), .B(a_bus[4]), .Z(n1276) );
  NAND U2252 ( .A(n887), .B(n863), .Z(n1275) );
  AND U2253 ( .A(n1278), .B(n1279), .Z(n1271) );
  NAND U2254 ( .A(n1280), .B(n865), .Z(n1268) );
  NAND U2255 ( .A(n1281), .B(n1282), .Z(n1280) );
  AND U2256 ( .A(n1283), .B(n1279), .Z(n1282) );
  NAND U2257 ( .A(n870), .B(n1127), .Z(n1279) );
  AND U2258 ( .A(n1278), .B(n1284), .Z(n1283) );
  NAND U2259 ( .A(n887), .B(n876), .Z(n1284) );
  NAND U2260 ( .A(n1133), .B(n874), .Z(n1278) );
  AND U2261 ( .A(n1274), .B(n1285), .Z(n1281) );
  NAND U2262 ( .A(n1286), .B(n1250), .Z(n1285) );
  NAND U2263 ( .A(n888), .B(n1287), .Z(n1274) );
  AND U2264 ( .A(n1288), .B(n1289), .Z(n1266) );
  NAND U2265 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][12] ), .Z(n1289) );
  NAND U2266 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N120 ), .Z(n1288) );
  AND U2267 ( .A(n1290), .B(n1291), .Z(n1264) );
  AND U2268 ( .A(n1292), .B(n1293), .Z(n1291) );
  NANDN U2269 ( .A(n891), .B(\ALU/N120 ), .Z(n1293) );
  NAND U2270 ( .A(n1294), .B(n1026), .Z(n1292) );
  XNOR U2271 ( .A(n965), .B(n2505), .Z(n1294) );
  AND U2272 ( .A(n1295), .B(n1296), .Z(n1290) );
  NAND U2273 ( .A(n1297), .B(n2505), .Z(n1296) );
  AND U2274 ( .A(n897), .B(b_bus[12]), .Z(n1297) );
  MUX U2275 ( .A(n1022), .B(n1023), .S(n1298), .Z(n1295) );
  NOR U2276 ( .A(b_bus[12]), .B(n2505), .Z(n1298) );
  ANDN U2277 ( .B(reg_source[12]), .A(n1015), .Z(n2505) );
  AND U2278 ( .A(n1299), .B(n1300), .Z(n1224) );
  IV U2279 ( .A(n359), .Z(n1300) );
  NAND U2280 ( .A(n1301), .B(n1302), .Z(n359) );
  AND U2281 ( .A(n1303), .B(n1304), .Z(n1302) );
  AND U2282 ( .A(n1305), .B(n1306), .Z(n1304) );
  NAND U2283 ( .A(n1307), .B(n852), .Z(n1306) );
  NAND U2284 ( .A(n1308), .B(n1309), .Z(n1307) );
  AND U2285 ( .A(n1310), .B(n1311), .Z(n1309) );
  AND U2286 ( .A(n1312), .B(n1313), .Z(n1310) );
  NAND U2287 ( .A(n1170), .B(n863), .Z(n1313) );
  AND U2288 ( .A(n1314), .B(n1315), .Z(n1308) );
  NAND U2289 ( .A(n888), .B(n1316), .Z(n1314) );
  NAND U2290 ( .A(n1317), .B(n865), .Z(n1305) );
  NAND U2291 ( .A(n1318), .B(n1319), .Z(n1317) );
  AND U2292 ( .A(n1320), .B(n1315), .Z(n1319) );
  NAND U2293 ( .A(n870), .B(n1175), .Z(n1315) );
  AND U2294 ( .A(n1311), .B(n1321), .Z(n1320) );
  NAND U2295 ( .A(n1170), .B(n876), .Z(n1321) );
  NAND U2296 ( .A(n1168), .B(n874), .Z(n1311) );
  AND U2297 ( .A(n1322), .B(n1323), .Z(n1318) );
  NANDN U2298 ( .A(n1324), .B(n1250), .Z(n1323) );
  NANDN U2299 ( .A(n1325), .B(n888), .Z(n1322) );
  AND U2300 ( .A(n1326), .B(n1327), .Z(n1303) );
  NAND U2301 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][15] ), .Z(n1327) );
  NAND U2302 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N123 ), .Z(n1326) );
  AND U2303 ( .A(n1328), .B(n1329), .Z(n1301) );
  AND U2304 ( .A(n1330), .B(n1331), .Z(n1329) );
  NANDN U2305 ( .A(n891), .B(\ALU/N123 ), .Z(n1331) );
  NAND U2306 ( .A(n1332), .B(n1026), .Z(n1330) );
  XNOR U2307 ( .A(n959), .B(n2502), .Z(n1332) );
  AND U2308 ( .A(n1333), .B(n1334), .Z(n1328) );
  NAND U2309 ( .A(n1335), .B(n2502), .Z(n1334) );
  AND U2310 ( .A(n897), .B(b_bus[15]), .Z(n1335) );
  MUX U2311 ( .A(n1022), .B(n1023), .S(n1336), .Z(n1333) );
  NOR U2312 ( .A(b_bus[15]), .B(n2502), .Z(n1336) );
  ANDN U2313 ( .B(reg_source[15]), .A(n1015), .Z(n2502) );
  IV U2314 ( .A(n364), .Z(n1299) );
  NAND U2315 ( .A(n1337), .B(n1338), .Z(n364) );
  AND U2316 ( .A(n1339), .B(n1340), .Z(n1338) );
  AND U2317 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U2318 ( .A(n1343), .B(n852), .Z(n1342) );
  NAND U2319 ( .A(n1344), .B(n1345), .Z(n1343) );
  AND U2320 ( .A(n1346), .B(n1347), .Z(n1345) );
  AND U2321 ( .A(n1348), .B(n1349), .Z(n1346) );
  NANDN U2322 ( .A(n1350), .B(a_bus[4]), .Z(n1349) );
  NAND U2323 ( .A(n1212), .B(n863), .Z(n1348) );
  AND U2324 ( .A(n1351), .B(n1352), .Z(n1344) );
  NAND U2325 ( .A(n1353), .B(n865), .Z(n1341) );
  NAND U2326 ( .A(n1354), .B(n1355), .Z(n1353) );
  AND U2327 ( .A(n1356), .B(n1352), .Z(n1355) );
  NAND U2328 ( .A(n870), .B(n1205), .Z(n1352) );
  AND U2329 ( .A(n1351), .B(n1357), .Z(n1356) );
  NAND U2330 ( .A(n1212), .B(n876), .Z(n1357) );
  NAND U2331 ( .A(n1211), .B(n874), .Z(n1351) );
  AND U2332 ( .A(n1347), .B(n1358), .Z(n1354) );
  NAND U2333 ( .A(n1250), .B(n1359), .Z(n1358) );
  ANDN U2334 ( .B(n1360), .A(n1361), .Z(n1250) );
  NAND U2335 ( .A(n888), .B(n1362), .Z(n1347) );
  AND U2336 ( .A(n1363), .B(n1364), .Z(n1339) );
  NAND U2337 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][14] ), .Z(n1364) );
  NAND U2338 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N122 ), .Z(n1363) );
  AND U2339 ( .A(n1365), .B(n1366), .Z(n1337) );
  AND U2340 ( .A(n1367), .B(n1368), .Z(n1366) );
  NANDN U2341 ( .A(n891), .B(\ALU/N122 ), .Z(n1368) );
  NAND U2342 ( .A(n1369), .B(n1026), .Z(n1367) );
  XNOR U2343 ( .A(n960), .B(n2503), .Z(n1369) );
  AND U2344 ( .A(n1370), .B(n1371), .Z(n1365) );
  NAND U2345 ( .A(n1372), .B(n2503), .Z(n1371) );
  AND U2346 ( .A(n897), .B(b_bus[14]), .Z(n1372) );
  MUX U2347 ( .A(n1022), .B(n1023), .S(n1373), .Z(n1370) );
  NOR U2348 ( .A(b_bus[14]), .B(n2503), .Z(n1373) );
  ANDN U2349 ( .B(reg_source[14]), .A(n1015), .Z(n2503) );
  AND U2350 ( .A(n1374), .B(n1375), .Z(n826) );
  AND U2351 ( .A(n1376), .B(n1377), .Z(n1375) );
  AND U2352 ( .A(n1378), .B(n1379), .Z(n1377) );
  AND U2353 ( .A(n1380), .B(n1381), .Z(n1379) );
  IV U2354 ( .A(n344), .Z(n1381) );
  NAND U2355 ( .A(n1382), .B(n1383), .Z(n344) );
  AND U2356 ( .A(n1384), .B(n1385), .Z(n1383) );
  AND U2357 ( .A(n1386), .B(n1387), .Z(n1385) );
  NAND U2358 ( .A(n1388), .B(n852), .Z(n1387) );
  NAND U2359 ( .A(n1389), .B(n1312), .Z(n1388) );
  NANDN U2360 ( .A(n1040), .B(n1361), .Z(n1389) );
  AND U2361 ( .A(n1390), .B(n1391), .Z(n1040) );
  AND U2362 ( .A(n1392), .B(n1393), .Z(n1391) );
  NAND U2363 ( .A(n1098), .B(n1394), .Z(n1393) );
  AND U2364 ( .A(n1395), .B(n1396), .Z(n1390) );
  NAND U2365 ( .A(n1397), .B(n1398), .Z(n1395) );
  NAND U2366 ( .A(n1399), .B(n865), .Z(n1386) );
  ANDN U2367 ( .B(n1361), .A(n1050), .Z(n1399) );
  AND U2368 ( .A(n1400), .B(n1401), .Z(n1050) );
  AND U2369 ( .A(n1392), .B(n1402), .Z(n1401) );
  NAND U2370 ( .A(n1360), .B(n1098), .Z(n1402) );
  NAND U2371 ( .A(n1092), .B(n1403), .Z(n1392) );
  AND U2372 ( .A(n1404), .B(n1396), .Z(n1400) );
  NAND U2373 ( .A(n1405), .B(n1252), .Z(n1396) );
  NAND U2374 ( .A(n1251), .B(n1397), .Z(n1404) );
  AND U2375 ( .A(n1406), .B(n1407), .Z(n1384) );
  NANDN U2376 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][17] ), .Z(n1407) );
  NAND U2377 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N125 ), .Z(n1406) );
  AND U2378 ( .A(n1409), .B(n1410), .Z(n1382) );
  AND U2379 ( .A(n1411), .B(n1412), .Z(n1410) );
  NANDN U2380 ( .A(n891), .B(\ALU/N125 ), .Z(n1412) );
  NAND U2381 ( .A(n1413), .B(n1026), .Z(n1411) );
  XNOR U2382 ( .A(n954), .B(n2500), .Z(n1413) );
  AND U2383 ( .A(n1414), .B(n1415), .Z(n1409) );
  NAND U2384 ( .A(n1416), .B(n2500), .Z(n1415) );
  AND U2385 ( .A(n897), .B(b_bus[17]), .Z(n1416) );
  MUX U2386 ( .A(n1022), .B(n1023), .S(n1417), .Z(n1414) );
  NOR U2387 ( .A(b_bus[17]), .B(n2500), .Z(n1417) );
  ANDN U2388 ( .B(reg_source[17]), .A(n1015), .Z(n2500) );
  IV U2389 ( .A(n351), .Z(n1380) );
  NAND U2390 ( .A(n1418), .B(n1419), .Z(n351) );
  AND U2391 ( .A(n1420), .B(n1421), .Z(n1419) );
  AND U2392 ( .A(n1422), .B(n1423), .Z(n1421) );
  NAND U2393 ( .A(n1424), .B(n852), .Z(n1423) );
  NAND U2394 ( .A(n1425), .B(n1312), .Z(n1424) );
  NANDN U2395 ( .A(n859), .B(n1361), .Z(n1425) );
  AND U2396 ( .A(n1426), .B(n1427), .Z(n859) );
  AND U2397 ( .A(n1428), .B(n1429), .Z(n1427) );
  NAND U2398 ( .A(n1133), .B(n1394), .Z(n1429) );
  NAND U2399 ( .A(n1430), .B(n865), .Z(n1422) );
  ANDN U2400 ( .B(n1361), .A(n872), .Z(n1430) );
  AND U2401 ( .A(n1426), .B(n1431), .Z(n872) );
  AND U2402 ( .A(n1428), .B(n1432), .Z(n1431) );
  NAND U2403 ( .A(n1360), .B(n1133), .Z(n1432) );
  NAND U2404 ( .A(n1127), .B(n1403), .Z(n1428) );
  AND U2405 ( .A(n1433), .B(n1434), .Z(n1426) );
  NAND U2406 ( .A(n1287), .B(n1405), .Z(n1434) );
  NAND U2407 ( .A(n1286), .B(n1397), .Z(n1433) );
  AND U2408 ( .A(n1435), .B(n1436), .Z(n1420) );
  NANDN U2409 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][16] ), .Z(n1436) );
  NAND U2410 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N124 ), .Z(n1435) );
  AND U2411 ( .A(n1437), .B(n1438), .Z(n1418) );
  AND U2412 ( .A(n1439), .B(n1440), .Z(n1438) );
  NANDN U2413 ( .A(n891), .B(\ALU/N124 ), .Z(n1440) );
  NAND U2414 ( .A(n1441), .B(n1026), .Z(n1439) );
  XNOR U2415 ( .A(n955), .B(n2501), .Z(n1441) );
  AND U2416 ( .A(n1442), .B(n1443), .Z(n1437) );
  NAND U2417 ( .A(n1444), .B(n2501), .Z(n1443) );
  AND U2418 ( .A(n897), .B(b_bus[16]), .Z(n1444) );
  MUX U2419 ( .A(n1022), .B(n1023), .S(n1445), .Z(n1442) );
  NOR U2420 ( .A(b_bus[16]), .B(n2501), .Z(n1445) );
  ANDN U2421 ( .B(reg_source[16]), .A(n1015), .Z(n2501) );
  AND U2422 ( .A(n1446), .B(n1447), .Z(n1378) );
  IV U2423 ( .A(n330), .Z(n1447) );
  NAND U2424 ( .A(n1448), .B(n1449), .Z(n330) );
  AND U2425 ( .A(n1450), .B(n1451), .Z(n1449) );
  AND U2426 ( .A(n1452), .B(n1453), .Z(n1451) );
  NAND U2427 ( .A(n1454), .B(n852), .Z(n1453) );
  NAND U2428 ( .A(n1455), .B(n1312), .Z(n1454) );
  NANDN U2429 ( .A(n1456), .B(n1361), .Z(n1455) );
  NAND U2430 ( .A(n1457), .B(n865), .Z(n1452) );
  ANDN U2431 ( .B(n1361), .A(n1458), .Z(n1457) );
  AND U2432 ( .A(n1459), .B(n1460), .Z(n1450) );
  NANDN U2433 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][19] ), .Z(n1460) );
  NAND U2434 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N127 ), .Z(n1459) );
  AND U2435 ( .A(n1461), .B(n1462), .Z(n1448) );
  AND U2436 ( .A(n1463), .B(n1464), .Z(n1462) );
  NANDN U2437 ( .A(n891), .B(\ALU/N127 ), .Z(n1464) );
  NAND U2438 ( .A(n1465), .B(n1026), .Z(n1463) );
  XNOR U2439 ( .A(n1466), .B(n2498), .Z(n1465) );
  AND U2440 ( .A(n1467), .B(n1468), .Z(n1461) );
  NAND U2441 ( .A(n1469), .B(n2498), .Z(n1468) );
  AND U2442 ( .A(n897), .B(b_bus[19]), .Z(n1469) );
  MUX U2443 ( .A(n1022), .B(n1023), .S(n1470), .Z(n1467) );
  NOR U2444 ( .A(b_bus[19]), .B(n2498), .Z(n1470) );
  ANDN U2445 ( .B(reg_source[19]), .A(n1015), .Z(n2498) );
  IV U2446 ( .A(n337), .Z(n1446) );
  NAND U2447 ( .A(n1471), .B(n1472), .Z(n337) );
  AND U2448 ( .A(n1473), .B(n1474), .Z(n1472) );
  AND U2449 ( .A(n1475), .B(n1476), .Z(n1474) );
  NAND U2450 ( .A(n1477), .B(n852), .Z(n1476) );
  NAND U2451 ( .A(n1478), .B(n1312), .Z(n1477) );
  NANDN U2452 ( .A(n1479), .B(n1361), .Z(n1478) );
  NAND U2453 ( .A(n1480), .B(n865), .Z(n1475) );
  ANDN U2454 ( .B(n1361), .A(n1481), .Z(n1480) );
  AND U2455 ( .A(n1482), .B(n1483), .Z(n1473) );
  NANDN U2456 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][18] ), .Z(n1483) );
  NAND U2457 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N126 ), .Z(n1482) );
  AND U2458 ( .A(n1484), .B(n1485), .Z(n1471) );
  AND U2459 ( .A(n1486), .B(n1487), .Z(n1485) );
  NANDN U2460 ( .A(n891), .B(\ALU/N126 ), .Z(n1487) );
  NAND U2461 ( .A(n1488), .B(n1026), .Z(n1486) );
  XNOR U2462 ( .A(n950), .B(n2499), .Z(n1488) );
  AND U2463 ( .A(n1489), .B(n1490), .Z(n1484) );
  NAND U2464 ( .A(n1491), .B(n2499), .Z(n1490) );
  AND U2465 ( .A(n897), .B(b_bus[18]), .Z(n1491) );
  MUX U2466 ( .A(n1022), .B(n1023), .S(n1492), .Z(n1489) );
  NOR U2467 ( .A(b_bus[18]), .B(n2499), .Z(n1492) );
  ANDN U2468 ( .B(reg_source[18]), .A(n1015), .Z(n2499) );
  AND U2469 ( .A(n1493), .B(n1494), .Z(n1376) );
  AND U2470 ( .A(n1495), .B(n1496), .Z(n1494) );
  IV U2471 ( .A(n316), .Z(n1496) );
  NAND U2472 ( .A(n1497), .B(n1498), .Z(n316) );
  AND U2473 ( .A(n1499), .B(n1500), .Z(n1498) );
  AND U2474 ( .A(n1501), .B(n1502), .Z(n1500) );
  NAND U2475 ( .A(n1503), .B(n852), .Z(n1502) );
  NAND U2476 ( .A(n1504), .B(n1312), .Z(n1503) );
  NANDN U2477 ( .A(n1505), .B(n1361), .Z(n1504) );
  NAND U2478 ( .A(n1506), .B(n865), .Z(n1501) );
  ANDN U2479 ( .B(n1361), .A(n1507), .Z(n1506) );
  AND U2480 ( .A(n1508), .B(n1509), .Z(n1499) );
  NANDN U2481 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][21] ), .Z(n1509) );
  NAND U2482 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N129 ), .Z(n1508) );
  AND U2483 ( .A(n1510), .B(n1511), .Z(n1497) );
  AND U2484 ( .A(n1512), .B(n1513), .Z(n1511) );
  NANDN U2485 ( .A(n891), .B(\ALU/N129 ), .Z(n1513) );
  NAND U2486 ( .A(n1514), .B(n1026), .Z(n1512) );
  XNOR U2487 ( .A(n1515), .B(n2496), .Z(n1514) );
  AND U2488 ( .A(n1516), .B(n1517), .Z(n1510) );
  NAND U2489 ( .A(n1518), .B(n2496), .Z(n1517) );
  AND U2490 ( .A(n897), .B(b_bus[21]), .Z(n1518) );
  MUX U2491 ( .A(n1022), .B(n1023), .S(n1519), .Z(n1516) );
  NOR U2492 ( .A(b_bus[21]), .B(n2496), .Z(n1519) );
  ANDN U2493 ( .B(reg_source[21]), .A(n1015), .Z(n2496) );
  IV U2494 ( .A(n323), .Z(n1495) );
  NAND U2495 ( .A(n1520), .B(n1521), .Z(n323) );
  AND U2496 ( .A(n1522), .B(n1523), .Z(n1521) );
  AND U2497 ( .A(n1524), .B(n1525), .Z(n1523) );
  NAND U2498 ( .A(n1526), .B(n852), .Z(n1525) );
  NAND U2499 ( .A(n1527), .B(n1312), .Z(n1526) );
  NANDN U2500 ( .A(n1528), .B(n1361), .Z(n1527) );
  NAND U2501 ( .A(n1529), .B(n865), .Z(n1524) );
  ANDN U2502 ( .B(n1361), .A(n1530), .Z(n1529) );
  AND U2503 ( .A(n1531), .B(n1532), .Z(n1522) );
  NANDN U2504 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][20] ), .Z(n1532) );
  NAND U2505 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N128 ), .Z(n1531) );
  AND U2506 ( .A(n1533), .B(n1534), .Z(n1520) );
  AND U2507 ( .A(n1535), .B(n1536), .Z(n1534) );
  NANDN U2508 ( .A(n891), .B(\ALU/N128 ), .Z(n1536) );
  NAND U2509 ( .A(n1537), .B(n1026), .Z(n1535) );
  XNOR U2510 ( .A(n944), .B(n2497), .Z(n1537) );
  AND U2511 ( .A(n1538), .B(n1539), .Z(n1533) );
  NAND U2512 ( .A(n1540), .B(n2497), .Z(n1539) );
  AND U2513 ( .A(n897), .B(b_bus[20]), .Z(n1540) );
  MUX U2514 ( .A(n1022), .B(n1023), .S(n1541), .Z(n1538) );
  NOR U2515 ( .A(b_bus[20]), .B(n2497), .Z(n1541) );
  ANDN U2516 ( .B(reg_source[20]), .A(n1015), .Z(n2497) );
  AND U2517 ( .A(n1542), .B(n1543), .Z(n1493) );
  IV U2518 ( .A(n302), .Z(n1543) );
  NAND U2519 ( .A(n1544), .B(n1545), .Z(n302) );
  AND U2520 ( .A(n1546), .B(n1547), .Z(n1545) );
  AND U2521 ( .A(n1548), .B(n1549), .Z(n1547) );
  NAND U2522 ( .A(n1550), .B(n852), .Z(n1549) );
  NAND U2523 ( .A(n1551), .B(n1312), .Z(n1550) );
  NANDN U2524 ( .A(n1552), .B(n1361), .Z(n1551) );
  NAND U2525 ( .A(n1553), .B(n865), .Z(n1548) );
  ANDN U2526 ( .B(n1361), .A(n1554), .Z(n1553) );
  AND U2527 ( .A(n1555), .B(n1556), .Z(n1546) );
  NANDN U2528 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][23] ), .Z(n1556) );
  NAND U2529 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N131 ), .Z(n1555) );
  AND U2530 ( .A(n1557), .B(n1558), .Z(n1544) );
  AND U2531 ( .A(n1559), .B(n1560), .Z(n1558) );
  NANDN U2532 ( .A(n891), .B(\ALU/N131 ), .Z(n1560) );
  NAND U2533 ( .A(n1561), .B(n1026), .Z(n1559) );
  XNOR U2534 ( .A(n1562), .B(n2494), .Z(n1561) );
  AND U2535 ( .A(n1563), .B(n1564), .Z(n1557) );
  NAND U2536 ( .A(n1565), .B(n2494), .Z(n1564) );
  AND U2537 ( .A(n897), .B(b_bus[23]), .Z(n1565) );
  MUX U2538 ( .A(n1022), .B(n1023), .S(n1566), .Z(n1563) );
  NOR U2539 ( .A(b_bus[23]), .B(n2494), .Z(n1566) );
  ANDN U2540 ( .B(reg_source[23]), .A(n1015), .Z(n2494) );
  IV U2541 ( .A(n309), .Z(n1542) );
  NAND U2542 ( .A(n1567), .B(n1568), .Z(n309) );
  AND U2543 ( .A(n1569), .B(n1570), .Z(n1568) );
  AND U2544 ( .A(n1571), .B(n1572), .Z(n1570) );
  NAND U2545 ( .A(n1573), .B(n852), .Z(n1572) );
  NAND U2546 ( .A(n1574), .B(n1312), .Z(n1573) );
  NANDN U2547 ( .A(n1575), .B(n1361), .Z(n1574) );
  NAND U2548 ( .A(n1576), .B(n865), .Z(n1571) );
  ANDN U2549 ( .B(n1361), .A(n1577), .Z(n1576) );
  AND U2550 ( .A(n1578), .B(n1579), .Z(n1569) );
  NANDN U2551 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][22] ), .Z(n1579) );
  NAND U2552 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N130 ), .Z(n1578) );
  AND U2553 ( .A(n1580), .B(n1581), .Z(n1567) );
  AND U2554 ( .A(n1582), .B(n1583), .Z(n1581) );
  NANDN U2555 ( .A(n891), .B(\ALU/N130 ), .Z(n1583) );
  NAND U2556 ( .A(n1584), .B(n1026), .Z(n1582) );
  XNOR U2557 ( .A(n938), .B(n2495), .Z(n1584) );
  AND U2558 ( .A(n1585), .B(n1586), .Z(n1580) );
  NAND U2559 ( .A(n1587), .B(n2495), .Z(n1586) );
  AND U2560 ( .A(n897), .B(b_bus[22]), .Z(n1587) );
  MUX U2561 ( .A(n1022), .B(n1023), .S(n1588), .Z(n1585) );
  NOR U2562 ( .A(b_bus[22]), .B(n2495), .Z(n1588) );
  ANDN U2563 ( .B(reg_source[22]), .A(n1015), .Z(n2495) );
  AND U2564 ( .A(n1589), .B(n1590), .Z(n1374) );
  AND U2565 ( .A(n1591), .B(n1592), .Z(n1590) );
  AND U2566 ( .A(n1593), .B(n1594), .Z(n1592) );
  IV U2567 ( .A(n288), .Z(n1594) );
  NAND U2568 ( .A(n1595), .B(n1596), .Z(n288) );
  AND U2569 ( .A(n1597), .B(n1598), .Z(n1596) );
  AND U2570 ( .A(n1599), .B(n1600), .Z(n1598) );
  NAND U2571 ( .A(n1601), .B(n852), .Z(n1600) );
  NAND U2572 ( .A(n1602), .B(n1312), .Z(n1601) );
  NANDN U2573 ( .A(n1088), .B(n1361), .Z(n1602) );
  AND U2574 ( .A(n1603), .B(n1604), .Z(n1088) );
  NAND U2575 ( .A(n1252), .B(n1394), .Z(n1604) );
  ANDN U2576 ( .B(n1605), .A(n1606), .Z(n1603) );
  NAND U2577 ( .A(n1398), .B(n1403), .Z(n1605) );
  NAND U2578 ( .A(n1607), .B(n865), .Z(n1599) );
  ANDN U2579 ( .B(n1361), .A(n1095), .Z(n1607) );
  AND U2580 ( .A(n1608), .B(n1609), .Z(n1095) );
  NAND U2581 ( .A(n1360), .B(n1252), .Z(n1609) );
  NAND U2582 ( .A(n1251), .B(n1403), .Z(n1608) );
  AND U2583 ( .A(n1610), .B(n1611), .Z(n1597) );
  NANDN U2584 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][25] ), .Z(n1611) );
  NAND U2585 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N133 ), .Z(n1610) );
  AND U2586 ( .A(n1612), .B(n1613), .Z(n1595) );
  AND U2587 ( .A(n1614), .B(n1615), .Z(n1613) );
  NANDN U2588 ( .A(n891), .B(\ALU/N133 ), .Z(n1615) );
  NAND U2589 ( .A(n1616), .B(n1026), .Z(n1614) );
  XNOR U2590 ( .A(n1617), .B(n2492), .Z(n1616) );
  AND U2591 ( .A(n1618), .B(n1619), .Z(n1612) );
  NAND U2592 ( .A(n1620), .B(n2492), .Z(n1619) );
  AND U2593 ( .A(n897), .B(b_bus[25]), .Z(n1620) );
  MUX U2594 ( .A(n1022), .B(n1023), .S(n1621), .Z(n1618) );
  NOR U2595 ( .A(b_bus[25]), .B(n2492), .Z(n1621) );
  ANDN U2596 ( .B(reg_source[25]), .A(n1015), .Z(n2492) );
  IV U2597 ( .A(n295), .Z(n1593) );
  NAND U2598 ( .A(n1622), .B(n1623), .Z(n295) );
  AND U2599 ( .A(n1624), .B(n1625), .Z(n1623) );
  AND U2600 ( .A(n1626), .B(n1627), .Z(n1625) );
  NAND U2601 ( .A(n1628), .B(n852), .Z(n1627) );
  NAND U2602 ( .A(n1629), .B(n1312), .Z(n1628) );
  NANDN U2603 ( .A(n1123), .B(n1361), .Z(n1629) );
  AND U2604 ( .A(n1630), .B(n1631), .Z(n1123) );
  NAND U2605 ( .A(n1287), .B(n1394), .Z(n1631) );
  ANDN U2606 ( .B(n1632), .A(n1606), .Z(n1630) );
  NAND U2607 ( .A(n1633), .B(n865), .Z(n1626) );
  ANDN U2608 ( .B(n1361), .A(n1130), .Z(n1633) );
  AND U2609 ( .A(n1632), .B(n1634), .Z(n1130) );
  NAND U2610 ( .A(n1360), .B(n1287), .Z(n1634) );
  NAND U2611 ( .A(n1286), .B(n1403), .Z(n1632) );
  AND U2612 ( .A(n1635), .B(n1636), .Z(n1624) );
  NANDN U2613 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][24] ), .Z(n1636) );
  NAND U2614 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N132 ), .Z(n1635) );
  AND U2615 ( .A(n1637), .B(n1638), .Z(n1622) );
  AND U2616 ( .A(n1639), .B(n1640), .Z(n1638) );
  NANDN U2617 ( .A(n891), .B(\ALU/N132 ), .Z(n1640) );
  NAND U2618 ( .A(n1641), .B(n1026), .Z(n1639) );
  XNOR U2619 ( .A(n932), .B(n2493), .Z(n1641) );
  AND U2620 ( .A(n1642), .B(n1643), .Z(n1637) );
  NAND U2621 ( .A(n1644), .B(n2493), .Z(n1643) );
  AND U2622 ( .A(n897), .B(b_bus[24]), .Z(n1644) );
  MUX U2623 ( .A(n1022), .B(n1023), .S(n1645), .Z(n1642) );
  NOR U2624 ( .A(b_bus[24]), .B(n2493), .Z(n1645) );
  ANDN U2625 ( .B(reg_source[24]), .A(n1015), .Z(n2493) );
  AND U2626 ( .A(n1646), .B(n1647), .Z(n1591) );
  IV U2627 ( .A(n274), .Z(n1647) );
  NAND U2628 ( .A(n1648), .B(n1649), .Z(n274) );
  AND U2629 ( .A(n1650), .B(n1651), .Z(n1649) );
  AND U2630 ( .A(n1652), .B(n1653), .Z(n1651) );
  NAND U2631 ( .A(n1654), .B(n852), .Z(n1653) );
  NAND U2632 ( .A(n1655), .B(n1312), .Z(n1654) );
  NAND U2633 ( .A(n1361), .B(n1160), .Z(n1655) );
  NAND U2634 ( .A(n1656), .B(n1657), .Z(n1160) );
  NAND U2635 ( .A(n1316), .B(n1394), .Z(n1656) );
  NAND U2636 ( .A(n1658), .B(n1659), .Z(n1652) );
  AND U2637 ( .A(n1361), .B(n1174), .Z(n1659) );
  AND U2638 ( .A(n865), .B(n1172), .Z(n1658) );
  AND U2639 ( .A(n1660), .B(n1661), .Z(n1650) );
  NANDN U2640 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][27] ), .Z(n1661) );
  NAND U2641 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N135 ), .Z(n1660) );
  AND U2642 ( .A(n1662), .B(n1663), .Z(n1648) );
  AND U2643 ( .A(n1664), .B(n1665), .Z(n1663) );
  NANDN U2644 ( .A(n891), .B(\ALU/N135 ), .Z(n1665) );
  NAND U2645 ( .A(n1666), .B(n1026), .Z(n1664) );
  XNOR U2646 ( .A(n1667), .B(n2490), .Z(n1666) );
  AND U2647 ( .A(n1668), .B(n1669), .Z(n1662) );
  NAND U2648 ( .A(n1670), .B(n2490), .Z(n1669) );
  AND U2649 ( .A(n897), .B(b_bus[27]), .Z(n1670) );
  MUX U2650 ( .A(n1022), .B(n1023), .S(n1671), .Z(n1668) );
  NOR U2651 ( .A(b_bus[27]), .B(n2490), .Z(n1671) );
  ANDN U2652 ( .B(reg_source[27]), .A(n1015), .Z(n2490) );
  IV U2653 ( .A(n281), .Z(n1646) );
  NAND U2654 ( .A(n1672), .B(n1673), .Z(n281) );
  AND U2655 ( .A(n1674), .B(n1675), .Z(n1673) );
  AND U2656 ( .A(n1676), .B(n1677), .Z(n1675) );
  NAND U2657 ( .A(n1678), .B(n852), .Z(n1677) );
  NAND U2658 ( .A(n1679), .B(n1312), .Z(n1678) );
  NANDN U2659 ( .A(n1200), .B(n1361), .Z(n1679) );
  AND U2660 ( .A(n1680), .B(n1681), .Z(n1200) );
  NAND U2661 ( .A(n1362), .B(n1394), .Z(n1681) );
  ANDN U2662 ( .B(n1682), .A(n1606), .Z(n1680) );
  NAND U2663 ( .A(n1683), .B(n1403), .Z(n1682) );
  NAND U2664 ( .A(n1684), .B(n865), .Z(n1676) );
  ANDN U2665 ( .B(n1361), .A(n1208), .Z(n1684) );
  AND U2666 ( .A(n1685), .B(n1686), .Z(n1208) );
  NAND U2667 ( .A(n1360), .B(n1362), .Z(n1686) );
  NAND U2668 ( .A(n1359), .B(n1403), .Z(n1685) );
  AND U2669 ( .A(n1687), .B(n1688), .Z(n1674) );
  NANDN U2670 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][26] ), .Z(n1688) );
  NAND U2671 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N134 ), .Z(n1687) );
  AND U2672 ( .A(n1689), .B(n1690), .Z(n1672) );
  AND U2673 ( .A(n1691), .B(n1692), .Z(n1690) );
  NANDN U2674 ( .A(n891), .B(\ALU/N134 ), .Z(n1692) );
  NAND U2675 ( .A(n1693), .B(n1026), .Z(n1691) );
  XNOR U2676 ( .A(n926), .B(n2491), .Z(n1693) );
  AND U2677 ( .A(n1694), .B(n1695), .Z(n1689) );
  NAND U2678 ( .A(n1696), .B(n2491), .Z(n1695) );
  AND U2679 ( .A(n897), .B(b_bus[26]), .Z(n1696) );
  MUX U2680 ( .A(n1022), .B(n1023), .S(n1697), .Z(n1694) );
  NOR U2681 ( .A(b_bus[26]), .B(n2491), .Z(n1697) );
  ANDN U2682 ( .B(reg_source[26]), .A(n1015), .Z(n2491) );
  AND U2683 ( .A(n1698), .B(n1699), .Z(n1589) );
  AND U2684 ( .A(n1700), .B(n1701), .Z(n1699) );
  IV U2685 ( .A(n260), .Z(n1701) );
  NAND U2686 ( .A(n1702), .B(n1703), .Z(n260) );
  AND U2687 ( .A(n1704), .B(n1705), .Z(n1703) );
  AND U2688 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U2689 ( .A(n1708), .B(n852), .Z(n1707) );
  NAND U2690 ( .A(n1709), .B(n1312), .Z(n1708) );
  NANDN U2691 ( .A(n1241), .B(n1361), .Z(n1709) );
  AND U2692 ( .A(n1710), .B(n1657), .Z(n1241) );
  NAND U2693 ( .A(n1398), .B(n1394), .Z(n1710) );
  NAND U2694 ( .A(n1711), .B(n865), .Z(n1706) );
  AND U2695 ( .A(n1251), .B(n876), .Z(n1711) );
  AND U2696 ( .A(n1712), .B(n1713), .Z(n1704) );
  NANDN U2697 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][29] ), .Z(n1713) );
  NAND U2698 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N137 ), .Z(n1712) );
  AND U2699 ( .A(n1714), .B(n1715), .Z(n1702) );
  AND U2700 ( .A(n1716), .B(n1717), .Z(n1715) );
  NANDN U2701 ( .A(n891), .B(\ALU/N137 ), .Z(n1717) );
  NAND U2702 ( .A(n1718), .B(n1026), .Z(n1716) );
  XNOR U2703 ( .A(n1719), .B(n2488), .Z(n1718) );
  AND U2704 ( .A(n1720), .B(n1721), .Z(n1714) );
  NAND U2705 ( .A(n1722), .B(n2488), .Z(n1721) );
  AND U2706 ( .A(n897), .B(b_bus[29]), .Z(n1722) );
  MUX U2707 ( .A(n1022), .B(n1023), .S(n1723), .Z(n1720) );
  NOR U2708 ( .A(b_bus[29]), .B(n2488), .Z(n1723) );
  ANDN U2709 ( .B(reg_source[29]), .A(n1015), .Z(n2488) );
  IV U2710 ( .A(n267), .Z(n1700) );
  NAND U2711 ( .A(n1724), .B(n1725), .Z(n267) );
  AND U2712 ( .A(n1726), .B(n1727), .Z(n1725) );
  AND U2713 ( .A(n1728), .B(n1729), .Z(n1727) );
  NAND U2714 ( .A(n1730), .B(n852), .Z(n1729) );
  NAND U2715 ( .A(n1731), .B(n1312), .Z(n1730) );
  NANDN U2716 ( .A(n1277), .B(n1361), .Z(n1731) );
  AND U2717 ( .A(n1657), .B(n1732), .Z(n1277) );
  NAND U2718 ( .A(n1286), .B(n1394), .Z(n1732) );
  NAND U2719 ( .A(n1733), .B(n865), .Z(n1728) );
  AND U2720 ( .A(n1286), .B(n876), .Z(n1733) );
  AND U2721 ( .A(n1734), .B(n1735), .Z(n1726) );
  NANDN U2722 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][28] ), .Z(n1735) );
  NAND U2723 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N136 ), .Z(n1734) );
  AND U2724 ( .A(n1736), .B(n1737), .Z(n1724) );
  AND U2725 ( .A(n1738), .B(n1739), .Z(n1737) );
  NANDN U2726 ( .A(n891), .B(\ALU/N136 ), .Z(n1739) );
  NAND U2727 ( .A(n1740), .B(n1026), .Z(n1738) );
  XNOR U2728 ( .A(n920), .B(n2489), .Z(n1740) );
  AND U2729 ( .A(n1741), .B(n1742), .Z(n1736) );
  NAND U2730 ( .A(n1743), .B(n2489), .Z(n1742) );
  AND U2731 ( .A(n897), .B(b_bus[28]), .Z(n1743) );
  MUX U2732 ( .A(n1022), .B(n1023), .S(n1744), .Z(n1741) );
  NOR U2733 ( .A(b_bus[28]), .B(n2489), .Z(n1744) );
  ANDN U2734 ( .B(reg_source[28]), .A(n1015), .Z(n2489) );
  AND U2735 ( .A(n1745), .B(n810), .Z(n1698) );
  IV U2736 ( .A(n243), .Z(n810) );
  IV U2737 ( .A(n253), .Z(n1745) );
  NAND U2738 ( .A(n1746), .B(n1747), .Z(n253) );
  AND U2739 ( .A(n1748), .B(n1749), .Z(n1747) );
  AND U2740 ( .A(n1750), .B(n1751), .Z(n1749) );
  NAND U2741 ( .A(n1752), .B(n852), .Z(n1751) );
  NAND U2742 ( .A(n1753), .B(n1312), .Z(n1752) );
  NANDN U2743 ( .A(n1361), .B(\Shifter/N75 ), .Z(n1312) );
  NANDN U2744 ( .A(n1350), .B(n1361), .Z(n1753) );
  AND U2745 ( .A(n1754), .B(n1657), .Z(n1350) );
  ANDN U2746 ( .B(n1755), .A(n1606), .Z(n1657) );
  NAND U2747 ( .A(\Shifter/N75 ), .B(a_bus[2]), .Z(n1755) );
  NAND U2748 ( .A(n1683), .B(n1394), .Z(n1754) );
  NAND U2749 ( .A(n1756), .B(n865), .Z(n1750) );
  AND U2750 ( .A(n1359), .B(n876), .Z(n1756) );
  AND U2751 ( .A(n1757), .B(n1758), .Z(n1748) );
  NANDN U2752 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][30] ), .Z(n1758) );
  NAND U2753 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N138 ), .Z(n1757) );
  AND U2754 ( .A(n1759), .B(n1760), .Z(n1746) );
  AND U2755 ( .A(n1761), .B(n1762), .Z(n1760) );
  NANDN U2756 ( .A(n891), .B(\ALU/N138 ), .Z(n1762) );
  NAND U2757 ( .A(n1763), .B(n1026), .Z(n1761) );
  XNOR U2758 ( .A(n1764), .B(n2487), .Z(n1763) );
  AND U2759 ( .A(n1765), .B(n1766), .Z(n1759) );
  NAND U2760 ( .A(n1767), .B(n2487), .Z(n1766) );
  AND U2761 ( .A(n897), .B(b_bus[30]), .Z(n1767) );
  MUX U2762 ( .A(n1022), .B(n1023), .S(n1768), .Z(n1765) );
  NOR U2763 ( .A(b_bus[30]), .B(n2487), .Z(n1768) );
  ANDN U2764 ( .B(reg_source[30]), .A(n1015), .Z(n2487) );
  XOR U2765 ( .A(pc_current[31]), .B(\PC_Next/add_30/carry[29] ), .Z(n247) );
  NAND U2766 ( .A(n243), .B(n584), .Z(n788) );
  AND U2767 ( .A(n1769), .B(n7), .Z(n584) );
  OR U2768 ( .A(n795), .B(n89), .Z(n1769) );
  ANDN U2769 ( .B(n10), .A(n1770), .Z(n795) );
  NAND U2770 ( .A(n1771), .B(n1772), .Z(n243) );
  AND U2771 ( .A(n1773), .B(n1774), .Z(n1772) );
  AND U2772 ( .A(n1775), .B(n1776), .Z(n1774) );
  NAND U2773 ( .A(\Shifter/N75 ), .B(n852), .Z(n1776) );
  NAND U2774 ( .A(n1777), .B(n865), .Z(n1775) );
  ANDN U2775 ( .B(n876), .A(n1324), .Z(n1777) );
  AND U2776 ( .A(n1778), .B(n1779), .Z(n1773) );
  NANDN U2777 ( .A(n1408), .B(\Shifter/sll_27/ML_int[5][31] ), .Z(n1779) );
  NAND U2778 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N139 ), .Z(n1778) );
  AND U2779 ( .A(n1780), .B(n1781), .Z(n1771) );
  AND U2780 ( .A(n1782), .B(n1783), .Z(n1781) );
  NANDN U2781 ( .A(n891), .B(\ALU/N139 ), .Z(n1783) );
  NAND U2782 ( .A(n1784), .B(n1026), .Z(n1782) );
  XOR U2783 ( .A(n907), .B(n909), .Z(n1784) );
  AND U2784 ( .A(n1785), .B(n1786), .Z(n1780) );
  NAND U2785 ( .A(n1787), .B(n897), .Z(n1786) );
  AND U2786 ( .A(\Shifter/N75 ), .B(n2486), .Z(n1787) );
  MUX U2787 ( .A(n1022), .B(n1023), .S(n1788), .Z(n1785) );
  AND U2788 ( .A(n909), .B(n907), .Z(n1788) );
  IV U2789 ( .A(n2486), .Z(n909) );
  ANDN U2790 ( .B(reg_source[31]), .A(n1015), .Z(n2486) );
  MUX U2791 ( .A(reg_target[31]), .B(data_mem_out_wire[31]), .S(n1789), .Z(
        \Data_Mem/n6263 ) );
  MUX U2792 ( .A(reg_target[30]), .B(data_mem_out_wire[30]), .S(n1789), .Z(
        \Data_Mem/n6262 ) );
  MUX U2793 ( .A(reg_target[29]), .B(data_mem_out_wire[29]), .S(n1789), .Z(
        \Data_Mem/n6261 ) );
  MUX U2794 ( .A(reg_target[28]), .B(data_mem_out_wire[28]), .S(n1789), .Z(
        \Data_Mem/n6260 ) );
  MUX U2795 ( .A(reg_target[27]), .B(data_mem_out_wire[27]), .S(n1789), .Z(
        \Data_Mem/n6259 ) );
  MUX U2796 ( .A(reg_target[26]), .B(data_mem_out_wire[26]), .S(n1789), .Z(
        \Data_Mem/n6258 ) );
  MUX U2797 ( .A(reg_target[25]), .B(data_mem_out_wire[25]), .S(n1789), .Z(
        \Data_Mem/n6257 ) );
  MUX U2798 ( .A(reg_target[24]), .B(data_mem_out_wire[24]), .S(n1789), .Z(
        \Data_Mem/n6256 ) );
  MUX U2799 ( .A(reg_target[23]), .B(data_mem_out_wire[23]), .S(n1789), .Z(
        \Data_Mem/n6255 ) );
  MUX U2800 ( .A(reg_target[22]), .B(data_mem_out_wire[22]), .S(n1789), .Z(
        \Data_Mem/n6254 ) );
  MUX U2801 ( .A(reg_target[21]), .B(data_mem_out_wire[21]), .S(n1789), .Z(
        \Data_Mem/n6253 ) );
  MUX U2802 ( .A(reg_target[20]), .B(data_mem_out_wire[20]), .S(n1789), .Z(
        \Data_Mem/n6252 ) );
  MUX U2803 ( .A(reg_target[19]), .B(data_mem_out_wire[19]), .S(n1789), .Z(
        \Data_Mem/n6251 ) );
  MUX U2804 ( .A(reg_target[18]), .B(data_mem_out_wire[18]), .S(n1789), .Z(
        \Data_Mem/n6250 ) );
  MUX U2805 ( .A(reg_target[17]), .B(data_mem_out_wire[17]), .S(n1789), .Z(
        \Data_Mem/n6249 ) );
  MUX U2806 ( .A(reg_target[16]), .B(data_mem_out_wire[16]), .S(n1789), .Z(
        \Data_Mem/n6248 ) );
  MUX U2807 ( .A(reg_target[15]), .B(data_mem_out_wire[15]), .S(n1789), .Z(
        \Data_Mem/n6247 ) );
  MUX U2808 ( .A(reg_target[14]), .B(data_mem_out_wire[14]), .S(n1789), .Z(
        \Data_Mem/n6246 ) );
  MUX U2809 ( .A(reg_target[13]), .B(data_mem_out_wire[13]), .S(n1789), .Z(
        \Data_Mem/n6245 ) );
  MUX U2810 ( .A(reg_target[12]), .B(data_mem_out_wire[12]), .S(n1789), .Z(
        \Data_Mem/n6244 ) );
  MUX U2811 ( .A(reg_target[11]), .B(data_mem_out_wire[11]), .S(n1789), .Z(
        \Data_Mem/n6243 ) );
  MUX U2812 ( .A(reg_target[10]), .B(data_mem_out_wire[10]), .S(n1789), .Z(
        \Data_Mem/n6242 ) );
  MUX U2813 ( .A(reg_target[9]), .B(data_mem_out_wire[9]), .S(n1789), .Z(
        \Data_Mem/n6241 ) );
  MUX U2814 ( .A(reg_target[8]), .B(data_mem_out_wire[8]), .S(n1789), .Z(
        \Data_Mem/n6240 ) );
  MUX U2815 ( .A(reg_target[7]), .B(data_mem_out_wire[7]), .S(n1789), .Z(
        \Data_Mem/n6239 ) );
  MUX U2816 ( .A(reg_target[6]), .B(data_mem_out_wire[6]), .S(n1789), .Z(
        \Data_Mem/n6238 ) );
  MUX U2817 ( .A(reg_target[5]), .B(data_mem_out_wire[5]), .S(n1789), .Z(
        \Data_Mem/n6237 ) );
  MUX U2818 ( .A(reg_target[4]), .B(data_mem_out_wire[4]), .S(n1789), .Z(
        \Data_Mem/n6236 ) );
  MUX U2819 ( .A(reg_target[3]), .B(data_mem_out_wire[3]), .S(n1789), .Z(
        \Data_Mem/n6235 ) );
  MUX U2820 ( .A(reg_target[2]), .B(data_mem_out_wire[2]), .S(n1789), .Z(
        \Data_Mem/n6234 ) );
  IV U2821 ( .A(n1790), .Z(n1789) );
  MUX U2822 ( .A(data_mem_out_wire[1]), .B(reg_target[1]), .S(n1790), .Z(
        \Data_Mem/n6233 ) );
  MUX U2823 ( .A(data_mem_out_wire[0]), .B(reg_target[0]), .S(n1790), .Z(
        \Data_Mem/n6232 ) );
  ANDN U2824 ( .B(n1791), .A(n1792), .Z(n1790) );
  MUX U2825 ( .A(reg_target[31]), .B(data_mem_out_wire[63]), .S(n1793), .Z(
        \Data_Mem/n6231 ) );
  MUX U2826 ( .A(reg_target[30]), .B(data_mem_out_wire[62]), .S(n1793), .Z(
        \Data_Mem/n6230 ) );
  MUX U2827 ( .A(reg_target[29]), .B(data_mem_out_wire[61]), .S(n1793), .Z(
        \Data_Mem/n6229 ) );
  MUX U2828 ( .A(reg_target[28]), .B(data_mem_out_wire[60]), .S(n1793), .Z(
        \Data_Mem/n6228 ) );
  MUX U2829 ( .A(reg_target[27]), .B(data_mem_out_wire[59]), .S(n1793), .Z(
        \Data_Mem/n6227 ) );
  MUX U2830 ( .A(reg_target[26]), .B(data_mem_out_wire[58]), .S(n1793), .Z(
        \Data_Mem/n6226 ) );
  MUX U2831 ( .A(reg_target[25]), .B(data_mem_out_wire[57]), .S(n1793), .Z(
        \Data_Mem/n6225 ) );
  MUX U2832 ( .A(reg_target[24]), .B(data_mem_out_wire[56]), .S(n1793), .Z(
        \Data_Mem/n6224 ) );
  MUX U2833 ( .A(reg_target[23]), .B(data_mem_out_wire[55]), .S(n1793), .Z(
        \Data_Mem/n6223 ) );
  MUX U2834 ( .A(reg_target[22]), .B(data_mem_out_wire[54]), .S(n1793), .Z(
        \Data_Mem/n6222 ) );
  MUX U2835 ( .A(reg_target[21]), .B(data_mem_out_wire[53]), .S(n1793), .Z(
        \Data_Mem/n6221 ) );
  MUX U2836 ( .A(reg_target[20]), .B(data_mem_out_wire[52]), .S(n1793), .Z(
        \Data_Mem/n6220 ) );
  MUX U2837 ( .A(reg_target[19]), .B(data_mem_out_wire[51]), .S(n1793), .Z(
        \Data_Mem/n6219 ) );
  MUX U2838 ( .A(reg_target[18]), .B(data_mem_out_wire[50]), .S(n1793), .Z(
        \Data_Mem/n6218 ) );
  MUX U2839 ( .A(reg_target[17]), .B(data_mem_out_wire[49]), .S(n1793), .Z(
        \Data_Mem/n6217 ) );
  MUX U2840 ( .A(reg_target[16]), .B(data_mem_out_wire[48]), .S(n1793), .Z(
        \Data_Mem/n6216 ) );
  MUX U2841 ( .A(reg_target[15]), .B(data_mem_out_wire[47]), .S(n1793), .Z(
        \Data_Mem/n6215 ) );
  MUX U2842 ( .A(reg_target[14]), .B(data_mem_out_wire[46]), .S(n1793), .Z(
        \Data_Mem/n6214 ) );
  MUX U2843 ( .A(reg_target[13]), .B(data_mem_out_wire[45]), .S(n1793), .Z(
        \Data_Mem/n6213 ) );
  MUX U2844 ( .A(reg_target[12]), .B(data_mem_out_wire[44]), .S(n1793), .Z(
        \Data_Mem/n6212 ) );
  MUX U2845 ( .A(reg_target[11]), .B(data_mem_out_wire[43]), .S(n1793), .Z(
        \Data_Mem/n6211 ) );
  MUX U2846 ( .A(reg_target[10]), .B(data_mem_out_wire[42]), .S(n1793), .Z(
        \Data_Mem/n6210 ) );
  MUX U2847 ( .A(reg_target[9]), .B(data_mem_out_wire[41]), .S(n1793), .Z(
        \Data_Mem/n6209 ) );
  MUX U2848 ( .A(reg_target[8]), .B(data_mem_out_wire[40]), .S(n1793), .Z(
        \Data_Mem/n6208 ) );
  MUX U2849 ( .A(reg_target[7]), .B(data_mem_out_wire[39]), .S(n1793), .Z(
        \Data_Mem/n6207 ) );
  MUX U2850 ( .A(reg_target[6]), .B(data_mem_out_wire[38]), .S(n1793), .Z(
        \Data_Mem/n6206 ) );
  MUX U2851 ( .A(reg_target[5]), .B(data_mem_out_wire[37]), .S(n1793), .Z(
        \Data_Mem/n6205 ) );
  MUX U2852 ( .A(reg_target[4]), .B(data_mem_out_wire[36]), .S(n1793), .Z(
        \Data_Mem/n6204 ) );
  MUX U2853 ( .A(reg_target[3]), .B(data_mem_out_wire[35]), .S(n1793), .Z(
        \Data_Mem/n6203 ) );
  MUX U2854 ( .A(reg_target[2]), .B(data_mem_out_wire[34]), .S(n1793), .Z(
        \Data_Mem/n6202 ) );
  IV U2855 ( .A(n1794), .Z(n1793) );
  MUX U2856 ( .A(data_mem_out_wire[33]), .B(reg_target[1]), .S(n1794), .Z(
        \Data_Mem/n6201 ) );
  MUX U2857 ( .A(data_mem_out_wire[32]), .B(reg_target[0]), .S(n1794), .Z(
        \Data_Mem/n6200 ) );
  ANDN U2858 ( .B(n1795), .A(n1792), .Z(n1794) );
  MUX U2859 ( .A(reg_target[31]), .B(data_mem_out_wire[95]), .S(n1796), .Z(
        \Data_Mem/n6199 ) );
  MUX U2860 ( .A(reg_target[30]), .B(data_mem_out_wire[94]), .S(n1796), .Z(
        \Data_Mem/n6198 ) );
  MUX U2861 ( .A(reg_target[29]), .B(data_mem_out_wire[93]), .S(n1796), .Z(
        \Data_Mem/n6197 ) );
  MUX U2862 ( .A(reg_target[28]), .B(data_mem_out_wire[92]), .S(n1796), .Z(
        \Data_Mem/n6196 ) );
  MUX U2863 ( .A(reg_target[27]), .B(data_mem_out_wire[91]), .S(n1796), .Z(
        \Data_Mem/n6195 ) );
  MUX U2864 ( .A(reg_target[26]), .B(data_mem_out_wire[90]), .S(n1796), .Z(
        \Data_Mem/n6194 ) );
  MUX U2865 ( .A(reg_target[25]), .B(data_mem_out_wire[89]), .S(n1796), .Z(
        \Data_Mem/n6193 ) );
  MUX U2866 ( .A(reg_target[24]), .B(data_mem_out_wire[88]), .S(n1796), .Z(
        \Data_Mem/n6192 ) );
  MUX U2867 ( .A(reg_target[23]), .B(data_mem_out_wire[87]), .S(n1796), .Z(
        \Data_Mem/n6191 ) );
  MUX U2868 ( .A(reg_target[22]), .B(data_mem_out_wire[86]), .S(n1796), .Z(
        \Data_Mem/n6190 ) );
  MUX U2869 ( .A(reg_target[21]), .B(data_mem_out_wire[85]), .S(n1796), .Z(
        \Data_Mem/n6189 ) );
  MUX U2870 ( .A(reg_target[20]), .B(data_mem_out_wire[84]), .S(n1796), .Z(
        \Data_Mem/n6188 ) );
  MUX U2871 ( .A(reg_target[19]), .B(data_mem_out_wire[83]), .S(n1796), .Z(
        \Data_Mem/n6187 ) );
  MUX U2872 ( .A(reg_target[18]), .B(data_mem_out_wire[82]), .S(n1796), .Z(
        \Data_Mem/n6186 ) );
  MUX U2873 ( .A(reg_target[17]), .B(data_mem_out_wire[81]), .S(n1796), .Z(
        \Data_Mem/n6185 ) );
  MUX U2874 ( .A(reg_target[16]), .B(data_mem_out_wire[80]), .S(n1796), .Z(
        \Data_Mem/n6184 ) );
  MUX U2875 ( .A(reg_target[15]), .B(data_mem_out_wire[79]), .S(n1796), .Z(
        \Data_Mem/n6183 ) );
  MUX U2876 ( .A(reg_target[14]), .B(data_mem_out_wire[78]), .S(n1796), .Z(
        \Data_Mem/n6182 ) );
  MUX U2877 ( .A(reg_target[13]), .B(data_mem_out_wire[77]), .S(n1796), .Z(
        \Data_Mem/n6181 ) );
  MUX U2878 ( .A(reg_target[12]), .B(data_mem_out_wire[76]), .S(n1796), .Z(
        \Data_Mem/n6180 ) );
  MUX U2879 ( .A(reg_target[11]), .B(data_mem_out_wire[75]), .S(n1796), .Z(
        \Data_Mem/n6179 ) );
  MUX U2880 ( .A(reg_target[10]), .B(data_mem_out_wire[74]), .S(n1796), .Z(
        \Data_Mem/n6178 ) );
  MUX U2881 ( .A(reg_target[9]), .B(data_mem_out_wire[73]), .S(n1796), .Z(
        \Data_Mem/n6177 ) );
  MUX U2882 ( .A(reg_target[8]), .B(data_mem_out_wire[72]), .S(n1796), .Z(
        \Data_Mem/n6176 ) );
  MUX U2883 ( .A(reg_target[7]), .B(data_mem_out_wire[71]), .S(n1796), .Z(
        \Data_Mem/n6175 ) );
  MUX U2884 ( .A(reg_target[6]), .B(data_mem_out_wire[70]), .S(n1796), .Z(
        \Data_Mem/n6174 ) );
  MUX U2885 ( .A(reg_target[5]), .B(data_mem_out_wire[69]), .S(n1796), .Z(
        \Data_Mem/n6173 ) );
  MUX U2886 ( .A(reg_target[4]), .B(data_mem_out_wire[68]), .S(n1796), .Z(
        \Data_Mem/n6172 ) );
  MUX U2887 ( .A(reg_target[3]), .B(data_mem_out_wire[67]), .S(n1796), .Z(
        \Data_Mem/n6171 ) );
  MUX U2888 ( .A(reg_target[2]), .B(data_mem_out_wire[66]), .S(n1796), .Z(
        \Data_Mem/n6170 ) );
  IV U2889 ( .A(n1797), .Z(n1796) );
  MUX U2890 ( .A(data_mem_out_wire[65]), .B(reg_target[1]), .S(n1797), .Z(
        \Data_Mem/n6169 ) );
  MUX U2891 ( .A(data_mem_out_wire[64]), .B(reg_target[0]), .S(n1797), .Z(
        \Data_Mem/n6168 ) );
  ANDN U2892 ( .B(n1798), .A(n1792), .Z(n1797) );
  MUX U2893 ( .A(reg_target[31]), .B(data_mem_out_wire[127]), .S(n1799), .Z(
        \Data_Mem/n6167 ) );
  MUX U2894 ( .A(reg_target[30]), .B(data_mem_out_wire[126]), .S(n1799), .Z(
        \Data_Mem/n6166 ) );
  MUX U2895 ( .A(reg_target[29]), .B(data_mem_out_wire[125]), .S(n1799), .Z(
        \Data_Mem/n6165 ) );
  MUX U2896 ( .A(reg_target[28]), .B(data_mem_out_wire[124]), .S(n1799), .Z(
        \Data_Mem/n6164 ) );
  MUX U2897 ( .A(reg_target[27]), .B(data_mem_out_wire[123]), .S(n1799), .Z(
        \Data_Mem/n6163 ) );
  MUX U2898 ( .A(reg_target[26]), .B(data_mem_out_wire[122]), .S(n1799), .Z(
        \Data_Mem/n6162 ) );
  MUX U2899 ( .A(reg_target[25]), .B(data_mem_out_wire[121]), .S(n1799), .Z(
        \Data_Mem/n6161 ) );
  MUX U2900 ( .A(reg_target[24]), .B(data_mem_out_wire[120]), .S(n1799), .Z(
        \Data_Mem/n6160 ) );
  MUX U2901 ( .A(reg_target[23]), .B(data_mem_out_wire[119]), .S(n1799), .Z(
        \Data_Mem/n6159 ) );
  MUX U2902 ( .A(reg_target[22]), .B(data_mem_out_wire[118]), .S(n1799), .Z(
        \Data_Mem/n6158 ) );
  MUX U2903 ( .A(reg_target[21]), .B(data_mem_out_wire[117]), .S(n1799), .Z(
        \Data_Mem/n6157 ) );
  MUX U2904 ( .A(reg_target[20]), .B(data_mem_out_wire[116]), .S(n1799), .Z(
        \Data_Mem/n6156 ) );
  MUX U2905 ( .A(reg_target[19]), .B(data_mem_out_wire[115]), .S(n1799), .Z(
        \Data_Mem/n6155 ) );
  MUX U2906 ( .A(reg_target[18]), .B(data_mem_out_wire[114]), .S(n1799), .Z(
        \Data_Mem/n6154 ) );
  MUX U2907 ( .A(reg_target[17]), .B(data_mem_out_wire[113]), .S(n1799), .Z(
        \Data_Mem/n6153 ) );
  MUX U2908 ( .A(reg_target[16]), .B(data_mem_out_wire[112]), .S(n1799), .Z(
        \Data_Mem/n6152 ) );
  MUX U2909 ( .A(reg_target[15]), .B(data_mem_out_wire[111]), .S(n1799), .Z(
        \Data_Mem/n6151 ) );
  MUX U2910 ( .A(reg_target[14]), .B(data_mem_out_wire[110]), .S(n1799), .Z(
        \Data_Mem/n6150 ) );
  MUX U2911 ( .A(reg_target[13]), .B(data_mem_out_wire[109]), .S(n1799), .Z(
        \Data_Mem/n6149 ) );
  MUX U2912 ( .A(reg_target[12]), .B(data_mem_out_wire[108]), .S(n1799), .Z(
        \Data_Mem/n6148 ) );
  MUX U2913 ( .A(reg_target[11]), .B(data_mem_out_wire[107]), .S(n1799), .Z(
        \Data_Mem/n6147 ) );
  MUX U2914 ( .A(reg_target[10]), .B(data_mem_out_wire[106]), .S(n1799), .Z(
        \Data_Mem/n6146 ) );
  MUX U2915 ( .A(reg_target[9]), .B(data_mem_out_wire[105]), .S(n1799), .Z(
        \Data_Mem/n6145 ) );
  MUX U2916 ( .A(reg_target[8]), .B(data_mem_out_wire[104]), .S(n1799), .Z(
        \Data_Mem/n6144 ) );
  MUX U2917 ( .A(reg_target[7]), .B(data_mem_out_wire[103]), .S(n1799), .Z(
        \Data_Mem/n6143 ) );
  MUX U2918 ( .A(reg_target[6]), .B(data_mem_out_wire[102]), .S(n1799), .Z(
        \Data_Mem/n6142 ) );
  MUX U2919 ( .A(reg_target[5]), .B(data_mem_out_wire[101]), .S(n1799), .Z(
        \Data_Mem/n6141 ) );
  MUX U2920 ( .A(reg_target[4]), .B(data_mem_out_wire[100]), .S(n1799), .Z(
        \Data_Mem/n6140 ) );
  MUX U2921 ( .A(reg_target[3]), .B(data_mem_out_wire[99]), .S(n1799), .Z(
        \Data_Mem/n6139 ) );
  MUX U2922 ( .A(reg_target[2]), .B(data_mem_out_wire[98]), .S(n1799), .Z(
        \Data_Mem/n6138 ) );
  IV U2923 ( .A(n1800), .Z(n1799) );
  MUX U2924 ( .A(data_mem_out_wire[97]), .B(reg_target[1]), .S(n1800), .Z(
        \Data_Mem/n6137 ) );
  MUX U2925 ( .A(data_mem_out_wire[96]), .B(reg_target[0]), .S(n1800), .Z(
        \Data_Mem/n6136 ) );
  ANDN U2926 ( .B(n1801), .A(n1792), .Z(n1800) );
  MUX U2927 ( .A(reg_target[31]), .B(data_mem_out_wire[159]), .S(n1802), .Z(
        \Data_Mem/n6135 ) );
  MUX U2928 ( .A(reg_target[30]), .B(data_mem_out_wire[158]), .S(n1802), .Z(
        \Data_Mem/n6134 ) );
  MUX U2929 ( .A(reg_target[29]), .B(data_mem_out_wire[157]), .S(n1802), .Z(
        \Data_Mem/n6133 ) );
  MUX U2930 ( .A(reg_target[28]), .B(data_mem_out_wire[156]), .S(n1802), .Z(
        \Data_Mem/n6132 ) );
  MUX U2931 ( .A(reg_target[27]), .B(data_mem_out_wire[155]), .S(n1802), .Z(
        \Data_Mem/n6131 ) );
  MUX U2932 ( .A(reg_target[26]), .B(data_mem_out_wire[154]), .S(n1802), .Z(
        \Data_Mem/n6130 ) );
  MUX U2933 ( .A(reg_target[25]), .B(data_mem_out_wire[153]), .S(n1802), .Z(
        \Data_Mem/n6129 ) );
  MUX U2934 ( .A(reg_target[24]), .B(data_mem_out_wire[152]), .S(n1802), .Z(
        \Data_Mem/n6128 ) );
  MUX U2935 ( .A(reg_target[23]), .B(data_mem_out_wire[151]), .S(n1802), .Z(
        \Data_Mem/n6127 ) );
  MUX U2936 ( .A(reg_target[22]), .B(data_mem_out_wire[150]), .S(n1802), .Z(
        \Data_Mem/n6126 ) );
  MUX U2937 ( .A(reg_target[21]), .B(data_mem_out_wire[149]), .S(n1802), .Z(
        \Data_Mem/n6125 ) );
  MUX U2938 ( .A(reg_target[20]), .B(data_mem_out_wire[148]), .S(n1802), .Z(
        \Data_Mem/n6124 ) );
  MUX U2939 ( .A(reg_target[19]), .B(data_mem_out_wire[147]), .S(n1802), .Z(
        \Data_Mem/n6123 ) );
  MUX U2940 ( .A(reg_target[18]), .B(data_mem_out_wire[146]), .S(n1802), .Z(
        \Data_Mem/n6122 ) );
  MUX U2941 ( .A(reg_target[17]), .B(data_mem_out_wire[145]), .S(n1802), .Z(
        \Data_Mem/n6121 ) );
  MUX U2942 ( .A(reg_target[16]), .B(data_mem_out_wire[144]), .S(n1802), .Z(
        \Data_Mem/n6120 ) );
  MUX U2943 ( .A(reg_target[15]), .B(data_mem_out_wire[143]), .S(n1802), .Z(
        \Data_Mem/n6119 ) );
  MUX U2944 ( .A(reg_target[14]), .B(data_mem_out_wire[142]), .S(n1802), .Z(
        \Data_Mem/n6118 ) );
  MUX U2945 ( .A(reg_target[13]), .B(data_mem_out_wire[141]), .S(n1802), .Z(
        \Data_Mem/n6117 ) );
  MUX U2946 ( .A(reg_target[12]), .B(data_mem_out_wire[140]), .S(n1802), .Z(
        \Data_Mem/n6116 ) );
  MUX U2947 ( .A(reg_target[11]), .B(data_mem_out_wire[139]), .S(n1802), .Z(
        \Data_Mem/n6115 ) );
  MUX U2948 ( .A(reg_target[10]), .B(data_mem_out_wire[138]), .S(n1802), .Z(
        \Data_Mem/n6114 ) );
  MUX U2949 ( .A(reg_target[9]), .B(data_mem_out_wire[137]), .S(n1802), .Z(
        \Data_Mem/n6113 ) );
  MUX U2950 ( .A(reg_target[8]), .B(data_mem_out_wire[136]), .S(n1802), .Z(
        \Data_Mem/n6112 ) );
  MUX U2951 ( .A(reg_target[7]), .B(data_mem_out_wire[135]), .S(n1802), .Z(
        \Data_Mem/n6111 ) );
  MUX U2952 ( .A(reg_target[6]), .B(data_mem_out_wire[134]), .S(n1802), .Z(
        \Data_Mem/n6110 ) );
  MUX U2953 ( .A(reg_target[5]), .B(data_mem_out_wire[133]), .S(n1802), .Z(
        \Data_Mem/n6109 ) );
  MUX U2954 ( .A(reg_target[4]), .B(data_mem_out_wire[132]), .S(n1802), .Z(
        \Data_Mem/n6108 ) );
  MUX U2955 ( .A(reg_target[3]), .B(data_mem_out_wire[131]), .S(n1802), .Z(
        \Data_Mem/n6107 ) );
  MUX U2956 ( .A(reg_target[2]), .B(data_mem_out_wire[130]), .S(n1802), .Z(
        \Data_Mem/n6106 ) );
  IV U2957 ( .A(n1803), .Z(n1802) );
  MUX U2958 ( .A(data_mem_out_wire[129]), .B(reg_target[1]), .S(n1803), .Z(
        \Data_Mem/n6105 ) );
  MUX U2959 ( .A(data_mem_out_wire[128]), .B(reg_target[0]), .S(n1803), .Z(
        \Data_Mem/n6104 ) );
  ANDN U2960 ( .B(n1804), .A(n1792), .Z(n1803) );
  MUX U2961 ( .A(reg_target[31]), .B(data_mem_out_wire[191]), .S(n1805), .Z(
        \Data_Mem/n6103 ) );
  MUX U2962 ( .A(reg_target[30]), .B(data_mem_out_wire[190]), .S(n1805), .Z(
        \Data_Mem/n6102 ) );
  MUX U2963 ( .A(reg_target[29]), .B(data_mem_out_wire[189]), .S(n1805), .Z(
        \Data_Mem/n6101 ) );
  MUX U2964 ( .A(reg_target[28]), .B(data_mem_out_wire[188]), .S(n1805), .Z(
        \Data_Mem/n6100 ) );
  MUX U2965 ( .A(reg_target[27]), .B(data_mem_out_wire[187]), .S(n1805), .Z(
        \Data_Mem/n6099 ) );
  MUX U2966 ( .A(reg_target[26]), .B(data_mem_out_wire[186]), .S(n1805), .Z(
        \Data_Mem/n6098 ) );
  MUX U2967 ( .A(reg_target[25]), .B(data_mem_out_wire[185]), .S(n1805), .Z(
        \Data_Mem/n6097 ) );
  MUX U2968 ( .A(reg_target[24]), .B(data_mem_out_wire[184]), .S(n1805), .Z(
        \Data_Mem/n6096 ) );
  MUX U2969 ( .A(reg_target[23]), .B(data_mem_out_wire[183]), .S(n1805), .Z(
        \Data_Mem/n6095 ) );
  MUX U2970 ( .A(reg_target[22]), .B(data_mem_out_wire[182]), .S(n1805), .Z(
        \Data_Mem/n6094 ) );
  MUX U2971 ( .A(reg_target[21]), .B(data_mem_out_wire[181]), .S(n1805), .Z(
        \Data_Mem/n6093 ) );
  MUX U2972 ( .A(reg_target[20]), .B(data_mem_out_wire[180]), .S(n1805), .Z(
        \Data_Mem/n6092 ) );
  MUX U2973 ( .A(reg_target[19]), .B(data_mem_out_wire[179]), .S(n1805), .Z(
        \Data_Mem/n6091 ) );
  MUX U2974 ( .A(reg_target[18]), .B(data_mem_out_wire[178]), .S(n1805), .Z(
        \Data_Mem/n6090 ) );
  MUX U2975 ( .A(reg_target[17]), .B(data_mem_out_wire[177]), .S(n1805), .Z(
        \Data_Mem/n6089 ) );
  MUX U2976 ( .A(reg_target[16]), .B(data_mem_out_wire[176]), .S(n1805), .Z(
        \Data_Mem/n6088 ) );
  MUX U2977 ( .A(reg_target[15]), .B(data_mem_out_wire[175]), .S(n1805), .Z(
        \Data_Mem/n6087 ) );
  MUX U2978 ( .A(reg_target[14]), .B(data_mem_out_wire[174]), .S(n1805), .Z(
        \Data_Mem/n6086 ) );
  MUX U2979 ( .A(reg_target[13]), .B(data_mem_out_wire[173]), .S(n1805), .Z(
        \Data_Mem/n6085 ) );
  MUX U2980 ( .A(reg_target[12]), .B(data_mem_out_wire[172]), .S(n1805), .Z(
        \Data_Mem/n6084 ) );
  MUX U2981 ( .A(reg_target[11]), .B(data_mem_out_wire[171]), .S(n1805), .Z(
        \Data_Mem/n6083 ) );
  MUX U2982 ( .A(reg_target[10]), .B(data_mem_out_wire[170]), .S(n1805), .Z(
        \Data_Mem/n6082 ) );
  MUX U2983 ( .A(reg_target[9]), .B(data_mem_out_wire[169]), .S(n1805), .Z(
        \Data_Mem/n6081 ) );
  MUX U2984 ( .A(reg_target[8]), .B(data_mem_out_wire[168]), .S(n1805), .Z(
        \Data_Mem/n6080 ) );
  MUX U2985 ( .A(reg_target[7]), .B(data_mem_out_wire[167]), .S(n1805), .Z(
        \Data_Mem/n6079 ) );
  MUX U2986 ( .A(reg_target[6]), .B(data_mem_out_wire[166]), .S(n1805), .Z(
        \Data_Mem/n6078 ) );
  MUX U2987 ( .A(reg_target[5]), .B(data_mem_out_wire[165]), .S(n1805), .Z(
        \Data_Mem/n6077 ) );
  MUX U2988 ( .A(reg_target[4]), .B(data_mem_out_wire[164]), .S(n1805), .Z(
        \Data_Mem/n6076 ) );
  MUX U2989 ( .A(reg_target[3]), .B(data_mem_out_wire[163]), .S(n1805), .Z(
        \Data_Mem/n6075 ) );
  MUX U2990 ( .A(reg_target[2]), .B(data_mem_out_wire[162]), .S(n1805), .Z(
        \Data_Mem/n6074 ) );
  IV U2991 ( .A(n1806), .Z(n1805) );
  MUX U2992 ( .A(data_mem_out_wire[161]), .B(reg_target[1]), .S(n1806), .Z(
        \Data_Mem/n6073 ) );
  MUX U2993 ( .A(data_mem_out_wire[160]), .B(reg_target[0]), .S(n1806), .Z(
        \Data_Mem/n6072 ) );
  ANDN U2994 ( .B(n1807), .A(n1792), .Z(n1806) );
  MUX U2995 ( .A(reg_target[31]), .B(data_mem_out_wire[223]), .S(n1808), .Z(
        \Data_Mem/n6071 ) );
  MUX U2996 ( .A(reg_target[30]), .B(data_mem_out_wire[222]), .S(n1808), .Z(
        \Data_Mem/n6070 ) );
  MUX U2997 ( .A(reg_target[29]), .B(data_mem_out_wire[221]), .S(n1808), .Z(
        \Data_Mem/n6069 ) );
  MUX U2998 ( .A(reg_target[28]), .B(data_mem_out_wire[220]), .S(n1808), .Z(
        \Data_Mem/n6068 ) );
  MUX U2999 ( .A(reg_target[27]), .B(data_mem_out_wire[219]), .S(n1808), .Z(
        \Data_Mem/n6067 ) );
  MUX U3000 ( .A(reg_target[26]), .B(data_mem_out_wire[218]), .S(n1808), .Z(
        \Data_Mem/n6066 ) );
  MUX U3001 ( .A(reg_target[25]), .B(data_mem_out_wire[217]), .S(n1808), .Z(
        \Data_Mem/n6065 ) );
  MUX U3002 ( .A(reg_target[24]), .B(data_mem_out_wire[216]), .S(n1808), .Z(
        \Data_Mem/n6064 ) );
  MUX U3003 ( .A(reg_target[23]), .B(data_mem_out_wire[215]), .S(n1808), .Z(
        \Data_Mem/n6063 ) );
  MUX U3004 ( .A(reg_target[22]), .B(data_mem_out_wire[214]), .S(n1808), .Z(
        \Data_Mem/n6062 ) );
  MUX U3005 ( .A(reg_target[21]), .B(data_mem_out_wire[213]), .S(n1808), .Z(
        \Data_Mem/n6061 ) );
  MUX U3006 ( .A(reg_target[20]), .B(data_mem_out_wire[212]), .S(n1808), .Z(
        \Data_Mem/n6060 ) );
  MUX U3007 ( .A(reg_target[19]), .B(data_mem_out_wire[211]), .S(n1808), .Z(
        \Data_Mem/n6059 ) );
  MUX U3008 ( .A(reg_target[18]), .B(data_mem_out_wire[210]), .S(n1808), .Z(
        \Data_Mem/n6058 ) );
  MUX U3009 ( .A(reg_target[17]), .B(data_mem_out_wire[209]), .S(n1808), .Z(
        \Data_Mem/n6057 ) );
  MUX U3010 ( .A(reg_target[16]), .B(data_mem_out_wire[208]), .S(n1808), .Z(
        \Data_Mem/n6056 ) );
  MUX U3011 ( .A(reg_target[15]), .B(data_mem_out_wire[207]), .S(n1808), .Z(
        \Data_Mem/n6055 ) );
  MUX U3012 ( .A(reg_target[14]), .B(data_mem_out_wire[206]), .S(n1808), .Z(
        \Data_Mem/n6054 ) );
  MUX U3013 ( .A(reg_target[13]), .B(data_mem_out_wire[205]), .S(n1808), .Z(
        \Data_Mem/n6053 ) );
  MUX U3014 ( .A(reg_target[12]), .B(data_mem_out_wire[204]), .S(n1808), .Z(
        \Data_Mem/n6052 ) );
  MUX U3015 ( .A(reg_target[11]), .B(data_mem_out_wire[203]), .S(n1808), .Z(
        \Data_Mem/n6051 ) );
  MUX U3016 ( .A(reg_target[10]), .B(data_mem_out_wire[202]), .S(n1808), .Z(
        \Data_Mem/n6050 ) );
  MUX U3017 ( .A(reg_target[9]), .B(data_mem_out_wire[201]), .S(n1808), .Z(
        \Data_Mem/n6049 ) );
  MUX U3018 ( .A(reg_target[8]), .B(data_mem_out_wire[200]), .S(n1808), .Z(
        \Data_Mem/n6048 ) );
  MUX U3019 ( .A(reg_target[7]), .B(data_mem_out_wire[199]), .S(n1808), .Z(
        \Data_Mem/n6047 ) );
  MUX U3020 ( .A(reg_target[6]), .B(data_mem_out_wire[198]), .S(n1808), .Z(
        \Data_Mem/n6046 ) );
  MUX U3021 ( .A(reg_target[5]), .B(data_mem_out_wire[197]), .S(n1808), .Z(
        \Data_Mem/n6045 ) );
  MUX U3022 ( .A(reg_target[4]), .B(data_mem_out_wire[196]), .S(n1808), .Z(
        \Data_Mem/n6044 ) );
  MUX U3023 ( .A(reg_target[3]), .B(data_mem_out_wire[195]), .S(n1808), .Z(
        \Data_Mem/n6043 ) );
  MUX U3024 ( .A(reg_target[2]), .B(data_mem_out_wire[194]), .S(n1808), .Z(
        \Data_Mem/n6042 ) );
  IV U3025 ( .A(n1809), .Z(n1808) );
  MUX U3026 ( .A(data_mem_out_wire[193]), .B(reg_target[1]), .S(n1809), .Z(
        \Data_Mem/n6041 ) );
  MUX U3027 ( .A(data_mem_out_wire[192]), .B(reg_target[0]), .S(n1809), .Z(
        \Data_Mem/n6040 ) );
  ANDN U3028 ( .B(n1810), .A(n1792), .Z(n1809) );
  MUX U3029 ( .A(data_mem_out_wire[255]), .B(reg_target[31]), .S(n1811), .Z(
        \Data_Mem/n6039 ) );
  MUX U3030 ( .A(data_mem_out_wire[254]), .B(reg_target[30]), .S(n1811), .Z(
        \Data_Mem/n6038 ) );
  MUX U3031 ( .A(data_mem_out_wire[253]), .B(reg_target[29]), .S(n1811), .Z(
        \Data_Mem/n6037 ) );
  MUX U3032 ( .A(data_mem_out_wire[252]), .B(reg_target[28]), .S(n1811), .Z(
        \Data_Mem/n6036 ) );
  MUX U3033 ( .A(data_mem_out_wire[251]), .B(reg_target[27]), .S(n1811), .Z(
        \Data_Mem/n6035 ) );
  MUX U3034 ( .A(data_mem_out_wire[250]), .B(reg_target[26]), .S(n1811), .Z(
        \Data_Mem/n6034 ) );
  MUX U3035 ( .A(data_mem_out_wire[249]), .B(reg_target[25]), .S(n1811), .Z(
        \Data_Mem/n6033 ) );
  MUX U3036 ( .A(data_mem_out_wire[248]), .B(reg_target[24]), .S(n1811), .Z(
        \Data_Mem/n6032 ) );
  MUX U3037 ( .A(data_mem_out_wire[247]), .B(reg_target[23]), .S(n1811), .Z(
        \Data_Mem/n6031 ) );
  MUX U3038 ( .A(data_mem_out_wire[246]), .B(reg_target[22]), .S(n1811), .Z(
        \Data_Mem/n6030 ) );
  MUX U3039 ( .A(data_mem_out_wire[245]), .B(reg_target[21]), .S(n1811), .Z(
        \Data_Mem/n6029 ) );
  MUX U3040 ( .A(data_mem_out_wire[244]), .B(reg_target[20]), .S(n1811), .Z(
        \Data_Mem/n6028 ) );
  MUX U3041 ( .A(data_mem_out_wire[243]), .B(reg_target[19]), .S(n1811), .Z(
        \Data_Mem/n6027 ) );
  MUX U3042 ( .A(data_mem_out_wire[242]), .B(reg_target[18]), .S(n1811), .Z(
        \Data_Mem/n6026 ) );
  MUX U3043 ( .A(data_mem_out_wire[241]), .B(reg_target[17]), .S(n1811), .Z(
        \Data_Mem/n6025 ) );
  MUX U3044 ( .A(data_mem_out_wire[240]), .B(reg_target[16]), .S(n1811), .Z(
        \Data_Mem/n6024 ) );
  MUX U3045 ( .A(data_mem_out_wire[239]), .B(reg_target[15]), .S(n1811), .Z(
        \Data_Mem/n6023 ) );
  MUX U3046 ( .A(data_mem_out_wire[238]), .B(reg_target[14]), .S(n1811), .Z(
        \Data_Mem/n6022 ) );
  MUX U3047 ( .A(data_mem_out_wire[237]), .B(reg_target[13]), .S(n1811), .Z(
        \Data_Mem/n6021 ) );
  MUX U3048 ( .A(data_mem_out_wire[236]), .B(reg_target[12]), .S(n1811), .Z(
        \Data_Mem/n6020 ) );
  MUX U3049 ( .A(data_mem_out_wire[235]), .B(reg_target[11]), .S(n1811), .Z(
        \Data_Mem/n6019 ) );
  MUX U3050 ( .A(data_mem_out_wire[234]), .B(reg_target[10]), .S(n1811), .Z(
        \Data_Mem/n6018 ) );
  MUX U3051 ( .A(data_mem_out_wire[233]), .B(reg_target[9]), .S(n1811), .Z(
        \Data_Mem/n6017 ) );
  MUX U3052 ( .A(data_mem_out_wire[232]), .B(reg_target[8]), .S(n1811), .Z(
        \Data_Mem/n6016 ) );
  MUX U3053 ( .A(data_mem_out_wire[231]), .B(reg_target[7]), .S(n1811), .Z(
        \Data_Mem/n6015 ) );
  MUX U3054 ( .A(data_mem_out_wire[230]), .B(reg_target[6]), .S(n1811), .Z(
        \Data_Mem/n6014 ) );
  MUX U3055 ( .A(data_mem_out_wire[229]), .B(reg_target[5]), .S(n1811), .Z(
        \Data_Mem/n6013 ) );
  MUX U3056 ( .A(data_mem_out_wire[228]), .B(reg_target[4]), .S(n1811), .Z(
        \Data_Mem/n6012 ) );
  MUX U3057 ( .A(data_mem_out_wire[227]), .B(reg_target[3]), .S(n1811), .Z(
        \Data_Mem/n6011 ) );
  MUX U3058 ( .A(data_mem_out_wire[226]), .B(reg_target[2]), .S(n1811), .Z(
        \Data_Mem/n6010 ) );
  MUX U3059 ( .A(data_mem_out_wire[225]), .B(reg_target[1]), .S(n1811), .Z(
        \Data_Mem/n6009 ) );
  MUX U3060 ( .A(data_mem_out_wire[224]), .B(reg_target[0]), .S(n1811), .Z(
        \Data_Mem/n6008 ) );
  NOR U3061 ( .A(n1812), .B(n1792), .Z(n1811) );
  NANDN U3062 ( .A(N24), .B(n1813), .Z(n1792) );
  MUX U3063 ( .A(reg_target[31]), .B(data_mem_out_wire[287]), .S(n1814), .Z(
        \Data_Mem/n6007 ) );
  MUX U3064 ( .A(reg_target[30]), .B(data_mem_out_wire[286]), .S(n1814), .Z(
        \Data_Mem/n6006 ) );
  MUX U3065 ( .A(reg_target[29]), .B(data_mem_out_wire[285]), .S(n1814), .Z(
        \Data_Mem/n6005 ) );
  MUX U3066 ( .A(reg_target[28]), .B(data_mem_out_wire[284]), .S(n1814), .Z(
        \Data_Mem/n6004 ) );
  MUX U3067 ( .A(reg_target[27]), .B(data_mem_out_wire[283]), .S(n1814), .Z(
        \Data_Mem/n6003 ) );
  MUX U3068 ( .A(reg_target[26]), .B(data_mem_out_wire[282]), .S(n1814), .Z(
        \Data_Mem/n6002 ) );
  MUX U3069 ( .A(reg_target[25]), .B(data_mem_out_wire[281]), .S(n1814), .Z(
        \Data_Mem/n6001 ) );
  MUX U3070 ( .A(reg_target[24]), .B(data_mem_out_wire[280]), .S(n1814), .Z(
        \Data_Mem/n6000 ) );
  MUX U3071 ( .A(reg_target[23]), .B(data_mem_out_wire[279]), .S(n1814), .Z(
        \Data_Mem/n5999 ) );
  MUX U3072 ( .A(reg_target[22]), .B(data_mem_out_wire[278]), .S(n1814), .Z(
        \Data_Mem/n5998 ) );
  MUX U3073 ( .A(reg_target[21]), .B(data_mem_out_wire[277]), .S(n1814), .Z(
        \Data_Mem/n5997 ) );
  MUX U3074 ( .A(reg_target[20]), .B(data_mem_out_wire[276]), .S(n1814), .Z(
        \Data_Mem/n5996 ) );
  MUX U3075 ( .A(reg_target[19]), .B(data_mem_out_wire[275]), .S(n1814), .Z(
        \Data_Mem/n5995 ) );
  MUX U3076 ( .A(reg_target[18]), .B(data_mem_out_wire[274]), .S(n1814), .Z(
        \Data_Mem/n5994 ) );
  MUX U3077 ( .A(reg_target[17]), .B(data_mem_out_wire[273]), .S(n1814), .Z(
        \Data_Mem/n5993 ) );
  MUX U3078 ( .A(reg_target[16]), .B(data_mem_out_wire[272]), .S(n1814), .Z(
        \Data_Mem/n5992 ) );
  MUX U3079 ( .A(reg_target[15]), .B(data_mem_out_wire[271]), .S(n1814), .Z(
        \Data_Mem/n5991 ) );
  MUX U3080 ( .A(reg_target[14]), .B(data_mem_out_wire[270]), .S(n1814), .Z(
        \Data_Mem/n5990 ) );
  MUX U3081 ( .A(reg_target[13]), .B(data_mem_out_wire[269]), .S(n1814), .Z(
        \Data_Mem/n5989 ) );
  MUX U3082 ( .A(reg_target[12]), .B(data_mem_out_wire[268]), .S(n1814), .Z(
        \Data_Mem/n5988 ) );
  MUX U3083 ( .A(reg_target[11]), .B(data_mem_out_wire[267]), .S(n1814), .Z(
        \Data_Mem/n5987 ) );
  MUX U3084 ( .A(reg_target[10]), .B(data_mem_out_wire[266]), .S(n1814), .Z(
        \Data_Mem/n5986 ) );
  MUX U3085 ( .A(reg_target[9]), .B(data_mem_out_wire[265]), .S(n1814), .Z(
        \Data_Mem/n5985 ) );
  MUX U3086 ( .A(reg_target[8]), .B(data_mem_out_wire[264]), .S(n1814), .Z(
        \Data_Mem/n5984 ) );
  MUX U3087 ( .A(reg_target[7]), .B(data_mem_out_wire[263]), .S(n1814), .Z(
        \Data_Mem/n5983 ) );
  MUX U3088 ( .A(reg_target[6]), .B(data_mem_out_wire[262]), .S(n1814), .Z(
        \Data_Mem/n5982 ) );
  MUX U3089 ( .A(reg_target[5]), .B(data_mem_out_wire[261]), .S(n1814), .Z(
        \Data_Mem/n5981 ) );
  MUX U3090 ( .A(reg_target[4]), .B(data_mem_out_wire[260]), .S(n1814), .Z(
        \Data_Mem/n5980 ) );
  MUX U3091 ( .A(reg_target[3]), .B(data_mem_out_wire[259]), .S(n1814), .Z(
        \Data_Mem/n5979 ) );
  MUX U3092 ( .A(reg_target[2]), .B(data_mem_out_wire[258]), .S(n1814), .Z(
        \Data_Mem/n5978 ) );
  IV U3093 ( .A(n1815), .Z(n1814) );
  MUX U3094 ( .A(data_mem_out_wire[257]), .B(reg_target[1]), .S(n1815), .Z(
        \Data_Mem/n5977 ) );
  MUX U3095 ( .A(data_mem_out_wire[256]), .B(reg_target[0]), .S(n1815), .Z(
        \Data_Mem/n5976 ) );
  AND U3096 ( .A(n1791), .B(n1816), .Z(n1815) );
  MUX U3097 ( .A(reg_target[31]), .B(data_mem_out_wire[319]), .S(n1817), .Z(
        \Data_Mem/n5975 ) );
  MUX U3098 ( .A(reg_target[30]), .B(data_mem_out_wire[318]), .S(n1817), .Z(
        \Data_Mem/n5974 ) );
  MUX U3099 ( .A(reg_target[29]), .B(data_mem_out_wire[317]), .S(n1817), .Z(
        \Data_Mem/n5973 ) );
  MUX U3100 ( .A(reg_target[28]), .B(data_mem_out_wire[316]), .S(n1817), .Z(
        \Data_Mem/n5972 ) );
  MUX U3101 ( .A(reg_target[27]), .B(data_mem_out_wire[315]), .S(n1817), .Z(
        \Data_Mem/n5971 ) );
  MUX U3102 ( .A(reg_target[26]), .B(data_mem_out_wire[314]), .S(n1817), .Z(
        \Data_Mem/n5970 ) );
  MUX U3103 ( .A(reg_target[25]), .B(data_mem_out_wire[313]), .S(n1817), .Z(
        \Data_Mem/n5969 ) );
  MUX U3104 ( .A(reg_target[24]), .B(data_mem_out_wire[312]), .S(n1817), .Z(
        \Data_Mem/n5968 ) );
  MUX U3105 ( .A(reg_target[23]), .B(data_mem_out_wire[311]), .S(n1817), .Z(
        \Data_Mem/n5967 ) );
  MUX U3106 ( .A(reg_target[22]), .B(data_mem_out_wire[310]), .S(n1817), .Z(
        \Data_Mem/n5966 ) );
  MUX U3107 ( .A(reg_target[21]), .B(data_mem_out_wire[309]), .S(n1817), .Z(
        \Data_Mem/n5965 ) );
  MUX U3108 ( .A(reg_target[20]), .B(data_mem_out_wire[308]), .S(n1817), .Z(
        \Data_Mem/n5964 ) );
  MUX U3109 ( .A(reg_target[19]), .B(data_mem_out_wire[307]), .S(n1817), .Z(
        \Data_Mem/n5963 ) );
  MUX U3110 ( .A(reg_target[18]), .B(data_mem_out_wire[306]), .S(n1817), .Z(
        \Data_Mem/n5962 ) );
  MUX U3111 ( .A(reg_target[17]), .B(data_mem_out_wire[305]), .S(n1817), .Z(
        \Data_Mem/n5961 ) );
  MUX U3112 ( .A(reg_target[16]), .B(data_mem_out_wire[304]), .S(n1817), .Z(
        \Data_Mem/n5960 ) );
  MUX U3113 ( .A(reg_target[15]), .B(data_mem_out_wire[303]), .S(n1817), .Z(
        \Data_Mem/n5959 ) );
  MUX U3114 ( .A(reg_target[14]), .B(data_mem_out_wire[302]), .S(n1817), .Z(
        \Data_Mem/n5958 ) );
  MUX U3115 ( .A(reg_target[13]), .B(data_mem_out_wire[301]), .S(n1817), .Z(
        \Data_Mem/n5957 ) );
  MUX U3116 ( .A(reg_target[12]), .B(data_mem_out_wire[300]), .S(n1817), .Z(
        \Data_Mem/n5956 ) );
  MUX U3117 ( .A(reg_target[11]), .B(data_mem_out_wire[299]), .S(n1817), .Z(
        \Data_Mem/n5955 ) );
  MUX U3118 ( .A(reg_target[10]), .B(data_mem_out_wire[298]), .S(n1817), .Z(
        \Data_Mem/n5954 ) );
  MUX U3119 ( .A(reg_target[9]), .B(data_mem_out_wire[297]), .S(n1817), .Z(
        \Data_Mem/n5953 ) );
  MUX U3120 ( .A(reg_target[8]), .B(data_mem_out_wire[296]), .S(n1817), .Z(
        \Data_Mem/n5952 ) );
  MUX U3121 ( .A(reg_target[7]), .B(data_mem_out_wire[295]), .S(n1817), .Z(
        \Data_Mem/n5951 ) );
  MUX U3122 ( .A(reg_target[6]), .B(data_mem_out_wire[294]), .S(n1817), .Z(
        \Data_Mem/n5950 ) );
  MUX U3123 ( .A(reg_target[5]), .B(data_mem_out_wire[293]), .S(n1817), .Z(
        \Data_Mem/n5949 ) );
  MUX U3124 ( .A(reg_target[4]), .B(data_mem_out_wire[292]), .S(n1817), .Z(
        \Data_Mem/n5948 ) );
  MUX U3125 ( .A(reg_target[3]), .B(data_mem_out_wire[291]), .S(n1817), .Z(
        \Data_Mem/n5947 ) );
  MUX U3126 ( .A(reg_target[2]), .B(data_mem_out_wire[290]), .S(n1817), .Z(
        \Data_Mem/n5946 ) );
  IV U3127 ( .A(n1818), .Z(n1817) );
  MUX U3128 ( .A(data_mem_out_wire[289]), .B(reg_target[1]), .S(n1818), .Z(
        \Data_Mem/n5945 ) );
  MUX U3129 ( .A(data_mem_out_wire[288]), .B(reg_target[0]), .S(n1818), .Z(
        \Data_Mem/n5944 ) );
  AND U3130 ( .A(n1795), .B(n1816), .Z(n1818) );
  MUX U3131 ( .A(reg_target[31]), .B(data_mem_out_wire[351]), .S(n1819), .Z(
        \Data_Mem/n5943 ) );
  MUX U3132 ( .A(reg_target[30]), .B(data_mem_out_wire[350]), .S(n1819), .Z(
        \Data_Mem/n5942 ) );
  MUX U3133 ( .A(reg_target[29]), .B(data_mem_out_wire[349]), .S(n1819), .Z(
        \Data_Mem/n5941 ) );
  MUX U3134 ( .A(reg_target[28]), .B(data_mem_out_wire[348]), .S(n1819), .Z(
        \Data_Mem/n5940 ) );
  MUX U3135 ( .A(reg_target[27]), .B(data_mem_out_wire[347]), .S(n1819), .Z(
        \Data_Mem/n5939 ) );
  MUX U3136 ( .A(reg_target[26]), .B(data_mem_out_wire[346]), .S(n1819), .Z(
        \Data_Mem/n5938 ) );
  MUX U3137 ( .A(reg_target[25]), .B(data_mem_out_wire[345]), .S(n1819), .Z(
        \Data_Mem/n5937 ) );
  MUX U3138 ( .A(reg_target[24]), .B(data_mem_out_wire[344]), .S(n1819), .Z(
        \Data_Mem/n5936 ) );
  MUX U3139 ( .A(reg_target[23]), .B(data_mem_out_wire[343]), .S(n1819), .Z(
        \Data_Mem/n5935 ) );
  MUX U3140 ( .A(reg_target[22]), .B(data_mem_out_wire[342]), .S(n1819), .Z(
        \Data_Mem/n5934 ) );
  MUX U3141 ( .A(reg_target[21]), .B(data_mem_out_wire[341]), .S(n1819), .Z(
        \Data_Mem/n5933 ) );
  MUX U3142 ( .A(reg_target[20]), .B(data_mem_out_wire[340]), .S(n1819), .Z(
        \Data_Mem/n5932 ) );
  MUX U3143 ( .A(reg_target[19]), .B(data_mem_out_wire[339]), .S(n1819), .Z(
        \Data_Mem/n5931 ) );
  MUX U3144 ( .A(reg_target[18]), .B(data_mem_out_wire[338]), .S(n1819), .Z(
        \Data_Mem/n5930 ) );
  MUX U3145 ( .A(reg_target[17]), .B(data_mem_out_wire[337]), .S(n1819), .Z(
        \Data_Mem/n5929 ) );
  MUX U3146 ( .A(reg_target[16]), .B(data_mem_out_wire[336]), .S(n1819), .Z(
        \Data_Mem/n5928 ) );
  MUX U3147 ( .A(reg_target[15]), .B(data_mem_out_wire[335]), .S(n1819), .Z(
        \Data_Mem/n5927 ) );
  MUX U3148 ( .A(reg_target[14]), .B(data_mem_out_wire[334]), .S(n1819), .Z(
        \Data_Mem/n5926 ) );
  MUX U3149 ( .A(reg_target[13]), .B(data_mem_out_wire[333]), .S(n1819), .Z(
        \Data_Mem/n5925 ) );
  MUX U3150 ( .A(reg_target[12]), .B(data_mem_out_wire[332]), .S(n1819), .Z(
        \Data_Mem/n5924 ) );
  MUX U3151 ( .A(reg_target[11]), .B(data_mem_out_wire[331]), .S(n1819), .Z(
        \Data_Mem/n5923 ) );
  MUX U3152 ( .A(reg_target[10]), .B(data_mem_out_wire[330]), .S(n1819), .Z(
        \Data_Mem/n5922 ) );
  MUX U3153 ( .A(reg_target[9]), .B(data_mem_out_wire[329]), .S(n1819), .Z(
        \Data_Mem/n5921 ) );
  MUX U3154 ( .A(reg_target[8]), .B(data_mem_out_wire[328]), .S(n1819), .Z(
        \Data_Mem/n5920 ) );
  MUX U3155 ( .A(reg_target[7]), .B(data_mem_out_wire[327]), .S(n1819), .Z(
        \Data_Mem/n5919 ) );
  MUX U3156 ( .A(reg_target[6]), .B(data_mem_out_wire[326]), .S(n1819), .Z(
        \Data_Mem/n5918 ) );
  MUX U3157 ( .A(reg_target[5]), .B(data_mem_out_wire[325]), .S(n1819), .Z(
        \Data_Mem/n5917 ) );
  MUX U3158 ( .A(reg_target[4]), .B(data_mem_out_wire[324]), .S(n1819), .Z(
        \Data_Mem/n5916 ) );
  MUX U3159 ( .A(reg_target[3]), .B(data_mem_out_wire[323]), .S(n1819), .Z(
        \Data_Mem/n5915 ) );
  MUX U3160 ( .A(reg_target[2]), .B(data_mem_out_wire[322]), .S(n1819), .Z(
        \Data_Mem/n5914 ) );
  IV U3161 ( .A(n1820), .Z(n1819) );
  MUX U3162 ( .A(data_mem_out_wire[321]), .B(reg_target[1]), .S(n1820), .Z(
        \Data_Mem/n5913 ) );
  MUX U3163 ( .A(data_mem_out_wire[320]), .B(reg_target[0]), .S(n1820), .Z(
        \Data_Mem/n5912 ) );
  AND U3164 ( .A(n1798), .B(n1816), .Z(n1820) );
  MUX U3165 ( .A(reg_target[31]), .B(data_mem_out_wire[383]), .S(n1821), .Z(
        \Data_Mem/n5911 ) );
  MUX U3166 ( .A(reg_target[30]), .B(data_mem_out_wire[382]), .S(n1821), .Z(
        \Data_Mem/n5910 ) );
  MUX U3167 ( .A(reg_target[29]), .B(data_mem_out_wire[381]), .S(n1821), .Z(
        \Data_Mem/n5909 ) );
  MUX U3168 ( .A(reg_target[28]), .B(data_mem_out_wire[380]), .S(n1821), .Z(
        \Data_Mem/n5908 ) );
  MUX U3169 ( .A(reg_target[27]), .B(data_mem_out_wire[379]), .S(n1821), .Z(
        \Data_Mem/n5907 ) );
  MUX U3170 ( .A(reg_target[26]), .B(data_mem_out_wire[378]), .S(n1821), .Z(
        \Data_Mem/n5906 ) );
  MUX U3171 ( .A(reg_target[25]), .B(data_mem_out_wire[377]), .S(n1821), .Z(
        \Data_Mem/n5905 ) );
  MUX U3172 ( .A(reg_target[24]), .B(data_mem_out_wire[376]), .S(n1821), .Z(
        \Data_Mem/n5904 ) );
  MUX U3173 ( .A(reg_target[23]), .B(data_mem_out_wire[375]), .S(n1821), .Z(
        \Data_Mem/n5903 ) );
  MUX U3174 ( .A(reg_target[22]), .B(data_mem_out_wire[374]), .S(n1821), .Z(
        \Data_Mem/n5902 ) );
  MUX U3175 ( .A(reg_target[21]), .B(data_mem_out_wire[373]), .S(n1821), .Z(
        \Data_Mem/n5901 ) );
  MUX U3176 ( .A(reg_target[20]), .B(data_mem_out_wire[372]), .S(n1821), .Z(
        \Data_Mem/n5900 ) );
  MUX U3177 ( .A(reg_target[19]), .B(data_mem_out_wire[371]), .S(n1821), .Z(
        \Data_Mem/n5899 ) );
  MUX U3178 ( .A(reg_target[18]), .B(data_mem_out_wire[370]), .S(n1821), .Z(
        \Data_Mem/n5898 ) );
  MUX U3179 ( .A(reg_target[17]), .B(data_mem_out_wire[369]), .S(n1821), .Z(
        \Data_Mem/n5897 ) );
  MUX U3180 ( .A(reg_target[16]), .B(data_mem_out_wire[368]), .S(n1821), .Z(
        \Data_Mem/n5896 ) );
  MUX U3181 ( .A(reg_target[15]), .B(data_mem_out_wire[367]), .S(n1821), .Z(
        \Data_Mem/n5895 ) );
  MUX U3182 ( .A(reg_target[14]), .B(data_mem_out_wire[366]), .S(n1821), .Z(
        \Data_Mem/n5894 ) );
  MUX U3183 ( .A(reg_target[13]), .B(data_mem_out_wire[365]), .S(n1821), .Z(
        \Data_Mem/n5893 ) );
  MUX U3184 ( .A(reg_target[12]), .B(data_mem_out_wire[364]), .S(n1821), .Z(
        \Data_Mem/n5892 ) );
  MUX U3185 ( .A(reg_target[11]), .B(data_mem_out_wire[363]), .S(n1821), .Z(
        \Data_Mem/n5891 ) );
  MUX U3186 ( .A(reg_target[10]), .B(data_mem_out_wire[362]), .S(n1821), .Z(
        \Data_Mem/n5890 ) );
  MUX U3187 ( .A(reg_target[9]), .B(data_mem_out_wire[361]), .S(n1821), .Z(
        \Data_Mem/n5889 ) );
  MUX U3188 ( .A(reg_target[8]), .B(data_mem_out_wire[360]), .S(n1821), .Z(
        \Data_Mem/n5888 ) );
  MUX U3189 ( .A(reg_target[7]), .B(data_mem_out_wire[359]), .S(n1821), .Z(
        \Data_Mem/n5887 ) );
  MUX U3190 ( .A(reg_target[6]), .B(data_mem_out_wire[358]), .S(n1821), .Z(
        \Data_Mem/n5886 ) );
  MUX U3191 ( .A(reg_target[5]), .B(data_mem_out_wire[357]), .S(n1821), .Z(
        \Data_Mem/n5885 ) );
  MUX U3192 ( .A(reg_target[4]), .B(data_mem_out_wire[356]), .S(n1821), .Z(
        \Data_Mem/n5884 ) );
  MUX U3193 ( .A(reg_target[3]), .B(data_mem_out_wire[355]), .S(n1821), .Z(
        \Data_Mem/n5883 ) );
  MUX U3194 ( .A(reg_target[2]), .B(data_mem_out_wire[354]), .S(n1821), .Z(
        \Data_Mem/n5882 ) );
  IV U3195 ( .A(n1822), .Z(n1821) );
  MUX U3196 ( .A(data_mem_out_wire[353]), .B(reg_target[1]), .S(n1822), .Z(
        \Data_Mem/n5881 ) );
  MUX U3197 ( .A(data_mem_out_wire[352]), .B(reg_target[0]), .S(n1822), .Z(
        \Data_Mem/n5880 ) );
  AND U3198 ( .A(n1801), .B(n1816), .Z(n1822) );
  MUX U3199 ( .A(reg_target[31]), .B(data_mem_out_wire[415]), .S(n1823), .Z(
        \Data_Mem/n5879 ) );
  MUX U3200 ( .A(reg_target[30]), .B(data_mem_out_wire[414]), .S(n1823), .Z(
        \Data_Mem/n5878 ) );
  MUX U3201 ( .A(reg_target[29]), .B(data_mem_out_wire[413]), .S(n1823), .Z(
        \Data_Mem/n5877 ) );
  MUX U3202 ( .A(reg_target[28]), .B(data_mem_out_wire[412]), .S(n1823), .Z(
        \Data_Mem/n5876 ) );
  MUX U3203 ( .A(reg_target[27]), .B(data_mem_out_wire[411]), .S(n1823), .Z(
        \Data_Mem/n5875 ) );
  MUX U3204 ( .A(reg_target[26]), .B(data_mem_out_wire[410]), .S(n1823), .Z(
        \Data_Mem/n5874 ) );
  MUX U3205 ( .A(reg_target[25]), .B(data_mem_out_wire[409]), .S(n1823), .Z(
        \Data_Mem/n5873 ) );
  MUX U3206 ( .A(reg_target[24]), .B(data_mem_out_wire[408]), .S(n1823), .Z(
        \Data_Mem/n5872 ) );
  MUX U3207 ( .A(reg_target[23]), .B(data_mem_out_wire[407]), .S(n1823), .Z(
        \Data_Mem/n5871 ) );
  MUX U3208 ( .A(reg_target[22]), .B(data_mem_out_wire[406]), .S(n1823), .Z(
        \Data_Mem/n5870 ) );
  MUX U3209 ( .A(reg_target[21]), .B(data_mem_out_wire[405]), .S(n1823), .Z(
        \Data_Mem/n5869 ) );
  MUX U3210 ( .A(reg_target[20]), .B(data_mem_out_wire[404]), .S(n1823), .Z(
        \Data_Mem/n5868 ) );
  MUX U3211 ( .A(reg_target[19]), .B(data_mem_out_wire[403]), .S(n1823), .Z(
        \Data_Mem/n5867 ) );
  MUX U3212 ( .A(reg_target[18]), .B(data_mem_out_wire[402]), .S(n1823), .Z(
        \Data_Mem/n5866 ) );
  MUX U3213 ( .A(reg_target[17]), .B(data_mem_out_wire[401]), .S(n1823), .Z(
        \Data_Mem/n5865 ) );
  MUX U3214 ( .A(reg_target[16]), .B(data_mem_out_wire[400]), .S(n1823), .Z(
        \Data_Mem/n5864 ) );
  MUX U3215 ( .A(reg_target[15]), .B(data_mem_out_wire[399]), .S(n1823), .Z(
        \Data_Mem/n5863 ) );
  MUX U3216 ( .A(reg_target[14]), .B(data_mem_out_wire[398]), .S(n1823), .Z(
        \Data_Mem/n5862 ) );
  MUX U3217 ( .A(reg_target[13]), .B(data_mem_out_wire[397]), .S(n1823), .Z(
        \Data_Mem/n5861 ) );
  MUX U3218 ( .A(reg_target[12]), .B(data_mem_out_wire[396]), .S(n1823), .Z(
        \Data_Mem/n5860 ) );
  MUX U3219 ( .A(reg_target[11]), .B(data_mem_out_wire[395]), .S(n1823), .Z(
        \Data_Mem/n5859 ) );
  MUX U3220 ( .A(reg_target[10]), .B(data_mem_out_wire[394]), .S(n1823), .Z(
        \Data_Mem/n5858 ) );
  MUX U3221 ( .A(reg_target[9]), .B(data_mem_out_wire[393]), .S(n1823), .Z(
        \Data_Mem/n5857 ) );
  MUX U3222 ( .A(reg_target[8]), .B(data_mem_out_wire[392]), .S(n1823), .Z(
        \Data_Mem/n5856 ) );
  MUX U3223 ( .A(reg_target[7]), .B(data_mem_out_wire[391]), .S(n1823), .Z(
        \Data_Mem/n5855 ) );
  MUX U3224 ( .A(reg_target[6]), .B(data_mem_out_wire[390]), .S(n1823), .Z(
        \Data_Mem/n5854 ) );
  MUX U3225 ( .A(reg_target[5]), .B(data_mem_out_wire[389]), .S(n1823), .Z(
        \Data_Mem/n5853 ) );
  MUX U3226 ( .A(reg_target[4]), .B(data_mem_out_wire[388]), .S(n1823), .Z(
        \Data_Mem/n5852 ) );
  MUX U3227 ( .A(reg_target[3]), .B(data_mem_out_wire[387]), .S(n1823), .Z(
        \Data_Mem/n5851 ) );
  MUX U3228 ( .A(reg_target[2]), .B(data_mem_out_wire[386]), .S(n1823), .Z(
        \Data_Mem/n5850 ) );
  IV U3229 ( .A(n1824), .Z(n1823) );
  MUX U3230 ( .A(data_mem_out_wire[385]), .B(reg_target[1]), .S(n1824), .Z(
        \Data_Mem/n5849 ) );
  MUX U3231 ( .A(data_mem_out_wire[384]), .B(reg_target[0]), .S(n1824), .Z(
        \Data_Mem/n5848 ) );
  AND U3232 ( .A(n1804), .B(n1816), .Z(n1824) );
  MUX U3233 ( .A(reg_target[31]), .B(data_mem_out_wire[447]), .S(n1825), .Z(
        \Data_Mem/n5847 ) );
  MUX U3234 ( .A(reg_target[30]), .B(data_mem_out_wire[446]), .S(n1825), .Z(
        \Data_Mem/n5846 ) );
  MUX U3235 ( .A(reg_target[29]), .B(data_mem_out_wire[445]), .S(n1825), .Z(
        \Data_Mem/n5845 ) );
  MUX U3236 ( .A(reg_target[28]), .B(data_mem_out_wire[444]), .S(n1825), .Z(
        \Data_Mem/n5844 ) );
  MUX U3237 ( .A(reg_target[27]), .B(data_mem_out_wire[443]), .S(n1825), .Z(
        \Data_Mem/n5843 ) );
  MUX U3238 ( .A(reg_target[26]), .B(data_mem_out_wire[442]), .S(n1825), .Z(
        \Data_Mem/n5842 ) );
  MUX U3239 ( .A(reg_target[25]), .B(data_mem_out_wire[441]), .S(n1825), .Z(
        \Data_Mem/n5841 ) );
  MUX U3240 ( .A(reg_target[24]), .B(data_mem_out_wire[440]), .S(n1825), .Z(
        \Data_Mem/n5840 ) );
  MUX U3241 ( .A(reg_target[23]), .B(data_mem_out_wire[439]), .S(n1825), .Z(
        \Data_Mem/n5839 ) );
  MUX U3242 ( .A(reg_target[22]), .B(data_mem_out_wire[438]), .S(n1825), .Z(
        \Data_Mem/n5838 ) );
  MUX U3243 ( .A(reg_target[21]), .B(data_mem_out_wire[437]), .S(n1825), .Z(
        \Data_Mem/n5837 ) );
  MUX U3244 ( .A(reg_target[20]), .B(data_mem_out_wire[436]), .S(n1825), .Z(
        \Data_Mem/n5836 ) );
  MUX U3245 ( .A(reg_target[19]), .B(data_mem_out_wire[435]), .S(n1825), .Z(
        \Data_Mem/n5835 ) );
  MUX U3246 ( .A(reg_target[18]), .B(data_mem_out_wire[434]), .S(n1825), .Z(
        \Data_Mem/n5834 ) );
  MUX U3247 ( .A(reg_target[17]), .B(data_mem_out_wire[433]), .S(n1825), .Z(
        \Data_Mem/n5833 ) );
  MUX U3248 ( .A(reg_target[16]), .B(data_mem_out_wire[432]), .S(n1825), .Z(
        \Data_Mem/n5832 ) );
  MUX U3249 ( .A(reg_target[15]), .B(data_mem_out_wire[431]), .S(n1825), .Z(
        \Data_Mem/n5831 ) );
  MUX U3250 ( .A(reg_target[14]), .B(data_mem_out_wire[430]), .S(n1825), .Z(
        \Data_Mem/n5830 ) );
  MUX U3251 ( .A(reg_target[13]), .B(data_mem_out_wire[429]), .S(n1825), .Z(
        \Data_Mem/n5829 ) );
  MUX U3252 ( .A(reg_target[12]), .B(data_mem_out_wire[428]), .S(n1825), .Z(
        \Data_Mem/n5828 ) );
  MUX U3253 ( .A(reg_target[11]), .B(data_mem_out_wire[427]), .S(n1825), .Z(
        \Data_Mem/n5827 ) );
  MUX U3254 ( .A(reg_target[10]), .B(data_mem_out_wire[426]), .S(n1825), .Z(
        \Data_Mem/n5826 ) );
  MUX U3255 ( .A(reg_target[9]), .B(data_mem_out_wire[425]), .S(n1825), .Z(
        \Data_Mem/n5825 ) );
  MUX U3256 ( .A(reg_target[8]), .B(data_mem_out_wire[424]), .S(n1825), .Z(
        \Data_Mem/n5824 ) );
  MUX U3257 ( .A(reg_target[7]), .B(data_mem_out_wire[423]), .S(n1825), .Z(
        \Data_Mem/n5823 ) );
  MUX U3258 ( .A(reg_target[6]), .B(data_mem_out_wire[422]), .S(n1825), .Z(
        \Data_Mem/n5822 ) );
  MUX U3259 ( .A(reg_target[5]), .B(data_mem_out_wire[421]), .S(n1825), .Z(
        \Data_Mem/n5821 ) );
  MUX U3260 ( .A(reg_target[4]), .B(data_mem_out_wire[420]), .S(n1825), .Z(
        \Data_Mem/n5820 ) );
  MUX U3261 ( .A(reg_target[3]), .B(data_mem_out_wire[419]), .S(n1825), .Z(
        \Data_Mem/n5819 ) );
  MUX U3262 ( .A(reg_target[2]), .B(data_mem_out_wire[418]), .S(n1825), .Z(
        \Data_Mem/n5818 ) );
  IV U3263 ( .A(n1826), .Z(n1825) );
  MUX U3264 ( .A(data_mem_out_wire[417]), .B(reg_target[1]), .S(n1826), .Z(
        \Data_Mem/n5817 ) );
  MUX U3265 ( .A(data_mem_out_wire[416]), .B(reg_target[0]), .S(n1826), .Z(
        \Data_Mem/n5816 ) );
  AND U3266 ( .A(n1807), .B(n1816), .Z(n1826) );
  MUX U3267 ( .A(reg_target[31]), .B(data_mem_out_wire[479]), .S(n1827), .Z(
        \Data_Mem/n5815 ) );
  MUX U3268 ( .A(reg_target[30]), .B(data_mem_out_wire[478]), .S(n1827), .Z(
        \Data_Mem/n5814 ) );
  MUX U3269 ( .A(reg_target[29]), .B(data_mem_out_wire[477]), .S(n1827), .Z(
        \Data_Mem/n5813 ) );
  MUX U3270 ( .A(reg_target[28]), .B(data_mem_out_wire[476]), .S(n1827), .Z(
        \Data_Mem/n5812 ) );
  MUX U3271 ( .A(reg_target[27]), .B(data_mem_out_wire[475]), .S(n1827), .Z(
        \Data_Mem/n5811 ) );
  MUX U3272 ( .A(reg_target[26]), .B(data_mem_out_wire[474]), .S(n1827), .Z(
        \Data_Mem/n5810 ) );
  MUX U3273 ( .A(reg_target[25]), .B(data_mem_out_wire[473]), .S(n1827), .Z(
        \Data_Mem/n5809 ) );
  MUX U3274 ( .A(reg_target[24]), .B(data_mem_out_wire[472]), .S(n1827), .Z(
        \Data_Mem/n5808 ) );
  MUX U3275 ( .A(reg_target[23]), .B(data_mem_out_wire[471]), .S(n1827), .Z(
        \Data_Mem/n5807 ) );
  MUX U3276 ( .A(reg_target[22]), .B(data_mem_out_wire[470]), .S(n1827), .Z(
        \Data_Mem/n5806 ) );
  MUX U3277 ( .A(reg_target[21]), .B(data_mem_out_wire[469]), .S(n1827), .Z(
        \Data_Mem/n5805 ) );
  MUX U3278 ( .A(reg_target[20]), .B(data_mem_out_wire[468]), .S(n1827), .Z(
        \Data_Mem/n5804 ) );
  MUX U3279 ( .A(reg_target[19]), .B(data_mem_out_wire[467]), .S(n1827), .Z(
        \Data_Mem/n5803 ) );
  MUX U3280 ( .A(reg_target[18]), .B(data_mem_out_wire[466]), .S(n1827), .Z(
        \Data_Mem/n5802 ) );
  MUX U3281 ( .A(reg_target[17]), .B(data_mem_out_wire[465]), .S(n1827), .Z(
        \Data_Mem/n5801 ) );
  MUX U3282 ( .A(reg_target[16]), .B(data_mem_out_wire[464]), .S(n1827), .Z(
        \Data_Mem/n5800 ) );
  MUX U3283 ( .A(reg_target[15]), .B(data_mem_out_wire[463]), .S(n1827), .Z(
        \Data_Mem/n5799 ) );
  MUX U3284 ( .A(reg_target[14]), .B(data_mem_out_wire[462]), .S(n1827), .Z(
        \Data_Mem/n5798 ) );
  MUX U3285 ( .A(reg_target[13]), .B(data_mem_out_wire[461]), .S(n1827), .Z(
        \Data_Mem/n5797 ) );
  MUX U3286 ( .A(reg_target[12]), .B(data_mem_out_wire[460]), .S(n1827), .Z(
        \Data_Mem/n5796 ) );
  MUX U3287 ( .A(reg_target[11]), .B(data_mem_out_wire[459]), .S(n1827), .Z(
        \Data_Mem/n5795 ) );
  MUX U3288 ( .A(reg_target[10]), .B(data_mem_out_wire[458]), .S(n1827), .Z(
        \Data_Mem/n5794 ) );
  MUX U3289 ( .A(reg_target[9]), .B(data_mem_out_wire[457]), .S(n1827), .Z(
        \Data_Mem/n5793 ) );
  MUX U3290 ( .A(reg_target[8]), .B(data_mem_out_wire[456]), .S(n1827), .Z(
        \Data_Mem/n5792 ) );
  MUX U3291 ( .A(reg_target[7]), .B(data_mem_out_wire[455]), .S(n1827), .Z(
        \Data_Mem/n5791 ) );
  MUX U3292 ( .A(reg_target[6]), .B(data_mem_out_wire[454]), .S(n1827), .Z(
        \Data_Mem/n5790 ) );
  MUX U3293 ( .A(reg_target[5]), .B(data_mem_out_wire[453]), .S(n1827), .Z(
        \Data_Mem/n5789 ) );
  MUX U3294 ( .A(reg_target[4]), .B(data_mem_out_wire[452]), .S(n1827), .Z(
        \Data_Mem/n5788 ) );
  MUX U3295 ( .A(reg_target[3]), .B(data_mem_out_wire[451]), .S(n1827), .Z(
        \Data_Mem/n5787 ) );
  MUX U3296 ( .A(reg_target[2]), .B(data_mem_out_wire[450]), .S(n1827), .Z(
        \Data_Mem/n5786 ) );
  IV U3297 ( .A(n1828), .Z(n1827) );
  MUX U3298 ( .A(data_mem_out_wire[449]), .B(reg_target[1]), .S(n1828), .Z(
        \Data_Mem/n5785 ) );
  MUX U3299 ( .A(data_mem_out_wire[448]), .B(reg_target[0]), .S(n1828), .Z(
        \Data_Mem/n5784 ) );
  AND U3300 ( .A(n1810), .B(n1816), .Z(n1828) );
  MUX U3301 ( .A(data_mem_out_wire[511]), .B(reg_target[31]), .S(n1829), .Z(
        \Data_Mem/n5783 ) );
  MUX U3302 ( .A(data_mem_out_wire[510]), .B(reg_target[30]), .S(n1829), .Z(
        \Data_Mem/n5782 ) );
  MUX U3303 ( .A(data_mem_out_wire[509]), .B(reg_target[29]), .S(n1829), .Z(
        \Data_Mem/n5781 ) );
  MUX U3304 ( .A(data_mem_out_wire[508]), .B(reg_target[28]), .S(n1829), .Z(
        \Data_Mem/n5780 ) );
  MUX U3305 ( .A(data_mem_out_wire[507]), .B(reg_target[27]), .S(n1829), .Z(
        \Data_Mem/n5779 ) );
  MUX U3306 ( .A(data_mem_out_wire[506]), .B(reg_target[26]), .S(n1829), .Z(
        \Data_Mem/n5778 ) );
  MUX U3307 ( .A(data_mem_out_wire[505]), .B(reg_target[25]), .S(n1829), .Z(
        \Data_Mem/n5777 ) );
  MUX U3308 ( .A(data_mem_out_wire[504]), .B(reg_target[24]), .S(n1829), .Z(
        \Data_Mem/n5776 ) );
  MUX U3309 ( .A(data_mem_out_wire[503]), .B(reg_target[23]), .S(n1829), .Z(
        \Data_Mem/n5775 ) );
  MUX U3310 ( .A(data_mem_out_wire[502]), .B(reg_target[22]), .S(n1829), .Z(
        \Data_Mem/n5774 ) );
  MUX U3311 ( .A(data_mem_out_wire[501]), .B(reg_target[21]), .S(n1829), .Z(
        \Data_Mem/n5773 ) );
  MUX U3312 ( .A(data_mem_out_wire[500]), .B(reg_target[20]), .S(n1829), .Z(
        \Data_Mem/n5772 ) );
  MUX U3313 ( .A(data_mem_out_wire[499]), .B(reg_target[19]), .S(n1829), .Z(
        \Data_Mem/n5771 ) );
  MUX U3314 ( .A(data_mem_out_wire[498]), .B(reg_target[18]), .S(n1829), .Z(
        \Data_Mem/n5770 ) );
  MUX U3315 ( .A(data_mem_out_wire[497]), .B(reg_target[17]), .S(n1829), .Z(
        \Data_Mem/n5769 ) );
  MUX U3316 ( .A(data_mem_out_wire[496]), .B(reg_target[16]), .S(n1829), .Z(
        \Data_Mem/n5768 ) );
  MUX U3317 ( .A(data_mem_out_wire[495]), .B(reg_target[15]), .S(n1829), .Z(
        \Data_Mem/n5767 ) );
  MUX U3318 ( .A(data_mem_out_wire[494]), .B(reg_target[14]), .S(n1829), .Z(
        \Data_Mem/n5766 ) );
  MUX U3319 ( .A(data_mem_out_wire[493]), .B(reg_target[13]), .S(n1829), .Z(
        \Data_Mem/n5765 ) );
  MUX U3320 ( .A(data_mem_out_wire[492]), .B(reg_target[12]), .S(n1829), .Z(
        \Data_Mem/n5764 ) );
  MUX U3321 ( .A(data_mem_out_wire[491]), .B(reg_target[11]), .S(n1829), .Z(
        \Data_Mem/n5763 ) );
  MUX U3322 ( .A(data_mem_out_wire[490]), .B(reg_target[10]), .S(n1829), .Z(
        \Data_Mem/n5762 ) );
  MUX U3323 ( .A(data_mem_out_wire[489]), .B(reg_target[9]), .S(n1829), .Z(
        \Data_Mem/n5761 ) );
  MUX U3324 ( .A(data_mem_out_wire[488]), .B(reg_target[8]), .S(n1829), .Z(
        \Data_Mem/n5760 ) );
  MUX U3325 ( .A(data_mem_out_wire[487]), .B(reg_target[7]), .S(n1829), .Z(
        \Data_Mem/n5759 ) );
  MUX U3326 ( .A(data_mem_out_wire[486]), .B(reg_target[6]), .S(n1829), .Z(
        \Data_Mem/n5758 ) );
  MUX U3327 ( .A(data_mem_out_wire[485]), .B(reg_target[5]), .S(n1829), .Z(
        \Data_Mem/n5757 ) );
  MUX U3328 ( .A(data_mem_out_wire[484]), .B(reg_target[4]), .S(n1829), .Z(
        \Data_Mem/n5756 ) );
  MUX U3329 ( .A(data_mem_out_wire[483]), .B(reg_target[3]), .S(n1829), .Z(
        \Data_Mem/n5755 ) );
  MUX U3330 ( .A(data_mem_out_wire[482]), .B(reg_target[2]), .S(n1829), .Z(
        \Data_Mem/n5754 ) );
  MUX U3331 ( .A(data_mem_out_wire[481]), .B(reg_target[1]), .S(n1829), .Z(
        \Data_Mem/n5753 ) );
  MUX U3332 ( .A(data_mem_out_wire[480]), .B(reg_target[0]), .S(n1829), .Z(
        \Data_Mem/n5752 ) );
  AND U3333 ( .A(n1816), .B(n1830), .Z(n1829) );
  ANDN U3334 ( .B(n1831), .A(N24), .Z(n1816) );
  MUX U3335 ( .A(reg_target[31]), .B(data_mem_out_wire[543]), .S(n1832), .Z(
        \Data_Mem/n5751 ) );
  MUX U3336 ( .A(reg_target[30]), .B(data_mem_out_wire[542]), .S(n1832), .Z(
        \Data_Mem/n5750 ) );
  MUX U3337 ( .A(reg_target[29]), .B(data_mem_out_wire[541]), .S(n1832), .Z(
        \Data_Mem/n5749 ) );
  MUX U3338 ( .A(reg_target[28]), .B(data_mem_out_wire[540]), .S(n1832), .Z(
        \Data_Mem/n5748 ) );
  MUX U3339 ( .A(reg_target[27]), .B(data_mem_out_wire[539]), .S(n1832), .Z(
        \Data_Mem/n5747 ) );
  MUX U3340 ( .A(reg_target[26]), .B(data_mem_out_wire[538]), .S(n1832), .Z(
        \Data_Mem/n5746 ) );
  MUX U3341 ( .A(reg_target[25]), .B(data_mem_out_wire[537]), .S(n1832), .Z(
        \Data_Mem/n5745 ) );
  MUX U3342 ( .A(reg_target[24]), .B(data_mem_out_wire[536]), .S(n1832), .Z(
        \Data_Mem/n5744 ) );
  MUX U3343 ( .A(reg_target[23]), .B(data_mem_out_wire[535]), .S(n1832), .Z(
        \Data_Mem/n5743 ) );
  MUX U3344 ( .A(reg_target[22]), .B(data_mem_out_wire[534]), .S(n1832), .Z(
        \Data_Mem/n5742 ) );
  MUX U3345 ( .A(reg_target[21]), .B(data_mem_out_wire[533]), .S(n1832), .Z(
        \Data_Mem/n5741 ) );
  MUX U3346 ( .A(reg_target[20]), .B(data_mem_out_wire[532]), .S(n1832), .Z(
        \Data_Mem/n5740 ) );
  MUX U3347 ( .A(reg_target[19]), .B(data_mem_out_wire[531]), .S(n1832), .Z(
        \Data_Mem/n5739 ) );
  MUX U3348 ( .A(reg_target[18]), .B(data_mem_out_wire[530]), .S(n1832), .Z(
        \Data_Mem/n5738 ) );
  MUX U3349 ( .A(reg_target[17]), .B(data_mem_out_wire[529]), .S(n1832), .Z(
        \Data_Mem/n5737 ) );
  MUX U3350 ( .A(reg_target[16]), .B(data_mem_out_wire[528]), .S(n1832), .Z(
        \Data_Mem/n5736 ) );
  MUX U3351 ( .A(reg_target[15]), .B(data_mem_out_wire[527]), .S(n1832), .Z(
        \Data_Mem/n5735 ) );
  MUX U3352 ( .A(reg_target[14]), .B(data_mem_out_wire[526]), .S(n1832), .Z(
        \Data_Mem/n5734 ) );
  MUX U3353 ( .A(reg_target[13]), .B(data_mem_out_wire[525]), .S(n1832), .Z(
        \Data_Mem/n5733 ) );
  MUX U3354 ( .A(reg_target[12]), .B(data_mem_out_wire[524]), .S(n1832), .Z(
        \Data_Mem/n5732 ) );
  MUX U3355 ( .A(reg_target[11]), .B(data_mem_out_wire[523]), .S(n1832), .Z(
        \Data_Mem/n5731 ) );
  MUX U3356 ( .A(reg_target[10]), .B(data_mem_out_wire[522]), .S(n1832), .Z(
        \Data_Mem/n5730 ) );
  MUX U3357 ( .A(reg_target[9]), .B(data_mem_out_wire[521]), .S(n1832), .Z(
        \Data_Mem/n5729 ) );
  MUX U3358 ( .A(reg_target[8]), .B(data_mem_out_wire[520]), .S(n1832), .Z(
        \Data_Mem/n5728 ) );
  MUX U3359 ( .A(reg_target[7]), .B(data_mem_out_wire[519]), .S(n1832), .Z(
        \Data_Mem/n5727 ) );
  MUX U3360 ( .A(reg_target[6]), .B(data_mem_out_wire[518]), .S(n1832), .Z(
        \Data_Mem/n5726 ) );
  MUX U3361 ( .A(reg_target[5]), .B(data_mem_out_wire[517]), .S(n1832), .Z(
        \Data_Mem/n5725 ) );
  MUX U3362 ( .A(reg_target[4]), .B(data_mem_out_wire[516]), .S(n1832), .Z(
        \Data_Mem/n5724 ) );
  MUX U3363 ( .A(reg_target[3]), .B(data_mem_out_wire[515]), .S(n1832), .Z(
        \Data_Mem/n5723 ) );
  MUX U3364 ( .A(reg_target[2]), .B(data_mem_out_wire[514]), .S(n1832), .Z(
        \Data_Mem/n5722 ) );
  IV U3365 ( .A(n1833), .Z(n1832) );
  MUX U3366 ( .A(data_mem_out_wire[513]), .B(reg_target[1]), .S(n1833), .Z(
        \Data_Mem/n5721 ) );
  MUX U3367 ( .A(data_mem_out_wire[512]), .B(reg_target[0]), .S(n1833), .Z(
        \Data_Mem/n5720 ) );
  AND U3368 ( .A(n1791), .B(n1834), .Z(n1833) );
  MUX U3369 ( .A(reg_target[31]), .B(data_mem_out_wire[575]), .S(n1835), .Z(
        \Data_Mem/n5719 ) );
  MUX U3370 ( .A(reg_target[30]), .B(data_mem_out_wire[574]), .S(n1835), .Z(
        \Data_Mem/n5718 ) );
  MUX U3371 ( .A(reg_target[29]), .B(data_mem_out_wire[573]), .S(n1835), .Z(
        \Data_Mem/n5717 ) );
  MUX U3372 ( .A(reg_target[28]), .B(data_mem_out_wire[572]), .S(n1835), .Z(
        \Data_Mem/n5716 ) );
  MUX U3373 ( .A(reg_target[27]), .B(data_mem_out_wire[571]), .S(n1835), .Z(
        \Data_Mem/n5715 ) );
  MUX U3374 ( .A(reg_target[26]), .B(data_mem_out_wire[570]), .S(n1835), .Z(
        \Data_Mem/n5714 ) );
  MUX U3375 ( .A(reg_target[25]), .B(data_mem_out_wire[569]), .S(n1835), .Z(
        \Data_Mem/n5713 ) );
  MUX U3376 ( .A(reg_target[24]), .B(data_mem_out_wire[568]), .S(n1835), .Z(
        \Data_Mem/n5712 ) );
  MUX U3377 ( .A(reg_target[23]), .B(data_mem_out_wire[567]), .S(n1835), .Z(
        \Data_Mem/n5711 ) );
  MUX U3378 ( .A(reg_target[22]), .B(data_mem_out_wire[566]), .S(n1835), .Z(
        \Data_Mem/n5710 ) );
  MUX U3379 ( .A(reg_target[21]), .B(data_mem_out_wire[565]), .S(n1835), .Z(
        \Data_Mem/n5709 ) );
  MUX U3380 ( .A(reg_target[20]), .B(data_mem_out_wire[564]), .S(n1835), .Z(
        \Data_Mem/n5708 ) );
  MUX U3381 ( .A(reg_target[19]), .B(data_mem_out_wire[563]), .S(n1835), .Z(
        \Data_Mem/n5707 ) );
  MUX U3382 ( .A(reg_target[18]), .B(data_mem_out_wire[562]), .S(n1835), .Z(
        \Data_Mem/n5706 ) );
  MUX U3383 ( .A(reg_target[17]), .B(data_mem_out_wire[561]), .S(n1835), .Z(
        \Data_Mem/n5705 ) );
  MUX U3384 ( .A(reg_target[16]), .B(data_mem_out_wire[560]), .S(n1835), .Z(
        \Data_Mem/n5704 ) );
  MUX U3385 ( .A(reg_target[15]), .B(data_mem_out_wire[559]), .S(n1835), .Z(
        \Data_Mem/n5703 ) );
  MUX U3386 ( .A(reg_target[14]), .B(data_mem_out_wire[558]), .S(n1835), .Z(
        \Data_Mem/n5702 ) );
  MUX U3387 ( .A(reg_target[13]), .B(data_mem_out_wire[557]), .S(n1835), .Z(
        \Data_Mem/n5701 ) );
  MUX U3388 ( .A(reg_target[12]), .B(data_mem_out_wire[556]), .S(n1835), .Z(
        \Data_Mem/n5700 ) );
  MUX U3389 ( .A(reg_target[11]), .B(data_mem_out_wire[555]), .S(n1835), .Z(
        \Data_Mem/n5699 ) );
  MUX U3390 ( .A(reg_target[10]), .B(data_mem_out_wire[554]), .S(n1835), .Z(
        \Data_Mem/n5698 ) );
  MUX U3391 ( .A(reg_target[9]), .B(data_mem_out_wire[553]), .S(n1835), .Z(
        \Data_Mem/n5697 ) );
  MUX U3392 ( .A(reg_target[8]), .B(data_mem_out_wire[552]), .S(n1835), .Z(
        \Data_Mem/n5696 ) );
  MUX U3393 ( .A(reg_target[7]), .B(data_mem_out_wire[551]), .S(n1835), .Z(
        \Data_Mem/n5695 ) );
  MUX U3394 ( .A(reg_target[6]), .B(data_mem_out_wire[550]), .S(n1835), .Z(
        \Data_Mem/n5694 ) );
  MUX U3395 ( .A(reg_target[5]), .B(data_mem_out_wire[549]), .S(n1835), .Z(
        \Data_Mem/n5693 ) );
  MUX U3396 ( .A(reg_target[4]), .B(data_mem_out_wire[548]), .S(n1835), .Z(
        \Data_Mem/n5692 ) );
  MUX U3397 ( .A(reg_target[3]), .B(data_mem_out_wire[547]), .S(n1835), .Z(
        \Data_Mem/n5691 ) );
  MUX U3398 ( .A(reg_target[2]), .B(data_mem_out_wire[546]), .S(n1835), .Z(
        \Data_Mem/n5690 ) );
  IV U3399 ( .A(n1836), .Z(n1835) );
  MUX U3400 ( .A(data_mem_out_wire[545]), .B(reg_target[1]), .S(n1836), .Z(
        \Data_Mem/n5689 ) );
  MUX U3401 ( .A(data_mem_out_wire[544]), .B(reg_target[0]), .S(n1836), .Z(
        \Data_Mem/n5688 ) );
  AND U3402 ( .A(n1795), .B(n1834), .Z(n1836) );
  MUX U3403 ( .A(reg_target[31]), .B(data_mem_out_wire[607]), .S(n1837), .Z(
        \Data_Mem/n5687 ) );
  MUX U3404 ( .A(reg_target[30]), .B(data_mem_out_wire[606]), .S(n1837), .Z(
        \Data_Mem/n5686 ) );
  MUX U3405 ( .A(reg_target[29]), .B(data_mem_out_wire[605]), .S(n1837), .Z(
        \Data_Mem/n5685 ) );
  MUX U3406 ( .A(reg_target[28]), .B(data_mem_out_wire[604]), .S(n1837), .Z(
        \Data_Mem/n5684 ) );
  MUX U3407 ( .A(reg_target[27]), .B(data_mem_out_wire[603]), .S(n1837), .Z(
        \Data_Mem/n5683 ) );
  MUX U3408 ( .A(reg_target[26]), .B(data_mem_out_wire[602]), .S(n1837), .Z(
        \Data_Mem/n5682 ) );
  MUX U3409 ( .A(reg_target[25]), .B(data_mem_out_wire[601]), .S(n1837), .Z(
        \Data_Mem/n5681 ) );
  MUX U3410 ( .A(reg_target[24]), .B(data_mem_out_wire[600]), .S(n1837), .Z(
        \Data_Mem/n5680 ) );
  MUX U3411 ( .A(reg_target[23]), .B(data_mem_out_wire[599]), .S(n1837), .Z(
        \Data_Mem/n5679 ) );
  MUX U3412 ( .A(reg_target[22]), .B(data_mem_out_wire[598]), .S(n1837), .Z(
        \Data_Mem/n5678 ) );
  MUX U3413 ( .A(reg_target[21]), .B(data_mem_out_wire[597]), .S(n1837), .Z(
        \Data_Mem/n5677 ) );
  MUX U3414 ( .A(reg_target[20]), .B(data_mem_out_wire[596]), .S(n1837), .Z(
        \Data_Mem/n5676 ) );
  MUX U3415 ( .A(reg_target[19]), .B(data_mem_out_wire[595]), .S(n1837), .Z(
        \Data_Mem/n5675 ) );
  MUX U3416 ( .A(reg_target[18]), .B(data_mem_out_wire[594]), .S(n1837), .Z(
        \Data_Mem/n5674 ) );
  MUX U3417 ( .A(reg_target[17]), .B(data_mem_out_wire[593]), .S(n1837), .Z(
        \Data_Mem/n5673 ) );
  MUX U3418 ( .A(reg_target[16]), .B(data_mem_out_wire[592]), .S(n1837), .Z(
        \Data_Mem/n5672 ) );
  MUX U3419 ( .A(reg_target[15]), .B(data_mem_out_wire[591]), .S(n1837), .Z(
        \Data_Mem/n5671 ) );
  MUX U3420 ( .A(reg_target[14]), .B(data_mem_out_wire[590]), .S(n1837), .Z(
        \Data_Mem/n5670 ) );
  MUX U3421 ( .A(reg_target[13]), .B(data_mem_out_wire[589]), .S(n1837), .Z(
        \Data_Mem/n5669 ) );
  MUX U3422 ( .A(reg_target[12]), .B(data_mem_out_wire[588]), .S(n1837), .Z(
        \Data_Mem/n5668 ) );
  MUX U3423 ( .A(reg_target[11]), .B(data_mem_out_wire[587]), .S(n1837), .Z(
        \Data_Mem/n5667 ) );
  MUX U3424 ( .A(reg_target[10]), .B(data_mem_out_wire[586]), .S(n1837), .Z(
        \Data_Mem/n5666 ) );
  MUX U3425 ( .A(reg_target[9]), .B(data_mem_out_wire[585]), .S(n1837), .Z(
        \Data_Mem/n5665 ) );
  MUX U3426 ( .A(reg_target[8]), .B(data_mem_out_wire[584]), .S(n1837), .Z(
        \Data_Mem/n5664 ) );
  MUX U3427 ( .A(reg_target[7]), .B(data_mem_out_wire[583]), .S(n1837), .Z(
        \Data_Mem/n5663 ) );
  MUX U3428 ( .A(reg_target[6]), .B(data_mem_out_wire[582]), .S(n1837), .Z(
        \Data_Mem/n5662 ) );
  MUX U3429 ( .A(reg_target[5]), .B(data_mem_out_wire[581]), .S(n1837), .Z(
        \Data_Mem/n5661 ) );
  MUX U3430 ( .A(reg_target[4]), .B(data_mem_out_wire[580]), .S(n1837), .Z(
        \Data_Mem/n5660 ) );
  MUX U3431 ( .A(reg_target[3]), .B(data_mem_out_wire[579]), .S(n1837), .Z(
        \Data_Mem/n5659 ) );
  MUX U3432 ( .A(reg_target[2]), .B(data_mem_out_wire[578]), .S(n1837), .Z(
        \Data_Mem/n5658 ) );
  IV U3433 ( .A(n1838), .Z(n1837) );
  MUX U3434 ( .A(data_mem_out_wire[577]), .B(reg_target[1]), .S(n1838), .Z(
        \Data_Mem/n5657 ) );
  MUX U3435 ( .A(data_mem_out_wire[576]), .B(reg_target[0]), .S(n1838), .Z(
        \Data_Mem/n5656 ) );
  AND U3436 ( .A(n1798), .B(n1834), .Z(n1838) );
  MUX U3437 ( .A(reg_target[31]), .B(data_mem_out_wire[639]), .S(n1839), .Z(
        \Data_Mem/n5655 ) );
  MUX U3438 ( .A(reg_target[30]), .B(data_mem_out_wire[638]), .S(n1839), .Z(
        \Data_Mem/n5654 ) );
  MUX U3439 ( .A(reg_target[29]), .B(data_mem_out_wire[637]), .S(n1839), .Z(
        \Data_Mem/n5653 ) );
  MUX U3440 ( .A(reg_target[28]), .B(data_mem_out_wire[636]), .S(n1839), .Z(
        \Data_Mem/n5652 ) );
  MUX U3441 ( .A(reg_target[27]), .B(data_mem_out_wire[635]), .S(n1839), .Z(
        \Data_Mem/n5651 ) );
  MUX U3442 ( .A(reg_target[26]), .B(data_mem_out_wire[634]), .S(n1839), .Z(
        \Data_Mem/n5650 ) );
  MUX U3443 ( .A(reg_target[25]), .B(data_mem_out_wire[633]), .S(n1839), .Z(
        \Data_Mem/n5649 ) );
  MUX U3444 ( .A(reg_target[24]), .B(data_mem_out_wire[632]), .S(n1839), .Z(
        \Data_Mem/n5648 ) );
  MUX U3445 ( .A(reg_target[23]), .B(data_mem_out_wire[631]), .S(n1839), .Z(
        \Data_Mem/n5647 ) );
  MUX U3446 ( .A(reg_target[22]), .B(data_mem_out_wire[630]), .S(n1839), .Z(
        \Data_Mem/n5646 ) );
  MUX U3447 ( .A(reg_target[21]), .B(data_mem_out_wire[629]), .S(n1839), .Z(
        \Data_Mem/n5645 ) );
  MUX U3448 ( .A(reg_target[20]), .B(data_mem_out_wire[628]), .S(n1839), .Z(
        \Data_Mem/n5644 ) );
  MUX U3449 ( .A(reg_target[19]), .B(data_mem_out_wire[627]), .S(n1839), .Z(
        \Data_Mem/n5643 ) );
  MUX U3450 ( .A(reg_target[18]), .B(data_mem_out_wire[626]), .S(n1839), .Z(
        \Data_Mem/n5642 ) );
  MUX U3451 ( .A(reg_target[17]), .B(data_mem_out_wire[625]), .S(n1839), .Z(
        \Data_Mem/n5641 ) );
  MUX U3452 ( .A(reg_target[16]), .B(data_mem_out_wire[624]), .S(n1839), .Z(
        \Data_Mem/n5640 ) );
  MUX U3453 ( .A(reg_target[15]), .B(data_mem_out_wire[623]), .S(n1839), .Z(
        \Data_Mem/n5639 ) );
  MUX U3454 ( .A(reg_target[14]), .B(data_mem_out_wire[622]), .S(n1839), .Z(
        \Data_Mem/n5638 ) );
  MUX U3455 ( .A(reg_target[13]), .B(data_mem_out_wire[621]), .S(n1839), .Z(
        \Data_Mem/n5637 ) );
  MUX U3456 ( .A(reg_target[12]), .B(data_mem_out_wire[620]), .S(n1839), .Z(
        \Data_Mem/n5636 ) );
  MUX U3457 ( .A(reg_target[11]), .B(data_mem_out_wire[619]), .S(n1839), .Z(
        \Data_Mem/n5635 ) );
  MUX U3458 ( .A(reg_target[10]), .B(data_mem_out_wire[618]), .S(n1839), .Z(
        \Data_Mem/n5634 ) );
  MUX U3459 ( .A(reg_target[9]), .B(data_mem_out_wire[617]), .S(n1839), .Z(
        \Data_Mem/n5633 ) );
  MUX U3460 ( .A(reg_target[8]), .B(data_mem_out_wire[616]), .S(n1839), .Z(
        \Data_Mem/n5632 ) );
  MUX U3461 ( .A(reg_target[7]), .B(data_mem_out_wire[615]), .S(n1839), .Z(
        \Data_Mem/n5631 ) );
  MUX U3462 ( .A(reg_target[6]), .B(data_mem_out_wire[614]), .S(n1839), .Z(
        \Data_Mem/n5630 ) );
  MUX U3463 ( .A(reg_target[5]), .B(data_mem_out_wire[613]), .S(n1839), .Z(
        \Data_Mem/n5629 ) );
  MUX U3464 ( .A(reg_target[4]), .B(data_mem_out_wire[612]), .S(n1839), .Z(
        \Data_Mem/n5628 ) );
  MUX U3465 ( .A(reg_target[3]), .B(data_mem_out_wire[611]), .S(n1839), .Z(
        \Data_Mem/n5627 ) );
  MUX U3466 ( .A(reg_target[2]), .B(data_mem_out_wire[610]), .S(n1839), .Z(
        \Data_Mem/n5626 ) );
  IV U3467 ( .A(n1840), .Z(n1839) );
  MUX U3468 ( .A(data_mem_out_wire[609]), .B(reg_target[1]), .S(n1840), .Z(
        \Data_Mem/n5625 ) );
  MUX U3469 ( .A(data_mem_out_wire[608]), .B(reg_target[0]), .S(n1840), .Z(
        \Data_Mem/n5624 ) );
  AND U3470 ( .A(n1801), .B(n1834), .Z(n1840) );
  MUX U3471 ( .A(reg_target[31]), .B(data_mem_out_wire[671]), .S(n1841), .Z(
        \Data_Mem/n5623 ) );
  MUX U3472 ( .A(reg_target[30]), .B(data_mem_out_wire[670]), .S(n1841), .Z(
        \Data_Mem/n5622 ) );
  MUX U3473 ( .A(reg_target[29]), .B(data_mem_out_wire[669]), .S(n1841), .Z(
        \Data_Mem/n5621 ) );
  MUX U3474 ( .A(reg_target[28]), .B(data_mem_out_wire[668]), .S(n1841), .Z(
        \Data_Mem/n5620 ) );
  MUX U3475 ( .A(reg_target[27]), .B(data_mem_out_wire[667]), .S(n1841), .Z(
        \Data_Mem/n5619 ) );
  MUX U3476 ( .A(reg_target[26]), .B(data_mem_out_wire[666]), .S(n1841), .Z(
        \Data_Mem/n5618 ) );
  MUX U3477 ( .A(reg_target[25]), .B(data_mem_out_wire[665]), .S(n1841), .Z(
        \Data_Mem/n5617 ) );
  MUX U3478 ( .A(reg_target[24]), .B(data_mem_out_wire[664]), .S(n1841), .Z(
        \Data_Mem/n5616 ) );
  MUX U3479 ( .A(reg_target[23]), .B(data_mem_out_wire[663]), .S(n1841), .Z(
        \Data_Mem/n5615 ) );
  MUX U3480 ( .A(reg_target[22]), .B(data_mem_out_wire[662]), .S(n1841), .Z(
        \Data_Mem/n5614 ) );
  MUX U3481 ( .A(reg_target[21]), .B(data_mem_out_wire[661]), .S(n1841), .Z(
        \Data_Mem/n5613 ) );
  MUX U3482 ( .A(reg_target[20]), .B(data_mem_out_wire[660]), .S(n1841), .Z(
        \Data_Mem/n5612 ) );
  MUX U3483 ( .A(reg_target[19]), .B(data_mem_out_wire[659]), .S(n1841), .Z(
        \Data_Mem/n5611 ) );
  MUX U3484 ( .A(reg_target[18]), .B(data_mem_out_wire[658]), .S(n1841), .Z(
        \Data_Mem/n5610 ) );
  MUX U3485 ( .A(reg_target[17]), .B(data_mem_out_wire[657]), .S(n1841), .Z(
        \Data_Mem/n5609 ) );
  MUX U3486 ( .A(reg_target[16]), .B(data_mem_out_wire[656]), .S(n1841), .Z(
        \Data_Mem/n5608 ) );
  MUX U3487 ( .A(reg_target[15]), .B(data_mem_out_wire[655]), .S(n1841), .Z(
        \Data_Mem/n5607 ) );
  MUX U3488 ( .A(reg_target[14]), .B(data_mem_out_wire[654]), .S(n1841), .Z(
        \Data_Mem/n5606 ) );
  MUX U3489 ( .A(reg_target[13]), .B(data_mem_out_wire[653]), .S(n1841), .Z(
        \Data_Mem/n5605 ) );
  MUX U3490 ( .A(reg_target[12]), .B(data_mem_out_wire[652]), .S(n1841), .Z(
        \Data_Mem/n5604 ) );
  MUX U3491 ( .A(reg_target[11]), .B(data_mem_out_wire[651]), .S(n1841), .Z(
        \Data_Mem/n5603 ) );
  MUX U3492 ( .A(reg_target[10]), .B(data_mem_out_wire[650]), .S(n1841), .Z(
        \Data_Mem/n5602 ) );
  MUX U3493 ( .A(reg_target[9]), .B(data_mem_out_wire[649]), .S(n1841), .Z(
        \Data_Mem/n5601 ) );
  MUX U3494 ( .A(reg_target[8]), .B(data_mem_out_wire[648]), .S(n1841), .Z(
        \Data_Mem/n5600 ) );
  MUX U3495 ( .A(reg_target[7]), .B(data_mem_out_wire[647]), .S(n1841), .Z(
        \Data_Mem/n5599 ) );
  MUX U3496 ( .A(reg_target[6]), .B(data_mem_out_wire[646]), .S(n1841), .Z(
        \Data_Mem/n5598 ) );
  MUX U3497 ( .A(reg_target[5]), .B(data_mem_out_wire[645]), .S(n1841), .Z(
        \Data_Mem/n5597 ) );
  MUX U3498 ( .A(reg_target[4]), .B(data_mem_out_wire[644]), .S(n1841), .Z(
        \Data_Mem/n5596 ) );
  MUX U3499 ( .A(reg_target[3]), .B(data_mem_out_wire[643]), .S(n1841), .Z(
        \Data_Mem/n5595 ) );
  MUX U3500 ( .A(reg_target[2]), .B(data_mem_out_wire[642]), .S(n1841), .Z(
        \Data_Mem/n5594 ) );
  IV U3501 ( .A(n1842), .Z(n1841) );
  MUX U3502 ( .A(data_mem_out_wire[641]), .B(reg_target[1]), .S(n1842), .Z(
        \Data_Mem/n5593 ) );
  MUX U3503 ( .A(data_mem_out_wire[640]), .B(reg_target[0]), .S(n1842), .Z(
        \Data_Mem/n5592 ) );
  AND U3504 ( .A(n1804), .B(n1834), .Z(n1842) );
  MUX U3505 ( .A(reg_target[31]), .B(data_mem_out_wire[703]), .S(n1843), .Z(
        \Data_Mem/n5591 ) );
  MUX U3506 ( .A(reg_target[30]), .B(data_mem_out_wire[702]), .S(n1843), .Z(
        \Data_Mem/n5590 ) );
  MUX U3507 ( .A(reg_target[29]), .B(data_mem_out_wire[701]), .S(n1843), .Z(
        \Data_Mem/n5589 ) );
  MUX U3508 ( .A(reg_target[28]), .B(data_mem_out_wire[700]), .S(n1843), .Z(
        \Data_Mem/n5588 ) );
  MUX U3509 ( .A(reg_target[27]), .B(data_mem_out_wire[699]), .S(n1843), .Z(
        \Data_Mem/n5587 ) );
  MUX U3510 ( .A(reg_target[26]), .B(data_mem_out_wire[698]), .S(n1843), .Z(
        \Data_Mem/n5586 ) );
  MUX U3511 ( .A(reg_target[25]), .B(data_mem_out_wire[697]), .S(n1843), .Z(
        \Data_Mem/n5585 ) );
  MUX U3512 ( .A(reg_target[24]), .B(data_mem_out_wire[696]), .S(n1843), .Z(
        \Data_Mem/n5584 ) );
  MUX U3513 ( .A(reg_target[23]), .B(data_mem_out_wire[695]), .S(n1843), .Z(
        \Data_Mem/n5583 ) );
  MUX U3514 ( .A(reg_target[22]), .B(data_mem_out_wire[694]), .S(n1843), .Z(
        \Data_Mem/n5582 ) );
  MUX U3515 ( .A(reg_target[21]), .B(data_mem_out_wire[693]), .S(n1843), .Z(
        \Data_Mem/n5581 ) );
  MUX U3516 ( .A(reg_target[20]), .B(data_mem_out_wire[692]), .S(n1843), .Z(
        \Data_Mem/n5580 ) );
  MUX U3517 ( .A(reg_target[19]), .B(data_mem_out_wire[691]), .S(n1843), .Z(
        \Data_Mem/n5579 ) );
  MUX U3518 ( .A(reg_target[18]), .B(data_mem_out_wire[690]), .S(n1843), .Z(
        \Data_Mem/n5578 ) );
  MUX U3519 ( .A(reg_target[17]), .B(data_mem_out_wire[689]), .S(n1843), .Z(
        \Data_Mem/n5577 ) );
  MUX U3520 ( .A(reg_target[16]), .B(data_mem_out_wire[688]), .S(n1843), .Z(
        \Data_Mem/n5576 ) );
  MUX U3521 ( .A(reg_target[15]), .B(data_mem_out_wire[687]), .S(n1843), .Z(
        \Data_Mem/n5575 ) );
  MUX U3522 ( .A(reg_target[14]), .B(data_mem_out_wire[686]), .S(n1843), .Z(
        \Data_Mem/n5574 ) );
  MUX U3523 ( .A(reg_target[13]), .B(data_mem_out_wire[685]), .S(n1843), .Z(
        \Data_Mem/n5573 ) );
  MUX U3524 ( .A(reg_target[12]), .B(data_mem_out_wire[684]), .S(n1843), .Z(
        \Data_Mem/n5572 ) );
  MUX U3525 ( .A(reg_target[11]), .B(data_mem_out_wire[683]), .S(n1843), .Z(
        \Data_Mem/n5571 ) );
  MUX U3526 ( .A(reg_target[10]), .B(data_mem_out_wire[682]), .S(n1843), .Z(
        \Data_Mem/n5570 ) );
  MUX U3527 ( .A(reg_target[9]), .B(data_mem_out_wire[681]), .S(n1843), .Z(
        \Data_Mem/n5569 ) );
  MUX U3528 ( .A(reg_target[8]), .B(data_mem_out_wire[680]), .S(n1843), .Z(
        \Data_Mem/n5568 ) );
  MUX U3529 ( .A(reg_target[7]), .B(data_mem_out_wire[679]), .S(n1843), .Z(
        \Data_Mem/n5567 ) );
  MUX U3530 ( .A(reg_target[6]), .B(data_mem_out_wire[678]), .S(n1843), .Z(
        \Data_Mem/n5566 ) );
  MUX U3531 ( .A(reg_target[5]), .B(data_mem_out_wire[677]), .S(n1843), .Z(
        \Data_Mem/n5565 ) );
  MUX U3532 ( .A(reg_target[4]), .B(data_mem_out_wire[676]), .S(n1843), .Z(
        \Data_Mem/n5564 ) );
  MUX U3533 ( .A(reg_target[3]), .B(data_mem_out_wire[675]), .S(n1843), .Z(
        \Data_Mem/n5563 ) );
  MUX U3534 ( .A(reg_target[2]), .B(data_mem_out_wire[674]), .S(n1843), .Z(
        \Data_Mem/n5562 ) );
  IV U3535 ( .A(n1844), .Z(n1843) );
  MUX U3536 ( .A(data_mem_out_wire[673]), .B(reg_target[1]), .S(n1844), .Z(
        \Data_Mem/n5561 ) );
  MUX U3537 ( .A(data_mem_out_wire[672]), .B(reg_target[0]), .S(n1844), .Z(
        \Data_Mem/n5560 ) );
  AND U3538 ( .A(n1807), .B(n1834), .Z(n1844) );
  MUX U3539 ( .A(reg_target[31]), .B(data_mem_out_wire[735]), .S(n1845), .Z(
        \Data_Mem/n5559 ) );
  MUX U3540 ( .A(reg_target[30]), .B(data_mem_out_wire[734]), .S(n1845), .Z(
        \Data_Mem/n5558 ) );
  MUX U3541 ( .A(reg_target[29]), .B(data_mem_out_wire[733]), .S(n1845), .Z(
        \Data_Mem/n5557 ) );
  MUX U3542 ( .A(reg_target[28]), .B(data_mem_out_wire[732]), .S(n1845), .Z(
        \Data_Mem/n5556 ) );
  MUX U3543 ( .A(reg_target[27]), .B(data_mem_out_wire[731]), .S(n1845), .Z(
        \Data_Mem/n5555 ) );
  MUX U3544 ( .A(reg_target[26]), .B(data_mem_out_wire[730]), .S(n1845), .Z(
        \Data_Mem/n5554 ) );
  MUX U3545 ( .A(reg_target[25]), .B(data_mem_out_wire[729]), .S(n1845), .Z(
        \Data_Mem/n5553 ) );
  MUX U3546 ( .A(reg_target[24]), .B(data_mem_out_wire[728]), .S(n1845), .Z(
        \Data_Mem/n5552 ) );
  MUX U3547 ( .A(reg_target[23]), .B(data_mem_out_wire[727]), .S(n1845), .Z(
        \Data_Mem/n5551 ) );
  MUX U3548 ( .A(reg_target[22]), .B(data_mem_out_wire[726]), .S(n1845), .Z(
        \Data_Mem/n5550 ) );
  MUX U3549 ( .A(reg_target[21]), .B(data_mem_out_wire[725]), .S(n1845), .Z(
        \Data_Mem/n5549 ) );
  MUX U3550 ( .A(reg_target[20]), .B(data_mem_out_wire[724]), .S(n1845), .Z(
        \Data_Mem/n5548 ) );
  MUX U3551 ( .A(reg_target[19]), .B(data_mem_out_wire[723]), .S(n1845), .Z(
        \Data_Mem/n5547 ) );
  MUX U3552 ( .A(reg_target[18]), .B(data_mem_out_wire[722]), .S(n1845), .Z(
        \Data_Mem/n5546 ) );
  MUX U3553 ( .A(reg_target[17]), .B(data_mem_out_wire[721]), .S(n1845), .Z(
        \Data_Mem/n5545 ) );
  MUX U3554 ( .A(reg_target[16]), .B(data_mem_out_wire[720]), .S(n1845), .Z(
        \Data_Mem/n5544 ) );
  MUX U3555 ( .A(reg_target[15]), .B(data_mem_out_wire[719]), .S(n1845), .Z(
        \Data_Mem/n5543 ) );
  MUX U3556 ( .A(reg_target[14]), .B(data_mem_out_wire[718]), .S(n1845), .Z(
        \Data_Mem/n5542 ) );
  MUX U3557 ( .A(reg_target[13]), .B(data_mem_out_wire[717]), .S(n1845), .Z(
        \Data_Mem/n5541 ) );
  MUX U3558 ( .A(reg_target[12]), .B(data_mem_out_wire[716]), .S(n1845), .Z(
        \Data_Mem/n5540 ) );
  MUX U3559 ( .A(reg_target[11]), .B(data_mem_out_wire[715]), .S(n1845), .Z(
        \Data_Mem/n5539 ) );
  MUX U3560 ( .A(reg_target[10]), .B(data_mem_out_wire[714]), .S(n1845), .Z(
        \Data_Mem/n5538 ) );
  MUX U3561 ( .A(reg_target[9]), .B(data_mem_out_wire[713]), .S(n1845), .Z(
        \Data_Mem/n5537 ) );
  MUX U3562 ( .A(reg_target[8]), .B(data_mem_out_wire[712]), .S(n1845), .Z(
        \Data_Mem/n5536 ) );
  MUX U3563 ( .A(reg_target[7]), .B(data_mem_out_wire[711]), .S(n1845), .Z(
        \Data_Mem/n5535 ) );
  MUX U3564 ( .A(reg_target[6]), .B(data_mem_out_wire[710]), .S(n1845), .Z(
        \Data_Mem/n5534 ) );
  MUX U3565 ( .A(reg_target[5]), .B(data_mem_out_wire[709]), .S(n1845), .Z(
        \Data_Mem/n5533 ) );
  MUX U3566 ( .A(reg_target[4]), .B(data_mem_out_wire[708]), .S(n1845), .Z(
        \Data_Mem/n5532 ) );
  MUX U3567 ( .A(reg_target[3]), .B(data_mem_out_wire[707]), .S(n1845), .Z(
        \Data_Mem/n5531 ) );
  MUX U3568 ( .A(reg_target[2]), .B(data_mem_out_wire[706]), .S(n1845), .Z(
        \Data_Mem/n5530 ) );
  IV U3569 ( .A(n1846), .Z(n1845) );
  MUX U3570 ( .A(data_mem_out_wire[705]), .B(reg_target[1]), .S(n1846), .Z(
        \Data_Mem/n5529 ) );
  MUX U3571 ( .A(data_mem_out_wire[704]), .B(reg_target[0]), .S(n1846), .Z(
        \Data_Mem/n5528 ) );
  AND U3572 ( .A(n1810), .B(n1834), .Z(n1846) );
  MUX U3573 ( .A(data_mem_out_wire[767]), .B(reg_target[31]), .S(n1847), .Z(
        \Data_Mem/n5527 ) );
  MUX U3574 ( .A(data_mem_out_wire[766]), .B(reg_target[30]), .S(n1847), .Z(
        \Data_Mem/n5526 ) );
  MUX U3575 ( .A(data_mem_out_wire[765]), .B(reg_target[29]), .S(n1847), .Z(
        \Data_Mem/n5525 ) );
  MUX U3576 ( .A(data_mem_out_wire[764]), .B(reg_target[28]), .S(n1847), .Z(
        \Data_Mem/n5524 ) );
  MUX U3577 ( .A(data_mem_out_wire[763]), .B(reg_target[27]), .S(n1847), .Z(
        \Data_Mem/n5523 ) );
  MUX U3578 ( .A(data_mem_out_wire[762]), .B(reg_target[26]), .S(n1847), .Z(
        \Data_Mem/n5522 ) );
  MUX U3579 ( .A(data_mem_out_wire[761]), .B(reg_target[25]), .S(n1847), .Z(
        \Data_Mem/n5521 ) );
  MUX U3580 ( .A(data_mem_out_wire[760]), .B(reg_target[24]), .S(n1847), .Z(
        \Data_Mem/n5520 ) );
  MUX U3581 ( .A(data_mem_out_wire[759]), .B(reg_target[23]), .S(n1847), .Z(
        \Data_Mem/n5519 ) );
  MUX U3582 ( .A(data_mem_out_wire[758]), .B(reg_target[22]), .S(n1847), .Z(
        \Data_Mem/n5518 ) );
  MUX U3583 ( .A(data_mem_out_wire[757]), .B(reg_target[21]), .S(n1847), .Z(
        \Data_Mem/n5517 ) );
  MUX U3584 ( .A(data_mem_out_wire[756]), .B(reg_target[20]), .S(n1847), .Z(
        \Data_Mem/n5516 ) );
  MUX U3585 ( .A(data_mem_out_wire[755]), .B(reg_target[19]), .S(n1847), .Z(
        \Data_Mem/n5515 ) );
  MUX U3586 ( .A(data_mem_out_wire[754]), .B(reg_target[18]), .S(n1847), .Z(
        \Data_Mem/n5514 ) );
  MUX U3587 ( .A(data_mem_out_wire[753]), .B(reg_target[17]), .S(n1847), .Z(
        \Data_Mem/n5513 ) );
  MUX U3588 ( .A(data_mem_out_wire[752]), .B(reg_target[16]), .S(n1847), .Z(
        \Data_Mem/n5512 ) );
  MUX U3589 ( .A(data_mem_out_wire[751]), .B(reg_target[15]), .S(n1847), .Z(
        \Data_Mem/n5511 ) );
  MUX U3590 ( .A(data_mem_out_wire[750]), .B(reg_target[14]), .S(n1847), .Z(
        \Data_Mem/n5510 ) );
  MUX U3591 ( .A(data_mem_out_wire[749]), .B(reg_target[13]), .S(n1847), .Z(
        \Data_Mem/n5509 ) );
  MUX U3592 ( .A(data_mem_out_wire[748]), .B(reg_target[12]), .S(n1847), .Z(
        \Data_Mem/n5508 ) );
  MUX U3593 ( .A(data_mem_out_wire[747]), .B(reg_target[11]), .S(n1847), .Z(
        \Data_Mem/n5507 ) );
  MUX U3594 ( .A(data_mem_out_wire[746]), .B(reg_target[10]), .S(n1847), .Z(
        \Data_Mem/n5506 ) );
  MUX U3595 ( .A(data_mem_out_wire[745]), .B(reg_target[9]), .S(n1847), .Z(
        \Data_Mem/n5505 ) );
  MUX U3596 ( .A(data_mem_out_wire[744]), .B(reg_target[8]), .S(n1847), .Z(
        \Data_Mem/n5504 ) );
  MUX U3597 ( .A(data_mem_out_wire[743]), .B(reg_target[7]), .S(n1847), .Z(
        \Data_Mem/n5503 ) );
  MUX U3598 ( .A(data_mem_out_wire[742]), .B(reg_target[6]), .S(n1847), .Z(
        \Data_Mem/n5502 ) );
  MUX U3599 ( .A(data_mem_out_wire[741]), .B(reg_target[5]), .S(n1847), .Z(
        \Data_Mem/n5501 ) );
  MUX U3600 ( .A(data_mem_out_wire[740]), .B(reg_target[4]), .S(n1847), .Z(
        \Data_Mem/n5500 ) );
  MUX U3601 ( .A(data_mem_out_wire[739]), .B(reg_target[3]), .S(n1847), .Z(
        \Data_Mem/n5499 ) );
  MUX U3602 ( .A(data_mem_out_wire[738]), .B(reg_target[2]), .S(n1847), .Z(
        \Data_Mem/n5498 ) );
  MUX U3603 ( .A(data_mem_out_wire[737]), .B(reg_target[1]), .S(n1847), .Z(
        \Data_Mem/n5497 ) );
  MUX U3604 ( .A(data_mem_out_wire[736]), .B(reg_target[0]), .S(n1847), .Z(
        \Data_Mem/n5496 ) );
  AND U3605 ( .A(n1834), .B(n1830), .Z(n1847) );
  ANDN U3606 ( .B(n1848), .A(N24), .Z(n1834) );
  MUX U3607 ( .A(reg_target[31]), .B(data_mem_out_wire[799]), .S(n1849), .Z(
        \Data_Mem/n5495 ) );
  MUX U3608 ( .A(reg_target[30]), .B(data_mem_out_wire[798]), .S(n1849), .Z(
        \Data_Mem/n5494 ) );
  MUX U3609 ( .A(reg_target[29]), .B(data_mem_out_wire[797]), .S(n1849), .Z(
        \Data_Mem/n5493 ) );
  MUX U3610 ( .A(reg_target[28]), .B(data_mem_out_wire[796]), .S(n1849), .Z(
        \Data_Mem/n5492 ) );
  MUX U3611 ( .A(reg_target[27]), .B(data_mem_out_wire[795]), .S(n1849), .Z(
        \Data_Mem/n5491 ) );
  MUX U3612 ( .A(reg_target[26]), .B(data_mem_out_wire[794]), .S(n1849), .Z(
        \Data_Mem/n5490 ) );
  MUX U3613 ( .A(reg_target[25]), .B(data_mem_out_wire[793]), .S(n1849), .Z(
        \Data_Mem/n5489 ) );
  MUX U3614 ( .A(reg_target[24]), .B(data_mem_out_wire[792]), .S(n1849), .Z(
        \Data_Mem/n5488 ) );
  MUX U3615 ( .A(reg_target[23]), .B(data_mem_out_wire[791]), .S(n1849), .Z(
        \Data_Mem/n5487 ) );
  MUX U3616 ( .A(reg_target[22]), .B(data_mem_out_wire[790]), .S(n1849), .Z(
        \Data_Mem/n5486 ) );
  MUX U3617 ( .A(reg_target[21]), .B(data_mem_out_wire[789]), .S(n1849), .Z(
        \Data_Mem/n5485 ) );
  MUX U3618 ( .A(reg_target[20]), .B(data_mem_out_wire[788]), .S(n1849), .Z(
        \Data_Mem/n5484 ) );
  MUX U3619 ( .A(reg_target[19]), .B(data_mem_out_wire[787]), .S(n1849), .Z(
        \Data_Mem/n5483 ) );
  MUX U3620 ( .A(reg_target[18]), .B(data_mem_out_wire[786]), .S(n1849), .Z(
        \Data_Mem/n5482 ) );
  MUX U3621 ( .A(reg_target[17]), .B(data_mem_out_wire[785]), .S(n1849), .Z(
        \Data_Mem/n5481 ) );
  MUX U3622 ( .A(reg_target[16]), .B(data_mem_out_wire[784]), .S(n1849), .Z(
        \Data_Mem/n5480 ) );
  MUX U3623 ( .A(reg_target[15]), .B(data_mem_out_wire[783]), .S(n1849), .Z(
        \Data_Mem/n5479 ) );
  MUX U3624 ( .A(reg_target[14]), .B(data_mem_out_wire[782]), .S(n1849), .Z(
        \Data_Mem/n5478 ) );
  MUX U3625 ( .A(reg_target[13]), .B(data_mem_out_wire[781]), .S(n1849), .Z(
        \Data_Mem/n5477 ) );
  MUX U3626 ( .A(reg_target[12]), .B(data_mem_out_wire[780]), .S(n1849), .Z(
        \Data_Mem/n5476 ) );
  MUX U3627 ( .A(reg_target[11]), .B(data_mem_out_wire[779]), .S(n1849), .Z(
        \Data_Mem/n5475 ) );
  MUX U3628 ( .A(reg_target[10]), .B(data_mem_out_wire[778]), .S(n1849), .Z(
        \Data_Mem/n5474 ) );
  MUX U3629 ( .A(reg_target[9]), .B(data_mem_out_wire[777]), .S(n1849), .Z(
        \Data_Mem/n5473 ) );
  MUX U3630 ( .A(reg_target[8]), .B(data_mem_out_wire[776]), .S(n1849), .Z(
        \Data_Mem/n5472 ) );
  MUX U3631 ( .A(reg_target[7]), .B(data_mem_out_wire[775]), .S(n1849), .Z(
        \Data_Mem/n5471 ) );
  MUX U3632 ( .A(reg_target[6]), .B(data_mem_out_wire[774]), .S(n1849), .Z(
        \Data_Mem/n5470 ) );
  MUX U3633 ( .A(reg_target[5]), .B(data_mem_out_wire[773]), .S(n1849), .Z(
        \Data_Mem/n5469 ) );
  MUX U3634 ( .A(reg_target[4]), .B(data_mem_out_wire[772]), .S(n1849), .Z(
        \Data_Mem/n5468 ) );
  MUX U3635 ( .A(reg_target[3]), .B(data_mem_out_wire[771]), .S(n1849), .Z(
        \Data_Mem/n5467 ) );
  MUX U3636 ( .A(reg_target[2]), .B(data_mem_out_wire[770]), .S(n1849), .Z(
        \Data_Mem/n5466 ) );
  IV U3637 ( .A(n1850), .Z(n1849) );
  MUX U3638 ( .A(data_mem_out_wire[769]), .B(reg_target[1]), .S(n1850), .Z(
        \Data_Mem/n5465 ) );
  MUX U3639 ( .A(data_mem_out_wire[768]), .B(reg_target[0]), .S(n1850), .Z(
        \Data_Mem/n5464 ) );
  AND U3640 ( .A(n1791), .B(n1851), .Z(n1850) );
  MUX U3641 ( .A(reg_target[31]), .B(data_mem_out_wire[831]), .S(n1852), .Z(
        \Data_Mem/n5463 ) );
  MUX U3642 ( .A(reg_target[30]), .B(data_mem_out_wire[830]), .S(n1852), .Z(
        \Data_Mem/n5462 ) );
  MUX U3643 ( .A(reg_target[29]), .B(data_mem_out_wire[829]), .S(n1852), .Z(
        \Data_Mem/n5461 ) );
  MUX U3644 ( .A(reg_target[28]), .B(data_mem_out_wire[828]), .S(n1852), .Z(
        \Data_Mem/n5460 ) );
  MUX U3645 ( .A(reg_target[27]), .B(data_mem_out_wire[827]), .S(n1852), .Z(
        \Data_Mem/n5459 ) );
  MUX U3646 ( .A(reg_target[26]), .B(data_mem_out_wire[826]), .S(n1852), .Z(
        \Data_Mem/n5458 ) );
  MUX U3647 ( .A(reg_target[25]), .B(data_mem_out_wire[825]), .S(n1852), .Z(
        \Data_Mem/n5457 ) );
  MUX U3648 ( .A(reg_target[24]), .B(data_mem_out_wire[824]), .S(n1852), .Z(
        \Data_Mem/n5456 ) );
  MUX U3649 ( .A(reg_target[23]), .B(data_mem_out_wire[823]), .S(n1852), .Z(
        \Data_Mem/n5455 ) );
  MUX U3650 ( .A(reg_target[22]), .B(data_mem_out_wire[822]), .S(n1852), .Z(
        \Data_Mem/n5454 ) );
  MUX U3651 ( .A(reg_target[21]), .B(data_mem_out_wire[821]), .S(n1852), .Z(
        \Data_Mem/n5453 ) );
  MUX U3652 ( .A(reg_target[20]), .B(data_mem_out_wire[820]), .S(n1852), .Z(
        \Data_Mem/n5452 ) );
  MUX U3653 ( .A(reg_target[19]), .B(data_mem_out_wire[819]), .S(n1852), .Z(
        \Data_Mem/n5451 ) );
  MUX U3654 ( .A(reg_target[18]), .B(data_mem_out_wire[818]), .S(n1852), .Z(
        \Data_Mem/n5450 ) );
  MUX U3655 ( .A(reg_target[17]), .B(data_mem_out_wire[817]), .S(n1852), .Z(
        \Data_Mem/n5449 ) );
  MUX U3656 ( .A(reg_target[16]), .B(data_mem_out_wire[816]), .S(n1852), .Z(
        \Data_Mem/n5448 ) );
  MUX U3657 ( .A(reg_target[15]), .B(data_mem_out_wire[815]), .S(n1852), .Z(
        \Data_Mem/n5447 ) );
  MUX U3658 ( .A(reg_target[14]), .B(data_mem_out_wire[814]), .S(n1852), .Z(
        \Data_Mem/n5446 ) );
  MUX U3659 ( .A(reg_target[13]), .B(data_mem_out_wire[813]), .S(n1852), .Z(
        \Data_Mem/n5445 ) );
  MUX U3660 ( .A(reg_target[12]), .B(data_mem_out_wire[812]), .S(n1852), .Z(
        \Data_Mem/n5444 ) );
  MUX U3661 ( .A(reg_target[11]), .B(data_mem_out_wire[811]), .S(n1852), .Z(
        \Data_Mem/n5443 ) );
  MUX U3662 ( .A(reg_target[10]), .B(data_mem_out_wire[810]), .S(n1852), .Z(
        \Data_Mem/n5442 ) );
  MUX U3663 ( .A(reg_target[9]), .B(data_mem_out_wire[809]), .S(n1852), .Z(
        \Data_Mem/n5441 ) );
  MUX U3664 ( .A(reg_target[8]), .B(data_mem_out_wire[808]), .S(n1852), .Z(
        \Data_Mem/n5440 ) );
  MUX U3665 ( .A(reg_target[7]), .B(data_mem_out_wire[807]), .S(n1852), .Z(
        \Data_Mem/n5439 ) );
  MUX U3666 ( .A(reg_target[6]), .B(data_mem_out_wire[806]), .S(n1852), .Z(
        \Data_Mem/n5438 ) );
  MUX U3667 ( .A(reg_target[5]), .B(data_mem_out_wire[805]), .S(n1852), .Z(
        \Data_Mem/n5437 ) );
  MUX U3668 ( .A(reg_target[4]), .B(data_mem_out_wire[804]), .S(n1852), .Z(
        \Data_Mem/n5436 ) );
  MUX U3669 ( .A(reg_target[3]), .B(data_mem_out_wire[803]), .S(n1852), .Z(
        \Data_Mem/n5435 ) );
  MUX U3670 ( .A(reg_target[2]), .B(data_mem_out_wire[802]), .S(n1852), .Z(
        \Data_Mem/n5434 ) );
  IV U3671 ( .A(n1853), .Z(n1852) );
  MUX U3672 ( .A(data_mem_out_wire[801]), .B(reg_target[1]), .S(n1853), .Z(
        \Data_Mem/n5433 ) );
  MUX U3673 ( .A(data_mem_out_wire[800]), .B(reg_target[0]), .S(n1853), .Z(
        \Data_Mem/n5432 ) );
  AND U3674 ( .A(n1795), .B(n1851), .Z(n1853) );
  MUX U3675 ( .A(reg_target[31]), .B(data_mem_out_wire[863]), .S(n1854), .Z(
        \Data_Mem/n5431 ) );
  MUX U3676 ( .A(reg_target[30]), .B(data_mem_out_wire[862]), .S(n1854), .Z(
        \Data_Mem/n5430 ) );
  MUX U3677 ( .A(reg_target[29]), .B(data_mem_out_wire[861]), .S(n1854), .Z(
        \Data_Mem/n5429 ) );
  MUX U3678 ( .A(reg_target[28]), .B(data_mem_out_wire[860]), .S(n1854), .Z(
        \Data_Mem/n5428 ) );
  MUX U3679 ( .A(reg_target[27]), .B(data_mem_out_wire[859]), .S(n1854), .Z(
        \Data_Mem/n5427 ) );
  MUX U3680 ( .A(reg_target[26]), .B(data_mem_out_wire[858]), .S(n1854), .Z(
        \Data_Mem/n5426 ) );
  MUX U3681 ( .A(reg_target[25]), .B(data_mem_out_wire[857]), .S(n1854), .Z(
        \Data_Mem/n5425 ) );
  MUX U3682 ( .A(reg_target[24]), .B(data_mem_out_wire[856]), .S(n1854), .Z(
        \Data_Mem/n5424 ) );
  MUX U3683 ( .A(reg_target[23]), .B(data_mem_out_wire[855]), .S(n1854), .Z(
        \Data_Mem/n5423 ) );
  MUX U3684 ( .A(reg_target[22]), .B(data_mem_out_wire[854]), .S(n1854), .Z(
        \Data_Mem/n5422 ) );
  MUX U3685 ( .A(reg_target[21]), .B(data_mem_out_wire[853]), .S(n1854), .Z(
        \Data_Mem/n5421 ) );
  MUX U3686 ( .A(reg_target[20]), .B(data_mem_out_wire[852]), .S(n1854), .Z(
        \Data_Mem/n5420 ) );
  MUX U3687 ( .A(reg_target[19]), .B(data_mem_out_wire[851]), .S(n1854), .Z(
        \Data_Mem/n5419 ) );
  MUX U3688 ( .A(reg_target[18]), .B(data_mem_out_wire[850]), .S(n1854), .Z(
        \Data_Mem/n5418 ) );
  MUX U3689 ( .A(reg_target[17]), .B(data_mem_out_wire[849]), .S(n1854), .Z(
        \Data_Mem/n5417 ) );
  MUX U3690 ( .A(reg_target[16]), .B(data_mem_out_wire[848]), .S(n1854), .Z(
        \Data_Mem/n5416 ) );
  MUX U3691 ( .A(reg_target[15]), .B(data_mem_out_wire[847]), .S(n1854), .Z(
        \Data_Mem/n5415 ) );
  MUX U3692 ( .A(reg_target[14]), .B(data_mem_out_wire[846]), .S(n1854), .Z(
        \Data_Mem/n5414 ) );
  MUX U3693 ( .A(reg_target[13]), .B(data_mem_out_wire[845]), .S(n1854), .Z(
        \Data_Mem/n5413 ) );
  MUX U3694 ( .A(reg_target[12]), .B(data_mem_out_wire[844]), .S(n1854), .Z(
        \Data_Mem/n5412 ) );
  MUX U3695 ( .A(reg_target[11]), .B(data_mem_out_wire[843]), .S(n1854), .Z(
        \Data_Mem/n5411 ) );
  MUX U3696 ( .A(reg_target[10]), .B(data_mem_out_wire[842]), .S(n1854), .Z(
        \Data_Mem/n5410 ) );
  MUX U3697 ( .A(reg_target[9]), .B(data_mem_out_wire[841]), .S(n1854), .Z(
        \Data_Mem/n5409 ) );
  MUX U3698 ( .A(reg_target[8]), .B(data_mem_out_wire[840]), .S(n1854), .Z(
        \Data_Mem/n5408 ) );
  MUX U3699 ( .A(reg_target[7]), .B(data_mem_out_wire[839]), .S(n1854), .Z(
        \Data_Mem/n5407 ) );
  MUX U3700 ( .A(reg_target[6]), .B(data_mem_out_wire[838]), .S(n1854), .Z(
        \Data_Mem/n5406 ) );
  MUX U3701 ( .A(reg_target[5]), .B(data_mem_out_wire[837]), .S(n1854), .Z(
        \Data_Mem/n5405 ) );
  MUX U3702 ( .A(reg_target[4]), .B(data_mem_out_wire[836]), .S(n1854), .Z(
        \Data_Mem/n5404 ) );
  MUX U3703 ( .A(reg_target[3]), .B(data_mem_out_wire[835]), .S(n1854), .Z(
        \Data_Mem/n5403 ) );
  MUX U3704 ( .A(reg_target[2]), .B(data_mem_out_wire[834]), .S(n1854), .Z(
        \Data_Mem/n5402 ) );
  IV U3705 ( .A(n1855), .Z(n1854) );
  MUX U3706 ( .A(data_mem_out_wire[833]), .B(reg_target[1]), .S(n1855), .Z(
        \Data_Mem/n5401 ) );
  MUX U3707 ( .A(data_mem_out_wire[832]), .B(reg_target[0]), .S(n1855), .Z(
        \Data_Mem/n5400 ) );
  AND U3708 ( .A(n1798), .B(n1851), .Z(n1855) );
  MUX U3709 ( .A(reg_target[31]), .B(data_mem_out_wire[895]), .S(n1856), .Z(
        \Data_Mem/n5399 ) );
  MUX U3710 ( .A(reg_target[30]), .B(data_mem_out_wire[894]), .S(n1856), .Z(
        \Data_Mem/n5398 ) );
  MUX U3711 ( .A(reg_target[29]), .B(data_mem_out_wire[893]), .S(n1856), .Z(
        \Data_Mem/n5397 ) );
  MUX U3712 ( .A(reg_target[28]), .B(data_mem_out_wire[892]), .S(n1856), .Z(
        \Data_Mem/n5396 ) );
  MUX U3713 ( .A(reg_target[27]), .B(data_mem_out_wire[891]), .S(n1856), .Z(
        \Data_Mem/n5395 ) );
  MUX U3714 ( .A(reg_target[26]), .B(data_mem_out_wire[890]), .S(n1856), .Z(
        \Data_Mem/n5394 ) );
  MUX U3715 ( .A(reg_target[25]), .B(data_mem_out_wire[889]), .S(n1856), .Z(
        \Data_Mem/n5393 ) );
  MUX U3716 ( .A(reg_target[24]), .B(data_mem_out_wire[888]), .S(n1856), .Z(
        \Data_Mem/n5392 ) );
  MUX U3717 ( .A(reg_target[23]), .B(data_mem_out_wire[887]), .S(n1856), .Z(
        \Data_Mem/n5391 ) );
  MUX U3718 ( .A(reg_target[22]), .B(data_mem_out_wire[886]), .S(n1856), .Z(
        \Data_Mem/n5390 ) );
  MUX U3719 ( .A(reg_target[21]), .B(data_mem_out_wire[885]), .S(n1856), .Z(
        \Data_Mem/n5389 ) );
  MUX U3720 ( .A(reg_target[20]), .B(data_mem_out_wire[884]), .S(n1856), .Z(
        \Data_Mem/n5388 ) );
  MUX U3721 ( .A(reg_target[19]), .B(data_mem_out_wire[883]), .S(n1856), .Z(
        \Data_Mem/n5387 ) );
  MUX U3722 ( .A(reg_target[18]), .B(data_mem_out_wire[882]), .S(n1856), .Z(
        \Data_Mem/n5386 ) );
  MUX U3723 ( .A(reg_target[17]), .B(data_mem_out_wire[881]), .S(n1856), .Z(
        \Data_Mem/n5385 ) );
  MUX U3724 ( .A(reg_target[16]), .B(data_mem_out_wire[880]), .S(n1856), .Z(
        \Data_Mem/n5384 ) );
  MUX U3725 ( .A(reg_target[15]), .B(data_mem_out_wire[879]), .S(n1856), .Z(
        \Data_Mem/n5383 ) );
  MUX U3726 ( .A(reg_target[14]), .B(data_mem_out_wire[878]), .S(n1856), .Z(
        \Data_Mem/n5382 ) );
  MUX U3727 ( .A(reg_target[13]), .B(data_mem_out_wire[877]), .S(n1856), .Z(
        \Data_Mem/n5381 ) );
  MUX U3728 ( .A(reg_target[12]), .B(data_mem_out_wire[876]), .S(n1856), .Z(
        \Data_Mem/n5380 ) );
  MUX U3729 ( .A(reg_target[11]), .B(data_mem_out_wire[875]), .S(n1856), .Z(
        \Data_Mem/n5379 ) );
  MUX U3730 ( .A(reg_target[10]), .B(data_mem_out_wire[874]), .S(n1856), .Z(
        \Data_Mem/n5378 ) );
  MUX U3731 ( .A(reg_target[9]), .B(data_mem_out_wire[873]), .S(n1856), .Z(
        \Data_Mem/n5377 ) );
  MUX U3732 ( .A(reg_target[8]), .B(data_mem_out_wire[872]), .S(n1856), .Z(
        \Data_Mem/n5376 ) );
  MUX U3733 ( .A(reg_target[7]), .B(data_mem_out_wire[871]), .S(n1856), .Z(
        \Data_Mem/n5375 ) );
  MUX U3734 ( .A(reg_target[6]), .B(data_mem_out_wire[870]), .S(n1856), .Z(
        \Data_Mem/n5374 ) );
  MUX U3735 ( .A(reg_target[5]), .B(data_mem_out_wire[869]), .S(n1856), .Z(
        \Data_Mem/n5373 ) );
  MUX U3736 ( .A(reg_target[4]), .B(data_mem_out_wire[868]), .S(n1856), .Z(
        \Data_Mem/n5372 ) );
  MUX U3737 ( .A(reg_target[3]), .B(data_mem_out_wire[867]), .S(n1856), .Z(
        \Data_Mem/n5371 ) );
  MUX U3738 ( .A(reg_target[2]), .B(data_mem_out_wire[866]), .S(n1856), .Z(
        \Data_Mem/n5370 ) );
  IV U3739 ( .A(n1857), .Z(n1856) );
  MUX U3740 ( .A(data_mem_out_wire[865]), .B(reg_target[1]), .S(n1857), .Z(
        \Data_Mem/n5369 ) );
  MUX U3741 ( .A(data_mem_out_wire[864]), .B(reg_target[0]), .S(n1857), .Z(
        \Data_Mem/n5368 ) );
  AND U3742 ( .A(n1801), .B(n1851), .Z(n1857) );
  MUX U3743 ( .A(reg_target[31]), .B(data_mem_out_wire[927]), .S(n1858), .Z(
        \Data_Mem/n5367 ) );
  MUX U3744 ( .A(reg_target[30]), .B(data_mem_out_wire[926]), .S(n1858), .Z(
        \Data_Mem/n5366 ) );
  MUX U3745 ( .A(reg_target[29]), .B(data_mem_out_wire[925]), .S(n1858), .Z(
        \Data_Mem/n5365 ) );
  MUX U3746 ( .A(reg_target[28]), .B(data_mem_out_wire[924]), .S(n1858), .Z(
        \Data_Mem/n5364 ) );
  MUX U3747 ( .A(reg_target[27]), .B(data_mem_out_wire[923]), .S(n1858), .Z(
        \Data_Mem/n5363 ) );
  MUX U3748 ( .A(reg_target[26]), .B(data_mem_out_wire[922]), .S(n1858), .Z(
        \Data_Mem/n5362 ) );
  MUX U3749 ( .A(reg_target[25]), .B(data_mem_out_wire[921]), .S(n1858), .Z(
        \Data_Mem/n5361 ) );
  MUX U3750 ( .A(reg_target[24]), .B(data_mem_out_wire[920]), .S(n1858), .Z(
        \Data_Mem/n5360 ) );
  MUX U3751 ( .A(reg_target[23]), .B(data_mem_out_wire[919]), .S(n1858), .Z(
        \Data_Mem/n5359 ) );
  MUX U3752 ( .A(reg_target[22]), .B(data_mem_out_wire[918]), .S(n1858), .Z(
        \Data_Mem/n5358 ) );
  MUX U3753 ( .A(reg_target[21]), .B(data_mem_out_wire[917]), .S(n1858), .Z(
        \Data_Mem/n5357 ) );
  MUX U3754 ( .A(reg_target[20]), .B(data_mem_out_wire[916]), .S(n1858), .Z(
        \Data_Mem/n5356 ) );
  MUX U3755 ( .A(reg_target[19]), .B(data_mem_out_wire[915]), .S(n1858), .Z(
        \Data_Mem/n5355 ) );
  MUX U3756 ( .A(reg_target[18]), .B(data_mem_out_wire[914]), .S(n1858), .Z(
        \Data_Mem/n5354 ) );
  MUX U3757 ( .A(reg_target[17]), .B(data_mem_out_wire[913]), .S(n1858), .Z(
        \Data_Mem/n5353 ) );
  MUX U3758 ( .A(reg_target[16]), .B(data_mem_out_wire[912]), .S(n1858), .Z(
        \Data_Mem/n5352 ) );
  MUX U3759 ( .A(reg_target[15]), .B(data_mem_out_wire[911]), .S(n1858), .Z(
        \Data_Mem/n5351 ) );
  MUX U3760 ( .A(reg_target[14]), .B(data_mem_out_wire[910]), .S(n1858), .Z(
        \Data_Mem/n5350 ) );
  MUX U3761 ( .A(reg_target[13]), .B(data_mem_out_wire[909]), .S(n1858), .Z(
        \Data_Mem/n5349 ) );
  MUX U3762 ( .A(reg_target[12]), .B(data_mem_out_wire[908]), .S(n1858), .Z(
        \Data_Mem/n5348 ) );
  MUX U3763 ( .A(reg_target[11]), .B(data_mem_out_wire[907]), .S(n1858), .Z(
        \Data_Mem/n5347 ) );
  MUX U3764 ( .A(reg_target[10]), .B(data_mem_out_wire[906]), .S(n1858), .Z(
        \Data_Mem/n5346 ) );
  MUX U3765 ( .A(reg_target[9]), .B(data_mem_out_wire[905]), .S(n1858), .Z(
        \Data_Mem/n5345 ) );
  MUX U3766 ( .A(reg_target[8]), .B(data_mem_out_wire[904]), .S(n1858), .Z(
        \Data_Mem/n5344 ) );
  MUX U3767 ( .A(reg_target[7]), .B(data_mem_out_wire[903]), .S(n1858), .Z(
        \Data_Mem/n5343 ) );
  MUX U3768 ( .A(reg_target[6]), .B(data_mem_out_wire[902]), .S(n1858), .Z(
        \Data_Mem/n5342 ) );
  MUX U3769 ( .A(reg_target[5]), .B(data_mem_out_wire[901]), .S(n1858), .Z(
        \Data_Mem/n5341 ) );
  MUX U3770 ( .A(reg_target[4]), .B(data_mem_out_wire[900]), .S(n1858), .Z(
        \Data_Mem/n5340 ) );
  MUX U3771 ( .A(reg_target[3]), .B(data_mem_out_wire[899]), .S(n1858), .Z(
        \Data_Mem/n5339 ) );
  MUX U3772 ( .A(reg_target[2]), .B(data_mem_out_wire[898]), .S(n1858), .Z(
        \Data_Mem/n5338 ) );
  IV U3773 ( .A(n1859), .Z(n1858) );
  MUX U3774 ( .A(data_mem_out_wire[897]), .B(reg_target[1]), .S(n1859), .Z(
        \Data_Mem/n5337 ) );
  MUX U3775 ( .A(data_mem_out_wire[896]), .B(reg_target[0]), .S(n1859), .Z(
        \Data_Mem/n5336 ) );
  AND U3776 ( .A(n1804), .B(n1851), .Z(n1859) );
  MUX U3777 ( .A(reg_target[31]), .B(data_mem_out_wire[959]), .S(n1860), .Z(
        \Data_Mem/n5335 ) );
  MUX U3778 ( .A(reg_target[30]), .B(data_mem_out_wire[958]), .S(n1860), .Z(
        \Data_Mem/n5334 ) );
  MUX U3779 ( .A(reg_target[29]), .B(data_mem_out_wire[957]), .S(n1860), .Z(
        \Data_Mem/n5333 ) );
  MUX U3780 ( .A(reg_target[28]), .B(data_mem_out_wire[956]), .S(n1860), .Z(
        \Data_Mem/n5332 ) );
  MUX U3781 ( .A(reg_target[27]), .B(data_mem_out_wire[955]), .S(n1860), .Z(
        \Data_Mem/n5331 ) );
  MUX U3782 ( .A(reg_target[26]), .B(data_mem_out_wire[954]), .S(n1860), .Z(
        \Data_Mem/n5330 ) );
  MUX U3783 ( .A(reg_target[25]), .B(data_mem_out_wire[953]), .S(n1860), .Z(
        \Data_Mem/n5329 ) );
  MUX U3784 ( .A(reg_target[24]), .B(data_mem_out_wire[952]), .S(n1860), .Z(
        \Data_Mem/n5328 ) );
  MUX U3785 ( .A(reg_target[23]), .B(data_mem_out_wire[951]), .S(n1860), .Z(
        \Data_Mem/n5327 ) );
  MUX U3786 ( .A(reg_target[22]), .B(data_mem_out_wire[950]), .S(n1860), .Z(
        \Data_Mem/n5326 ) );
  MUX U3787 ( .A(reg_target[21]), .B(data_mem_out_wire[949]), .S(n1860), .Z(
        \Data_Mem/n5325 ) );
  MUX U3788 ( .A(reg_target[20]), .B(data_mem_out_wire[948]), .S(n1860), .Z(
        \Data_Mem/n5324 ) );
  MUX U3789 ( .A(reg_target[19]), .B(data_mem_out_wire[947]), .S(n1860), .Z(
        \Data_Mem/n5323 ) );
  MUX U3790 ( .A(reg_target[18]), .B(data_mem_out_wire[946]), .S(n1860), .Z(
        \Data_Mem/n5322 ) );
  MUX U3791 ( .A(reg_target[17]), .B(data_mem_out_wire[945]), .S(n1860), .Z(
        \Data_Mem/n5321 ) );
  MUX U3792 ( .A(reg_target[16]), .B(data_mem_out_wire[944]), .S(n1860), .Z(
        \Data_Mem/n5320 ) );
  MUX U3793 ( .A(reg_target[15]), .B(data_mem_out_wire[943]), .S(n1860), .Z(
        \Data_Mem/n5319 ) );
  MUX U3794 ( .A(reg_target[14]), .B(data_mem_out_wire[942]), .S(n1860), .Z(
        \Data_Mem/n5318 ) );
  MUX U3795 ( .A(reg_target[13]), .B(data_mem_out_wire[941]), .S(n1860), .Z(
        \Data_Mem/n5317 ) );
  MUX U3796 ( .A(reg_target[12]), .B(data_mem_out_wire[940]), .S(n1860), .Z(
        \Data_Mem/n5316 ) );
  MUX U3797 ( .A(reg_target[11]), .B(data_mem_out_wire[939]), .S(n1860), .Z(
        \Data_Mem/n5315 ) );
  MUX U3798 ( .A(reg_target[10]), .B(data_mem_out_wire[938]), .S(n1860), .Z(
        \Data_Mem/n5314 ) );
  MUX U3799 ( .A(reg_target[9]), .B(data_mem_out_wire[937]), .S(n1860), .Z(
        \Data_Mem/n5313 ) );
  MUX U3800 ( .A(reg_target[8]), .B(data_mem_out_wire[936]), .S(n1860), .Z(
        \Data_Mem/n5312 ) );
  MUX U3801 ( .A(reg_target[7]), .B(data_mem_out_wire[935]), .S(n1860), .Z(
        \Data_Mem/n5311 ) );
  MUX U3802 ( .A(reg_target[6]), .B(data_mem_out_wire[934]), .S(n1860), .Z(
        \Data_Mem/n5310 ) );
  MUX U3803 ( .A(reg_target[5]), .B(data_mem_out_wire[933]), .S(n1860), .Z(
        \Data_Mem/n5309 ) );
  MUX U3804 ( .A(reg_target[4]), .B(data_mem_out_wire[932]), .S(n1860), .Z(
        \Data_Mem/n5308 ) );
  MUX U3805 ( .A(reg_target[3]), .B(data_mem_out_wire[931]), .S(n1860), .Z(
        \Data_Mem/n5307 ) );
  MUX U3806 ( .A(reg_target[2]), .B(data_mem_out_wire[930]), .S(n1860), .Z(
        \Data_Mem/n5306 ) );
  IV U3807 ( .A(n1861), .Z(n1860) );
  MUX U3808 ( .A(data_mem_out_wire[929]), .B(reg_target[1]), .S(n1861), .Z(
        \Data_Mem/n5305 ) );
  MUX U3809 ( .A(data_mem_out_wire[928]), .B(reg_target[0]), .S(n1861), .Z(
        \Data_Mem/n5304 ) );
  AND U3810 ( .A(n1807), .B(n1851), .Z(n1861) );
  MUX U3811 ( .A(reg_target[31]), .B(data_mem_out_wire[991]), .S(n1862), .Z(
        \Data_Mem/n5303 ) );
  MUX U3812 ( .A(reg_target[30]), .B(data_mem_out_wire[990]), .S(n1862), .Z(
        \Data_Mem/n5302 ) );
  MUX U3813 ( .A(reg_target[29]), .B(data_mem_out_wire[989]), .S(n1862), .Z(
        \Data_Mem/n5301 ) );
  MUX U3814 ( .A(reg_target[28]), .B(data_mem_out_wire[988]), .S(n1862), .Z(
        \Data_Mem/n5300 ) );
  MUX U3815 ( .A(reg_target[27]), .B(data_mem_out_wire[987]), .S(n1862), .Z(
        \Data_Mem/n5299 ) );
  MUX U3816 ( .A(reg_target[26]), .B(data_mem_out_wire[986]), .S(n1862), .Z(
        \Data_Mem/n5298 ) );
  MUX U3817 ( .A(reg_target[25]), .B(data_mem_out_wire[985]), .S(n1862), .Z(
        \Data_Mem/n5297 ) );
  MUX U3818 ( .A(reg_target[24]), .B(data_mem_out_wire[984]), .S(n1862), .Z(
        \Data_Mem/n5296 ) );
  MUX U3819 ( .A(reg_target[23]), .B(data_mem_out_wire[983]), .S(n1862), .Z(
        \Data_Mem/n5295 ) );
  MUX U3820 ( .A(reg_target[22]), .B(data_mem_out_wire[982]), .S(n1862), .Z(
        \Data_Mem/n5294 ) );
  MUX U3821 ( .A(reg_target[21]), .B(data_mem_out_wire[981]), .S(n1862), .Z(
        \Data_Mem/n5293 ) );
  MUX U3822 ( .A(reg_target[20]), .B(data_mem_out_wire[980]), .S(n1862), .Z(
        \Data_Mem/n5292 ) );
  MUX U3823 ( .A(reg_target[19]), .B(data_mem_out_wire[979]), .S(n1862), .Z(
        \Data_Mem/n5291 ) );
  MUX U3824 ( .A(reg_target[18]), .B(data_mem_out_wire[978]), .S(n1862), .Z(
        \Data_Mem/n5290 ) );
  MUX U3825 ( .A(reg_target[17]), .B(data_mem_out_wire[977]), .S(n1862), .Z(
        \Data_Mem/n5289 ) );
  MUX U3826 ( .A(reg_target[16]), .B(data_mem_out_wire[976]), .S(n1862), .Z(
        \Data_Mem/n5288 ) );
  MUX U3827 ( .A(reg_target[15]), .B(data_mem_out_wire[975]), .S(n1862), .Z(
        \Data_Mem/n5287 ) );
  MUX U3828 ( .A(reg_target[14]), .B(data_mem_out_wire[974]), .S(n1862), .Z(
        \Data_Mem/n5286 ) );
  MUX U3829 ( .A(reg_target[13]), .B(data_mem_out_wire[973]), .S(n1862), .Z(
        \Data_Mem/n5285 ) );
  MUX U3830 ( .A(reg_target[12]), .B(data_mem_out_wire[972]), .S(n1862), .Z(
        \Data_Mem/n5284 ) );
  MUX U3831 ( .A(reg_target[11]), .B(data_mem_out_wire[971]), .S(n1862), .Z(
        \Data_Mem/n5283 ) );
  MUX U3832 ( .A(reg_target[10]), .B(data_mem_out_wire[970]), .S(n1862), .Z(
        \Data_Mem/n5282 ) );
  MUX U3833 ( .A(reg_target[9]), .B(data_mem_out_wire[969]), .S(n1862), .Z(
        \Data_Mem/n5281 ) );
  MUX U3834 ( .A(reg_target[8]), .B(data_mem_out_wire[968]), .S(n1862), .Z(
        \Data_Mem/n5280 ) );
  MUX U3835 ( .A(reg_target[7]), .B(data_mem_out_wire[967]), .S(n1862), .Z(
        \Data_Mem/n5279 ) );
  MUX U3836 ( .A(reg_target[6]), .B(data_mem_out_wire[966]), .S(n1862), .Z(
        \Data_Mem/n5278 ) );
  MUX U3837 ( .A(reg_target[5]), .B(data_mem_out_wire[965]), .S(n1862), .Z(
        \Data_Mem/n5277 ) );
  MUX U3838 ( .A(reg_target[4]), .B(data_mem_out_wire[964]), .S(n1862), .Z(
        \Data_Mem/n5276 ) );
  MUX U3839 ( .A(reg_target[3]), .B(data_mem_out_wire[963]), .S(n1862), .Z(
        \Data_Mem/n5275 ) );
  MUX U3840 ( .A(reg_target[2]), .B(data_mem_out_wire[962]), .S(n1862), .Z(
        \Data_Mem/n5274 ) );
  IV U3841 ( .A(n1863), .Z(n1862) );
  MUX U3842 ( .A(data_mem_out_wire[961]), .B(reg_target[1]), .S(n1863), .Z(
        \Data_Mem/n5273 ) );
  MUX U3843 ( .A(data_mem_out_wire[960]), .B(reg_target[0]), .S(n1863), .Z(
        \Data_Mem/n5272 ) );
  AND U3844 ( .A(n1810), .B(n1851), .Z(n1863) );
  MUX U3845 ( .A(data_mem_out_wire[1023]), .B(reg_target[31]), .S(n1864), .Z(
        \Data_Mem/n5271 ) );
  MUX U3846 ( .A(data_mem_out_wire[1022]), .B(reg_target[30]), .S(n1864), .Z(
        \Data_Mem/n5270 ) );
  MUX U3847 ( .A(data_mem_out_wire[1021]), .B(reg_target[29]), .S(n1864), .Z(
        \Data_Mem/n5269 ) );
  MUX U3848 ( .A(data_mem_out_wire[1020]), .B(reg_target[28]), .S(n1864), .Z(
        \Data_Mem/n5268 ) );
  MUX U3849 ( .A(data_mem_out_wire[1019]), .B(reg_target[27]), .S(n1864), .Z(
        \Data_Mem/n5267 ) );
  MUX U3850 ( .A(data_mem_out_wire[1018]), .B(reg_target[26]), .S(n1864), .Z(
        \Data_Mem/n5266 ) );
  MUX U3851 ( .A(data_mem_out_wire[1017]), .B(reg_target[25]), .S(n1864), .Z(
        \Data_Mem/n5265 ) );
  MUX U3852 ( .A(data_mem_out_wire[1016]), .B(reg_target[24]), .S(n1864), .Z(
        \Data_Mem/n5264 ) );
  MUX U3853 ( .A(data_mem_out_wire[1015]), .B(reg_target[23]), .S(n1864), .Z(
        \Data_Mem/n5263 ) );
  MUX U3854 ( .A(data_mem_out_wire[1014]), .B(reg_target[22]), .S(n1864), .Z(
        \Data_Mem/n5262 ) );
  MUX U3855 ( .A(data_mem_out_wire[1013]), .B(reg_target[21]), .S(n1864), .Z(
        \Data_Mem/n5261 ) );
  MUX U3856 ( .A(data_mem_out_wire[1012]), .B(reg_target[20]), .S(n1864), .Z(
        \Data_Mem/n5260 ) );
  MUX U3857 ( .A(data_mem_out_wire[1011]), .B(reg_target[19]), .S(n1864), .Z(
        \Data_Mem/n5259 ) );
  MUX U3858 ( .A(data_mem_out_wire[1010]), .B(reg_target[18]), .S(n1864), .Z(
        \Data_Mem/n5258 ) );
  MUX U3859 ( .A(data_mem_out_wire[1009]), .B(reg_target[17]), .S(n1864), .Z(
        \Data_Mem/n5257 ) );
  MUX U3860 ( .A(data_mem_out_wire[1008]), .B(reg_target[16]), .S(n1864), .Z(
        \Data_Mem/n5256 ) );
  MUX U3861 ( .A(data_mem_out_wire[1007]), .B(reg_target[15]), .S(n1864), .Z(
        \Data_Mem/n5255 ) );
  MUX U3862 ( .A(data_mem_out_wire[1006]), .B(reg_target[14]), .S(n1864), .Z(
        \Data_Mem/n5254 ) );
  MUX U3863 ( .A(data_mem_out_wire[1005]), .B(reg_target[13]), .S(n1864), .Z(
        \Data_Mem/n5253 ) );
  MUX U3864 ( .A(data_mem_out_wire[1004]), .B(reg_target[12]), .S(n1864), .Z(
        \Data_Mem/n5252 ) );
  MUX U3865 ( .A(data_mem_out_wire[1003]), .B(reg_target[11]), .S(n1864), .Z(
        \Data_Mem/n5251 ) );
  MUX U3866 ( .A(data_mem_out_wire[1002]), .B(reg_target[10]), .S(n1864), .Z(
        \Data_Mem/n5250 ) );
  MUX U3867 ( .A(data_mem_out_wire[1001]), .B(reg_target[9]), .S(n1864), .Z(
        \Data_Mem/n5249 ) );
  MUX U3868 ( .A(data_mem_out_wire[1000]), .B(reg_target[8]), .S(n1864), .Z(
        \Data_Mem/n5248 ) );
  MUX U3869 ( .A(data_mem_out_wire[999]), .B(reg_target[7]), .S(n1864), .Z(
        \Data_Mem/n5247 ) );
  MUX U3870 ( .A(data_mem_out_wire[998]), .B(reg_target[6]), .S(n1864), .Z(
        \Data_Mem/n5246 ) );
  MUX U3871 ( .A(data_mem_out_wire[997]), .B(reg_target[5]), .S(n1864), .Z(
        \Data_Mem/n5245 ) );
  MUX U3872 ( .A(data_mem_out_wire[996]), .B(reg_target[4]), .S(n1864), .Z(
        \Data_Mem/n5244 ) );
  MUX U3873 ( .A(data_mem_out_wire[995]), .B(reg_target[3]), .S(n1864), .Z(
        \Data_Mem/n5243 ) );
  MUX U3874 ( .A(data_mem_out_wire[994]), .B(reg_target[2]), .S(n1864), .Z(
        \Data_Mem/n5242 ) );
  MUX U3875 ( .A(data_mem_out_wire[993]), .B(reg_target[1]), .S(n1864), .Z(
        \Data_Mem/n5241 ) );
  MUX U3876 ( .A(data_mem_out_wire[992]), .B(reg_target[0]), .S(n1864), .Z(
        \Data_Mem/n5240 ) );
  AND U3877 ( .A(n1851), .B(n1830), .Z(n1864) );
  ANDN U3878 ( .B(n1865), .A(N24), .Z(n1851) );
  MUX U3879 ( .A(reg_target[31]), .B(data_mem_out_wire[1055]), .S(n1866), .Z(
        \Data_Mem/n5239 ) );
  MUX U3880 ( .A(reg_target[30]), .B(data_mem_out_wire[1054]), .S(n1866), .Z(
        \Data_Mem/n5238 ) );
  MUX U3881 ( .A(reg_target[29]), .B(data_mem_out_wire[1053]), .S(n1866), .Z(
        \Data_Mem/n5237 ) );
  MUX U3882 ( .A(reg_target[28]), .B(data_mem_out_wire[1052]), .S(n1866), .Z(
        \Data_Mem/n5236 ) );
  MUX U3883 ( .A(reg_target[27]), .B(data_mem_out_wire[1051]), .S(n1866), .Z(
        \Data_Mem/n5235 ) );
  MUX U3884 ( .A(reg_target[26]), .B(data_mem_out_wire[1050]), .S(n1866), .Z(
        \Data_Mem/n5234 ) );
  MUX U3885 ( .A(reg_target[25]), .B(data_mem_out_wire[1049]), .S(n1866), .Z(
        \Data_Mem/n5233 ) );
  MUX U3886 ( .A(reg_target[24]), .B(data_mem_out_wire[1048]), .S(n1866), .Z(
        \Data_Mem/n5232 ) );
  MUX U3887 ( .A(reg_target[23]), .B(data_mem_out_wire[1047]), .S(n1866), .Z(
        \Data_Mem/n5231 ) );
  MUX U3888 ( .A(reg_target[22]), .B(data_mem_out_wire[1046]), .S(n1866), .Z(
        \Data_Mem/n5230 ) );
  MUX U3889 ( .A(reg_target[21]), .B(data_mem_out_wire[1045]), .S(n1866), .Z(
        \Data_Mem/n5229 ) );
  MUX U3890 ( .A(reg_target[20]), .B(data_mem_out_wire[1044]), .S(n1866), .Z(
        \Data_Mem/n5228 ) );
  MUX U3891 ( .A(reg_target[19]), .B(data_mem_out_wire[1043]), .S(n1866), .Z(
        \Data_Mem/n5227 ) );
  MUX U3892 ( .A(reg_target[18]), .B(data_mem_out_wire[1042]), .S(n1866), .Z(
        \Data_Mem/n5226 ) );
  MUX U3893 ( .A(reg_target[17]), .B(data_mem_out_wire[1041]), .S(n1866), .Z(
        \Data_Mem/n5225 ) );
  MUX U3894 ( .A(reg_target[16]), .B(data_mem_out_wire[1040]), .S(n1866), .Z(
        \Data_Mem/n5224 ) );
  MUX U3895 ( .A(reg_target[15]), .B(data_mem_out_wire[1039]), .S(n1866), .Z(
        \Data_Mem/n5223 ) );
  MUX U3896 ( .A(reg_target[14]), .B(data_mem_out_wire[1038]), .S(n1866), .Z(
        \Data_Mem/n5222 ) );
  MUX U3897 ( .A(reg_target[13]), .B(data_mem_out_wire[1037]), .S(n1866), .Z(
        \Data_Mem/n5221 ) );
  MUX U3898 ( .A(reg_target[12]), .B(data_mem_out_wire[1036]), .S(n1866), .Z(
        \Data_Mem/n5220 ) );
  MUX U3899 ( .A(reg_target[11]), .B(data_mem_out_wire[1035]), .S(n1866), .Z(
        \Data_Mem/n5219 ) );
  MUX U3900 ( .A(reg_target[10]), .B(data_mem_out_wire[1034]), .S(n1866), .Z(
        \Data_Mem/n5218 ) );
  MUX U3901 ( .A(reg_target[9]), .B(data_mem_out_wire[1033]), .S(n1866), .Z(
        \Data_Mem/n5217 ) );
  MUX U3902 ( .A(reg_target[8]), .B(data_mem_out_wire[1032]), .S(n1866), .Z(
        \Data_Mem/n5216 ) );
  MUX U3903 ( .A(reg_target[7]), .B(data_mem_out_wire[1031]), .S(n1866), .Z(
        \Data_Mem/n5215 ) );
  MUX U3904 ( .A(reg_target[6]), .B(data_mem_out_wire[1030]), .S(n1866), .Z(
        \Data_Mem/n5214 ) );
  MUX U3905 ( .A(reg_target[5]), .B(data_mem_out_wire[1029]), .S(n1866), .Z(
        \Data_Mem/n5213 ) );
  MUX U3906 ( .A(reg_target[4]), .B(data_mem_out_wire[1028]), .S(n1866), .Z(
        \Data_Mem/n5212 ) );
  MUX U3907 ( .A(reg_target[3]), .B(data_mem_out_wire[1027]), .S(n1866), .Z(
        \Data_Mem/n5211 ) );
  MUX U3908 ( .A(reg_target[2]), .B(data_mem_out_wire[1026]), .S(n1866), .Z(
        \Data_Mem/n5210 ) );
  IV U3909 ( .A(n1867), .Z(n1866) );
  MUX U3910 ( .A(data_mem_out_wire[1025]), .B(reg_target[1]), .S(n1867), .Z(
        \Data_Mem/n5209 ) );
  MUX U3911 ( .A(data_mem_out_wire[1024]), .B(reg_target[0]), .S(n1867), .Z(
        \Data_Mem/n5208 ) );
  AND U3912 ( .A(n1791), .B(n1868), .Z(n1867) );
  MUX U3913 ( .A(reg_target[31]), .B(data_mem_out_wire[1087]), .S(n1869), .Z(
        \Data_Mem/n5207 ) );
  MUX U3914 ( .A(reg_target[30]), .B(data_mem_out_wire[1086]), .S(n1869), .Z(
        \Data_Mem/n5206 ) );
  MUX U3915 ( .A(reg_target[29]), .B(data_mem_out_wire[1085]), .S(n1869), .Z(
        \Data_Mem/n5205 ) );
  MUX U3916 ( .A(reg_target[28]), .B(data_mem_out_wire[1084]), .S(n1869), .Z(
        \Data_Mem/n5204 ) );
  MUX U3917 ( .A(reg_target[27]), .B(data_mem_out_wire[1083]), .S(n1869), .Z(
        \Data_Mem/n5203 ) );
  MUX U3918 ( .A(reg_target[26]), .B(data_mem_out_wire[1082]), .S(n1869), .Z(
        \Data_Mem/n5202 ) );
  MUX U3919 ( .A(reg_target[25]), .B(data_mem_out_wire[1081]), .S(n1869), .Z(
        \Data_Mem/n5201 ) );
  MUX U3920 ( .A(reg_target[24]), .B(data_mem_out_wire[1080]), .S(n1869), .Z(
        \Data_Mem/n5200 ) );
  MUX U3921 ( .A(reg_target[23]), .B(data_mem_out_wire[1079]), .S(n1869), .Z(
        \Data_Mem/n5199 ) );
  MUX U3922 ( .A(reg_target[22]), .B(data_mem_out_wire[1078]), .S(n1869), .Z(
        \Data_Mem/n5198 ) );
  MUX U3923 ( .A(reg_target[21]), .B(data_mem_out_wire[1077]), .S(n1869), .Z(
        \Data_Mem/n5197 ) );
  MUX U3924 ( .A(reg_target[20]), .B(data_mem_out_wire[1076]), .S(n1869), .Z(
        \Data_Mem/n5196 ) );
  MUX U3925 ( .A(reg_target[19]), .B(data_mem_out_wire[1075]), .S(n1869), .Z(
        \Data_Mem/n5195 ) );
  MUX U3926 ( .A(reg_target[18]), .B(data_mem_out_wire[1074]), .S(n1869), .Z(
        \Data_Mem/n5194 ) );
  MUX U3927 ( .A(reg_target[17]), .B(data_mem_out_wire[1073]), .S(n1869), .Z(
        \Data_Mem/n5193 ) );
  MUX U3928 ( .A(reg_target[16]), .B(data_mem_out_wire[1072]), .S(n1869), .Z(
        \Data_Mem/n5192 ) );
  MUX U3929 ( .A(reg_target[15]), .B(data_mem_out_wire[1071]), .S(n1869), .Z(
        \Data_Mem/n5191 ) );
  MUX U3930 ( .A(reg_target[14]), .B(data_mem_out_wire[1070]), .S(n1869), .Z(
        \Data_Mem/n5190 ) );
  MUX U3931 ( .A(reg_target[13]), .B(data_mem_out_wire[1069]), .S(n1869), .Z(
        \Data_Mem/n5189 ) );
  MUX U3932 ( .A(reg_target[12]), .B(data_mem_out_wire[1068]), .S(n1869), .Z(
        \Data_Mem/n5188 ) );
  MUX U3933 ( .A(reg_target[11]), .B(data_mem_out_wire[1067]), .S(n1869), .Z(
        \Data_Mem/n5187 ) );
  MUX U3934 ( .A(reg_target[10]), .B(data_mem_out_wire[1066]), .S(n1869), .Z(
        \Data_Mem/n5186 ) );
  MUX U3935 ( .A(reg_target[9]), .B(data_mem_out_wire[1065]), .S(n1869), .Z(
        \Data_Mem/n5185 ) );
  MUX U3936 ( .A(reg_target[8]), .B(data_mem_out_wire[1064]), .S(n1869), .Z(
        \Data_Mem/n5184 ) );
  MUX U3937 ( .A(reg_target[7]), .B(data_mem_out_wire[1063]), .S(n1869), .Z(
        \Data_Mem/n5183 ) );
  MUX U3938 ( .A(reg_target[6]), .B(data_mem_out_wire[1062]), .S(n1869), .Z(
        \Data_Mem/n5182 ) );
  MUX U3939 ( .A(reg_target[5]), .B(data_mem_out_wire[1061]), .S(n1869), .Z(
        \Data_Mem/n5181 ) );
  MUX U3940 ( .A(reg_target[4]), .B(data_mem_out_wire[1060]), .S(n1869), .Z(
        \Data_Mem/n5180 ) );
  MUX U3941 ( .A(reg_target[3]), .B(data_mem_out_wire[1059]), .S(n1869), .Z(
        \Data_Mem/n5179 ) );
  MUX U3942 ( .A(reg_target[2]), .B(data_mem_out_wire[1058]), .S(n1869), .Z(
        \Data_Mem/n5178 ) );
  IV U3943 ( .A(n1870), .Z(n1869) );
  MUX U3944 ( .A(data_mem_out_wire[1057]), .B(reg_target[1]), .S(n1870), .Z(
        \Data_Mem/n5177 ) );
  MUX U3945 ( .A(data_mem_out_wire[1056]), .B(reg_target[0]), .S(n1870), .Z(
        \Data_Mem/n5176 ) );
  AND U3946 ( .A(n1795), .B(n1868), .Z(n1870) );
  MUX U3947 ( .A(reg_target[31]), .B(data_mem_out_wire[1119]), .S(n1871), .Z(
        \Data_Mem/n5175 ) );
  MUX U3948 ( .A(reg_target[30]), .B(data_mem_out_wire[1118]), .S(n1871), .Z(
        \Data_Mem/n5174 ) );
  MUX U3949 ( .A(reg_target[29]), .B(data_mem_out_wire[1117]), .S(n1871), .Z(
        \Data_Mem/n5173 ) );
  MUX U3950 ( .A(reg_target[28]), .B(data_mem_out_wire[1116]), .S(n1871), .Z(
        \Data_Mem/n5172 ) );
  MUX U3951 ( .A(reg_target[27]), .B(data_mem_out_wire[1115]), .S(n1871), .Z(
        \Data_Mem/n5171 ) );
  MUX U3952 ( .A(reg_target[26]), .B(data_mem_out_wire[1114]), .S(n1871), .Z(
        \Data_Mem/n5170 ) );
  MUX U3953 ( .A(reg_target[25]), .B(data_mem_out_wire[1113]), .S(n1871), .Z(
        \Data_Mem/n5169 ) );
  MUX U3954 ( .A(reg_target[24]), .B(data_mem_out_wire[1112]), .S(n1871), .Z(
        \Data_Mem/n5168 ) );
  MUX U3955 ( .A(reg_target[23]), .B(data_mem_out_wire[1111]), .S(n1871), .Z(
        \Data_Mem/n5167 ) );
  MUX U3956 ( .A(reg_target[22]), .B(data_mem_out_wire[1110]), .S(n1871), .Z(
        \Data_Mem/n5166 ) );
  MUX U3957 ( .A(reg_target[21]), .B(data_mem_out_wire[1109]), .S(n1871), .Z(
        \Data_Mem/n5165 ) );
  MUX U3958 ( .A(reg_target[20]), .B(data_mem_out_wire[1108]), .S(n1871), .Z(
        \Data_Mem/n5164 ) );
  MUX U3959 ( .A(reg_target[19]), .B(data_mem_out_wire[1107]), .S(n1871), .Z(
        \Data_Mem/n5163 ) );
  MUX U3960 ( .A(reg_target[18]), .B(data_mem_out_wire[1106]), .S(n1871), .Z(
        \Data_Mem/n5162 ) );
  MUX U3961 ( .A(reg_target[17]), .B(data_mem_out_wire[1105]), .S(n1871), .Z(
        \Data_Mem/n5161 ) );
  MUX U3962 ( .A(reg_target[16]), .B(data_mem_out_wire[1104]), .S(n1871), .Z(
        \Data_Mem/n5160 ) );
  MUX U3963 ( .A(reg_target[15]), .B(data_mem_out_wire[1103]), .S(n1871), .Z(
        \Data_Mem/n5159 ) );
  MUX U3964 ( .A(reg_target[14]), .B(data_mem_out_wire[1102]), .S(n1871), .Z(
        \Data_Mem/n5158 ) );
  MUX U3965 ( .A(reg_target[13]), .B(data_mem_out_wire[1101]), .S(n1871), .Z(
        \Data_Mem/n5157 ) );
  MUX U3966 ( .A(reg_target[12]), .B(data_mem_out_wire[1100]), .S(n1871), .Z(
        \Data_Mem/n5156 ) );
  MUX U3967 ( .A(reg_target[11]), .B(data_mem_out_wire[1099]), .S(n1871), .Z(
        \Data_Mem/n5155 ) );
  MUX U3968 ( .A(reg_target[10]), .B(data_mem_out_wire[1098]), .S(n1871), .Z(
        \Data_Mem/n5154 ) );
  MUX U3969 ( .A(reg_target[9]), .B(data_mem_out_wire[1097]), .S(n1871), .Z(
        \Data_Mem/n5153 ) );
  MUX U3970 ( .A(reg_target[8]), .B(data_mem_out_wire[1096]), .S(n1871), .Z(
        \Data_Mem/n5152 ) );
  MUX U3971 ( .A(reg_target[7]), .B(data_mem_out_wire[1095]), .S(n1871), .Z(
        \Data_Mem/n5151 ) );
  MUX U3972 ( .A(reg_target[6]), .B(data_mem_out_wire[1094]), .S(n1871), .Z(
        \Data_Mem/n5150 ) );
  MUX U3973 ( .A(reg_target[5]), .B(data_mem_out_wire[1093]), .S(n1871), .Z(
        \Data_Mem/n5149 ) );
  MUX U3974 ( .A(reg_target[4]), .B(data_mem_out_wire[1092]), .S(n1871), .Z(
        \Data_Mem/n5148 ) );
  MUX U3975 ( .A(reg_target[3]), .B(data_mem_out_wire[1091]), .S(n1871), .Z(
        \Data_Mem/n5147 ) );
  MUX U3976 ( .A(reg_target[2]), .B(data_mem_out_wire[1090]), .S(n1871), .Z(
        \Data_Mem/n5146 ) );
  IV U3977 ( .A(n1872), .Z(n1871) );
  MUX U3978 ( .A(data_mem_out_wire[1089]), .B(reg_target[1]), .S(n1872), .Z(
        \Data_Mem/n5145 ) );
  MUX U3979 ( .A(data_mem_out_wire[1088]), .B(reg_target[0]), .S(n1872), .Z(
        \Data_Mem/n5144 ) );
  AND U3980 ( .A(n1798), .B(n1868), .Z(n1872) );
  MUX U3981 ( .A(reg_target[31]), .B(data_mem_out_wire[1151]), .S(n1873), .Z(
        \Data_Mem/n5143 ) );
  MUX U3982 ( .A(reg_target[30]), .B(data_mem_out_wire[1150]), .S(n1873), .Z(
        \Data_Mem/n5142 ) );
  MUX U3983 ( .A(reg_target[29]), .B(data_mem_out_wire[1149]), .S(n1873), .Z(
        \Data_Mem/n5141 ) );
  MUX U3984 ( .A(reg_target[28]), .B(data_mem_out_wire[1148]), .S(n1873), .Z(
        \Data_Mem/n5140 ) );
  MUX U3985 ( .A(reg_target[27]), .B(data_mem_out_wire[1147]), .S(n1873), .Z(
        \Data_Mem/n5139 ) );
  MUX U3986 ( .A(reg_target[26]), .B(data_mem_out_wire[1146]), .S(n1873), .Z(
        \Data_Mem/n5138 ) );
  MUX U3987 ( .A(reg_target[25]), .B(data_mem_out_wire[1145]), .S(n1873), .Z(
        \Data_Mem/n5137 ) );
  MUX U3988 ( .A(reg_target[24]), .B(data_mem_out_wire[1144]), .S(n1873), .Z(
        \Data_Mem/n5136 ) );
  MUX U3989 ( .A(reg_target[23]), .B(data_mem_out_wire[1143]), .S(n1873), .Z(
        \Data_Mem/n5135 ) );
  MUX U3990 ( .A(reg_target[22]), .B(data_mem_out_wire[1142]), .S(n1873), .Z(
        \Data_Mem/n5134 ) );
  MUX U3991 ( .A(reg_target[21]), .B(data_mem_out_wire[1141]), .S(n1873), .Z(
        \Data_Mem/n5133 ) );
  MUX U3992 ( .A(reg_target[20]), .B(data_mem_out_wire[1140]), .S(n1873), .Z(
        \Data_Mem/n5132 ) );
  MUX U3993 ( .A(reg_target[19]), .B(data_mem_out_wire[1139]), .S(n1873), .Z(
        \Data_Mem/n5131 ) );
  MUX U3994 ( .A(reg_target[18]), .B(data_mem_out_wire[1138]), .S(n1873), .Z(
        \Data_Mem/n5130 ) );
  MUX U3995 ( .A(reg_target[17]), .B(data_mem_out_wire[1137]), .S(n1873), .Z(
        \Data_Mem/n5129 ) );
  MUX U3996 ( .A(reg_target[16]), .B(data_mem_out_wire[1136]), .S(n1873), .Z(
        \Data_Mem/n5128 ) );
  MUX U3997 ( .A(reg_target[15]), .B(data_mem_out_wire[1135]), .S(n1873), .Z(
        \Data_Mem/n5127 ) );
  MUX U3998 ( .A(reg_target[14]), .B(data_mem_out_wire[1134]), .S(n1873), .Z(
        \Data_Mem/n5126 ) );
  MUX U3999 ( .A(reg_target[13]), .B(data_mem_out_wire[1133]), .S(n1873), .Z(
        \Data_Mem/n5125 ) );
  MUX U4000 ( .A(reg_target[12]), .B(data_mem_out_wire[1132]), .S(n1873), .Z(
        \Data_Mem/n5124 ) );
  MUX U4001 ( .A(reg_target[11]), .B(data_mem_out_wire[1131]), .S(n1873), .Z(
        \Data_Mem/n5123 ) );
  MUX U4002 ( .A(reg_target[10]), .B(data_mem_out_wire[1130]), .S(n1873), .Z(
        \Data_Mem/n5122 ) );
  MUX U4003 ( .A(reg_target[9]), .B(data_mem_out_wire[1129]), .S(n1873), .Z(
        \Data_Mem/n5121 ) );
  MUX U4004 ( .A(reg_target[8]), .B(data_mem_out_wire[1128]), .S(n1873), .Z(
        \Data_Mem/n5120 ) );
  MUX U4005 ( .A(reg_target[7]), .B(data_mem_out_wire[1127]), .S(n1873), .Z(
        \Data_Mem/n5119 ) );
  MUX U4006 ( .A(reg_target[6]), .B(data_mem_out_wire[1126]), .S(n1873), .Z(
        \Data_Mem/n5118 ) );
  MUX U4007 ( .A(reg_target[5]), .B(data_mem_out_wire[1125]), .S(n1873), .Z(
        \Data_Mem/n5117 ) );
  MUX U4008 ( .A(reg_target[4]), .B(data_mem_out_wire[1124]), .S(n1873), .Z(
        \Data_Mem/n5116 ) );
  MUX U4009 ( .A(reg_target[3]), .B(data_mem_out_wire[1123]), .S(n1873), .Z(
        \Data_Mem/n5115 ) );
  MUX U4010 ( .A(reg_target[2]), .B(data_mem_out_wire[1122]), .S(n1873), .Z(
        \Data_Mem/n5114 ) );
  IV U4011 ( .A(n1874), .Z(n1873) );
  MUX U4012 ( .A(data_mem_out_wire[1121]), .B(reg_target[1]), .S(n1874), .Z(
        \Data_Mem/n5113 ) );
  MUX U4013 ( .A(data_mem_out_wire[1120]), .B(reg_target[0]), .S(n1874), .Z(
        \Data_Mem/n5112 ) );
  AND U4014 ( .A(n1801), .B(n1868), .Z(n1874) );
  MUX U4015 ( .A(reg_target[31]), .B(data_mem_out_wire[1183]), .S(n1875), .Z(
        \Data_Mem/n5111 ) );
  MUX U4016 ( .A(reg_target[30]), .B(data_mem_out_wire[1182]), .S(n1875), .Z(
        \Data_Mem/n5110 ) );
  MUX U4017 ( .A(reg_target[29]), .B(data_mem_out_wire[1181]), .S(n1875), .Z(
        \Data_Mem/n5109 ) );
  MUX U4018 ( .A(reg_target[28]), .B(data_mem_out_wire[1180]), .S(n1875), .Z(
        \Data_Mem/n5108 ) );
  MUX U4019 ( .A(reg_target[27]), .B(data_mem_out_wire[1179]), .S(n1875), .Z(
        \Data_Mem/n5107 ) );
  MUX U4020 ( .A(reg_target[26]), .B(data_mem_out_wire[1178]), .S(n1875), .Z(
        \Data_Mem/n5106 ) );
  MUX U4021 ( .A(reg_target[25]), .B(data_mem_out_wire[1177]), .S(n1875), .Z(
        \Data_Mem/n5105 ) );
  MUX U4022 ( .A(reg_target[24]), .B(data_mem_out_wire[1176]), .S(n1875), .Z(
        \Data_Mem/n5104 ) );
  MUX U4023 ( .A(reg_target[23]), .B(data_mem_out_wire[1175]), .S(n1875), .Z(
        \Data_Mem/n5103 ) );
  MUX U4024 ( .A(reg_target[22]), .B(data_mem_out_wire[1174]), .S(n1875), .Z(
        \Data_Mem/n5102 ) );
  MUX U4025 ( .A(reg_target[21]), .B(data_mem_out_wire[1173]), .S(n1875), .Z(
        \Data_Mem/n5101 ) );
  MUX U4026 ( .A(reg_target[20]), .B(data_mem_out_wire[1172]), .S(n1875), .Z(
        \Data_Mem/n5100 ) );
  MUX U4027 ( .A(reg_target[19]), .B(data_mem_out_wire[1171]), .S(n1875), .Z(
        \Data_Mem/n5099 ) );
  MUX U4028 ( .A(reg_target[18]), .B(data_mem_out_wire[1170]), .S(n1875), .Z(
        \Data_Mem/n5098 ) );
  MUX U4029 ( .A(reg_target[17]), .B(data_mem_out_wire[1169]), .S(n1875), .Z(
        \Data_Mem/n5097 ) );
  MUX U4030 ( .A(reg_target[16]), .B(data_mem_out_wire[1168]), .S(n1875), .Z(
        \Data_Mem/n5096 ) );
  MUX U4031 ( .A(reg_target[15]), .B(data_mem_out_wire[1167]), .S(n1875), .Z(
        \Data_Mem/n5095 ) );
  MUX U4032 ( .A(reg_target[14]), .B(data_mem_out_wire[1166]), .S(n1875), .Z(
        \Data_Mem/n5094 ) );
  MUX U4033 ( .A(reg_target[13]), .B(data_mem_out_wire[1165]), .S(n1875), .Z(
        \Data_Mem/n5093 ) );
  MUX U4034 ( .A(reg_target[12]), .B(data_mem_out_wire[1164]), .S(n1875), .Z(
        \Data_Mem/n5092 ) );
  MUX U4035 ( .A(reg_target[11]), .B(data_mem_out_wire[1163]), .S(n1875), .Z(
        \Data_Mem/n5091 ) );
  MUX U4036 ( .A(reg_target[10]), .B(data_mem_out_wire[1162]), .S(n1875), .Z(
        \Data_Mem/n5090 ) );
  MUX U4037 ( .A(reg_target[9]), .B(data_mem_out_wire[1161]), .S(n1875), .Z(
        \Data_Mem/n5089 ) );
  MUX U4038 ( .A(reg_target[8]), .B(data_mem_out_wire[1160]), .S(n1875), .Z(
        \Data_Mem/n5088 ) );
  MUX U4039 ( .A(reg_target[7]), .B(data_mem_out_wire[1159]), .S(n1875), .Z(
        \Data_Mem/n5087 ) );
  MUX U4040 ( .A(reg_target[6]), .B(data_mem_out_wire[1158]), .S(n1875), .Z(
        \Data_Mem/n5086 ) );
  MUX U4041 ( .A(reg_target[5]), .B(data_mem_out_wire[1157]), .S(n1875), .Z(
        \Data_Mem/n5085 ) );
  MUX U4042 ( .A(reg_target[4]), .B(data_mem_out_wire[1156]), .S(n1875), .Z(
        \Data_Mem/n5084 ) );
  MUX U4043 ( .A(reg_target[3]), .B(data_mem_out_wire[1155]), .S(n1875), .Z(
        \Data_Mem/n5083 ) );
  MUX U4044 ( .A(reg_target[2]), .B(data_mem_out_wire[1154]), .S(n1875), .Z(
        \Data_Mem/n5082 ) );
  IV U4045 ( .A(n1876), .Z(n1875) );
  MUX U4046 ( .A(data_mem_out_wire[1153]), .B(reg_target[1]), .S(n1876), .Z(
        \Data_Mem/n5081 ) );
  MUX U4047 ( .A(data_mem_out_wire[1152]), .B(reg_target[0]), .S(n1876), .Z(
        \Data_Mem/n5080 ) );
  AND U4048 ( .A(n1804), .B(n1868), .Z(n1876) );
  MUX U4049 ( .A(reg_target[31]), .B(data_mem_out_wire[1215]), .S(n1877), .Z(
        \Data_Mem/n5079 ) );
  MUX U4050 ( .A(reg_target[30]), .B(data_mem_out_wire[1214]), .S(n1877), .Z(
        \Data_Mem/n5078 ) );
  MUX U4051 ( .A(reg_target[29]), .B(data_mem_out_wire[1213]), .S(n1877), .Z(
        \Data_Mem/n5077 ) );
  MUX U4052 ( .A(reg_target[28]), .B(data_mem_out_wire[1212]), .S(n1877), .Z(
        \Data_Mem/n5076 ) );
  MUX U4053 ( .A(reg_target[27]), .B(data_mem_out_wire[1211]), .S(n1877), .Z(
        \Data_Mem/n5075 ) );
  MUX U4054 ( .A(reg_target[26]), .B(data_mem_out_wire[1210]), .S(n1877), .Z(
        \Data_Mem/n5074 ) );
  MUX U4055 ( .A(reg_target[25]), .B(data_mem_out_wire[1209]), .S(n1877), .Z(
        \Data_Mem/n5073 ) );
  MUX U4056 ( .A(reg_target[24]), .B(data_mem_out_wire[1208]), .S(n1877), .Z(
        \Data_Mem/n5072 ) );
  MUX U4057 ( .A(reg_target[23]), .B(data_mem_out_wire[1207]), .S(n1877), .Z(
        \Data_Mem/n5071 ) );
  MUX U4058 ( .A(reg_target[22]), .B(data_mem_out_wire[1206]), .S(n1877), .Z(
        \Data_Mem/n5070 ) );
  MUX U4059 ( .A(reg_target[21]), .B(data_mem_out_wire[1205]), .S(n1877), .Z(
        \Data_Mem/n5069 ) );
  MUX U4060 ( .A(reg_target[20]), .B(data_mem_out_wire[1204]), .S(n1877), .Z(
        \Data_Mem/n5068 ) );
  MUX U4061 ( .A(reg_target[19]), .B(data_mem_out_wire[1203]), .S(n1877), .Z(
        \Data_Mem/n5067 ) );
  MUX U4062 ( .A(reg_target[18]), .B(data_mem_out_wire[1202]), .S(n1877), .Z(
        \Data_Mem/n5066 ) );
  MUX U4063 ( .A(reg_target[17]), .B(data_mem_out_wire[1201]), .S(n1877), .Z(
        \Data_Mem/n5065 ) );
  MUX U4064 ( .A(reg_target[16]), .B(data_mem_out_wire[1200]), .S(n1877), .Z(
        \Data_Mem/n5064 ) );
  MUX U4065 ( .A(reg_target[15]), .B(data_mem_out_wire[1199]), .S(n1877), .Z(
        \Data_Mem/n5063 ) );
  MUX U4066 ( .A(reg_target[14]), .B(data_mem_out_wire[1198]), .S(n1877), .Z(
        \Data_Mem/n5062 ) );
  MUX U4067 ( .A(reg_target[13]), .B(data_mem_out_wire[1197]), .S(n1877), .Z(
        \Data_Mem/n5061 ) );
  MUX U4068 ( .A(reg_target[12]), .B(data_mem_out_wire[1196]), .S(n1877), .Z(
        \Data_Mem/n5060 ) );
  MUX U4069 ( .A(reg_target[11]), .B(data_mem_out_wire[1195]), .S(n1877), .Z(
        \Data_Mem/n5059 ) );
  MUX U4070 ( .A(reg_target[10]), .B(data_mem_out_wire[1194]), .S(n1877), .Z(
        \Data_Mem/n5058 ) );
  MUX U4071 ( .A(reg_target[9]), .B(data_mem_out_wire[1193]), .S(n1877), .Z(
        \Data_Mem/n5057 ) );
  MUX U4072 ( .A(reg_target[8]), .B(data_mem_out_wire[1192]), .S(n1877), .Z(
        \Data_Mem/n5056 ) );
  MUX U4073 ( .A(reg_target[7]), .B(data_mem_out_wire[1191]), .S(n1877), .Z(
        \Data_Mem/n5055 ) );
  MUX U4074 ( .A(reg_target[6]), .B(data_mem_out_wire[1190]), .S(n1877), .Z(
        \Data_Mem/n5054 ) );
  MUX U4075 ( .A(reg_target[5]), .B(data_mem_out_wire[1189]), .S(n1877), .Z(
        \Data_Mem/n5053 ) );
  MUX U4076 ( .A(reg_target[4]), .B(data_mem_out_wire[1188]), .S(n1877), .Z(
        \Data_Mem/n5052 ) );
  MUX U4077 ( .A(reg_target[3]), .B(data_mem_out_wire[1187]), .S(n1877), .Z(
        \Data_Mem/n5051 ) );
  MUX U4078 ( .A(reg_target[2]), .B(data_mem_out_wire[1186]), .S(n1877), .Z(
        \Data_Mem/n5050 ) );
  IV U4079 ( .A(n1878), .Z(n1877) );
  MUX U4080 ( .A(data_mem_out_wire[1185]), .B(reg_target[1]), .S(n1878), .Z(
        \Data_Mem/n5049 ) );
  MUX U4081 ( .A(data_mem_out_wire[1184]), .B(reg_target[0]), .S(n1878), .Z(
        \Data_Mem/n5048 ) );
  AND U4082 ( .A(n1807), .B(n1868), .Z(n1878) );
  MUX U4083 ( .A(reg_target[31]), .B(data_mem_out_wire[1247]), .S(n1879), .Z(
        \Data_Mem/n5047 ) );
  MUX U4084 ( .A(reg_target[30]), .B(data_mem_out_wire[1246]), .S(n1879), .Z(
        \Data_Mem/n5046 ) );
  MUX U4085 ( .A(reg_target[29]), .B(data_mem_out_wire[1245]), .S(n1879), .Z(
        \Data_Mem/n5045 ) );
  MUX U4086 ( .A(reg_target[28]), .B(data_mem_out_wire[1244]), .S(n1879), .Z(
        \Data_Mem/n5044 ) );
  MUX U4087 ( .A(reg_target[27]), .B(data_mem_out_wire[1243]), .S(n1879), .Z(
        \Data_Mem/n5043 ) );
  MUX U4088 ( .A(reg_target[26]), .B(data_mem_out_wire[1242]), .S(n1879), .Z(
        \Data_Mem/n5042 ) );
  MUX U4089 ( .A(reg_target[25]), .B(data_mem_out_wire[1241]), .S(n1879), .Z(
        \Data_Mem/n5041 ) );
  MUX U4090 ( .A(reg_target[24]), .B(data_mem_out_wire[1240]), .S(n1879), .Z(
        \Data_Mem/n5040 ) );
  MUX U4091 ( .A(reg_target[23]), .B(data_mem_out_wire[1239]), .S(n1879), .Z(
        \Data_Mem/n5039 ) );
  MUX U4092 ( .A(reg_target[22]), .B(data_mem_out_wire[1238]), .S(n1879), .Z(
        \Data_Mem/n5038 ) );
  MUX U4093 ( .A(reg_target[21]), .B(data_mem_out_wire[1237]), .S(n1879), .Z(
        \Data_Mem/n5037 ) );
  MUX U4094 ( .A(reg_target[20]), .B(data_mem_out_wire[1236]), .S(n1879), .Z(
        \Data_Mem/n5036 ) );
  MUX U4095 ( .A(reg_target[19]), .B(data_mem_out_wire[1235]), .S(n1879), .Z(
        \Data_Mem/n5035 ) );
  MUX U4096 ( .A(reg_target[18]), .B(data_mem_out_wire[1234]), .S(n1879), .Z(
        \Data_Mem/n5034 ) );
  MUX U4097 ( .A(reg_target[17]), .B(data_mem_out_wire[1233]), .S(n1879), .Z(
        \Data_Mem/n5033 ) );
  MUX U4098 ( .A(reg_target[16]), .B(data_mem_out_wire[1232]), .S(n1879), .Z(
        \Data_Mem/n5032 ) );
  MUX U4099 ( .A(reg_target[15]), .B(data_mem_out_wire[1231]), .S(n1879), .Z(
        \Data_Mem/n5031 ) );
  MUX U4100 ( .A(reg_target[14]), .B(data_mem_out_wire[1230]), .S(n1879), .Z(
        \Data_Mem/n5030 ) );
  MUX U4101 ( .A(reg_target[13]), .B(data_mem_out_wire[1229]), .S(n1879), .Z(
        \Data_Mem/n5029 ) );
  MUX U4102 ( .A(reg_target[12]), .B(data_mem_out_wire[1228]), .S(n1879), .Z(
        \Data_Mem/n5028 ) );
  MUX U4103 ( .A(reg_target[11]), .B(data_mem_out_wire[1227]), .S(n1879), .Z(
        \Data_Mem/n5027 ) );
  MUX U4104 ( .A(reg_target[10]), .B(data_mem_out_wire[1226]), .S(n1879), .Z(
        \Data_Mem/n5026 ) );
  MUX U4105 ( .A(reg_target[9]), .B(data_mem_out_wire[1225]), .S(n1879), .Z(
        \Data_Mem/n5025 ) );
  MUX U4106 ( .A(reg_target[8]), .B(data_mem_out_wire[1224]), .S(n1879), .Z(
        \Data_Mem/n5024 ) );
  MUX U4107 ( .A(reg_target[7]), .B(data_mem_out_wire[1223]), .S(n1879), .Z(
        \Data_Mem/n5023 ) );
  MUX U4108 ( .A(reg_target[6]), .B(data_mem_out_wire[1222]), .S(n1879), .Z(
        \Data_Mem/n5022 ) );
  MUX U4109 ( .A(reg_target[5]), .B(data_mem_out_wire[1221]), .S(n1879), .Z(
        \Data_Mem/n5021 ) );
  MUX U4110 ( .A(reg_target[4]), .B(data_mem_out_wire[1220]), .S(n1879), .Z(
        \Data_Mem/n5020 ) );
  MUX U4111 ( .A(reg_target[3]), .B(data_mem_out_wire[1219]), .S(n1879), .Z(
        \Data_Mem/n5019 ) );
  MUX U4112 ( .A(reg_target[2]), .B(data_mem_out_wire[1218]), .S(n1879), .Z(
        \Data_Mem/n5018 ) );
  IV U4113 ( .A(n1880), .Z(n1879) );
  MUX U4114 ( .A(data_mem_out_wire[1217]), .B(reg_target[1]), .S(n1880), .Z(
        \Data_Mem/n5017 ) );
  MUX U4115 ( .A(data_mem_out_wire[1216]), .B(reg_target[0]), .S(n1880), .Z(
        \Data_Mem/n5016 ) );
  AND U4116 ( .A(n1810), .B(n1868), .Z(n1880) );
  MUX U4117 ( .A(data_mem_out_wire[1279]), .B(reg_target[31]), .S(n1881), .Z(
        \Data_Mem/n5015 ) );
  MUX U4118 ( .A(data_mem_out_wire[1278]), .B(reg_target[30]), .S(n1881), .Z(
        \Data_Mem/n5014 ) );
  MUX U4119 ( .A(data_mem_out_wire[1277]), .B(reg_target[29]), .S(n1881), .Z(
        \Data_Mem/n5013 ) );
  MUX U4120 ( .A(data_mem_out_wire[1276]), .B(reg_target[28]), .S(n1881), .Z(
        \Data_Mem/n5012 ) );
  MUX U4121 ( .A(data_mem_out_wire[1275]), .B(reg_target[27]), .S(n1881), .Z(
        \Data_Mem/n5011 ) );
  MUX U4122 ( .A(data_mem_out_wire[1274]), .B(reg_target[26]), .S(n1881), .Z(
        \Data_Mem/n5010 ) );
  MUX U4123 ( .A(data_mem_out_wire[1273]), .B(reg_target[25]), .S(n1881), .Z(
        \Data_Mem/n5009 ) );
  MUX U4124 ( .A(data_mem_out_wire[1272]), .B(reg_target[24]), .S(n1881), .Z(
        \Data_Mem/n5008 ) );
  MUX U4125 ( .A(data_mem_out_wire[1271]), .B(reg_target[23]), .S(n1881), .Z(
        \Data_Mem/n5007 ) );
  MUX U4126 ( .A(data_mem_out_wire[1270]), .B(reg_target[22]), .S(n1881), .Z(
        \Data_Mem/n5006 ) );
  MUX U4127 ( .A(data_mem_out_wire[1269]), .B(reg_target[21]), .S(n1881), .Z(
        \Data_Mem/n5005 ) );
  MUX U4128 ( .A(data_mem_out_wire[1268]), .B(reg_target[20]), .S(n1881), .Z(
        \Data_Mem/n5004 ) );
  MUX U4129 ( .A(data_mem_out_wire[1267]), .B(reg_target[19]), .S(n1881), .Z(
        \Data_Mem/n5003 ) );
  MUX U4130 ( .A(data_mem_out_wire[1266]), .B(reg_target[18]), .S(n1881), .Z(
        \Data_Mem/n5002 ) );
  MUX U4131 ( .A(data_mem_out_wire[1265]), .B(reg_target[17]), .S(n1881), .Z(
        \Data_Mem/n5001 ) );
  MUX U4132 ( .A(data_mem_out_wire[1264]), .B(reg_target[16]), .S(n1881), .Z(
        \Data_Mem/n5000 ) );
  MUX U4133 ( .A(data_mem_out_wire[1263]), .B(reg_target[15]), .S(n1881), .Z(
        \Data_Mem/n4999 ) );
  MUX U4134 ( .A(data_mem_out_wire[1262]), .B(reg_target[14]), .S(n1881), .Z(
        \Data_Mem/n4998 ) );
  MUX U4135 ( .A(data_mem_out_wire[1261]), .B(reg_target[13]), .S(n1881), .Z(
        \Data_Mem/n4997 ) );
  MUX U4136 ( .A(data_mem_out_wire[1260]), .B(reg_target[12]), .S(n1881), .Z(
        \Data_Mem/n4996 ) );
  MUX U4137 ( .A(data_mem_out_wire[1259]), .B(reg_target[11]), .S(n1881), .Z(
        \Data_Mem/n4995 ) );
  MUX U4138 ( .A(data_mem_out_wire[1258]), .B(reg_target[10]), .S(n1881), .Z(
        \Data_Mem/n4994 ) );
  MUX U4139 ( .A(data_mem_out_wire[1257]), .B(reg_target[9]), .S(n1881), .Z(
        \Data_Mem/n4993 ) );
  MUX U4140 ( .A(data_mem_out_wire[1256]), .B(reg_target[8]), .S(n1881), .Z(
        \Data_Mem/n4992 ) );
  MUX U4141 ( .A(data_mem_out_wire[1255]), .B(reg_target[7]), .S(n1881), .Z(
        \Data_Mem/n4991 ) );
  MUX U4142 ( .A(data_mem_out_wire[1254]), .B(reg_target[6]), .S(n1881), .Z(
        \Data_Mem/n4990 ) );
  MUX U4143 ( .A(data_mem_out_wire[1253]), .B(reg_target[5]), .S(n1881), .Z(
        \Data_Mem/n4989 ) );
  MUX U4144 ( .A(data_mem_out_wire[1252]), .B(reg_target[4]), .S(n1881), .Z(
        \Data_Mem/n4988 ) );
  MUX U4145 ( .A(data_mem_out_wire[1251]), .B(reg_target[3]), .S(n1881), .Z(
        \Data_Mem/n4987 ) );
  MUX U4146 ( .A(data_mem_out_wire[1250]), .B(reg_target[2]), .S(n1881), .Z(
        \Data_Mem/n4986 ) );
  MUX U4147 ( .A(data_mem_out_wire[1249]), .B(reg_target[1]), .S(n1881), .Z(
        \Data_Mem/n4985 ) );
  MUX U4148 ( .A(data_mem_out_wire[1248]), .B(reg_target[0]), .S(n1881), .Z(
        \Data_Mem/n4984 ) );
  AND U4149 ( .A(n1868), .B(n1830), .Z(n1881) );
  AND U4150 ( .A(n1813), .B(N24), .Z(n1868) );
  ANDN U4151 ( .B(n837), .A(N25), .Z(n1813) );
  MUX U4152 ( .A(reg_target[31]), .B(data_mem_out_wire[1311]), .S(n1882), .Z(
        \Data_Mem/n4983 ) );
  MUX U4153 ( .A(reg_target[30]), .B(data_mem_out_wire[1310]), .S(n1882), .Z(
        \Data_Mem/n4982 ) );
  MUX U4154 ( .A(reg_target[29]), .B(data_mem_out_wire[1309]), .S(n1882), .Z(
        \Data_Mem/n4981 ) );
  MUX U4155 ( .A(reg_target[28]), .B(data_mem_out_wire[1308]), .S(n1882), .Z(
        \Data_Mem/n4980 ) );
  MUX U4156 ( .A(reg_target[27]), .B(data_mem_out_wire[1307]), .S(n1882), .Z(
        \Data_Mem/n4979 ) );
  MUX U4157 ( .A(reg_target[26]), .B(data_mem_out_wire[1306]), .S(n1882), .Z(
        \Data_Mem/n4978 ) );
  MUX U4158 ( .A(reg_target[25]), .B(data_mem_out_wire[1305]), .S(n1882), .Z(
        \Data_Mem/n4977 ) );
  MUX U4159 ( .A(reg_target[24]), .B(data_mem_out_wire[1304]), .S(n1882), .Z(
        \Data_Mem/n4976 ) );
  MUX U4160 ( .A(reg_target[23]), .B(data_mem_out_wire[1303]), .S(n1882), .Z(
        \Data_Mem/n4975 ) );
  MUX U4161 ( .A(reg_target[22]), .B(data_mem_out_wire[1302]), .S(n1882), .Z(
        \Data_Mem/n4974 ) );
  MUX U4162 ( .A(reg_target[21]), .B(data_mem_out_wire[1301]), .S(n1882), .Z(
        \Data_Mem/n4973 ) );
  MUX U4163 ( .A(reg_target[20]), .B(data_mem_out_wire[1300]), .S(n1882), .Z(
        \Data_Mem/n4972 ) );
  MUX U4164 ( .A(reg_target[19]), .B(data_mem_out_wire[1299]), .S(n1882), .Z(
        \Data_Mem/n4971 ) );
  MUX U4165 ( .A(reg_target[18]), .B(data_mem_out_wire[1298]), .S(n1882), .Z(
        \Data_Mem/n4970 ) );
  MUX U4166 ( .A(reg_target[17]), .B(data_mem_out_wire[1297]), .S(n1882), .Z(
        \Data_Mem/n4969 ) );
  MUX U4167 ( .A(reg_target[16]), .B(data_mem_out_wire[1296]), .S(n1882), .Z(
        \Data_Mem/n4968 ) );
  MUX U4168 ( .A(reg_target[15]), .B(data_mem_out_wire[1295]), .S(n1882), .Z(
        \Data_Mem/n4967 ) );
  MUX U4169 ( .A(reg_target[14]), .B(data_mem_out_wire[1294]), .S(n1882), .Z(
        \Data_Mem/n4966 ) );
  MUX U4170 ( .A(reg_target[13]), .B(data_mem_out_wire[1293]), .S(n1882), .Z(
        \Data_Mem/n4965 ) );
  MUX U4171 ( .A(reg_target[12]), .B(data_mem_out_wire[1292]), .S(n1882), .Z(
        \Data_Mem/n4964 ) );
  MUX U4172 ( .A(reg_target[11]), .B(data_mem_out_wire[1291]), .S(n1882), .Z(
        \Data_Mem/n4963 ) );
  MUX U4173 ( .A(reg_target[10]), .B(data_mem_out_wire[1290]), .S(n1882), .Z(
        \Data_Mem/n4962 ) );
  MUX U4174 ( .A(reg_target[9]), .B(data_mem_out_wire[1289]), .S(n1882), .Z(
        \Data_Mem/n4961 ) );
  MUX U4175 ( .A(reg_target[8]), .B(data_mem_out_wire[1288]), .S(n1882), .Z(
        \Data_Mem/n4960 ) );
  MUX U4176 ( .A(reg_target[7]), .B(data_mem_out_wire[1287]), .S(n1882), .Z(
        \Data_Mem/n4959 ) );
  MUX U4177 ( .A(reg_target[6]), .B(data_mem_out_wire[1286]), .S(n1882), .Z(
        \Data_Mem/n4958 ) );
  MUX U4178 ( .A(reg_target[5]), .B(data_mem_out_wire[1285]), .S(n1882), .Z(
        \Data_Mem/n4957 ) );
  MUX U4179 ( .A(reg_target[4]), .B(data_mem_out_wire[1284]), .S(n1882), .Z(
        \Data_Mem/n4956 ) );
  MUX U4180 ( .A(reg_target[3]), .B(data_mem_out_wire[1283]), .S(n1882), .Z(
        \Data_Mem/n4955 ) );
  MUX U4181 ( .A(reg_target[2]), .B(data_mem_out_wire[1282]), .S(n1882), .Z(
        \Data_Mem/n4954 ) );
  IV U4182 ( .A(n1883), .Z(n1882) );
  MUX U4183 ( .A(data_mem_out_wire[1281]), .B(reg_target[1]), .S(n1883), .Z(
        \Data_Mem/n4953 ) );
  MUX U4184 ( .A(data_mem_out_wire[1280]), .B(reg_target[0]), .S(n1883), .Z(
        \Data_Mem/n4952 ) );
  AND U4185 ( .A(n1791), .B(n1884), .Z(n1883) );
  MUX U4186 ( .A(reg_target[31]), .B(data_mem_out_wire[1343]), .S(n1885), .Z(
        \Data_Mem/n4951 ) );
  MUX U4187 ( .A(reg_target[30]), .B(data_mem_out_wire[1342]), .S(n1885), .Z(
        \Data_Mem/n4950 ) );
  MUX U4188 ( .A(reg_target[29]), .B(data_mem_out_wire[1341]), .S(n1885), .Z(
        \Data_Mem/n4949 ) );
  MUX U4189 ( .A(reg_target[28]), .B(data_mem_out_wire[1340]), .S(n1885), .Z(
        \Data_Mem/n4948 ) );
  MUX U4190 ( .A(reg_target[27]), .B(data_mem_out_wire[1339]), .S(n1885), .Z(
        \Data_Mem/n4947 ) );
  MUX U4191 ( .A(reg_target[26]), .B(data_mem_out_wire[1338]), .S(n1885), .Z(
        \Data_Mem/n4946 ) );
  MUX U4192 ( .A(reg_target[25]), .B(data_mem_out_wire[1337]), .S(n1885), .Z(
        \Data_Mem/n4945 ) );
  MUX U4193 ( .A(reg_target[24]), .B(data_mem_out_wire[1336]), .S(n1885), .Z(
        \Data_Mem/n4944 ) );
  MUX U4194 ( .A(reg_target[23]), .B(data_mem_out_wire[1335]), .S(n1885), .Z(
        \Data_Mem/n4943 ) );
  MUX U4195 ( .A(reg_target[22]), .B(data_mem_out_wire[1334]), .S(n1885), .Z(
        \Data_Mem/n4942 ) );
  MUX U4196 ( .A(reg_target[21]), .B(data_mem_out_wire[1333]), .S(n1885), .Z(
        \Data_Mem/n4941 ) );
  MUX U4197 ( .A(reg_target[20]), .B(data_mem_out_wire[1332]), .S(n1885), .Z(
        \Data_Mem/n4940 ) );
  MUX U4198 ( .A(reg_target[19]), .B(data_mem_out_wire[1331]), .S(n1885), .Z(
        \Data_Mem/n4939 ) );
  MUX U4199 ( .A(reg_target[18]), .B(data_mem_out_wire[1330]), .S(n1885), .Z(
        \Data_Mem/n4938 ) );
  MUX U4200 ( .A(reg_target[17]), .B(data_mem_out_wire[1329]), .S(n1885), .Z(
        \Data_Mem/n4937 ) );
  MUX U4201 ( .A(reg_target[16]), .B(data_mem_out_wire[1328]), .S(n1885), .Z(
        \Data_Mem/n4936 ) );
  MUX U4202 ( .A(reg_target[15]), .B(data_mem_out_wire[1327]), .S(n1885), .Z(
        \Data_Mem/n4935 ) );
  MUX U4203 ( .A(reg_target[14]), .B(data_mem_out_wire[1326]), .S(n1885), .Z(
        \Data_Mem/n4934 ) );
  MUX U4204 ( .A(reg_target[13]), .B(data_mem_out_wire[1325]), .S(n1885), .Z(
        \Data_Mem/n4933 ) );
  MUX U4205 ( .A(reg_target[12]), .B(data_mem_out_wire[1324]), .S(n1885), .Z(
        \Data_Mem/n4932 ) );
  MUX U4206 ( .A(reg_target[11]), .B(data_mem_out_wire[1323]), .S(n1885), .Z(
        \Data_Mem/n4931 ) );
  MUX U4207 ( .A(reg_target[10]), .B(data_mem_out_wire[1322]), .S(n1885), .Z(
        \Data_Mem/n4930 ) );
  MUX U4208 ( .A(reg_target[9]), .B(data_mem_out_wire[1321]), .S(n1885), .Z(
        \Data_Mem/n4929 ) );
  MUX U4209 ( .A(reg_target[8]), .B(data_mem_out_wire[1320]), .S(n1885), .Z(
        \Data_Mem/n4928 ) );
  MUX U4210 ( .A(reg_target[7]), .B(data_mem_out_wire[1319]), .S(n1885), .Z(
        \Data_Mem/n4927 ) );
  MUX U4211 ( .A(reg_target[6]), .B(data_mem_out_wire[1318]), .S(n1885), .Z(
        \Data_Mem/n4926 ) );
  MUX U4212 ( .A(reg_target[5]), .B(data_mem_out_wire[1317]), .S(n1885), .Z(
        \Data_Mem/n4925 ) );
  MUX U4213 ( .A(reg_target[4]), .B(data_mem_out_wire[1316]), .S(n1885), .Z(
        \Data_Mem/n4924 ) );
  MUX U4214 ( .A(reg_target[3]), .B(data_mem_out_wire[1315]), .S(n1885), .Z(
        \Data_Mem/n4923 ) );
  MUX U4215 ( .A(reg_target[2]), .B(data_mem_out_wire[1314]), .S(n1885), .Z(
        \Data_Mem/n4922 ) );
  IV U4216 ( .A(n1886), .Z(n1885) );
  MUX U4217 ( .A(data_mem_out_wire[1313]), .B(reg_target[1]), .S(n1886), .Z(
        \Data_Mem/n4921 ) );
  MUX U4218 ( .A(data_mem_out_wire[1312]), .B(reg_target[0]), .S(n1886), .Z(
        \Data_Mem/n4920 ) );
  AND U4219 ( .A(n1795), .B(n1884), .Z(n1886) );
  MUX U4220 ( .A(reg_target[31]), .B(data_mem_out_wire[1375]), .S(n1887), .Z(
        \Data_Mem/n4919 ) );
  MUX U4221 ( .A(reg_target[30]), .B(data_mem_out_wire[1374]), .S(n1887), .Z(
        \Data_Mem/n4918 ) );
  MUX U4222 ( .A(reg_target[29]), .B(data_mem_out_wire[1373]), .S(n1887), .Z(
        \Data_Mem/n4917 ) );
  MUX U4223 ( .A(reg_target[28]), .B(data_mem_out_wire[1372]), .S(n1887), .Z(
        \Data_Mem/n4916 ) );
  MUX U4224 ( .A(reg_target[27]), .B(data_mem_out_wire[1371]), .S(n1887), .Z(
        \Data_Mem/n4915 ) );
  MUX U4225 ( .A(reg_target[26]), .B(data_mem_out_wire[1370]), .S(n1887), .Z(
        \Data_Mem/n4914 ) );
  MUX U4226 ( .A(reg_target[25]), .B(data_mem_out_wire[1369]), .S(n1887), .Z(
        \Data_Mem/n4913 ) );
  MUX U4227 ( .A(reg_target[24]), .B(data_mem_out_wire[1368]), .S(n1887), .Z(
        \Data_Mem/n4912 ) );
  MUX U4228 ( .A(reg_target[23]), .B(data_mem_out_wire[1367]), .S(n1887), .Z(
        \Data_Mem/n4911 ) );
  MUX U4229 ( .A(reg_target[22]), .B(data_mem_out_wire[1366]), .S(n1887), .Z(
        \Data_Mem/n4910 ) );
  MUX U4230 ( .A(reg_target[21]), .B(data_mem_out_wire[1365]), .S(n1887), .Z(
        \Data_Mem/n4909 ) );
  MUX U4231 ( .A(reg_target[20]), .B(data_mem_out_wire[1364]), .S(n1887), .Z(
        \Data_Mem/n4908 ) );
  MUX U4232 ( .A(reg_target[19]), .B(data_mem_out_wire[1363]), .S(n1887), .Z(
        \Data_Mem/n4907 ) );
  MUX U4233 ( .A(reg_target[18]), .B(data_mem_out_wire[1362]), .S(n1887), .Z(
        \Data_Mem/n4906 ) );
  MUX U4234 ( .A(reg_target[17]), .B(data_mem_out_wire[1361]), .S(n1887), .Z(
        \Data_Mem/n4905 ) );
  MUX U4235 ( .A(reg_target[16]), .B(data_mem_out_wire[1360]), .S(n1887), .Z(
        \Data_Mem/n4904 ) );
  MUX U4236 ( .A(reg_target[15]), .B(data_mem_out_wire[1359]), .S(n1887), .Z(
        \Data_Mem/n4903 ) );
  MUX U4237 ( .A(reg_target[14]), .B(data_mem_out_wire[1358]), .S(n1887), .Z(
        \Data_Mem/n4902 ) );
  MUX U4238 ( .A(reg_target[13]), .B(data_mem_out_wire[1357]), .S(n1887), .Z(
        \Data_Mem/n4901 ) );
  MUX U4239 ( .A(reg_target[12]), .B(data_mem_out_wire[1356]), .S(n1887), .Z(
        \Data_Mem/n4900 ) );
  MUX U4240 ( .A(reg_target[11]), .B(data_mem_out_wire[1355]), .S(n1887), .Z(
        \Data_Mem/n4899 ) );
  MUX U4241 ( .A(reg_target[10]), .B(data_mem_out_wire[1354]), .S(n1887), .Z(
        \Data_Mem/n4898 ) );
  MUX U4242 ( .A(reg_target[9]), .B(data_mem_out_wire[1353]), .S(n1887), .Z(
        \Data_Mem/n4897 ) );
  MUX U4243 ( .A(reg_target[8]), .B(data_mem_out_wire[1352]), .S(n1887), .Z(
        \Data_Mem/n4896 ) );
  MUX U4244 ( .A(reg_target[7]), .B(data_mem_out_wire[1351]), .S(n1887), .Z(
        \Data_Mem/n4895 ) );
  MUX U4245 ( .A(reg_target[6]), .B(data_mem_out_wire[1350]), .S(n1887), .Z(
        \Data_Mem/n4894 ) );
  MUX U4246 ( .A(reg_target[5]), .B(data_mem_out_wire[1349]), .S(n1887), .Z(
        \Data_Mem/n4893 ) );
  MUX U4247 ( .A(reg_target[4]), .B(data_mem_out_wire[1348]), .S(n1887), .Z(
        \Data_Mem/n4892 ) );
  MUX U4248 ( .A(reg_target[3]), .B(data_mem_out_wire[1347]), .S(n1887), .Z(
        \Data_Mem/n4891 ) );
  MUX U4249 ( .A(reg_target[2]), .B(data_mem_out_wire[1346]), .S(n1887), .Z(
        \Data_Mem/n4890 ) );
  IV U4250 ( .A(n1888), .Z(n1887) );
  MUX U4251 ( .A(data_mem_out_wire[1345]), .B(reg_target[1]), .S(n1888), .Z(
        \Data_Mem/n4889 ) );
  MUX U4252 ( .A(data_mem_out_wire[1344]), .B(reg_target[0]), .S(n1888), .Z(
        \Data_Mem/n4888 ) );
  AND U4253 ( .A(n1798), .B(n1884), .Z(n1888) );
  MUX U4254 ( .A(reg_target[31]), .B(data_mem_out_wire[1407]), .S(n1889), .Z(
        \Data_Mem/n4887 ) );
  MUX U4255 ( .A(reg_target[30]), .B(data_mem_out_wire[1406]), .S(n1889), .Z(
        \Data_Mem/n4886 ) );
  MUX U4256 ( .A(reg_target[29]), .B(data_mem_out_wire[1405]), .S(n1889), .Z(
        \Data_Mem/n4885 ) );
  MUX U4257 ( .A(reg_target[28]), .B(data_mem_out_wire[1404]), .S(n1889), .Z(
        \Data_Mem/n4884 ) );
  MUX U4258 ( .A(reg_target[27]), .B(data_mem_out_wire[1403]), .S(n1889), .Z(
        \Data_Mem/n4883 ) );
  MUX U4259 ( .A(reg_target[26]), .B(data_mem_out_wire[1402]), .S(n1889), .Z(
        \Data_Mem/n4882 ) );
  MUX U4260 ( .A(reg_target[25]), .B(data_mem_out_wire[1401]), .S(n1889), .Z(
        \Data_Mem/n4881 ) );
  MUX U4261 ( .A(reg_target[24]), .B(data_mem_out_wire[1400]), .S(n1889), .Z(
        \Data_Mem/n4880 ) );
  MUX U4262 ( .A(reg_target[23]), .B(data_mem_out_wire[1399]), .S(n1889), .Z(
        \Data_Mem/n4879 ) );
  MUX U4263 ( .A(reg_target[22]), .B(data_mem_out_wire[1398]), .S(n1889), .Z(
        \Data_Mem/n4878 ) );
  MUX U4264 ( .A(reg_target[21]), .B(data_mem_out_wire[1397]), .S(n1889), .Z(
        \Data_Mem/n4877 ) );
  MUX U4265 ( .A(reg_target[20]), .B(data_mem_out_wire[1396]), .S(n1889), .Z(
        \Data_Mem/n4876 ) );
  MUX U4266 ( .A(reg_target[19]), .B(data_mem_out_wire[1395]), .S(n1889), .Z(
        \Data_Mem/n4875 ) );
  MUX U4267 ( .A(reg_target[18]), .B(data_mem_out_wire[1394]), .S(n1889), .Z(
        \Data_Mem/n4874 ) );
  MUX U4268 ( .A(reg_target[17]), .B(data_mem_out_wire[1393]), .S(n1889), .Z(
        \Data_Mem/n4873 ) );
  MUX U4269 ( .A(reg_target[16]), .B(data_mem_out_wire[1392]), .S(n1889), .Z(
        \Data_Mem/n4872 ) );
  MUX U4270 ( .A(reg_target[15]), .B(data_mem_out_wire[1391]), .S(n1889), .Z(
        \Data_Mem/n4871 ) );
  MUX U4271 ( .A(reg_target[14]), .B(data_mem_out_wire[1390]), .S(n1889), .Z(
        \Data_Mem/n4870 ) );
  MUX U4272 ( .A(reg_target[13]), .B(data_mem_out_wire[1389]), .S(n1889), .Z(
        \Data_Mem/n4869 ) );
  MUX U4273 ( .A(reg_target[12]), .B(data_mem_out_wire[1388]), .S(n1889), .Z(
        \Data_Mem/n4868 ) );
  MUX U4274 ( .A(reg_target[11]), .B(data_mem_out_wire[1387]), .S(n1889), .Z(
        \Data_Mem/n4867 ) );
  MUX U4275 ( .A(reg_target[10]), .B(data_mem_out_wire[1386]), .S(n1889), .Z(
        \Data_Mem/n4866 ) );
  MUX U4276 ( .A(reg_target[9]), .B(data_mem_out_wire[1385]), .S(n1889), .Z(
        \Data_Mem/n4865 ) );
  MUX U4277 ( .A(reg_target[8]), .B(data_mem_out_wire[1384]), .S(n1889), .Z(
        \Data_Mem/n4864 ) );
  MUX U4278 ( .A(reg_target[7]), .B(data_mem_out_wire[1383]), .S(n1889), .Z(
        \Data_Mem/n4863 ) );
  MUX U4279 ( .A(reg_target[6]), .B(data_mem_out_wire[1382]), .S(n1889), .Z(
        \Data_Mem/n4862 ) );
  MUX U4280 ( .A(reg_target[5]), .B(data_mem_out_wire[1381]), .S(n1889), .Z(
        \Data_Mem/n4861 ) );
  MUX U4281 ( .A(reg_target[4]), .B(data_mem_out_wire[1380]), .S(n1889), .Z(
        \Data_Mem/n4860 ) );
  MUX U4282 ( .A(reg_target[3]), .B(data_mem_out_wire[1379]), .S(n1889), .Z(
        \Data_Mem/n4859 ) );
  MUX U4283 ( .A(reg_target[2]), .B(data_mem_out_wire[1378]), .S(n1889), .Z(
        \Data_Mem/n4858 ) );
  IV U4284 ( .A(n1890), .Z(n1889) );
  MUX U4285 ( .A(data_mem_out_wire[1377]), .B(reg_target[1]), .S(n1890), .Z(
        \Data_Mem/n4857 ) );
  MUX U4286 ( .A(data_mem_out_wire[1376]), .B(reg_target[0]), .S(n1890), .Z(
        \Data_Mem/n4856 ) );
  AND U4287 ( .A(n1801), .B(n1884), .Z(n1890) );
  MUX U4288 ( .A(reg_target[31]), .B(data_mem_out_wire[1439]), .S(n1891), .Z(
        \Data_Mem/n4855 ) );
  MUX U4289 ( .A(reg_target[30]), .B(data_mem_out_wire[1438]), .S(n1891), .Z(
        \Data_Mem/n4854 ) );
  MUX U4290 ( .A(reg_target[29]), .B(data_mem_out_wire[1437]), .S(n1891), .Z(
        \Data_Mem/n4853 ) );
  MUX U4291 ( .A(reg_target[28]), .B(data_mem_out_wire[1436]), .S(n1891), .Z(
        \Data_Mem/n4852 ) );
  MUX U4292 ( .A(reg_target[27]), .B(data_mem_out_wire[1435]), .S(n1891), .Z(
        \Data_Mem/n4851 ) );
  MUX U4293 ( .A(reg_target[26]), .B(data_mem_out_wire[1434]), .S(n1891), .Z(
        \Data_Mem/n4850 ) );
  MUX U4294 ( .A(reg_target[25]), .B(data_mem_out_wire[1433]), .S(n1891), .Z(
        \Data_Mem/n4849 ) );
  MUX U4295 ( .A(reg_target[24]), .B(data_mem_out_wire[1432]), .S(n1891), .Z(
        \Data_Mem/n4848 ) );
  MUX U4296 ( .A(reg_target[23]), .B(data_mem_out_wire[1431]), .S(n1891), .Z(
        \Data_Mem/n4847 ) );
  MUX U4297 ( .A(reg_target[22]), .B(data_mem_out_wire[1430]), .S(n1891), .Z(
        \Data_Mem/n4846 ) );
  MUX U4298 ( .A(reg_target[21]), .B(data_mem_out_wire[1429]), .S(n1891), .Z(
        \Data_Mem/n4845 ) );
  MUX U4299 ( .A(reg_target[20]), .B(data_mem_out_wire[1428]), .S(n1891), .Z(
        \Data_Mem/n4844 ) );
  MUX U4300 ( .A(reg_target[19]), .B(data_mem_out_wire[1427]), .S(n1891), .Z(
        \Data_Mem/n4843 ) );
  MUX U4301 ( .A(reg_target[18]), .B(data_mem_out_wire[1426]), .S(n1891), .Z(
        \Data_Mem/n4842 ) );
  MUX U4302 ( .A(reg_target[17]), .B(data_mem_out_wire[1425]), .S(n1891), .Z(
        \Data_Mem/n4841 ) );
  MUX U4303 ( .A(reg_target[16]), .B(data_mem_out_wire[1424]), .S(n1891), .Z(
        \Data_Mem/n4840 ) );
  MUX U4304 ( .A(reg_target[15]), .B(data_mem_out_wire[1423]), .S(n1891), .Z(
        \Data_Mem/n4839 ) );
  MUX U4305 ( .A(reg_target[14]), .B(data_mem_out_wire[1422]), .S(n1891), .Z(
        \Data_Mem/n4838 ) );
  MUX U4306 ( .A(reg_target[13]), .B(data_mem_out_wire[1421]), .S(n1891), .Z(
        \Data_Mem/n4837 ) );
  MUX U4307 ( .A(reg_target[12]), .B(data_mem_out_wire[1420]), .S(n1891), .Z(
        \Data_Mem/n4836 ) );
  MUX U4308 ( .A(reg_target[11]), .B(data_mem_out_wire[1419]), .S(n1891), .Z(
        \Data_Mem/n4835 ) );
  MUX U4309 ( .A(reg_target[10]), .B(data_mem_out_wire[1418]), .S(n1891), .Z(
        \Data_Mem/n4834 ) );
  MUX U4310 ( .A(reg_target[9]), .B(data_mem_out_wire[1417]), .S(n1891), .Z(
        \Data_Mem/n4833 ) );
  MUX U4311 ( .A(reg_target[8]), .B(data_mem_out_wire[1416]), .S(n1891), .Z(
        \Data_Mem/n4832 ) );
  MUX U4312 ( .A(reg_target[7]), .B(data_mem_out_wire[1415]), .S(n1891), .Z(
        \Data_Mem/n4831 ) );
  MUX U4313 ( .A(reg_target[6]), .B(data_mem_out_wire[1414]), .S(n1891), .Z(
        \Data_Mem/n4830 ) );
  MUX U4314 ( .A(reg_target[5]), .B(data_mem_out_wire[1413]), .S(n1891), .Z(
        \Data_Mem/n4829 ) );
  MUX U4315 ( .A(reg_target[4]), .B(data_mem_out_wire[1412]), .S(n1891), .Z(
        \Data_Mem/n4828 ) );
  MUX U4316 ( .A(reg_target[3]), .B(data_mem_out_wire[1411]), .S(n1891), .Z(
        \Data_Mem/n4827 ) );
  MUX U4317 ( .A(reg_target[2]), .B(data_mem_out_wire[1410]), .S(n1891), .Z(
        \Data_Mem/n4826 ) );
  IV U4318 ( .A(n1892), .Z(n1891) );
  MUX U4319 ( .A(data_mem_out_wire[1409]), .B(reg_target[1]), .S(n1892), .Z(
        \Data_Mem/n4825 ) );
  MUX U4320 ( .A(data_mem_out_wire[1408]), .B(reg_target[0]), .S(n1892), .Z(
        \Data_Mem/n4824 ) );
  AND U4321 ( .A(n1804), .B(n1884), .Z(n1892) );
  MUX U4322 ( .A(reg_target[31]), .B(data_mem_out_wire[1471]), .S(n1893), .Z(
        \Data_Mem/n4823 ) );
  MUX U4323 ( .A(reg_target[30]), .B(data_mem_out_wire[1470]), .S(n1893), .Z(
        \Data_Mem/n4822 ) );
  MUX U4324 ( .A(reg_target[29]), .B(data_mem_out_wire[1469]), .S(n1893), .Z(
        \Data_Mem/n4821 ) );
  MUX U4325 ( .A(reg_target[28]), .B(data_mem_out_wire[1468]), .S(n1893), .Z(
        \Data_Mem/n4820 ) );
  MUX U4326 ( .A(reg_target[27]), .B(data_mem_out_wire[1467]), .S(n1893), .Z(
        \Data_Mem/n4819 ) );
  MUX U4327 ( .A(reg_target[26]), .B(data_mem_out_wire[1466]), .S(n1893), .Z(
        \Data_Mem/n4818 ) );
  MUX U4328 ( .A(reg_target[25]), .B(data_mem_out_wire[1465]), .S(n1893), .Z(
        \Data_Mem/n4817 ) );
  MUX U4329 ( .A(reg_target[24]), .B(data_mem_out_wire[1464]), .S(n1893), .Z(
        \Data_Mem/n4816 ) );
  MUX U4330 ( .A(reg_target[23]), .B(data_mem_out_wire[1463]), .S(n1893), .Z(
        \Data_Mem/n4815 ) );
  MUX U4331 ( .A(reg_target[22]), .B(data_mem_out_wire[1462]), .S(n1893), .Z(
        \Data_Mem/n4814 ) );
  MUX U4332 ( .A(reg_target[21]), .B(data_mem_out_wire[1461]), .S(n1893), .Z(
        \Data_Mem/n4813 ) );
  MUX U4333 ( .A(reg_target[20]), .B(data_mem_out_wire[1460]), .S(n1893), .Z(
        \Data_Mem/n4812 ) );
  MUX U4334 ( .A(reg_target[19]), .B(data_mem_out_wire[1459]), .S(n1893), .Z(
        \Data_Mem/n4811 ) );
  MUX U4335 ( .A(reg_target[18]), .B(data_mem_out_wire[1458]), .S(n1893), .Z(
        \Data_Mem/n4810 ) );
  MUX U4336 ( .A(reg_target[17]), .B(data_mem_out_wire[1457]), .S(n1893), .Z(
        \Data_Mem/n4809 ) );
  MUX U4337 ( .A(reg_target[16]), .B(data_mem_out_wire[1456]), .S(n1893), .Z(
        \Data_Mem/n4808 ) );
  MUX U4338 ( .A(reg_target[15]), .B(data_mem_out_wire[1455]), .S(n1893), .Z(
        \Data_Mem/n4807 ) );
  MUX U4339 ( .A(reg_target[14]), .B(data_mem_out_wire[1454]), .S(n1893), .Z(
        \Data_Mem/n4806 ) );
  MUX U4340 ( .A(reg_target[13]), .B(data_mem_out_wire[1453]), .S(n1893), .Z(
        \Data_Mem/n4805 ) );
  MUX U4341 ( .A(reg_target[12]), .B(data_mem_out_wire[1452]), .S(n1893), .Z(
        \Data_Mem/n4804 ) );
  MUX U4342 ( .A(reg_target[11]), .B(data_mem_out_wire[1451]), .S(n1893), .Z(
        \Data_Mem/n4803 ) );
  MUX U4343 ( .A(reg_target[10]), .B(data_mem_out_wire[1450]), .S(n1893), .Z(
        \Data_Mem/n4802 ) );
  MUX U4344 ( .A(reg_target[9]), .B(data_mem_out_wire[1449]), .S(n1893), .Z(
        \Data_Mem/n4801 ) );
  MUX U4345 ( .A(reg_target[8]), .B(data_mem_out_wire[1448]), .S(n1893), .Z(
        \Data_Mem/n4800 ) );
  MUX U4346 ( .A(reg_target[7]), .B(data_mem_out_wire[1447]), .S(n1893), .Z(
        \Data_Mem/n4799 ) );
  MUX U4347 ( .A(reg_target[6]), .B(data_mem_out_wire[1446]), .S(n1893), .Z(
        \Data_Mem/n4798 ) );
  MUX U4348 ( .A(reg_target[5]), .B(data_mem_out_wire[1445]), .S(n1893), .Z(
        \Data_Mem/n4797 ) );
  MUX U4349 ( .A(reg_target[4]), .B(data_mem_out_wire[1444]), .S(n1893), .Z(
        \Data_Mem/n4796 ) );
  MUX U4350 ( .A(reg_target[3]), .B(data_mem_out_wire[1443]), .S(n1893), .Z(
        \Data_Mem/n4795 ) );
  MUX U4351 ( .A(reg_target[2]), .B(data_mem_out_wire[1442]), .S(n1893), .Z(
        \Data_Mem/n4794 ) );
  IV U4352 ( .A(n1894), .Z(n1893) );
  MUX U4353 ( .A(data_mem_out_wire[1441]), .B(reg_target[1]), .S(n1894), .Z(
        \Data_Mem/n4793 ) );
  MUX U4354 ( .A(data_mem_out_wire[1440]), .B(reg_target[0]), .S(n1894), .Z(
        \Data_Mem/n4792 ) );
  AND U4355 ( .A(n1807), .B(n1884), .Z(n1894) );
  MUX U4356 ( .A(reg_target[31]), .B(data_mem_out_wire[1503]), .S(n1895), .Z(
        \Data_Mem/n4791 ) );
  MUX U4357 ( .A(reg_target[30]), .B(data_mem_out_wire[1502]), .S(n1895), .Z(
        \Data_Mem/n4790 ) );
  MUX U4358 ( .A(reg_target[29]), .B(data_mem_out_wire[1501]), .S(n1895), .Z(
        \Data_Mem/n4789 ) );
  MUX U4359 ( .A(reg_target[28]), .B(data_mem_out_wire[1500]), .S(n1895), .Z(
        \Data_Mem/n4788 ) );
  MUX U4360 ( .A(reg_target[27]), .B(data_mem_out_wire[1499]), .S(n1895), .Z(
        \Data_Mem/n4787 ) );
  MUX U4361 ( .A(reg_target[26]), .B(data_mem_out_wire[1498]), .S(n1895), .Z(
        \Data_Mem/n4786 ) );
  MUX U4362 ( .A(reg_target[25]), .B(data_mem_out_wire[1497]), .S(n1895), .Z(
        \Data_Mem/n4785 ) );
  MUX U4363 ( .A(reg_target[24]), .B(data_mem_out_wire[1496]), .S(n1895), .Z(
        \Data_Mem/n4784 ) );
  MUX U4364 ( .A(reg_target[23]), .B(data_mem_out_wire[1495]), .S(n1895), .Z(
        \Data_Mem/n4783 ) );
  MUX U4365 ( .A(reg_target[22]), .B(data_mem_out_wire[1494]), .S(n1895), .Z(
        \Data_Mem/n4782 ) );
  MUX U4366 ( .A(reg_target[21]), .B(data_mem_out_wire[1493]), .S(n1895), .Z(
        \Data_Mem/n4781 ) );
  MUX U4367 ( .A(reg_target[20]), .B(data_mem_out_wire[1492]), .S(n1895), .Z(
        \Data_Mem/n4780 ) );
  MUX U4368 ( .A(reg_target[19]), .B(data_mem_out_wire[1491]), .S(n1895), .Z(
        \Data_Mem/n4779 ) );
  MUX U4369 ( .A(reg_target[18]), .B(data_mem_out_wire[1490]), .S(n1895), .Z(
        \Data_Mem/n4778 ) );
  MUX U4370 ( .A(reg_target[17]), .B(data_mem_out_wire[1489]), .S(n1895), .Z(
        \Data_Mem/n4777 ) );
  MUX U4371 ( .A(reg_target[16]), .B(data_mem_out_wire[1488]), .S(n1895), .Z(
        \Data_Mem/n4776 ) );
  MUX U4372 ( .A(reg_target[15]), .B(data_mem_out_wire[1487]), .S(n1895), .Z(
        \Data_Mem/n4775 ) );
  MUX U4373 ( .A(reg_target[14]), .B(data_mem_out_wire[1486]), .S(n1895), .Z(
        \Data_Mem/n4774 ) );
  MUX U4374 ( .A(reg_target[13]), .B(data_mem_out_wire[1485]), .S(n1895), .Z(
        \Data_Mem/n4773 ) );
  MUX U4375 ( .A(reg_target[12]), .B(data_mem_out_wire[1484]), .S(n1895), .Z(
        \Data_Mem/n4772 ) );
  MUX U4376 ( .A(reg_target[11]), .B(data_mem_out_wire[1483]), .S(n1895), .Z(
        \Data_Mem/n4771 ) );
  MUX U4377 ( .A(reg_target[10]), .B(data_mem_out_wire[1482]), .S(n1895), .Z(
        \Data_Mem/n4770 ) );
  MUX U4378 ( .A(reg_target[9]), .B(data_mem_out_wire[1481]), .S(n1895), .Z(
        \Data_Mem/n4769 ) );
  MUX U4379 ( .A(reg_target[8]), .B(data_mem_out_wire[1480]), .S(n1895), .Z(
        \Data_Mem/n4768 ) );
  MUX U4380 ( .A(reg_target[7]), .B(data_mem_out_wire[1479]), .S(n1895), .Z(
        \Data_Mem/n4767 ) );
  MUX U4381 ( .A(reg_target[6]), .B(data_mem_out_wire[1478]), .S(n1895), .Z(
        \Data_Mem/n4766 ) );
  MUX U4382 ( .A(reg_target[5]), .B(data_mem_out_wire[1477]), .S(n1895), .Z(
        \Data_Mem/n4765 ) );
  MUX U4383 ( .A(reg_target[4]), .B(data_mem_out_wire[1476]), .S(n1895), .Z(
        \Data_Mem/n4764 ) );
  MUX U4384 ( .A(reg_target[3]), .B(data_mem_out_wire[1475]), .S(n1895), .Z(
        \Data_Mem/n4763 ) );
  MUX U4385 ( .A(reg_target[2]), .B(data_mem_out_wire[1474]), .S(n1895), .Z(
        \Data_Mem/n4762 ) );
  IV U4386 ( .A(n1896), .Z(n1895) );
  MUX U4387 ( .A(data_mem_out_wire[1473]), .B(reg_target[1]), .S(n1896), .Z(
        \Data_Mem/n4761 ) );
  MUX U4388 ( .A(data_mem_out_wire[1472]), .B(reg_target[0]), .S(n1896), .Z(
        \Data_Mem/n4760 ) );
  AND U4389 ( .A(n1810), .B(n1884), .Z(n1896) );
  MUX U4390 ( .A(data_mem_out_wire[1535]), .B(reg_target[31]), .S(n1897), .Z(
        \Data_Mem/n4759 ) );
  MUX U4391 ( .A(data_mem_out_wire[1534]), .B(reg_target[30]), .S(n1897), .Z(
        \Data_Mem/n4758 ) );
  MUX U4392 ( .A(data_mem_out_wire[1533]), .B(reg_target[29]), .S(n1897), .Z(
        \Data_Mem/n4757 ) );
  MUX U4393 ( .A(data_mem_out_wire[1532]), .B(reg_target[28]), .S(n1897), .Z(
        \Data_Mem/n4756 ) );
  MUX U4394 ( .A(data_mem_out_wire[1531]), .B(reg_target[27]), .S(n1897), .Z(
        \Data_Mem/n4755 ) );
  MUX U4395 ( .A(data_mem_out_wire[1530]), .B(reg_target[26]), .S(n1897), .Z(
        \Data_Mem/n4754 ) );
  MUX U4396 ( .A(data_mem_out_wire[1529]), .B(reg_target[25]), .S(n1897), .Z(
        \Data_Mem/n4753 ) );
  MUX U4397 ( .A(data_mem_out_wire[1528]), .B(reg_target[24]), .S(n1897), .Z(
        \Data_Mem/n4752 ) );
  MUX U4398 ( .A(data_mem_out_wire[1527]), .B(reg_target[23]), .S(n1897), .Z(
        \Data_Mem/n4751 ) );
  MUX U4399 ( .A(data_mem_out_wire[1526]), .B(reg_target[22]), .S(n1897), .Z(
        \Data_Mem/n4750 ) );
  MUX U4400 ( .A(data_mem_out_wire[1525]), .B(reg_target[21]), .S(n1897), .Z(
        \Data_Mem/n4749 ) );
  MUX U4401 ( .A(data_mem_out_wire[1524]), .B(reg_target[20]), .S(n1897), .Z(
        \Data_Mem/n4748 ) );
  MUX U4402 ( .A(data_mem_out_wire[1523]), .B(reg_target[19]), .S(n1897), .Z(
        \Data_Mem/n4747 ) );
  MUX U4403 ( .A(data_mem_out_wire[1522]), .B(reg_target[18]), .S(n1897), .Z(
        \Data_Mem/n4746 ) );
  MUX U4404 ( .A(data_mem_out_wire[1521]), .B(reg_target[17]), .S(n1897), .Z(
        \Data_Mem/n4745 ) );
  MUX U4405 ( .A(data_mem_out_wire[1520]), .B(reg_target[16]), .S(n1897), .Z(
        \Data_Mem/n4744 ) );
  MUX U4406 ( .A(data_mem_out_wire[1519]), .B(reg_target[15]), .S(n1897), .Z(
        \Data_Mem/n4743 ) );
  MUX U4407 ( .A(data_mem_out_wire[1518]), .B(reg_target[14]), .S(n1897), .Z(
        \Data_Mem/n4742 ) );
  MUX U4408 ( .A(data_mem_out_wire[1517]), .B(reg_target[13]), .S(n1897), .Z(
        \Data_Mem/n4741 ) );
  MUX U4409 ( .A(data_mem_out_wire[1516]), .B(reg_target[12]), .S(n1897), .Z(
        \Data_Mem/n4740 ) );
  MUX U4410 ( .A(data_mem_out_wire[1515]), .B(reg_target[11]), .S(n1897), .Z(
        \Data_Mem/n4739 ) );
  MUX U4411 ( .A(data_mem_out_wire[1514]), .B(reg_target[10]), .S(n1897), .Z(
        \Data_Mem/n4738 ) );
  MUX U4412 ( .A(data_mem_out_wire[1513]), .B(reg_target[9]), .S(n1897), .Z(
        \Data_Mem/n4737 ) );
  MUX U4413 ( .A(data_mem_out_wire[1512]), .B(reg_target[8]), .S(n1897), .Z(
        \Data_Mem/n4736 ) );
  MUX U4414 ( .A(data_mem_out_wire[1511]), .B(reg_target[7]), .S(n1897), .Z(
        \Data_Mem/n4735 ) );
  MUX U4415 ( .A(data_mem_out_wire[1510]), .B(reg_target[6]), .S(n1897), .Z(
        \Data_Mem/n4734 ) );
  MUX U4416 ( .A(data_mem_out_wire[1509]), .B(reg_target[5]), .S(n1897), .Z(
        \Data_Mem/n4733 ) );
  MUX U4417 ( .A(data_mem_out_wire[1508]), .B(reg_target[4]), .S(n1897), .Z(
        \Data_Mem/n4732 ) );
  MUX U4418 ( .A(data_mem_out_wire[1507]), .B(reg_target[3]), .S(n1897), .Z(
        \Data_Mem/n4731 ) );
  MUX U4419 ( .A(data_mem_out_wire[1506]), .B(reg_target[2]), .S(n1897), .Z(
        \Data_Mem/n4730 ) );
  MUX U4420 ( .A(data_mem_out_wire[1505]), .B(reg_target[1]), .S(n1897), .Z(
        \Data_Mem/n4729 ) );
  MUX U4421 ( .A(data_mem_out_wire[1504]), .B(reg_target[0]), .S(n1897), .Z(
        \Data_Mem/n4728 ) );
  AND U4422 ( .A(n1884), .B(n1830), .Z(n1897) );
  AND U4423 ( .A(n1831), .B(N24), .Z(n1884) );
  ANDN U4424 ( .B(n840), .A(n837), .Z(n1831) );
  MUX U4425 ( .A(data_mem_out_wire[1567]), .B(reg_target[31]), .S(n1898), .Z(
        \Data_Mem/n4727 ) );
  MUX U4426 ( .A(data_mem_out_wire[1566]), .B(reg_target[30]), .S(n1898), .Z(
        \Data_Mem/n4726 ) );
  MUX U4427 ( .A(data_mem_out_wire[1565]), .B(reg_target[29]), .S(n1898), .Z(
        \Data_Mem/n4725 ) );
  MUX U4428 ( .A(data_mem_out_wire[1564]), .B(reg_target[28]), .S(n1898), .Z(
        \Data_Mem/n4724 ) );
  MUX U4429 ( .A(data_mem_out_wire[1563]), .B(reg_target[27]), .S(n1898), .Z(
        \Data_Mem/n4723 ) );
  MUX U4430 ( .A(data_mem_out_wire[1562]), .B(reg_target[26]), .S(n1898), .Z(
        \Data_Mem/n4722 ) );
  MUX U4431 ( .A(data_mem_out_wire[1561]), .B(reg_target[25]), .S(n1898), .Z(
        \Data_Mem/n4721 ) );
  MUX U4432 ( .A(data_mem_out_wire[1560]), .B(reg_target[24]), .S(n1898), .Z(
        \Data_Mem/n4720 ) );
  MUX U4433 ( .A(data_mem_out_wire[1559]), .B(reg_target[23]), .S(n1898), .Z(
        \Data_Mem/n4719 ) );
  MUX U4434 ( .A(data_mem_out_wire[1558]), .B(reg_target[22]), .S(n1898), .Z(
        \Data_Mem/n4718 ) );
  MUX U4435 ( .A(data_mem_out_wire[1557]), .B(reg_target[21]), .S(n1898), .Z(
        \Data_Mem/n4717 ) );
  MUX U4436 ( .A(data_mem_out_wire[1556]), .B(reg_target[20]), .S(n1898), .Z(
        \Data_Mem/n4716 ) );
  MUX U4437 ( .A(data_mem_out_wire[1555]), .B(reg_target[19]), .S(n1898), .Z(
        \Data_Mem/n4715 ) );
  MUX U4438 ( .A(data_mem_out_wire[1554]), .B(reg_target[18]), .S(n1898), .Z(
        \Data_Mem/n4714 ) );
  MUX U4439 ( .A(data_mem_out_wire[1553]), .B(reg_target[17]), .S(n1898), .Z(
        \Data_Mem/n4713 ) );
  MUX U4440 ( .A(data_mem_out_wire[1552]), .B(reg_target[16]), .S(n1898), .Z(
        \Data_Mem/n4712 ) );
  MUX U4441 ( .A(data_mem_out_wire[1551]), .B(reg_target[15]), .S(n1898), .Z(
        \Data_Mem/n4711 ) );
  MUX U4442 ( .A(data_mem_out_wire[1550]), .B(reg_target[14]), .S(n1898), .Z(
        \Data_Mem/n4710 ) );
  MUX U4443 ( .A(data_mem_out_wire[1549]), .B(reg_target[13]), .S(n1898), .Z(
        \Data_Mem/n4709 ) );
  MUX U4444 ( .A(data_mem_out_wire[1548]), .B(reg_target[12]), .S(n1898), .Z(
        \Data_Mem/n4708 ) );
  MUX U4445 ( .A(data_mem_out_wire[1547]), .B(reg_target[11]), .S(n1898), .Z(
        \Data_Mem/n4707 ) );
  MUX U4446 ( .A(data_mem_out_wire[1546]), .B(reg_target[10]), .S(n1898), .Z(
        \Data_Mem/n4706 ) );
  MUX U4447 ( .A(data_mem_out_wire[1545]), .B(reg_target[9]), .S(n1898), .Z(
        \Data_Mem/n4705 ) );
  MUX U4448 ( .A(data_mem_out_wire[1544]), .B(reg_target[8]), .S(n1898), .Z(
        \Data_Mem/n4704 ) );
  MUX U4449 ( .A(data_mem_out_wire[1543]), .B(reg_target[7]), .S(n1898), .Z(
        \Data_Mem/n4703 ) );
  MUX U4450 ( .A(data_mem_out_wire[1542]), .B(reg_target[6]), .S(n1898), .Z(
        \Data_Mem/n4702 ) );
  MUX U4451 ( .A(data_mem_out_wire[1541]), .B(reg_target[5]), .S(n1898), .Z(
        \Data_Mem/n4701 ) );
  MUX U4452 ( .A(data_mem_out_wire[1540]), .B(reg_target[4]), .S(n1898), .Z(
        \Data_Mem/n4700 ) );
  MUX U4453 ( .A(data_mem_out_wire[1539]), .B(reg_target[3]), .S(n1898), .Z(
        \Data_Mem/n4699 ) );
  MUX U4454 ( .A(data_mem_out_wire[1538]), .B(reg_target[2]), .S(n1898), .Z(
        \Data_Mem/n4698 ) );
  MUX U4455 ( .A(data_mem_out_wire[1537]), .B(reg_target[1]), .S(n1898), .Z(
        \Data_Mem/n4697 ) );
  MUX U4456 ( .A(data_mem_out_wire[1536]), .B(reg_target[0]), .S(n1898), .Z(
        \Data_Mem/n4696 ) );
  ANDN U4457 ( .B(n1791), .A(n1899), .Z(n1898) );
  ANDN U4458 ( .B(n1900), .A(n1901), .Z(n1791) );
  MUX U4459 ( .A(data_mem_out_wire[1599]), .B(reg_target[31]), .S(n1902), .Z(
        \Data_Mem/n4695 ) );
  MUX U4460 ( .A(data_mem_out_wire[1598]), .B(reg_target[30]), .S(n1902), .Z(
        \Data_Mem/n4694 ) );
  MUX U4461 ( .A(data_mem_out_wire[1597]), .B(reg_target[29]), .S(n1902), .Z(
        \Data_Mem/n4693 ) );
  MUX U4462 ( .A(data_mem_out_wire[1596]), .B(reg_target[28]), .S(n1902), .Z(
        \Data_Mem/n4692 ) );
  MUX U4463 ( .A(data_mem_out_wire[1595]), .B(reg_target[27]), .S(n1902), .Z(
        \Data_Mem/n4691 ) );
  MUX U4464 ( .A(data_mem_out_wire[1594]), .B(reg_target[26]), .S(n1902), .Z(
        \Data_Mem/n4690 ) );
  MUX U4465 ( .A(data_mem_out_wire[1593]), .B(reg_target[25]), .S(n1902), .Z(
        \Data_Mem/n4689 ) );
  MUX U4466 ( .A(data_mem_out_wire[1592]), .B(reg_target[24]), .S(n1902), .Z(
        \Data_Mem/n4688 ) );
  MUX U4467 ( .A(data_mem_out_wire[1591]), .B(reg_target[23]), .S(n1902), .Z(
        \Data_Mem/n4687 ) );
  MUX U4468 ( .A(data_mem_out_wire[1590]), .B(reg_target[22]), .S(n1902), .Z(
        \Data_Mem/n4686 ) );
  MUX U4469 ( .A(data_mem_out_wire[1589]), .B(reg_target[21]), .S(n1902), .Z(
        \Data_Mem/n4685 ) );
  MUX U4470 ( .A(data_mem_out_wire[1588]), .B(reg_target[20]), .S(n1902), .Z(
        \Data_Mem/n4684 ) );
  MUX U4471 ( .A(data_mem_out_wire[1587]), .B(reg_target[19]), .S(n1902), .Z(
        \Data_Mem/n4683 ) );
  MUX U4472 ( .A(data_mem_out_wire[1586]), .B(reg_target[18]), .S(n1902), .Z(
        \Data_Mem/n4682 ) );
  MUX U4473 ( .A(data_mem_out_wire[1585]), .B(reg_target[17]), .S(n1902), .Z(
        \Data_Mem/n4681 ) );
  MUX U4474 ( .A(data_mem_out_wire[1584]), .B(reg_target[16]), .S(n1902), .Z(
        \Data_Mem/n4680 ) );
  MUX U4475 ( .A(data_mem_out_wire[1583]), .B(reg_target[15]), .S(n1902), .Z(
        \Data_Mem/n4679 ) );
  MUX U4476 ( .A(data_mem_out_wire[1582]), .B(reg_target[14]), .S(n1902), .Z(
        \Data_Mem/n4678 ) );
  MUX U4477 ( .A(data_mem_out_wire[1581]), .B(reg_target[13]), .S(n1902), .Z(
        \Data_Mem/n4677 ) );
  MUX U4478 ( .A(data_mem_out_wire[1580]), .B(reg_target[12]), .S(n1902), .Z(
        \Data_Mem/n4676 ) );
  MUX U4479 ( .A(data_mem_out_wire[1579]), .B(reg_target[11]), .S(n1902), .Z(
        \Data_Mem/n4675 ) );
  MUX U4480 ( .A(data_mem_out_wire[1578]), .B(reg_target[10]), .S(n1902), .Z(
        \Data_Mem/n4674 ) );
  MUX U4481 ( .A(data_mem_out_wire[1577]), .B(reg_target[9]), .S(n1902), .Z(
        \Data_Mem/n4673 ) );
  MUX U4482 ( .A(data_mem_out_wire[1576]), .B(reg_target[8]), .S(n1902), .Z(
        \Data_Mem/n4672 ) );
  MUX U4483 ( .A(data_mem_out_wire[1575]), .B(reg_target[7]), .S(n1902), .Z(
        \Data_Mem/n4671 ) );
  MUX U4484 ( .A(data_mem_out_wire[1574]), .B(reg_target[6]), .S(n1902), .Z(
        \Data_Mem/n4670 ) );
  MUX U4485 ( .A(data_mem_out_wire[1573]), .B(reg_target[5]), .S(n1902), .Z(
        \Data_Mem/n4669 ) );
  MUX U4486 ( .A(data_mem_out_wire[1572]), .B(reg_target[4]), .S(n1902), .Z(
        \Data_Mem/n4668 ) );
  MUX U4487 ( .A(data_mem_out_wire[1571]), .B(reg_target[3]), .S(n1902), .Z(
        \Data_Mem/n4667 ) );
  MUX U4488 ( .A(data_mem_out_wire[1570]), .B(reg_target[2]), .S(n1902), .Z(
        \Data_Mem/n4666 ) );
  MUX U4489 ( .A(data_mem_out_wire[1569]), .B(reg_target[1]), .S(n1902), .Z(
        \Data_Mem/n4665 ) );
  MUX U4490 ( .A(data_mem_out_wire[1568]), .B(reg_target[0]), .S(n1902), .Z(
        \Data_Mem/n4664 ) );
  ANDN U4491 ( .B(n1795), .A(n1899), .Z(n1902) );
  ANDN U4492 ( .B(n1903), .A(n1901), .Z(n1795) );
  MUX U4493 ( .A(data_mem_out_wire[1631]), .B(reg_target[31]), .S(n1904), .Z(
        \Data_Mem/n4663 ) );
  MUX U4494 ( .A(data_mem_out_wire[1630]), .B(reg_target[30]), .S(n1904), .Z(
        \Data_Mem/n4662 ) );
  MUX U4495 ( .A(data_mem_out_wire[1629]), .B(reg_target[29]), .S(n1904), .Z(
        \Data_Mem/n4661 ) );
  MUX U4496 ( .A(data_mem_out_wire[1628]), .B(reg_target[28]), .S(n1904), .Z(
        \Data_Mem/n4660 ) );
  MUX U4497 ( .A(data_mem_out_wire[1627]), .B(reg_target[27]), .S(n1904), .Z(
        \Data_Mem/n4659 ) );
  MUX U4498 ( .A(data_mem_out_wire[1626]), .B(reg_target[26]), .S(n1904), .Z(
        \Data_Mem/n4658 ) );
  MUX U4499 ( .A(data_mem_out_wire[1625]), .B(reg_target[25]), .S(n1904), .Z(
        \Data_Mem/n4657 ) );
  MUX U4500 ( .A(data_mem_out_wire[1624]), .B(reg_target[24]), .S(n1904), .Z(
        \Data_Mem/n4656 ) );
  MUX U4501 ( .A(data_mem_out_wire[1623]), .B(reg_target[23]), .S(n1904), .Z(
        \Data_Mem/n4655 ) );
  MUX U4502 ( .A(data_mem_out_wire[1622]), .B(reg_target[22]), .S(n1904), .Z(
        \Data_Mem/n4654 ) );
  MUX U4503 ( .A(data_mem_out_wire[1621]), .B(reg_target[21]), .S(n1904), .Z(
        \Data_Mem/n4653 ) );
  MUX U4504 ( .A(data_mem_out_wire[1620]), .B(reg_target[20]), .S(n1904), .Z(
        \Data_Mem/n4652 ) );
  MUX U4505 ( .A(data_mem_out_wire[1619]), .B(reg_target[19]), .S(n1904), .Z(
        \Data_Mem/n4651 ) );
  MUX U4506 ( .A(data_mem_out_wire[1618]), .B(reg_target[18]), .S(n1904), .Z(
        \Data_Mem/n4650 ) );
  MUX U4507 ( .A(data_mem_out_wire[1617]), .B(reg_target[17]), .S(n1904), .Z(
        \Data_Mem/n4649 ) );
  MUX U4508 ( .A(data_mem_out_wire[1616]), .B(reg_target[16]), .S(n1904), .Z(
        \Data_Mem/n4648 ) );
  MUX U4509 ( .A(data_mem_out_wire[1615]), .B(reg_target[15]), .S(n1904), .Z(
        \Data_Mem/n4647 ) );
  MUX U4510 ( .A(data_mem_out_wire[1614]), .B(reg_target[14]), .S(n1904), .Z(
        \Data_Mem/n4646 ) );
  MUX U4511 ( .A(data_mem_out_wire[1613]), .B(reg_target[13]), .S(n1904), .Z(
        \Data_Mem/n4645 ) );
  MUX U4512 ( .A(data_mem_out_wire[1612]), .B(reg_target[12]), .S(n1904), .Z(
        \Data_Mem/n4644 ) );
  MUX U4513 ( .A(data_mem_out_wire[1611]), .B(reg_target[11]), .S(n1904), .Z(
        \Data_Mem/n4643 ) );
  MUX U4514 ( .A(data_mem_out_wire[1610]), .B(reg_target[10]), .S(n1904), .Z(
        \Data_Mem/n4642 ) );
  MUX U4515 ( .A(data_mem_out_wire[1609]), .B(reg_target[9]), .S(n1904), .Z(
        \Data_Mem/n4641 ) );
  MUX U4516 ( .A(data_mem_out_wire[1608]), .B(reg_target[8]), .S(n1904), .Z(
        \Data_Mem/n4640 ) );
  MUX U4517 ( .A(data_mem_out_wire[1607]), .B(reg_target[7]), .S(n1904), .Z(
        \Data_Mem/n4639 ) );
  MUX U4518 ( .A(data_mem_out_wire[1606]), .B(reg_target[6]), .S(n1904), .Z(
        \Data_Mem/n4638 ) );
  MUX U4519 ( .A(data_mem_out_wire[1605]), .B(reg_target[5]), .S(n1904), .Z(
        \Data_Mem/n4637 ) );
  MUX U4520 ( .A(data_mem_out_wire[1604]), .B(reg_target[4]), .S(n1904), .Z(
        \Data_Mem/n4636 ) );
  MUX U4521 ( .A(data_mem_out_wire[1603]), .B(reg_target[3]), .S(n1904), .Z(
        \Data_Mem/n4635 ) );
  MUX U4522 ( .A(data_mem_out_wire[1602]), .B(reg_target[2]), .S(n1904), .Z(
        \Data_Mem/n4634 ) );
  MUX U4523 ( .A(data_mem_out_wire[1601]), .B(reg_target[1]), .S(n1904), .Z(
        \Data_Mem/n4633 ) );
  MUX U4524 ( .A(data_mem_out_wire[1600]), .B(reg_target[0]), .S(n1904), .Z(
        \Data_Mem/n4632 ) );
  ANDN U4525 ( .B(n1798), .A(n1899), .Z(n1904) );
  ANDN U4526 ( .B(n1905), .A(n1901), .Z(n1798) );
  MUX U4527 ( .A(data_mem_out_wire[1663]), .B(reg_target[31]), .S(n1906), .Z(
        \Data_Mem/n4631 ) );
  MUX U4528 ( .A(data_mem_out_wire[1662]), .B(reg_target[30]), .S(n1906), .Z(
        \Data_Mem/n4630 ) );
  MUX U4529 ( .A(data_mem_out_wire[1661]), .B(reg_target[29]), .S(n1906), .Z(
        \Data_Mem/n4629 ) );
  MUX U4530 ( .A(data_mem_out_wire[1660]), .B(reg_target[28]), .S(n1906), .Z(
        \Data_Mem/n4628 ) );
  MUX U4531 ( .A(data_mem_out_wire[1659]), .B(reg_target[27]), .S(n1906), .Z(
        \Data_Mem/n4627 ) );
  MUX U4532 ( .A(data_mem_out_wire[1658]), .B(reg_target[26]), .S(n1906), .Z(
        \Data_Mem/n4626 ) );
  MUX U4533 ( .A(data_mem_out_wire[1657]), .B(reg_target[25]), .S(n1906), .Z(
        \Data_Mem/n4625 ) );
  MUX U4534 ( .A(data_mem_out_wire[1656]), .B(reg_target[24]), .S(n1906), .Z(
        \Data_Mem/n4624 ) );
  MUX U4535 ( .A(data_mem_out_wire[1655]), .B(reg_target[23]), .S(n1906), .Z(
        \Data_Mem/n4623 ) );
  MUX U4536 ( .A(data_mem_out_wire[1654]), .B(reg_target[22]), .S(n1906), .Z(
        \Data_Mem/n4622 ) );
  MUX U4537 ( .A(data_mem_out_wire[1653]), .B(reg_target[21]), .S(n1906), .Z(
        \Data_Mem/n4621 ) );
  MUX U4538 ( .A(data_mem_out_wire[1652]), .B(reg_target[20]), .S(n1906), .Z(
        \Data_Mem/n4620 ) );
  MUX U4539 ( .A(data_mem_out_wire[1651]), .B(reg_target[19]), .S(n1906), .Z(
        \Data_Mem/n4619 ) );
  MUX U4540 ( .A(data_mem_out_wire[1650]), .B(reg_target[18]), .S(n1906), .Z(
        \Data_Mem/n4618 ) );
  MUX U4541 ( .A(data_mem_out_wire[1649]), .B(reg_target[17]), .S(n1906), .Z(
        \Data_Mem/n4617 ) );
  MUX U4542 ( .A(data_mem_out_wire[1648]), .B(reg_target[16]), .S(n1906), .Z(
        \Data_Mem/n4616 ) );
  MUX U4543 ( .A(data_mem_out_wire[1647]), .B(reg_target[15]), .S(n1906), .Z(
        \Data_Mem/n4615 ) );
  MUX U4544 ( .A(data_mem_out_wire[1646]), .B(reg_target[14]), .S(n1906), .Z(
        \Data_Mem/n4614 ) );
  MUX U4545 ( .A(data_mem_out_wire[1645]), .B(reg_target[13]), .S(n1906), .Z(
        \Data_Mem/n4613 ) );
  MUX U4546 ( .A(data_mem_out_wire[1644]), .B(reg_target[12]), .S(n1906), .Z(
        \Data_Mem/n4612 ) );
  MUX U4547 ( .A(data_mem_out_wire[1643]), .B(reg_target[11]), .S(n1906), .Z(
        \Data_Mem/n4611 ) );
  MUX U4548 ( .A(data_mem_out_wire[1642]), .B(reg_target[10]), .S(n1906), .Z(
        \Data_Mem/n4610 ) );
  MUX U4549 ( .A(data_mem_out_wire[1641]), .B(reg_target[9]), .S(n1906), .Z(
        \Data_Mem/n4609 ) );
  MUX U4550 ( .A(data_mem_out_wire[1640]), .B(reg_target[8]), .S(n1906), .Z(
        \Data_Mem/n4608 ) );
  MUX U4551 ( .A(data_mem_out_wire[1639]), .B(reg_target[7]), .S(n1906), .Z(
        \Data_Mem/n4607 ) );
  MUX U4552 ( .A(data_mem_out_wire[1638]), .B(reg_target[6]), .S(n1906), .Z(
        \Data_Mem/n4606 ) );
  MUX U4553 ( .A(data_mem_out_wire[1637]), .B(reg_target[5]), .S(n1906), .Z(
        \Data_Mem/n4605 ) );
  MUX U4554 ( .A(data_mem_out_wire[1636]), .B(reg_target[4]), .S(n1906), .Z(
        \Data_Mem/n4604 ) );
  MUX U4555 ( .A(data_mem_out_wire[1635]), .B(reg_target[3]), .S(n1906), .Z(
        \Data_Mem/n4603 ) );
  MUX U4556 ( .A(data_mem_out_wire[1634]), .B(reg_target[2]), .S(n1906), .Z(
        \Data_Mem/n4602 ) );
  MUX U4557 ( .A(data_mem_out_wire[1633]), .B(reg_target[1]), .S(n1906), .Z(
        \Data_Mem/n4601 ) );
  MUX U4558 ( .A(data_mem_out_wire[1632]), .B(reg_target[0]), .S(n1906), .Z(
        \Data_Mem/n4600 ) );
  ANDN U4559 ( .B(n1801), .A(n1899), .Z(n1906) );
  ANDN U4560 ( .B(n1907), .A(n1901), .Z(n1801) );
  MUX U4561 ( .A(data_mem_out_wire[1695]), .B(reg_target[31]), .S(n1908), .Z(
        \Data_Mem/n4599 ) );
  MUX U4562 ( .A(data_mem_out_wire[1694]), .B(reg_target[30]), .S(n1908), .Z(
        \Data_Mem/n4598 ) );
  MUX U4563 ( .A(data_mem_out_wire[1693]), .B(reg_target[29]), .S(n1908), .Z(
        \Data_Mem/n4597 ) );
  MUX U4564 ( .A(data_mem_out_wire[1692]), .B(reg_target[28]), .S(n1908), .Z(
        \Data_Mem/n4596 ) );
  MUX U4565 ( .A(data_mem_out_wire[1691]), .B(reg_target[27]), .S(n1908), .Z(
        \Data_Mem/n4595 ) );
  MUX U4566 ( .A(data_mem_out_wire[1690]), .B(reg_target[26]), .S(n1908), .Z(
        \Data_Mem/n4594 ) );
  MUX U4567 ( .A(data_mem_out_wire[1689]), .B(reg_target[25]), .S(n1908), .Z(
        \Data_Mem/n4593 ) );
  MUX U4568 ( .A(data_mem_out_wire[1688]), .B(reg_target[24]), .S(n1908), .Z(
        \Data_Mem/n4592 ) );
  MUX U4569 ( .A(data_mem_out_wire[1687]), .B(reg_target[23]), .S(n1908), .Z(
        \Data_Mem/n4591 ) );
  MUX U4570 ( .A(data_mem_out_wire[1686]), .B(reg_target[22]), .S(n1908), .Z(
        \Data_Mem/n4590 ) );
  MUX U4571 ( .A(data_mem_out_wire[1685]), .B(reg_target[21]), .S(n1908), .Z(
        \Data_Mem/n4589 ) );
  MUX U4572 ( .A(data_mem_out_wire[1684]), .B(reg_target[20]), .S(n1908), .Z(
        \Data_Mem/n4588 ) );
  MUX U4573 ( .A(data_mem_out_wire[1683]), .B(reg_target[19]), .S(n1908), .Z(
        \Data_Mem/n4587 ) );
  MUX U4574 ( .A(data_mem_out_wire[1682]), .B(reg_target[18]), .S(n1908), .Z(
        \Data_Mem/n4586 ) );
  MUX U4575 ( .A(data_mem_out_wire[1681]), .B(reg_target[17]), .S(n1908), .Z(
        \Data_Mem/n4585 ) );
  MUX U4576 ( .A(data_mem_out_wire[1680]), .B(reg_target[16]), .S(n1908), .Z(
        \Data_Mem/n4584 ) );
  MUX U4577 ( .A(data_mem_out_wire[1679]), .B(reg_target[15]), .S(n1908), .Z(
        \Data_Mem/n4583 ) );
  MUX U4578 ( .A(data_mem_out_wire[1678]), .B(reg_target[14]), .S(n1908), .Z(
        \Data_Mem/n4582 ) );
  MUX U4579 ( .A(data_mem_out_wire[1677]), .B(reg_target[13]), .S(n1908), .Z(
        \Data_Mem/n4581 ) );
  MUX U4580 ( .A(data_mem_out_wire[1676]), .B(reg_target[12]), .S(n1908), .Z(
        \Data_Mem/n4580 ) );
  MUX U4581 ( .A(data_mem_out_wire[1675]), .B(reg_target[11]), .S(n1908), .Z(
        \Data_Mem/n4579 ) );
  MUX U4582 ( .A(data_mem_out_wire[1674]), .B(reg_target[10]), .S(n1908), .Z(
        \Data_Mem/n4578 ) );
  MUX U4583 ( .A(data_mem_out_wire[1673]), .B(reg_target[9]), .S(n1908), .Z(
        \Data_Mem/n4577 ) );
  MUX U4584 ( .A(data_mem_out_wire[1672]), .B(reg_target[8]), .S(n1908), .Z(
        \Data_Mem/n4576 ) );
  MUX U4585 ( .A(data_mem_out_wire[1671]), .B(reg_target[7]), .S(n1908), .Z(
        \Data_Mem/n4575 ) );
  MUX U4586 ( .A(data_mem_out_wire[1670]), .B(reg_target[6]), .S(n1908), .Z(
        \Data_Mem/n4574 ) );
  MUX U4587 ( .A(data_mem_out_wire[1669]), .B(reg_target[5]), .S(n1908), .Z(
        \Data_Mem/n4573 ) );
  MUX U4588 ( .A(data_mem_out_wire[1668]), .B(reg_target[4]), .S(n1908), .Z(
        \Data_Mem/n4572 ) );
  MUX U4589 ( .A(data_mem_out_wire[1667]), .B(reg_target[3]), .S(n1908), .Z(
        \Data_Mem/n4571 ) );
  MUX U4590 ( .A(data_mem_out_wire[1666]), .B(reg_target[2]), .S(n1908), .Z(
        \Data_Mem/n4570 ) );
  MUX U4591 ( .A(data_mem_out_wire[1665]), .B(reg_target[1]), .S(n1908), .Z(
        \Data_Mem/n4569 ) );
  MUX U4592 ( .A(data_mem_out_wire[1664]), .B(reg_target[0]), .S(n1908), .Z(
        \Data_Mem/n4568 ) );
  ANDN U4593 ( .B(n1804), .A(n1899), .Z(n1908) );
  ANDN U4594 ( .B(n1909), .A(n1901), .Z(n1804) );
  MUX U4595 ( .A(data_mem_out_wire[1727]), .B(reg_target[31]), .S(n1910), .Z(
        \Data_Mem/n4567 ) );
  MUX U4596 ( .A(data_mem_out_wire[1726]), .B(reg_target[30]), .S(n1910), .Z(
        \Data_Mem/n4566 ) );
  MUX U4597 ( .A(data_mem_out_wire[1725]), .B(reg_target[29]), .S(n1910), .Z(
        \Data_Mem/n4565 ) );
  MUX U4598 ( .A(data_mem_out_wire[1724]), .B(reg_target[28]), .S(n1910), .Z(
        \Data_Mem/n4564 ) );
  MUX U4599 ( .A(data_mem_out_wire[1723]), .B(reg_target[27]), .S(n1910), .Z(
        \Data_Mem/n4563 ) );
  MUX U4600 ( .A(data_mem_out_wire[1722]), .B(reg_target[26]), .S(n1910), .Z(
        \Data_Mem/n4562 ) );
  MUX U4601 ( .A(data_mem_out_wire[1721]), .B(reg_target[25]), .S(n1910), .Z(
        \Data_Mem/n4561 ) );
  MUX U4602 ( .A(data_mem_out_wire[1720]), .B(reg_target[24]), .S(n1910), .Z(
        \Data_Mem/n4560 ) );
  MUX U4603 ( .A(data_mem_out_wire[1719]), .B(reg_target[23]), .S(n1910), .Z(
        \Data_Mem/n4559 ) );
  MUX U4604 ( .A(data_mem_out_wire[1718]), .B(reg_target[22]), .S(n1910), .Z(
        \Data_Mem/n4558 ) );
  MUX U4605 ( .A(data_mem_out_wire[1717]), .B(reg_target[21]), .S(n1910), .Z(
        \Data_Mem/n4557 ) );
  MUX U4606 ( .A(data_mem_out_wire[1716]), .B(reg_target[20]), .S(n1910), .Z(
        \Data_Mem/n4556 ) );
  MUX U4607 ( .A(data_mem_out_wire[1715]), .B(reg_target[19]), .S(n1910), .Z(
        \Data_Mem/n4555 ) );
  MUX U4608 ( .A(data_mem_out_wire[1714]), .B(reg_target[18]), .S(n1910), .Z(
        \Data_Mem/n4554 ) );
  MUX U4609 ( .A(data_mem_out_wire[1713]), .B(reg_target[17]), .S(n1910), .Z(
        \Data_Mem/n4553 ) );
  MUX U4610 ( .A(data_mem_out_wire[1712]), .B(reg_target[16]), .S(n1910), .Z(
        \Data_Mem/n4552 ) );
  MUX U4611 ( .A(data_mem_out_wire[1711]), .B(reg_target[15]), .S(n1910), .Z(
        \Data_Mem/n4551 ) );
  MUX U4612 ( .A(data_mem_out_wire[1710]), .B(reg_target[14]), .S(n1910), .Z(
        \Data_Mem/n4550 ) );
  MUX U4613 ( .A(data_mem_out_wire[1709]), .B(reg_target[13]), .S(n1910), .Z(
        \Data_Mem/n4549 ) );
  MUX U4614 ( .A(data_mem_out_wire[1708]), .B(reg_target[12]), .S(n1910), .Z(
        \Data_Mem/n4548 ) );
  MUX U4615 ( .A(data_mem_out_wire[1707]), .B(reg_target[11]), .S(n1910), .Z(
        \Data_Mem/n4547 ) );
  MUX U4616 ( .A(data_mem_out_wire[1706]), .B(reg_target[10]), .S(n1910), .Z(
        \Data_Mem/n4546 ) );
  MUX U4617 ( .A(data_mem_out_wire[1705]), .B(reg_target[9]), .S(n1910), .Z(
        \Data_Mem/n4545 ) );
  MUX U4618 ( .A(data_mem_out_wire[1704]), .B(reg_target[8]), .S(n1910), .Z(
        \Data_Mem/n4544 ) );
  MUX U4619 ( .A(data_mem_out_wire[1703]), .B(reg_target[7]), .S(n1910), .Z(
        \Data_Mem/n4543 ) );
  MUX U4620 ( .A(data_mem_out_wire[1702]), .B(reg_target[6]), .S(n1910), .Z(
        \Data_Mem/n4542 ) );
  MUX U4621 ( .A(data_mem_out_wire[1701]), .B(reg_target[5]), .S(n1910), .Z(
        \Data_Mem/n4541 ) );
  MUX U4622 ( .A(data_mem_out_wire[1700]), .B(reg_target[4]), .S(n1910), .Z(
        \Data_Mem/n4540 ) );
  MUX U4623 ( .A(data_mem_out_wire[1699]), .B(reg_target[3]), .S(n1910), .Z(
        \Data_Mem/n4539 ) );
  MUX U4624 ( .A(data_mem_out_wire[1698]), .B(reg_target[2]), .S(n1910), .Z(
        \Data_Mem/n4538 ) );
  MUX U4625 ( .A(data_mem_out_wire[1697]), .B(reg_target[1]), .S(n1910), .Z(
        \Data_Mem/n4537 ) );
  MUX U4626 ( .A(data_mem_out_wire[1696]), .B(reg_target[0]), .S(n1910), .Z(
        \Data_Mem/n4536 ) );
  ANDN U4627 ( .B(n1807), .A(n1899), .Z(n1910) );
  ANDN U4628 ( .B(n1911), .A(n1901), .Z(n1807) );
  MUX U4629 ( .A(data_mem_out_wire[1759]), .B(reg_target[31]), .S(n1912), .Z(
        \Data_Mem/n4535 ) );
  MUX U4630 ( .A(data_mem_out_wire[1758]), .B(reg_target[30]), .S(n1912), .Z(
        \Data_Mem/n4534 ) );
  MUX U4631 ( .A(data_mem_out_wire[1757]), .B(reg_target[29]), .S(n1912), .Z(
        \Data_Mem/n4533 ) );
  MUX U4632 ( .A(data_mem_out_wire[1756]), .B(reg_target[28]), .S(n1912), .Z(
        \Data_Mem/n4532 ) );
  MUX U4633 ( .A(data_mem_out_wire[1755]), .B(reg_target[27]), .S(n1912), .Z(
        \Data_Mem/n4531 ) );
  MUX U4634 ( .A(data_mem_out_wire[1754]), .B(reg_target[26]), .S(n1912), .Z(
        \Data_Mem/n4530 ) );
  MUX U4635 ( .A(data_mem_out_wire[1753]), .B(reg_target[25]), .S(n1912), .Z(
        \Data_Mem/n4529 ) );
  MUX U4636 ( .A(data_mem_out_wire[1752]), .B(reg_target[24]), .S(n1912), .Z(
        \Data_Mem/n4528 ) );
  MUX U4637 ( .A(data_mem_out_wire[1751]), .B(reg_target[23]), .S(n1912), .Z(
        \Data_Mem/n4527 ) );
  MUX U4638 ( .A(data_mem_out_wire[1750]), .B(reg_target[22]), .S(n1912), .Z(
        \Data_Mem/n4526 ) );
  MUX U4639 ( .A(data_mem_out_wire[1749]), .B(reg_target[21]), .S(n1912), .Z(
        \Data_Mem/n4525 ) );
  MUX U4640 ( .A(data_mem_out_wire[1748]), .B(reg_target[20]), .S(n1912), .Z(
        \Data_Mem/n4524 ) );
  MUX U4641 ( .A(data_mem_out_wire[1747]), .B(reg_target[19]), .S(n1912), .Z(
        \Data_Mem/n4523 ) );
  MUX U4642 ( .A(data_mem_out_wire[1746]), .B(reg_target[18]), .S(n1912), .Z(
        \Data_Mem/n4522 ) );
  MUX U4643 ( .A(data_mem_out_wire[1745]), .B(reg_target[17]), .S(n1912), .Z(
        \Data_Mem/n4521 ) );
  MUX U4644 ( .A(data_mem_out_wire[1744]), .B(reg_target[16]), .S(n1912), .Z(
        \Data_Mem/n4520 ) );
  MUX U4645 ( .A(data_mem_out_wire[1743]), .B(reg_target[15]), .S(n1912), .Z(
        \Data_Mem/n4519 ) );
  MUX U4646 ( .A(data_mem_out_wire[1742]), .B(reg_target[14]), .S(n1912), .Z(
        \Data_Mem/n4518 ) );
  MUX U4647 ( .A(data_mem_out_wire[1741]), .B(reg_target[13]), .S(n1912), .Z(
        \Data_Mem/n4517 ) );
  MUX U4648 ( .A(data_mem_out_wire[1740]), .B(reg_target[12]), .S(n1912), .Z(
        \Data_Mem/n4516 ) );
  MUX U4649 ( .A(data_mem_out_wire[1739]), .B(reg_target[11]), .S(n1912), .Z(
        \Data_Mem/n4515 ) );
  MUX U4650 ( .A(data_mem_out_wire[1738]), .B(reg_target[10]), .S(n1912), .Z(
        \Data_Mem/n4514 ) );
  MUX U4651 ( .A(data_mem_out_wire[1737]), .B(reg_target[9]), .S(n1912), .Z(
        \Data_Mem/n4513 ) );
  MUX U4652 ( .A(data_mem_out_wire[1736]), .B(reg_target[8]), .S(n1912), .Z(
        \Data_Mem/n4512 ) );
  MUX U4653 ( .A(data_mem_out_wire[1735]), .B(reg_target[7]), .S(n1912), .Z(
        \Data_Mem/n4511 ) );
  MUX U4654 ( .A(data_mem_out_wire[1734]), .B(reg_target[6]), .S(n1912), .Z(
        \Data_Mem/n4510 ) );
  MUX U4655 ( .A(data_mem_out_wire[1733]), .B(reg_target[5]), .S(n1912), .Z(
        \Data_Mem/n4509 ) );
  MUX U4656 ( .A(data_mem_out_wire[1732]), .B(reg_target[4]), .S(n1912), .Z(
        \Data_Mem/n4508 ) );
  MUX U4657 ( .A(data_mem_out_wire[1731]), .B(reg_target[3]), .S(n1912), .Z(
        \Data_Mem/n4507 ) );
  MUX U4658 ( .A(data_mem_out_wire[1730]), .B(reg_target[2]), .S(n1912), .Z(
        \Data_Mem/n4506 ) );
  MUX U4659 ( .A(data_mem_out_wire[1729]), .B(reg_target[1]), .S(n1912), .Z(
        \Data_Mem/n4505 ) );
  MUX U4660 ( .A(data_mem_out_wire[1728]), .B(reg_target[0]), .S(n1912), .Z(
        \Data_Mem/n4504 ) );
  ANDN U4661 ( .B(n1810), .A(n1899), .Z(n1912) );
  ANDN U4662 ( .B(n1913), .A(n1901), .Z(n1810) );
  MUX U4663 ( .A(data_mem_out_wire[1791]), .B(reg_target[31]), .S(n1914), .Z(
        \Data_Mem/n4503 ) );
  MUX U4664 ( .A(data_mem_out_wire[1790]), .B(reg_target[30]), .S(n1914), .Z(
        \Data_Mem/n4502 ) );
  MUX U4665 ( .A(data_mem_out_wire[1789]), .B(reg_target[29]), .S(n1914), .Z(
        \Data_Mem/n4501 ) );
  MUX U4666 ( .A(data_mem_out_wire[1788]), .B(reg_target[28]), .S(n1914), .Z(
        \Data_Mem/n4500 ) );
  MUX U4667 ( .A(data_mem_out_wire[1787]), .B(reg_target[27]), .S(n1914), .Z(
        \Data_Mem/n4499 ) );
  MUX U4668 ( .A(data_mem_out_wire[1786]), .B(reg_target[26]), .S(n1914), .Z(
        \Data_Mem/n4498 ) );
  MUX U4669 ( .A(data_mem_out_wire[1785]), .B(reg_target[25]), .S(n1914), .Z(
        \Data_Mem/n4497 ) );
  MUX U4670 ( .A(data_mem_out_wire[1784]), .B(reg_target[24]), .S(n1914), .Z(
        \Data_Mem/n4496 ) );
  MUX U4671 ( .A(data_mem_out_wire[1783]), .B(reg_target[23]), .S(n1914), .Z(
        \Data_Mem/n4495 ) );
  MUX U4672 ( .A(data_mem_out_wire[1782]), .B(reg_target[22]), .S(n1914), .Z(
        \Data_Mem/n4494 ) );
  MUX U4673 ( .A(data_mem_out_wire[1781]), .B(reg_target[21]), .S(n1914), .Z(
        \Data_Mem/n4493 ) );
  MUX U4674 ( .A(data_mem_out_wire[1780]), .B(reg_target[20]), .S(n1914), .Z(
        \Data_Mem/n4492 ) );
  MUX U4675 ( .A(data_mem_out_wire[1779]), .B(reg_target[19]), .S(n1914), .Z(
        \Data_Mem/n4491 ) );
  MUX U4676 ( .A(data_mem_out_wire[1778]), .B(reg_target[18]), .S(n1914), .Z(
        \Data_Mem/n4490 ) );
  MUX U4677 ( .A(data_mem_out_wire[1777]), .B(reg_target[17]), .S(n1914), .Z(
        \Data_Mem/n4489 ) );
  MUX U4678 ( .A(data_mem_out_wire[1776]), .B(reg_target[16]), .S(n1914), .Z(
        \Data_Mem/n4488 ) );
  MUX U4679 ( .A(data_mem_out_wire[1775]), .B(reg_target[15]), .S(n1914), .Z(
        \Data_Mem/n4487 ) );
  MUX U4680 ( .A(data_mem_out_wire[1774]), .B(reg_target[14]), .S(n1914), .Z(
        \Data_Mem/n4486 ) );
  MUX U4681 ( .A(data_mem_out_wire[1773]), .B(reg_target[13]), .S(n1914), .Z(
        \Data_Mem/n4485 ) );
  MUX U4682 ( .A(data_mem_out_wire[1772]), .B(reg_target[12]), .S(n1914), .Z(
        \Data_Mem/n4484 ) );
  MUX U4683 ( .A(data_mem_out_wire[1771]), .B(reg_target[11]), .S(n1914), .Z(
        \Data_Mem/n4483 ) );
  MUX U4684 ( .A(data_mem_out_wire[1770]), .B(reg_target[10]), .S(n1914), .Z(
        \Data_Mem/n4482 ) );
  MUX U4685 ( .A(data_mem_out_wire[1769]), .B(reg_target[9]), .S(n1914), .Z(
        \Data_Mem/n4481 ) );
  MUX U4686 ( .A(data_mem_out_wire[1768]), .B(reg_target[8]), .S(n1914), .Z(
        \Data_Mem/n4480 ) );
  MUX U4687 ( .A(data_mem_out_wire[1767]), .B(reg_target[7]), .S(n1914), .Z(
        \Data_Mem/n4479 ) );
  MUX U4688 ( .A(data_mem_out_wire[1766]), .B(reg_target[6]), .S(n1914), .Z(
        \Data_Mem/n4478 ) );
  MUX U4689 ( .A(data_mem_out_wire[1765]), .B(reg_target[5]), .S(n1914), .Z(
        \Data_Mem/n4477 ) );
  MUX U4690 ( .A(data_mem_out_wire[1764]), .B(reg_target[4]), .S(n1914), .Z(
        \Data_Mem/n4476 ) );
  MUX U4691 ( .A(data_mem_out_wire[1763]), .B(reg_target[3]), .S(n1914), .Z(
        \Data_Mem/n4475 ) );
  MUX U4692 ( .A(data_mem_out_wire[1762]), .B(reg_target[2]), .S(n1914), .Z(
        \Data_Mem/n4474 ) );
  MUX U4693 ( .A(data_mem_out_wire[1761]), .B(reg_target[1]), .S(n1914), .Z(
        \Data_Mem/n4473 ) );
  MUX U4694 ( .A(data_mem_out_wire[1760]), .B(reg_target[0]), .S(n1914), .Z(
        \Data_Mem/n4472 ) );
  NOR U4695 ( .A(n1812), .B(n1899), .Z(n1914) );
  NAND U4696 ( .A(N24), .B(n1848), .Z(n1899) );
  ANDN U4697 ( .B(n837), .A(n840), .Z(n1848) );
  IV U4698 ( .A(N25), .Z(n840) );
  IV U4699 ( .A(n1830), .Z(n1812) );
  ANDN U4700 ( .B(n1915), .A(n1901), .Z(n1830) );
  MUX U4701 ( .A(data_mem_out_wire[1823]), .B(reg_target[31]), .S(n1916), .Z(
        \Data_Mem/n4471 ) );
  MUX U4702 ( .A(data_mem_out_wire[1822]), .B(reg_target[30]), .S(n1916), .Z(
        \Data_Mem/n4470 ) );
  MUX U4703 ( .A(data_mem_out_wire[1821]), .B(reg_target[29]), .S(n1916), .Z(
        \Data_Mem/n4469 ) );
  MUX U4704 ( .A(data_mem_out_wire[1820]), .B(reg_target[28]), .S(n1916), .Z(
        \Data_Mem/n4468 ) );
  MUX U4705 ( .A(data_mem_out_wire[1819]), .B(reg_target[27]), .S(n1916), .Z(
        \Data_Mem/n4467 ) );
  MUX U4706 ( .A(data_mem_out_wire[1818]), .B(reg_target[26]), .S(n1916), .Z(
        \Data_Mem/n4466 ) );
  MUX U4707 ( .A(data_mem_out_wire[1817]), .B(reg_target[25]), .S(n1916), .Z(
        \Data_Mem/n4465 ) );
  MUX U4708 ( .A(data_mem_out_wire[1816]), .B(reg_target[24]), .S(n1916), .Z(
        \Data_Mem/n4464 ) );
  MUX U4709 ( .A(data_mem_out_wire[1815]), .B(reg_target[23]), .S(n1916), .Z(
        \Data_Mem/n4463 ) );
  MUX U4710 ( .A(data_mem_out_wire[1814]), .B(reg_target[22]), .S(n1916), .Z(
        \Data_Mem/n4462 ) );
  MUX U4711 ( .A(data_mem_out_wire[1813]), .B(reg_target[21]), .S(n1916), .Z(
        \Data_Mem/n4461 ) );
  MUX U4712 ( .A(data_mem_out_wire[1812]), .B(reg_target[20]), .S(n1916), .Z(
        \Data_Mem/n4460 ) );
  MUX U4713 ( .A(data_mem_out_wire[1811]), .B(reg_target[19]), .S(n1916), .Z(
        \Data_Mem/n4459 ) );
  MUX U4714 ( .A(data_mem_out_wire[1810]), .B(reg_target[18]), .S(n1916), .Z(
        \Data_Mem/n4458 ) );
  MUX U4715 ( .A(data_mem_out_wire[1809]), .B(reg_target[17]), .S(n1916), .Z(
        \Data_Mem/n4457 ) );
  MUX U4716 ( .A(data_mem_out_wire[1808]), .B(reg_target[16]), .S(n1916), .Z(
        \Data_Mem/n4456 ) );
  MUX U4717 ( .A(data_mem_out_wire[1807]), .B(reg_target[15]), .S(n1916), .Z(
        \Data_Mem/n4455 ) );
  MUX U4718 ( .A(data_mem_out_wire[1806]), .B(reg_target[14]), .S(n1916), .Z(
        \Data_Mem/n4454 ) );
  MUX U4719 ( .A(data_mem_out_wire[1805]), .B(reg_target[13]), .S(n1916), .Z(
        \Data_Mem/n4453 ) );
  MUX U4720 ( .A(data_mem_out_wire[1804]), .B(reg_target[12]), .S(n1916), .Z(
        \Data_Mem/n4452 ) );
  MUX U4721 ( .A(data_mem_out_wire[1803]), .B(reg_target[11]), .S(n1916), .Z(
        \Data_Mem/n4451 ) );
  MUX U4722 ( .A(data_mem_out_wire[1802]), .B(reg_target[10]), .S(n1916), .Z(
        \Data_Mem/n4450 ) );
  MUX U4723 ( .A(data_mem_out_wire[1801]), .B(reg_target[9]), .S(n1916), .Z(
        \Data_Mem/n4449 ) );
  MUX U4724 ( .A(data_mem_out_wire[1800]), .B(reg_target[8]), .S(n1916), .Z(
        \Data_Mem/n4448 ) );
  MUX U4725 ( .A(data_mem_out_wire[1799]), .B(reg_target[7]), .S(n1916), .Z(
        \Data_Mem/n4447 ) );
  MUX U4726 ( .A(data_mem_out_wire[1798]), .B(reg_target[6]), .S(n1916), .Z(
        \Data_Mem/n4446 ) );
  MUX U4727 ( .A(data_mem_out_wire[1797]), .B(reg_target[5]), .S(n1916), .Z(
        \Data_Mem/n4445 ) );
  MUX U4728 ( .A(data_mem_out_wire[1796]), .B(reg_target[4]), .S(n1916), .Z(
        \Data_Mem/n4444 ) );
  MUX U4729 ( .A(data_mem_out_wire[1795]), .B(reg_target[3]), .S(n1916), .Z(
        \Data_Mem/n4443 ) );
  MUX U4730 ( .A(data_mem_out_wire[1794]), .B(reg_target[2]), .S(n1916), .Z(
        \Data_Mem/n4442 ) );
  MUX U4731 ( .A(data_mem_out_wire[1793]), .B(reg_target[1]), .S(n1916), .Z(
        \Data_Mem/n4441 ) );
  MUX U4732 ( .A(data_mem_out_wire[1792]), .B(reg_target[0]), .S(n1916), .Z(
        \Data_Mem/n4440 ) );
  ANDN U4733 ( .B(n1900), .A(n1917), .Z(n1916) );
  ANDN U4734 ( .B(n1918), .A(N27), .Z(n1900) );
  MUX U4735 ( .A(data_mem_out_wire[1855]), .B(reg_target[31]), .S(n1919), .Z(
        \Data_Mem/n4439 ) );
  MUX U4736 ( .A(data_mem_out_wire[1854]), .B(reg_target[30]), .S(n1919), .Z(
        \Data_Mem/n4438 ) );
  MUX U4737 ( .A(data_mem_out_wire[1853]), .B(reg_target[29]), .S(n1919), .Z(
        \Data_Mem/n4437 ) );
  MUX U4738 ( .A(data_mem_out_wire[1852]), .B(reg_target[28]), .S(n1919), .Z(
        \Data_Mem/n4436 ) );
  MUX U4739 ( .A(data_mem_out_wire[1851]), .B(reg_target[27]), .S(n1919), .Z(
        \Data_Mem/n4435 ) );
  MUX U4740 ( .A(data_mem_out_wire[1850]), .B(reg_target[26]), .S(n1919), .Z(
        \Data_Mem/n4434 ) );
  MUX U4741 ( .A(data_mem_out_wire[1849]), .B(reg_target[25]), .S(n1919), .Z(
        \Data_Mem/n4433 ) );
  MUX U4742 ( .A(data_mem_out_wire[1848]), .B(reg_target[24]), .S(n1919), .Z(
        \Data_Mem/n4432 ) );
  MUX U4743 ( .A(data_mem_out_wire[1847]), .B(reg_target[23]), .S(n1919), .Z(
        \Data_Mem/n4431 ) );
  MUX U4744 ( .A(data_mem_out_wire[1846]), .B(reg_target[22]), .S(n1919), .Z(
        \Data_Mem/n4430 ) );
  MUX U4745 ( .A(data_mem_out_wire[1845]), .B(reg_target[21]), .S(n1919), .Z(
        \Data_Mem/n4429 ) );
  MUX U4746 ( .A(data_mem_out_wire[1844]), .B(reg_target[20]), .S(n1919), .Z(
        \Data_Mem/n4428 ) );
  MUX U4747 ( .A(data_mem_out_wire[1843]), .B(reg_target[19]), .S(n1919), .Z(
        \Data_Mem/n4427 ) );
  MUX U4748 ( .A(data_mem_out_wire[1842]), .B(reg_target[18]), .S(n1919), .Z(
        \Data_Mem/n4426 ) );
  MUX U4749 ( .A(data_mem_out_wire[1841]), .B(reg_target[17]), .S(n1919), .Z(
        \Data_Mem/n4425 ) );
  MUX U4750 ( .A(data_mem_out_wire[1840]), .B(reg_target[16]), .S(n1919), .Z(
        \Data_Mem/n4424 ) );
  MUX U4751 ( .A(data_mem_out_wire[1839]), .B(reg_target[15]), .S(n1919), .Z(
        \Data_Mem/n4423 ) );
  MUX U4752 ( .A(data_mem_out_wire[1838]), .B(reg_target[14]), .S(n1919), .Z(
        \Data_Mem/n4422 ) );
  MUX U4753 ( .A(data_mem_out_wire[1837]), .B(reg_target[13]), .S(n1919), .Z(
        \Data_Mem/n4421 ) );
  MUX U4754 ( .A(data_mem_out_wire[1836]), .B(reg_target[12]), .S(n1919), .Z(
        \Data_Mem/n4420 ) );
  MUX U4755 ( .A(data_mem_out_wire[1835]), .B(reg_target[11]), .S(n1919), .Z(
        \Data_Mem/n4419 ) );
  MUX U4756 ( .A(data_mem_out_wire[1834]), .B(reg_target[10]), .S(n1919), .Z(
        \Data_Mem/n4418 ) );
  MUX U4757 ( .A(data_mem_out_wire[1833]), .B(reg_target[9]), .S(n1919), .Z(
        \Data_Mem/n4417 ) );
  MUX U4758 ( .A(data_mem_out_wire[1832]), .B(reg_target[8]), .S(n1919), .Z(
        \Data_Mem/n4416 ) );
  MUX U4759 ( .A(data_mem_out_wire[1831]), .B(reg_target[7]), .S(n1919), .Z(
        \Data_Mem/n4415 ) );
  MUX U4760 ( .A(data_mem_out_wire[1830]), .B(reg_target[6]), .S(n1919), .Z(
        \Data_Mem/n4414 ) );
  MUX U4761 ( .A(data_mem_out_wire[1829]), .B(reg_target[5]), .S(n1919), .Z(
        \Data_Mem/n4413 ) );
  MUX U4762 ( .A(data_mem_out_wire[1828]), .B(reg_target[4]), .S(n1919), .Z(
        \Data_Mem/n4412 ) );
  MUX U4763 ( .A(data_mem_out_wire[1827]), .B(reg_target[3]), .S(n1919), .Z(
        \Data_Mem/n4411 ) );
  MUX U4764 ( .A(data_mem_out_wire[1826]), .B(reg_target[2]), .S(n1919), .Z(
        \Data_Mem/n4410 ) );
  MUX U4765 ( .A(data_mem_out_wire[1825]), .B(reg_target[1]), .S(n1919), .Z(
        \Data_Mem/n4409 ) );
  MUX U4766 ( .A(data_mem_out_wire[1824]), .B(reg_target[0]), .S(n1919), .Z(
        \Data_Mem/n4408 ) );
  ANDN U4767 ( .B(n1903), .A(n1917), .Z(n1919) );
  ANDN U4768 ( .B(n1920), .A(N27), .Z(n1903) );
  MUX U4769 ( .A(data_mem_out_wire[1887]), .B(reg_target[31]), .S(n1921), .Z(
        \Data_Mem/n4407 ) );
  MUX U4770 ( .A(data_mem_out_wire[1886]), .B(reg_target[30]), .S(n1921), .Z(
        \Data_Mem/n4406 ) );
  MUX U4771 ( .A(data_mem_out_wire[1885]), .B(reg_target[29]), .S(n1921), .Z(
        \Data_Mem/n4405 ) );
  MUX U4772 ( .A(data_mem_out_wire[1884]), .B(reg_target[28]), .S(n1921), .Z(
        \Data_Mem/n4404 ) );
  MUX U4773 ( .A(data_mem_out_wire[1883]), .B(reg_target[27]), .S(n1921), .Z(
        \Data_Mem/n4403 ) );
  MUX U4774 ( .A(data_mem_out_wire[1882]), .B(reg_target[26]), .S(n1921), .Z(
        \Data_Mem/n4402 ) );
  MUX U4775 ( .A(data_mem_out_wire[1881]), .B(reg_target[25]), .S(n1921), .Z(
        \Data_Mem/n4401 ) );
  MUX U4776 ( .A(data_mem_out_wire[1880]), .B(reg_target[24]), .S(n1921), .Z(
        \Data_Mem/n4400 ) );
  MUX U4777 ( .A(data_mem_out_wire[1879]), .B(reg_target[23]), .S(n1921), .Z(
        \Data_Mem/n4399 ) );
  MUX U4778 ( .A(data_mem_out_wire[1878]), .B(reg_target[22]), .S(n1921), .Z(
        \Data_Mem/n4398 ) );
  MUX U4779 ( .A(data_mem_out_wire[1877]), .B(reg_target[21]), .S(n1921), .Z(
        \Data_Mem/n4397 ) );
  MUX U4780 ( .A(data_mem_out_wire[1876]), .B(reg_target[20]), .S(n1921), .Z(
        \Data_Mem/n4396 ) );
  MUX U4781 ( .A(data_mem_out_wire[1875]), .B(reg_target[19]), .S(n1921), .Z(
        \Data_Mem/n4395 ) );
  MUX U4782 ( .A(data_mem_out_wire[1874]), .B(reg_target[18]), .S(n1921), .Z(
        \Data_Mem/n4394 ) );
  MUX U4783 ( .A(data_mem_out_wire[1873]), .B(reg_target[17]), .S(n1921), .Z(
        \Data_Mem/n4393 ) );
  MUX U4784 ( .A(data_mem_out_wire[1872]), .B(reg_target[16]), .S(n1921), .Z(
        \Data_Mem/n4392 ) );
  MUX U4785 ( .A(data_mem_out_wire[1871]), .B(reg_target[15]), .S(n1921), .Z(
        \Data_Mem/n4391 ) );
  MUX U4786 ( .A(data_mem_out_wire[1870]), .B(reg_target[14]), .S(n1921), .Z(
        \Data_Mem/n4390 ) );
  MUX U4787 ( .A(data_mem_out_wire[1869]), .B(reg_target[13]), .S(n1921), .Z(
        \Data_Mem/n4389 ) );
  MUX U4788 ( .A(data_mem_out_wire[1868]), .B(reg_target[12]), .S(n1921), .Z(
        \Data_Mem/n4388 ) );
  MUX U4789 ( .A(data_mem_out_wire[1867]), .B(reg_target[11]), .S(n1921), .Z(
        \Data_Mem/n4387 ) );
  MUX U4790 ( .A(data_mem_out_wire[1866]), .B(reg_target[10]), .S(n1921), .Z(
        \Data_Mem/n4386 ) );
  MUX U4791 ( .A(data_mem_out_wire[1865]), .B(reg_target[9]), .S(n1921), .Z(
        \Data_Mem/n4385 ) );
  MUX U4792 ( .A(data_mem_out_wire[1864]), .B(reg_target[8]), .S(n1921), .Z(
        \Data_Mem/n4384 ) );
  MUX U4793 ( .A(data_mem_out_wire[1863]), .B(reg_target[7]), .S(n1921), .Z(
        \Data_Mem/n4383 ) );
  MUX U4794 ( .A(data_mem_out_wire[1862]), .B(reg_target[6]), .S(n1921), .Z(
        \Data_Mem/n4382 ) );
  MUX U4795 ( .A(data_mem_out_wire[1861]), .B(reg_target[5]), .S(n1921), .Z(
        \Data_Mem/n4381 ) );
  MUX U4796 ( .A(data_mem_out_wire[1860]), .B(reg_target[4]), .S(n1921), .Z(
        \Data_Mem/n4380 ) );
  MUX U4797 ( .A(data_mem_out_wire[1859]), .B(reg_target[3]), .S(n1921), .Z(
        \Data_Mem/n4379 ) );
  MUX U4798 ( .A(data_mem_out_wire[1858]), .B(reg_target[2]), .S(n1921), .Z(
        \Data_Mem/n4378 ) );
  MUX U4799 ( .A(data_mem_out_wire[1857]), .B(reg_target[1]), .S(n1921), .Z(
        \Data_Mem/n4377 ) );
  MUX U4800 ( .A(data_mem_out_wire[1856]), .B(reg_target[0]), .S(n1921), .Z(
        \Data_Mem/n4376 ) );
  ANDN U4801 ( .B(n1905), .A(n1917), .Z(n1921) );
  ANDN U4802 ( .B(n1922), .A(N27), .Z(n1905) );
  MUX U4803 ( .A(data_mem_out_wire[1919]), .B(reg_target[31]), .S(n1923), .Z(
        \Data_Mem/n4375 ) );
  MUX U4804 ( .A(data_mem_out_wire[1918]), .B(reg_target[30]), .S(n1923), .Z(
        \Data_Mem/n4374 ) );
  MUX U4805 ( .A(data_mem_out_wire[1917]), .B(reg_target[29]), .S(n1923), .Z(
        \Data_Mem/n4373 ) );
  MUX U4806 ( .A(data_mem_out_wire[1916]), .B(reg_target[28]), .S(n1923), .Z(
        \Data_Mem/n4372 ) );
  MUX U4807 ( .A(data_mem_out_wire[1915]), .B(reg_target[27]), .S(n1923), .Z(
        \Data_Mem/n4371 ) );
  MUX U4808 ( .A(data_mem_out_wire[1914]), .B(reg_target[26]), .S(n1923), .Z(
        \Data_Mem/n4370 ) );
  MUX U4809 ( .A(data_mem_out_wire[1913]), .B(reg_target[25]), .S(n1923), .Z(
        \Data_Mem/n4369 ) );
  MUX U4810 ( .A(data_mem_out_wire[1912]), .B(reg_target[24]), .S(n1923), .Z(
        \Data_Mem/n4368 ) );
  MUX U4811 ( .A(data_mem_out_wire[1911]), .B(reg_target[23]), .S(n1923), .Z(
        \Data_Mem/n4367 ) );
  MUX U4812 ( .A(data_mem_out_wire[1910]), .B(reg_target[22]), .S(n1923), .Z(
        \Data_Mem/n4366 ) );
  MUX U4813 ( .A(data_mem_out_wire[1909]), .B(reg_target[21]), .S(n1923), .Z(
        \Data_Mem/n4365 ) );
  MUX U4814 ( .A(data_mem_out_wire[1908]), .B(reg_target[20]), .S(n1923), .Z(
        \Data_Mem/n4364 ) );
  MUX U4815 ( .A(data_mem_out_wire[1907]), .B(reg_target[19]), .S(n1923), .Z(
        \Data_Mem/n4363 ) );
  MUX U4816 ( .A(data_mem_out_wire[1906]), .B(reg_target[18]), .S(n1923), .Z(
        \Data_Mem/n4362 ) );
  MUX U4817 ( .A(data_mem_out_wire[1905]), .B(reg_target[17]), .S(n1923), .Z(
        \Data_Mem/n4361 ) );
  MUX U4818 ( .A(data_mem_out_wire[1904]), .B(reg_target[16]), .S(n1923), .Z(
        \Data_Mem/n4360 ) );
  MUX U4819 ( .A(data_mem_out_wire[1903]), .B(reg_target[15]), .S(n1923), .Z(
        \Data_Mem/n4359 ) );
  MUX U4820 ( .A(data_mem_out_wire[1902]), .B(reg_target[14]), .S(n1923), .Z(
        \Data_Mem/n4358 ) );
  MUX U4821 ( .A(data_mem_out_wire[1901]), .B(reg_target[13]), .S(n1923), .Z(
        \Data_Mem/n4357 ) );
  MUX U4822 ( .A(data_mem_out_wire[1900]), .B(reg_target[12]), .S(n1923), .Z(
        \Data_Mem/n4356 ) );
  MUX U4823 ( .A(data_mem_out_wire[1899]), .B(reg_target[11]), .S(n1923), .Z(
        \Data_Mem/n4355 ) );
  MUX U4824 ( .A(data_mem_out_wire[1898]), .B(reg_target[10]), .S(n1923), .Z(
        \Data_Mem/n4354 ) );
  MUX U4825 ( .A(data_mem_out_wire[1897]), .B(reg_target[9]), .S(n1923), .Z(
        \Data_Mem/n4353 ) );
  MUX U4826 ( .A(data_mem_out_wire[1896]), .B(reg_target[8]), .S(n1923), .Z(
        \Data_Mem/n4352 ) );
  MUX U4827 ( .A(data_mem_out_wire[1895]), .B(reg_target[7]), .S(n1923), .Z(
        \Data_Mem/n4351 ) );
  MUX U4828 ( .A(data_mem_out_wire[1894]), .B(reg_target[6]), .S(n1923), .Z(
        \Data_Mem/n4350 ) );
  MUX U4829 ( .A(data_mem_out_wire[1893]), .B(reg_target[5]), .S(n1923), .Z(
        \Data_Mem/n4349 ) );
  MUX U4830 ( .A(data_mem_out_wire[1892]), .B(reg_target[4]), .S(n1923), .Z(
        \Data_Mem/n4348 ) );
  MUX U4831 ( .A(data_mem_out_wire[1891]), .B(reg_target[3]), .S(n1923), .Z(
        \Data_Mem/n4347 ) );
  MUX U4832 ( .A(data_mem_out_wire[1890]), .B(reg_target[2]), .S(n1923), .Z(
        \Data_Mem/n4346 ) );
  MUX U4833 ( .A(data_mem_out_wire[1889]), .B(reg_target[1]), .S(n1923), .Z(
        \Data_Mem/n4345 ) );
  MUX U4834 ( .A(data_mem_out_wire[1888]), .B(reg_target[0]), .S(n1923), .Z(
        \Data_Mem/n4344 ) );
  ANDN U4835 ( .B(n1907), .A(n1917), .Z(n1923) );
  ANDN U4836 ( .B(n1924), .A(N27), .Z(n1907) );
  MUX U4837 ( .A(data_mem_out_wire[1951]), .B(reg_target[31]), .S(n1925), .Z(
        \Data_Mem/n4343 ) );
  MUX U4838 ( .A(data_mem_out_wire[1950]), .B(reg_target[30]), .S(n1925), .Z(
        \Data_Mem/n4342 ) );
  MUX U4839 ( .A(data_mem_out_wire[1949]), .B(reg_target[29]), .S(n1925), .Z(
        \Data_Mem/n4341 ) );
  MUX U4840 ( .A(data_mem_out_wire[1948]), .B(reg_target[28]), .S(n1925), .Z(
        \Data_Mem/n4340 ) );
  MUX U4841 ( .A(data_mem_out_wire[1947]), .B(reg_target[27]), .S(n1925), .Z(
        \Data_Mem/n4339 ) );
  MUX U4842 ( .A(data_mem_out_wire[1946]), .B(reg_target[26]), .S(n1925), .Z(
        \Data_Mem/n4338 ) );
  MUX U4843 ( .A(data_mem_out_wire[1945]), .B(reg_target[25]), .S(n1925), .Z(
        \Data_Mem/n4337 ) );
  MUX U4844 ( .A(data_mem_out_wire[1944]), .B(reg_target[24]), .S(n1925), .Z(
        \Data_Mem/n4336 ) );
  MUX U4845 ( .A(data_mem_out_wire[1943]), .B(reg_target[23]), .S(n1925), .Z(
        \Data_Mem/n4335 ) );
  MUX U4846 ( .A(data_mem_out_wire[1942]), .B(reg_target[22]), .S(n1925), .Z(
        \Data_Mem/n4334 ) );
  MUX U4847 ( .A(data_mem_out_wire[1941]), .B(reg_target[21]), .S(n1925), .Z(
        \Data_Mem/n4333 ) );
  MUX U4848 ( .A(data_mem_out_wire[1940]), .B(reg_target[20]), .S(n1925), .Z(
        \Data_Mem/n4332 ) );
  MUX U4849 ( .A(data_mem_out_wire[1939]), .B(reg_target[19]), .S(n1925), .Z(
        \Data_Mem/n4331 ) );
  MUX U4850 ( .A(data_mem_out_wire[1938]), .B(reg_target[18]), .S(n1925), .Z(
        \Data_Mem/n4330 ) );
  MUX U4851 ( .A(data_mem_out_wire[1937]), .B(reg_target[17]), .S(n1925), .Z(
        \Data_Mem/n4329 ) );
  MUX U4852 ( .A(data_mem_out_wire[1936]), .B(reg_target[16]), .S(n1925), .Z(
        \Data_Mem/n4328 ) );
  MUX U4853 ( .A(data_mem_out_wire[1935]), .B(reg_target[15]), .S(n1925), .Z(
        \Data_Mem/n4327 ) );
  MUX U4854 ( .A(data_mem_out_wire[1934]), .B(reg_target[14]), .S(n1925), .Z(
        \Data_Mem/n4326 ) );
  MUX U4855 ( .A(data_mem_out_wire[1933]), .B(reg_target[13]), .S(n1925), .Z(
        \Data_Mem/n4325 ) );
  MUX U4856 ( .A(data_mem_out_wire[1932]), .B(reg_target[12]), .S(n1925), .Z(
        \Data_Mem/n4324 ) );
  MUX U4857 ( .A(data_mem_out_wire[1931]), .B(reg_target[11]), .S(n1925), .Z(
        \Data_Mem/n4323 ) );
  MUX U4858 ( .A(data_mem_out_wire[1930]), .B(reg_target[10]), .S(n1925), .Z(
        \Data_Mem/n4322 ) );
  MUX U4859 ( .A(data_mem_out_wire[1929]), .B(reg_target[9]), .S(n1925), .Z(
        \Data_Mem/n4321 ) );
  MUX U4860 ( .A(data_mem_out_wire[1928]), .B(reg_target[8]), .S(n1925), .Z(
        \Data_Mem/n4320 ) );
  MUX U4861 ( .A(data_mem_out_wire[1927]), .B(reg_target[7]), .S(n1925), .Z(
        \Data_Mem/n4319 ) );
  MUX U4862 ( .A(data_mem_out_wire[1926]), .B(reg_target[6]), .S(n1925), .Z(
        \Data_Mem/n4318 ) );
  MUX U4863 ( .A(data_mem_out_wire[1925]), .B(reg_target[5]), .S(n1925), .Z(
        \Data_Mem/n4317 ) );
  MUX U4864 ( .A(data_mem_out_wire[1924]), .B(reg_target[4]), .S(n1925), .Z(
        \Data_Mem/n4316 ) );
  MUX U4865 ( .A(data_mem_out_wire[1923]), .B(reg_target[3]), .S(n1925), .Z(
        \Data_Mem/n4315 ) );
  MUX U4866 ( .A(data_mem_out_wire[1922]), .B(reg_target[2]), .S(n1925), .Z(
        \Data_Mem/n4314 ) );
  MUX U4867 ( .A(data_mem_out_wire[1921]), .B(reg_target[1]), .S(n1925), .Z(
        \Data_Mem/n4313 ) );
  MUX U4868 ( .A(data_mem_out_wire[1920]), .B(reg_target[0]), .S(n1925), .Z(
        \Data_Mem/n4312 ) );
  ANDN U4869 ( .B(n1909), .A(n1917), .Z(n1925) );
  AND U4870 ( .A(n1918), .B(N27), .Z(n1909) );
  ANDN U4871 ( .B(n834), .A(N28), .Z(n1918) );
  MUX U4872 ( .A(data_mem_out_wire[1983]), .B(reg_target[31]), .S(n1926), .Z(
        \Data_Mem/n4311 ) );
  MUX U4873 ( .A(data_mem_out_wire[1982]), .B(reg_target[30]), .S(n1926), .Z(
        \Data_Mem/n4310 ) );
  MUX U4874 ( .A(data_mem_out_wire[1981]), .B(reg_target[29]), .S(n1926), .Z(
        \Data_Mem/n4309 ) );
  MUX U4875 ( .A(data_mem_out_wire[1980]), .B(reg_target[28]), .S(n1926), .Z(
        \Data_Mem/n4308 ) );
  MUX U4876 ( .A(data_mem_out_wire[1979]), .B(reg_target[27]), .S(n1926), .Z(
        \Data_Mem/n4307 ) );
  MUX U4877 ( .A(data_mem_out_wire[1978]), .B(reg_target[26]), .S(n1926), .Z(
        \Data_Mem/n4306 ) );
  MUX U4878 ( .A(data_mem_out_wire[1977]), .B(reg_target[25]), .S(n1926), .Z(
        \Data_Mem/n4305 ) );
  MUX U4879 ( .A(data_mem_out_wire[1976]), .B(reg_target[24]), .S(n1926), .Z(
        \Data_Mem/n4304 ) );
  MUX U4880 ( .A(data_mem_out_wire[1975]), .B(reg_target[23]), .S(n1926), .Z(
        \Data_Mem/n4303 ) );
  MUX U4881 ( .A(data_mem_out_wire[1974]), .B(reg_target[22]), .S(n1926), .Z(
        \Data_Mem/n4302 ) );
  MUX U4882 ( .A(data_mem_out_wire[1973]), .B(reg_target[21]), .S(n1926), .Z(
        \Data_Mem/n4301 ) );
  MUX U4883 ( .A(data_mem_out_wire[1972]), .B(reg_target[20]), .S(n1926), .Z(
        \Data_Mem/n4300 ) );
  MUX U4884 ( .A(data_mem_out_wire[1971]), .B(reg_target[19]), .S(n1926), .Z(
        \Data_Mem/n4299 ) );
  MUX U4885 ( .A(data_mem_out_wire[1970]), .B(reg_target[18]), .S(n1926), .Z(
        \Data_Mem/n4298 ) );
  MUX U4886 ( .A(data_mem_out_wire[1969]), .B(reg_target[17]), .S(n1926), .Z(
        \Data_Mem/n4297 ) );
  MUX U4887 ( .A(data_mem_out_wire[1968]), .B(reg_target[16]), .S(n1926), .Z(
        \Data_Mem/n4296 ) );
  MUX U4888 ( .A(data_mem_out_wire[1967]), .B(reg_target[15]), .S(n1926), .Z(
        \Data_Mem/n4295 ) );
  MUX U4889 ( .A(data_mem_out_wire[1966]), .B(reg_target[14]), .S(n1926), .Z(
        \Data_Mem/n4294 ) );
  MUX U4890 ( .A(data_mem_out_wire[1965]), .B(reg_target[13]), .S(n1926), .Z(
        \Data_Mem/n4293 ) );
  MUX U4891 ( .A(data_mem_out_wire[1964]), .B(reg_target[12]), .S(n1926), .Z(
        \Data_Mem/n4292 ) );
  MUX U4892 ( .A(data_mem_out_wire[1963]), .B(reg_target[11]), .S(n1926), .Z(
        \Data_Mem/n4291 ) );
  MUX U4893 ( .A(data_mem_out_wire[1962]), .B(reg_target[10]), .S(n1926), .Z(
        \Data_Mem/n4290 ) );
  MUX U4894 ( .A(data_mem_out_wire[1961]), .B(reg_target[9]), .S(n1926), .Z(
        \Data_Mem/n4289 ) );
  MUX U4895 ( .A(data_mem_out_wire[1960]), .B(reg_target[8]), .S(n1926), .Z(
        \Data_Mem/n4288 ) );
  MUX U4896 ( .A(data_mem_out_wire[1959]), .B(reg_target[7]), .S(n1926), .Z(
        \Data_Mem/n4287 ) );
  MUX U4897 ( .A(data_mem_out_wire[1958]), .B(reg_target[6]), .S(n1926), .Z(
        \Data_Mem/n4286 ) );
  MUX U4898 ( .A(data_mem_out_wire[1957]), .B(reg_target[5]), .S(n1926), .Z(
        \Data_Mem/n4285 ) );
  MUX U4899 ( .A(data_mem_out_wire[1956]), .B(reg_target[4]), .S(n1926), .Z(
        \Data_Mem/n4284 ) );
  MUX U4900 ( .A(data_mem_out_wire[1955]), .B(reg_target[3]), .S(n1926), .Z(
        \Data_Mem/n4283 ) );
  MUX U4901 ( .A(data_mem_out_wire[1954]), .B(reg_target[2]), .S(n1926), .Z(
        \Data_Mem/n4282 ) );
  MUX U4902 ( .A(data_mem_out_wire[1953]), .B(reg_target[1]), .S(n1926), .Z(
        \Data_Mem/n4281 ) );
  MUX U4903 ( .A(data_mem_out_wire[1952]), .B(reg_target[0]), .S(n1926), .Z(
        \Data_Mem/n4280 ) );
  ANDN U4904 ( .B(n1911), .A(n1917), .Z(n1926) );
  AND U4905 ( .A(n1920), .B(N27), .Z(n1911) );
  ANDN U4906 ( .B(n835), .A(n834), .Z(n1920) );
  MUX U4907 ( .A(data_mem_out_wire[2015]), .B(reg_target[31]), .S(n1927), .Z(
        \Data_Mem/n4279 ) );
  MUX U4908 ( .A(data_mem_out_wire[2014]), .B(reg_target[30]), .S(n1927), .Z(
        \Data_Mem/n4278 ) );
  MUX U4909 ( .A(data_mem_out_wire[2013]), .B(reg_target[29]), .S(n1927), .Z(
        \Data_Mem/n4277 ) );
  MUX U4910 ( .A(data_mem_out_wire[2012]), .B(reg_target[28]), .S(n1927), .Z(
        \Data_Mem/n4276 ) );
  MUX U4911 ( .A(data_mem_out_wire[2011]), .B(reg_target[27]), .S(n1927), .Z(
        \Data_Mem/n4275 ) );
  MUX U4912 ( .A(data_mem_out_wire[2010]), .B(reg_target[26]), .S(n1927), .Z(
        \Data_Mem/n4274 ) );
  MUX U4913 ( .A(data_mem_out_wire[2009]), .B(reg_target[25]), .S(n1927), .Z(
        \Data_Mem/n4273 ) );
  MUX U4914 ( .A(data_mem_out_wire[2008]), .B(reg_target[24]), .S(n1927), .Z(
        \Data_Mem/n4272 ) );
  MUX U4915 ( .A(data_mem_out_wire[2007]), .B(reg_target[23]), .S(n1927), .Z(
        \Data_Mem/n4271 ) );
  MUX U4916 ( .A(data_mem_out_wire[2006]), .B(reg_target[22]), .S(n1927), .Z(
        \Data_Mem/n4270 ) );
  MUX U4917 ( .A(data_mem_out_wire[2005]), .B(reg_target[21]), .S(n1927), .Z(
        \Data_Mem/n4269 ) );
  MUX U4918 ( .A(data_mem_out_wire[2004]), .B(reg_target[20]), .S(n1927), .Z(
        \Data_Mem/n4268 ) );
  MUX U4919 ( .A(data_mem_out_wire[2003]), .B(reg_target[19]), .S(n1927), .Z(
        \Data_Mem/n4267 ) );
  MUX U4920 ( .A(data_mem_out_wire[2002]), .B(reg_target[18]), .S(n1927), .Z(
        \Data_Mem/n4266 ) );
  MUX U4921 ( .A(data_mem_out_wire[2001]), .B(reg_target[17]), .S(n1927), .Z(
        \Data_Mem/n4265 ) );
  MUX U4922 ( .A(data_mem_out_wire[2000]), .B(reg_target[16]), .S(n1927), .Z(
        \Data_Mem/n4264 ) );
  MUX U4923 ( .A(data_mem_out_wire[1999]), .B(reg_target[15]), .S(n1927), .Z(
        \Data_Mem/n4263 ) );
  MUX U4924 ( .A(data_mem_out_wire[1998]), .B(reg_target[14]), .S(n1927), .Z(
        \Data_Mem/n4262 ) );
  MUX U4925 ( .A(data_mem_out_wire[1997]), .B(reg_target[13]), .S(n1927), .Z(
        \Data_Mem/n4261 ) );
  MUX U4926 ( .A(data_mem_out_wire[1996]), .B(reg_target[12]), .S(n1927), .Z(
        \Data_Mem/n4260 ) );
  MUX U4927 ( .A(data_mem_out_wire[1995]), .B(reg_target[11]), .S(n1927), .Z(
        \Data_Mem/n4259 ) );
  MUX U4928 ( .A(data_mem_out_wire[1994]), .B(reg_target[10]), .S(n1927), .Z(
        \Data_Mem/n4258 ) );
  MUX U4929 ( .A(data_mem_out_wire[1993]), .B(reg_target[9]), .S(n1927), .Z(
        \Data_Mem/n4257 ) );
  MUX U4930 ( .A(data_mem_out_wire[1992]), .B(reg_target[8]), .S(n1927), .Z(
        \Data_Mem/n4256 ) );
  MUX U4931 ( .A(data_mem_out_wire[1991]), .B(reg_target[7]), .S(n1927), .Z(
        \Data_Mem/n4255 ) );
  MUX U4932 ( .A(data_mem_out_wire[1990]), .B(reg_target[6]), .S(n1927), .Z(
        \Data_Mem/n4254 ) );
  MUX U4933 ( .A(data_mem_out_wire[1989]), .B(reg_target[5]), .S(n1927), .Z(
        \Data_Mem/n4253 ) );
  MUX U4934 ( .A(data_mem_out_wire[1988]), .B(reg_target[4]), .S(n1927), .Z(
        \Data_Mem/n4252 ) );
  MUX U4935 ( .A(data_mem_out_wire[1987]), .B(reg_target[3]), .S(n1927), .Z(
        \Data_Mem/n4251 ) );
  MUX U4936 ( .A(data_mem_out_wire[1986]), .B(reg_target[2]), .S(n1927), .Z(
        \Data_Mem/n4250 ) );
  MUX U4937 ( .A(data_mem_out_wire[1985]), .B(reg_target[1]), .S(n1927), .Z(
        \Data_Mem/n4249 ) );
  MUX U4938 ( .A(data_mem_out_wire[1984]), .B(reg_target[0]), .S(n1927), .Z(
        \Data_Mem/n4248 ) );
  ANDN U4939 ( .B(n1913), .A(n1917), .Z(n1927) );
  AND U4940 ( .A(n1922), .B(N27), .Z(n1913) );
  ANDN U4941 ( .B(n834), .A(n835), .Z(n1922) );
  IV U4942 ( .A(N28), .Z(n835) );
  MUX U4943 ( .A(data_mem_out_wire[2047]), .B(reg_target[31]), .S(n1928), .Z(
        \Data_Mem/n4247 ) );
  MUX U4944 ( .A(data_mem_out_wire[2046]), .B(reg_target[30]), .S(n1928), .Z(
        \Data_Mem/n4246 ) );
  MUX U4945 ( .A(data_mem_out_wire[2045]), .B(reg_target[29]), .S(n1928), .Z(
        \Data_Mem/n4245 ) );
  MUX U4946 ( .A(data_mem_out_wire[2044]), .B(reg_target[28]), .S(n1928), .Z(
        \Data_Mem/n4244 ) );
  MUX U4947 ( .A(data_mem_out_wire[2043]), .B(reg_target[27]), .S(n1928), .Z(
        \Data_Mem/n4243 ) );
  MUX U4948 ( .A(data_mem_out_wire[2042]), .B(reg_target[26]), .S(n1928), .Z(
        \Data_Mem/n4242 ) );
  MUX U4949 ( .A(data_mem_out_wire[2041]), .B(reg_target[25]), .S(n1928), .Z(
        \Data_Mem/n4241 ) );
  MUX U4950 ( .A(data_mem_out_wire[2040]), .B(reg_target[24]), .S(n1928), .Z(
        \Data_Mem/n4240 ) );
  MUX U4951 ( .A(data_mem_out_wire[2039]), .B(reg_target[23]), .S(n1928), .Z(
        \Data_Mem/n4239 ) );
  MUX U4952 ( .A(data_mem_out_wire[2038]), .B(reg_target[22]), .S(n1928), .Z(
        \Data_Mem/n4238 ) );
  MUX U4953 ( .A(data_mem_out_wire[2037]), .B(reg_target[21]), .S(n1928), .Z(
        \Data_Mem/n4237 ) );
  MUX U4954 ( .A(data_mem_out_wire[2036]), .B(reg_target[20]), .S(n1928), .Z(
        \Data_Mem/n4236 ) );
  MUX U4955 ( .A(data_mem_out_wire[2035]), .B(reg_target[19]), .S(n1928), .Z(
        \Data_Mem/n4235 ) );
  MUX U4956 ( .A(data_mem_out_wire[2034]), .B(reg_target[18]), .S(n1928), .Z(
        \Data_Mem/n4234 ) );
  MUX U4957 ( .A(data_mem_out_wire[2033]), .B(reg_target[17]), .S(n1928), .Z(
        \Data_Mem/n4233 ) );
  MUX U4958 ( .A(data_mem_out_wire[2032]), .B(reg_target[16]), .S(n1928), .Z(
        \Data_Mem/n4232 ) );
  MUX U4959 ( .A(data_mem_out_wire[2031]), .B(reg_target[15]), .S(n1928), .Z(
        \Data_Mem/n4231 ) );
  MUX U4960 ( .A(data_mem_out_wire[2030]), .B(reg_target[14]), .S(n1928), .Z(
        \Data_Mem/n4230 ) );
  MUX U4961 ( .A(data_mem_out_wire[2029]), .B(reg_target[13]), .S(n1928), .Z(
        \Data_Mem/n4229 ) );
  MUX U4962 ( .A(data_mem_out_wire[2028]), .B(reg_target[12]), .S(n1928), .Z(
        \Data_Mem/n4228 ) );
  MUX U4963 ( .A(data_mem_out_wire[2027]), .B(reg_target[11]), .S(n1928), .Z(
        \Data_Mem/n4227 ) );
  MUX U4964 ( .A(data_mem_out_wire[2026]), .B(reg_target[10]), .S(n1928), .Z(
        \Data_Mem/n4226 ) );
  MUX U4965 ( .A(data_mem_out_wire[2025]), .B(reg_target[9]), .S(n1928), .Z(
        \Data_Mem/n4225 ) );
  MUX U4966 ( .A(data_mem_out_wire[2024]), .B(reg_target[8]), .S(n1928), .Z(
        \Data_Mem/n4224 ) );
  MUX U4967 ( .A(data_mem_out_wire[2023]), .B(reg_target[7]), .S(n1928), .Z(
        \Data_Mem/n4223 ) );
  MUX U4968 ( .A(data_mem_out_wire[2022]), .B(reg_target[6]), .S(n1928), .Z(
        \Data_Mem/n4222 ) );
  MUX U4969 ( .A(data_mem_out_wire[2021]), .B(reg_target[5]), .S(n1928), .Z(
        \Data_Mem/n4221 ) );
  MUX U4970 ( .A(data_mem_out_wire[2020]), .B(reg_target[4]), .S(n1928), .Z(
        \Data_Mem/n4220 ) );
  MUX U4971 ( .A(data_mem_out_wire[2019]), .B(reg_target[3]), .S(n1928), .Z(
        \Data_Mem/n4219 ) );
  MUX U4972 ( .A(data_mem_out_wire[2018]), .B(reg_target[2]), .S(n1928), .Z(
        \Data_Mem/n4218 ) );
  MUX U4973 ( .A(data_mem_out_wire[2017]), .B(reg_target[1]), .S(n1928), .Z(
        \Data_Mem/n4217 ) );
  MUX U4974 ( .A(data_mem_out_wire[2016]), .B(reg_target[0]), .S(n1928), .Z(
        \Data_Mem/n4216 ) );
  ANDN U4975 ( .B(n1915), .A(n1917), .Z(n1928) );
  NAND U4976 ( .A(n1929), .B(n1865), .Z(n1917) );
  ANDN U4977 ( .B(N25), .A(n837), .Z(n1865) );
  IV U4978 ( .A(N26), .Z(n837) );
  NAND U4979 ( .A(n1930), .B(n1931), .Z(N26) );
  AND U4980 ( .A(n1932), .B(n1933), .Z(n1931) );
  AND U4981 ( .A(n1934), .B(n1935), .Z(n1933) );
  NAND U4982 ( .A(n1936), .B(n852), .Z(n1935) );
  NAND U4983 ( .A(n1937), .B(n1938), .Z(n1936) );
  AND U4984 ( .A(n1939), .B(n1940), .Z(n1938) );
  AND U4985 ( .A(n1941), .B(n1942), .Z(n1939) );
  NANDN U4986 ( .A(n1505), .B(a_bus[4]), .Z(n1942) );
  AND U4987 ( .A(n1943), .B(n1944), .Z(n1505) );
  AND U4988 ( .A(n1945), .B(n1946), .Z(n1944) );
  NAND U4989 ( .A(n1092), .B(n1394), .Z(n1946) );
  AND U4990 ( .A(n1947), .B(n1948), .Z(n1943) );
  NAND U4991 ( .A(n1405), .B(n1398), .Z(n1947) );
  NAND U4992 ( .A(n1949), .B(n1950), .Z(n1398) );
  NAND U4993 ( .A(\Shifter/N75 ), .B(a_bus[1]), .Z(n1950) );
  AND U4994 ( .A(n1951), .B(n1952), .Z(n1949) );
  NANDN U4995 ( .A(n1051), .B(n863), .Z(n1941) );
  NAND U4996 ( .A(n1953), .B(n865), .Z(n1934) );
  NAND U4997 ( .A(n1937), .B(n1954), .Z(n1953) );
  AND U4998 ( .A(n1955), .B(n1940), .Z(n1954) );
  NAND U4999 ( .A(n888), .B(n1098), .Z(n1940) );
  NAND U5000 ( .A(n1956), .B(n1957), .Z(n1098) );
  AND U5001 ( .A(n1958), .B(n1959), .Z(n1957) );
  NANDN U5002 ( .A(n881), .B(b_bus[17]), .Z(n1959) );
  NANDN U5003 ( .A(n882), .B(b_bus[18]), .Z(n1958) );
  AND U5004 ( .A(n1960), .B(n1961), .Z(n1956) );
  NANDN U5005 ( .A(n885), .B(b_bus[20]), .Z(n1961) );
  NANDN U5006 ( .A(n886), .B(b_bus[19]), .Z(n1960) );
  AND U5007 ( .A(n1962), .B(n1963), .Z(n1955) );
  NANDN U5008 ( .A(n1507), .B(a_bus[4]), .Z(n1963) );
  AND U5009 ( .A(n1964), .B(n1965), .Z(n1507) );
  NAND U5010 ( .A(n1360), .B(n1092), .Z(n1965) );
  NAND U5011 ( .A(n1966), .B(n1967), .Z(n1092) );
  AND U5012 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U5013 ( .A(n881), .B(b_bus[21]), .Z(n1969) );
  NANDN U5014 ( .A(n882), .B(b_bus[22]), .Z(n1968) );
  AND U5015 ( .A(n1970), .B(n1971), .Z(n1966) );
  NANDN U5016 ( .A(n885), .B(b_bus[24]), .Z(n1971) );
  NANDN U5017 ( .A(n886), .B(b_bus[23]), .Z(n1970) );
  AND U5018 ( .A(n1972), .B(n1948), .Z(n1964) );
  NAND U5019 ( .A(n1252), .B(n1403), .Z(n1948) );
  NAND U5020 ( .A(n1973), .B(n1974), .Z(n1252) );
  AND U5021 ( .A(n1975), .B(n1976), .Z(n1974) );
  NANDN U5022 ( .A(n881), .B(b_bus[25]), .Z(n1976) );
  NANDN U5023 ( .A(n882), .B(b_bus[26]), .Z(n1975) );
  AND U5024 ( .A(n1977), .B(n1978), .Z(n1973) );
  NANDN U5025 ( .A(n885), .B(b_bus[28]), .Z(n1978) );
  NANDN U5026 ( .A(n886), .B(b_bus[27]), .Z(n1977) );
  NAND U5027 ( .A(n1251), .B(n1405), .Z(n1972) );
  NAND U5028 ( .A(n1979), .B(n1952), .Z(n1251) );
  NANDN U5029 ( .A(n881), .B(b_bus[29]), .Z(n1952) );
  AND U5030 ( .A(n1980), .B(n1951), .Z(n1979) );
  NANDN U5031 ( .A(n882), .B(b_bus[30]), .Z(n1951) );
  NANDN U5032 ( .A(n886), .B(\Shifter/N75 ), .Z(n1980) );
  NANDN U5033 ( .A(n1051), .B(n876), .Z(n1962) );
  AND U5034 ( .A(n1981), .B(n1982), .Z(n1051) );
  AND U5035 ( .A(n1983), .B(n1984), .Z(n1982) );
  NANDN U5036 ( .A(n881), .B(b_bus[5]), .Z(n1984) );
  NANDN U5037 ( .A(n882), .B(b_bus[6]), .Z(n1983) );
  AND U5038 ( .A(n1985), .B(n1986), .Z(n1981) );
  NANDN U5039 ( .A(n885), .B(b_bus[8]), .Z(n1986) );
  NANDN U5040 ( .A(n886), .B(b_bus[7]), .Z(n1985) );
  AND U5041 ( .A(n1987), .B(n1988), .Z(n1937) );
  NAND U5042 ( .A(n870), .B(n1059), .Z(n1988) );
  NAND U5043 ( .A(n1989), .B(n1990), .Z(n1059) );
  AND U5044 ( .A(n1991), .B(n1992), .Z(n1990) );
  NANDN U5045 ( .A(n881), .B(b_bus[13]), .Z(n1992) );
  NANDN U5046 ( .A(n882), .B(b_bus[14]), .Z(n1991) );
  AND U5047 ( .A(n1993), .B(n1994), .Z(n1989) );
  NANDN U5048 ( .A(n885), .B(b_bus[16]), .Z(n1994) );
  NANDN U5049 ( .A(n886), .B(b_bus[15]), .Z(n1993) );
  NAND U5050 ( .A(n874), .B(n1048), .Z(n1987) );
  NAND U5051 ( .A(n1995), .B(n1996), .Z(n1048) );
  AND U5052 ( .A(n1997), .B(n1998), .Z(n1996) );
  NANDN U5053 ( .A(n881), .B(b_bus[9]), .Z(n1998) );
  NANDN U5054 ( .A(n882), .B(b_bus[10]), .Z(n1997) );
  AND U5055 ( .A(n1999), .B(n2000), .Z(n1995) );
  NANDN U5056 ( .A(n885), .B(b_bus[12]), .Z(n2000) );
  NANDN U5057 ( .A(n886), .B(b_bus[11]), .Z(n1999) );
  AND U5058 ( .A(n2001), .B(n2002), .Z(n1932) );
  NAND U5059 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][5] ), .Z(n2002) );
  ANDN U5060 ( .B(\Shifter/sll_27/ML_int[3][5] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][5] ) );
  NAND U5061 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N113 ), .Z(n2001) );
  AND U5062 ( .A(n2003), .B(n2004), .Z(n1930) );
  AND U5063 ( .A(n2005), .B(n2006), .Z(n2004) );
  NANDN U5064 ( .A(n891), .B(\ALU/N113 ), .Z(n2006) );
  NAND U5065 ( .A(n2007), .B(n1026), .Z(n2005) );
  XNOR U5066 ( .A(n989), .B(n2485), .Z(n2007) );
  AND U5067 ( .A(n2008), .B(n2009), .Z(n2003) );
  NAND U5068 ( .A(n2010), .B(n2485), .Z(n2009) );
  AND U5069 ( .A(n897), .B(b_bus[5]), .Z(n2010) );
  MUX U5070 ( .A(n1022), .B(n1023), .S(n2011), .Z(n2008) );
  NOR U5071 ( .A(b_bus[5]), .B(n2485), .Z(n2011) );
  ANDN U5072 ( .B(reg_source[5]), .A(n1015), .Z(n2485) );
  NAND U5073 ( .A(n2012), .B(n2013), .Z(N25) );
  AND U5074 ( .A(n2014), .B(n2015), .Z(n2013) );
  AND U5075 ( .A(n2016), .B(n2017), .Z(n2015) );
  NAND U5076 ( .A(n2018), .B(n852), .Z(n2017) );
  NAND U5077 ( .A(n2019), .B(n2020), .Z(n2018) );
  AND U5078 ( .A(n2021), .B(n2022), .Z(n2020) );
  AND U5079 ( .A(n2023), .B(n2024), .Z(n2021) );
  NANDN U5080 ( .A(n1575), .B(a_bus[4]), .Z(n2024) );
  AND U5081 ( .A(n2025), .B(n2026), .Z(n1575) );
  AND U5082 ( .A(n2027), .B(n2028), .Z(n2026) );
  NAND U5083 ( .A(n1205), .B(n1394), .Z(n2028) );
  AND U5084 ( .A(n1945), .B(n2029), .Z(n2025) );
  NAND U5085 ( .A(n1683), .B(n1405), .Z(n2029) );
  NANDN U5086 ( .A(n2030), .B(n863), .Z(n2023) );
  NAND U5087 ( .A(n2031), .B(n865), .Z(n2016) );
  NAND U5088 ( .A(n2019), .B(n2032), .Z(n2031) );
  AND U5089 ( .A(n2033), .B(n2022), .Z(n2032) );
  NAND U5090 ( .A(n888), .B(n1211), .Z(n2022) );
  AND U5091 ( .A(n2034), .B(n2035), .Z(n2033) );
  NANDN U5092 ( .A(n1577), .B(a_bus[4]), .Z(n2035) );
  AND U5093 ( .A(n2036), .B(n2037), .Z(n1577) );
  NAND U5094 ( .A(n1360), .B(n1205), .Z(n2037) );
  AND U5095 ( .A(n2038), .B(n2027), .Z(n2036) );
  NAND U5096 ( .A(n1362), .B(n1403), .Z(n2027) );
  NAND U5097 ( .A(n1359), .B(n1405), .Z(n2038) );
  NANDN U5098 ( .A(n2030), .B(n876), .Z(n2034) );
  AND U5099 ( .A(n2039), .B(n2040), .Z(n2019) );
  NAND U5100 ( .A(n870), .B(n1212), .Z(n2040) );
  NAND U5101 ( .A(n874), .B(n1201), .Z(n2039) );
  AND U5102 ( .A(n2041), .B(n2042), .Z(n2014) );
  NAND U5103 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][6] ), .Z(n2042) );
  ANDN U5104 ( .B(\Shifter/sll_27/ML_int[3][6] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][6] ) );
  NAND U5105 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N114 ), .Z(n2041) );
  AND U5106 ( .A(n2043), .B(n2044), .Z(n2012) );
  AND U5107 ( .A(n2045), .B(n2046), .Z(n2044) );
  NANDN U5108 ( .A(n891), .B(\ALU/N114 ), .Z(n2046) );
  NAND U5109 ( .A(n2047), .B(n1026), .Z(n2045) );
  XNOR U5110 ( .A(n985), .B(n2484), .Z(n2047) );
  AND U5111 ( .A(n2048), .B(n2049), .Z(n2043) );
  NAND U5112 ( .A(n2050), .B(n2484), .Z(n2049) );
  AND U5113 ( .A(n897), .B(b_bus[6]), .Z(n2050) );
  MUX U5114 ( .A(n1022), .B(n1023), .S(n2051), .Z(n2048) );
  NOR U5115 ( .A(b_bus[6]), .B(n2484), .Z(n2051) );
  ANDN U5116 ( .B(reg_source[6]), .A(n1015), .Z(n2484) );
  ANDN U5117 ( .B(N24), .A(n1901), .Z(n1929) );
  AND U5118 ( .A(n2052), .B(n2053), .Z(n1901) );
  NAND U5119 ( .A(n17), .B(n2054), .Z(n2053) );
  NAND U5120 ( .A(n2055), .B(n2054), .Z(n2052) );
  NANDN U5121 ( .A(n824), .B(n130), .Z(n2055) );
  NAND U5122 ( .A(n821), .B(n125), .Z(n824) );
  NAND U5123 ( .A(n2056), .B(n2057), .Z(N24) );
  AND U5124 ( .A(n2058), .B(n2059), .Z(n2057) );
  AND U5125 ( .A(n2060), .B(n2061), .Z(n2059) );
  NAND U5126 ( .A(n2062), .B(n852), .Z(n2061) );
  NAND U5127 ( .A(n2063), .B(n2064), .Z(n2062) );
  AND U5128 ( .A(n2065), .B(n2066), .Z(n2064) );
  AND U5129 ( .A(n2067), .B(n2068), .Z(n2065) );
  NANDN U5130 ( .A(n1552), .B(a_bus[4]), .Z(n2068) );
  AND U5131 ( .A(n2069), .B(n2070), .Z(n1552) );
  NAND U5132 ( .A(n1175), .B(n1394), .Z(n2070) );
  ANDN U5133 ( .B(n2071), .A(n1606), .Z(n2069) );
  NAND U5134 ( .A(n1316), .B(n1403), .Z(n2071) );
  NANDN U5135 ( .A(n2072), .B(n863), .Z(n2067) );
  NAND U5136 ( .A(n2073), .B(n865), .Z(n2060) );
  NAND U5137 ( .A(n2063), .B(n2074), .Z(n2073) );
  AND U5138 ( .A(n2075), .B(n2066), .Z(n2074) );
  NAND U5139 ( .A(n888), .B(n1168), .Z(n2066) );
  AND U5140 ( .A(n2076), .B(n2077), .Z(n2075) );
  NANDN U5141 ( .A(n1554), .B(a_bus[4]), .Z(n2077) );
  AND U5142 ( .A(n2078), .B(n2079), .Z(n1554) );
  NAND U5143 ( .A(n1360), .B(n1175), .Z(n2079) );
  AND U5144 ( .A(n2080), .B(n2081), .Z(n2078) );
  NANDN U5145 ( .A(n1325), .B(n1403), .Z(n2081) );
  NANDN U5146 ( .A(n1324), .B(n1405), .Z(n2080) );
  NANDN U5147 ( .A(n2072), .B(n876), .Z(n2076) );
  AND U5148 ( .A(n2082), .B(n2083), .Z(n2063) );
  NAND U5149 ( .A(n870), .B(n1170), .Z(n2083) );
  NAND U5150 ( .A(n874), .B(n1161), .Z(n2082) );
  AND U5151 ( .A(n2084), .B(n2085), .Z(n2058) );
  NAND U5152 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][7] ), .Z(n2085) );
  ANDN U5153 ( .B(\Shifter/sll_27/ML_int[3][7] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][7] ) );
  NAND U5154 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N115 ), .Z(n2084) );
  AND U5155 ( .A(n2086), .B(n2087), .Z(n2056) );
  AND U5156 ( .A(n2088), .B(n2089), .Z(n2087) );
  NANDN U5157 ( .A(n891), .B(\ALU/N115 ), .Z(n2089) );
  NAND U5158 ( .A(n2090), .B(n1026), .Z(n2088) );
  XNOR U5159 ( .A(n984), .B(n2483), .Z(n2090) );
  AND U5160 ( .A(n2091), .B(n2092), .Z(n2086) );
  NAND U5161 ( .A(n2093), .B(n2483), .Z(n2092) );
  AND U5162 ( .A(n897), .B(b_bus[7]), .Z(n2093) );
  MUX U5163 ( .A(n1022), .B(n1023), .S(n2094), .Z(n2091) );
  NOR U5164 ( .A(b_bus[7]), .B(n2483), .Z(n2094) );
  ANDN U5165 ( .B(reg_source[7]), .A(n1015), .Z(n2483) );
  AND U5166 ( .A(n1924), .B(N27), .Z(n1915) );
  NAND U5167 ( .A(n2095), .B(n2096), .Z(N27) );
  AND U5168 ( .A(n2097), .B(n2098), .Z(n2096) );
  AND U5169 ( .A(n2099), .B(n2100), .Z(n2098) );
  NAND U5170 ( .A(n2101), .B(n852), .Z(n2100) );
  NAND U5171 ( .A(n2102), .B(n2103), .Z(n2101) );
  AND U5172 ( .A(n2104), .B(n2105), .Z(n2103) );
  AND U5173 ( .A(n2106), .B(n2107), .Z(n2104) );
  NANDN U5174 ( .A(n1528), .B(a_bus[4]), .Z(n2107) );
  AND U5175 ( .A(n2108), .B(n2109), .Z(n1528) );
  AND U5176 ( .A(n1945), .B(n2110), .Z(n2109) );
  NAND U5177 ( .A(n1127), .B(n1394), .Z(n2110) );
  NAND U5178 ( .A(n863), .B(n873), .Z(n2106) );
  NAND U5179 ( .A(n2111), .B(n865), .Z(n2099) );
  NAND U5180 ( .A(n2102), .B(n2112), .Z(n2111) );
  AND U5181 ( .A(n2113), .B(n2105), .Z(n2112) );
  NAND U5182 ( .A(n888), .B(n1133), .Z(n2105) );
  NAND U5183 ( .A(n2114), .B(n2115), .Z(n1133) );
  AND U5184 ( .A(n2116), .B(n2117), .Z(n2115) );
  NANDN U5185 ( .A(n881), .B(b_bus[16]), .Z(n2117) );
  NANDN U5186 ( .A(n882), .B(b_bus[17]), .Z(n2116) );
  AND U5187 ( .A(n2118), .B(n2119), .Z(n2114) );
  NANDN U5188 ( .A(n885), .B(b_bus[19]), .Z(n2119) );
  NANDN U5189 ( .A(n886), .B(b_bus[18]), .Z(n2118) );
  AND U5190 ( .A(n2120), .B(n2121), .Z(n2113) );
  NANDN U5191 ( .A(n1530), .B(a_bus[4]), .Z(n2121) );
  AND U5192 ( .A(n2108), .B(n2122), .Z(n1530) );
  NAND U5193 ( .A(n1360), .B(n1127), .Z(n2122) );
  NAND U5194 ( .A(n2123), .B(n2124), .Z(n1127) );
  AND U5195 ( .A(n2125), .B(n2126), .Z(n2124) );
  NANDN U5196 ( .A(n881), .B(b_bus[20]), .Z(n2126) );
  NANDN U5197 ( .A(n882), .B(b_bus[21]), .Z(n2125) );
  AND U5198 ( .A(n2127), .B(n2128), .Z(n2123) );
  NANDN U5199 ( .A(n885), .B(b_bus[23]), .Z(n2128) );
  NANDN U5200 ( .A(n886), .B(b_bus[22]), .Z(n2127) );
  AND U5201 ( .A(n2129), .B(n2130), .Z(n2108) );
  NAND U5202 ( .A(n1287), .B(n1403), .Z(n2130) );
  NAND U5203 ( .A(n2131), .B(n2132), .Z(n1287) );
  AND U5204 ( .A(n2133), .B(n2134), .Z(n2132) );
  NANDN U5205 ( .A(n881), .B(b_bus[24]), .Z(n2134) );
  NANDN U5206 ( .A(n882), .B(b_bus[25]), .Z(n2133) );
  AND U5207 ( .A(n2135), .B(n2136), .Z(n2131) );
  NANDN U5208 ( .A(n885), .B(b_bus[27]), .Z(n2136) );
  NANDN U5209 ( .A(n886), .B(b_bus[26]), .Z(n2135) );
  NAND U5210 ( .A(n1405), .B(n1286), .Z(n2129) );
  NAND U5211 ( .A(n2137), .B(n2138), .Z(n1286) );
  AND U5212 ( .A(n2139), .B(n2140), .Z(n2138) );
  NANDN U5213 ( .A(n881), .B(b_bus[28]), .Z(n2140) );
  NANDN U5214 ( .A(n882), .B(b_bus[29]), .Z(n2139) );
  AND U5215 ( .A(n2141), .B(n2142), .Z(n2137) );
  NANDN U5216 ( .A(n885), .B(\Shifter/N75 ), .Z(n2142) );
  NANDN U5217 ( .A(n886), .B(b_bus[30]), .Z(n2141) );
  NAND U5218 ( .A(n876), .B(n873), .Z(n2120) );
  NAND U5219 ( .A(n2143), .B(n2144), .Z(n873) );
  AND U5220 ( .A(n2145), .B(n2146), .Z(n2144) );
  NANDN U5221 ( .A(n881), .B(b_bus[4]), .Z(n2146) );
  NANDN U5222 ( .A(n882), .B(b_bus[5]), .Z(n2145) );
  AND U5223 ( .A(n2147), .B(n2148), .Z(n2143) );
  NANDN U5224 ( .A(n885), .B(b_bus[7]), .Z(n2148) );
  NANDN U5225 ( .A(n886), .B(b_bus[6]), .Z(n2147) );
  AND U5226 ( .A(n2149), .B(n2150), .Z(n2102) );
  NAND U5227 ( .A(n870), .B(n887), .Z(n2150) );
  NAND U5228 ( .A(n2151), .B(n2152), .Z(n887) );
  AND U5229 ( .A(n2153), .B(n2154), .Z(n2152) );
  NANDN U5230 ( .A(n881), .B(b_bus[12]), .Z(n2154) );
  NANDN U5231 ( .A(n882), .B(b_bus[13]), .Z(n2153) );
  AND U5232 ( .A(n2155), .B(n2156), .Z(n2151) );
  NANDN U5233 ( .A(n885), .B(b_bus[15]), .Z(n2156) );
  NANDN U5234 ( .A(n886), .B(b_bus[14]), .Z(n2155) );
  NAND U5235 ( .A(n874), .B(n869), .Z(n2149) );
  NAND U5236 ( .A(n2157), .B(n2158), .Z(n869) );
  AND U5237 ( .A(n2159), .B(n2160), .Z(n2158) );
  NANDN U5238 ( .A(n881), .B(b_bus[8]), .Z(n2160) );
  NANDN U5239 ( .A(n882), .B(b_bus[9]), .Z(n2159) );
  AND U5240 ( .A(n2161), .B(n2162), .Z(n2157) );
  NANDN U5241 ( .A(n885), .B(b_bus[11]), .Z(n2162) );
  NANDN U5242 ( .A(n886), .B(b_bus[10]), .Z(n2161) );
  AND U5243 ( .A(n2163), .B(n2164), .Z(n2097) );
  NAND U5244 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N112 ), .Z(n2164) );
  NANDN U5245 ( .A(n891), .B(\ALU/N112 ), .Z(n2163) );
  AND U5246 ( .A(n2165), .B(n2166), .Z(n2095) );
  AND U5247 ( .A(n2167), .B(n2168), .Z(n2166) );
  NAND U5248 ( .A(n2169), .B(n1026), .Z(n2168) );
  XOR U5249 ( .A(a_bus[4]), .B(b_bus[4]), .Z(n2169) );
  MUX U5250 ( .A(n1022), .B(n1023), .S(n2170), .Z(n2167) );
  AND U5251 ( .A(n990), .B(n1361), .Z(n2170) );
  MUX U5252 ( .A(n2171), .B(n2172), .S(a_bus[4]), .Z(n2165) );
  NAND U5253 ( .A(b_bus[4]), .B(n897), .Z(n2172) );
  NANDN U5254 ( .A(n1408), .B(\Shifter/sll_27/ML_int[4][4] ), .Z(n2171) );
  ANDN U5255 ( .B(\Shifter/sll_27/ML_int[3][4] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][4] ) );
  ANDN U5256 ( .B(N28), .A(n834), .Z(n1924) );
  IV U5257 ( .A(N29), .Z(n834) );
  NAND U5258 ( .A(n2173), .B(n2174), .Z(N29) );
  AND U5259 ( .A(n2175), .B(n2176), .Z(n2174) );
  AND U5260 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U5261 ( .A(n2179), .B(n852), .Z(n2178) );
  NAND U5262 ( .A(n2180), .B(n2181), .Z(n2179) );
  AND U5263 ( .A(n2182), .B(n2183), .Z(n2181) );
  AND U5264 ( .A(n2184), .B(n2185), .Z(n2182) );
  NANDN U5265 ( .A(n1479), .B(a_bus[4]), .Z(n2185) );
  AND U5266 ( .A(n2186), .B(n2187), .Z(n1479) );
  AND U5267 ( .A(n2188), .B(n2189), .Z(n2187) );
  NAND U5268 ( .A(n1211), .B(n1394), .Z(n2189) );
  AND U5269 ( .A(n2190), .B(n2191), .Z(n2186) );
  NAND U5270 ( .A(n1397), .B(n1683), .Z(n2190) );
  MUX U5271 ( .A(b_bus[30]), .B(\Shifter/N75 ), .S(n881), .Z(n1683) );
  AND U5272 ( .A(n2192), .B(n2193), .Z(n2180) );
  NAND U5273 ( .A(n2194), .B(n863), .Z(n2193) );
  NAND U5274 ( .A(n2195), .B(n865), .Z(n2177) );
  NAND U5275 ( .A(n2196), .B(n2197), .Z(n2195) );
  AND U5276 ( .A(n2198), .B(n2183), .Z(n2197) );
  NAND U5277 ( .A(n870), .B(n1201), .Z(n2183) );
  NAND U5278 ( .A(n2199), .B(n2200), .Z(n1201) );
  AND U5279 ( .A(n2201), .B(n2202), .Z(n2200) );
  NANDN U5280 ( .A(n881), .B(b_bus[10]), .Z(n2202) );
  NANDN U5281 ( .A(n882), .B(b_bus[11]), .Z(n2201) );
  AND U5282 ( .A(n2203), .B(n2204), .Z(n2199) );
  NANDN U5283 ( .A(n885), .B(b_bus[13]), .Z(n2204) );
  NANDN U5284 ( .A(n886), .B(b_bus[12]), .Z(n2203) );
  AND U5285 ( .A(n2184), .B(n2205), .Z(n2198) );
  NANDN U5286 ( .A(n1481), .B(a_bus[4]), .Z(n2205) );
  AND U5287 ( .A(n2206), .B(n2207), .Z(n1481) );
  AND U5288 ( .A(n2188), .B(n2208), .Z(n2207) );
  NAND U5289 ( .A(n1360), .B(n1211), .Z(n2208) );
  NAND U5290 ( .A(n2209), .B(n2210), .Z(n1211) );
  AND U5291 ( .A(n2211), .B(n2212), .Z(n2210) );
  NANDN U5292 ( .A(n881), .B(b_bus[18]), .Z(n2212) );
  NANDN U5293 ( .A(n882), .B(b_bus[19]), .Z(n2211) );
  AND U5294 ( .A(n2213), .B(n2214), .Z(n2209) );
  NANDN U5295 ( .A(n885), .B(b_bus[21]), .Z(n2214) );
  NANDN U5296 ( .A(n886), .B(b_bus[20]), .Z(n2213) );
  NAND U5297 ( .A(n1205), .B(n1403), .Z(n2188) );
  NAND U5298 ( .A(n2215), .B(n2216), .Z(n1205) );
  AND U5299 ( .A(n2217), .B(n2218), .Z(n2216) );
  NANDN U5300 ( .A(n881), .B(b_bus[22]), .Z(n2218) );
  NANDN U5301 ( .A(n882), .B(b_bus[23]), .Z(n2217) );
  AND U5302 ( .A(n2219), .B(n2220), .Z(n2215) );
  NANDN U5303 ( .A(n885), .B(b_bus[25]), .Z(n2220) );
  NANDN U5304 ( .A(n886), .B(b_bus[24]), .Z(n2219) );
  AND U5305 ( .A(n2221), .B(n2191), .Z(n2206) );
  NAND U5306 ( .A(n1405), .B(n1362), .Z(n2191) );
  NAND U5307 ( .A(n2222), .B(n2223), .Z(n1362) );
  AND U5308 ( .A(n2224), .B(n2225), .Z(n2223) );
  NANDN U5309 ( .A(n881), .B(b_bus[26]), .Z(n2225) );
  NANDN U5310 ( .A(n882), .B(b_bus[27]), .Z(n2224) );
  AND U5311 ( .A(n2226), .B(n2227), .Z(n2222) );
  NANDN U5312 ( .A(n885), .B(b_bus[29]), .Z(n2227) );
  NANDN U5313 ( .A(n886), .B(b_bus[28]), .Z(n2226) );
  NAND U5314 ( .A(n1359), .B(n1397), .Z(n2221) );
  ANDN U5315 ( .B(a_bus[3]), .A(n2228), .Z(n1397) );
  NAND U5316 ( .A(n2229), .B(n2230), .Z(n1359) );
  NANDN U5317 ( .A(n882), .B(\Shifter/N75 ), .Z(n2230) );
  NANDN U5318 ( .A(n881), .B(b_bus[30]), .Z(n2229) );
  NANDN U5319 ( .A(n2030), .B(n874), .Z(n2184) );
  AND U5320 ( .A(n2231), .B(n2232), .Z(n2030) );
  AND U5321 ( .A(n2233), .B(n2234), .Z(n2232) );
  NANDN U5322 ( .A(n881), .B(b_bus[6]), .Z(n2234) );
  NANDN U5323 ( .A(n882), .B(b_bus[7]), .Z(n2233) );
  AND U5324 ( .A(n2235), .B(n2236), .Z(n2231) );
  NANDN U5325 ( .A(n885), .B(b_bus[9]), .Z(n2236) );
  NANDN U5326 ( .A(n886), .B(b_bus[8]), .Z(n2235) );
  AND U5327 ( .A(n2192), .B(n2237), .Z(n2196) );
  NAND U5328 ( .A(n2194), .B(n876), .Z(n2237) );
  NAND U5329 ( .A(n2238), .B(n2239), .Z(n2194) );
  AND U5330 ( .A(n2240), .B(n2241), .Z(n2239) );
  NANDN U5331 ( .A(n881), .B(b_bus[2]), .Z(n2241) );
  NANDN U5332 ( .A(n882), .B(b_bus[3]), .Z(n2240) );
  AND U5333 ( .A(n2242), .B(n2243), .Z(n2238) );
  NANDN U5334 ( .A(n885), .B(b_bus[5]), .Z(n2243) );
  NANDN U5335 ( .A(n886), .B(b_bus[4]), .Z(n2242) );
  NAND U5336 ( .A(n888), .B(n1212), .Z(n2192) );
  NAND U5337 ( .A(n2244), .B(n2245), .Z(n1212) );
  AND U5338 ( .A(n2246), .B(n2247), .Z(n2245) );
  NANDN U5339 ( .A(n881), .B(b_bus[14]), .Z(n2247) );
  NANDN U5340 ( .A(n882), .B(b_bus[15]), .Z(n2246) );
  AND U5341 ( .A(n2248), .B(n2249), .Z(n2244) );
  NANDN U5342 ( .A(n885), .B(b_bus[17]), .Z(n2249) );
  NANDN U5343 ( .A(n886), .B(b_bus[16]), .Z(n2248) );
  AND U5344 ( .A(n2250), .B(n2251), .Z(n2175) );
  NAND U5345 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][2] ), .Z(n2251) );
  ANDN U5346 ( .B(\Shifter/sll_27/ML_int[3][2] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][2] ) );
  ANDN U5347 ( .B(\Shifter/sll_27/ML_int[2][2] ), .A(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][2] ) );
  NAND U5348 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N110 ), .Z(n2250) );
  AND U5349 ( .A(n2252), .B(n2253), .Z(n2173) );
  AND U5350 ( .A(n2254), .B(n2255), .Z(n2253) );
  NANDN U5351 ( .A(n891), .B(\ALU/N110 ), .Z(n2255) );
  NAND U5352 ( .A(n2256), .B(n1026), .Z(n2254) );
  XOR U5353 ( .A(a_bus[2]), .B(b_bus[2]), .Z(n2256) );
  AND U5354 ( .A(n2257), .B(n2258), .Z(n2252) );
  NAND U5355 ( .A(n2259), .B(n897), .Z(n2258) );
  AND U5356 ( .A(b_bus[2]), .B(a_bus[2]), .Z(n2259) );
  IV U5357 ( .A(n995), .Z(b_bus[2]) );
  MUX U5358 ( .A(n1022), .B(n1023), .S(n2260), .Z(n2257) );
  AND U5359 ( .A(n995), .B(n2228), .Z(n2260) );
  NAND U5360 ( .A(n2261), .B(n2262), .Z(N28) );
  AND U5361 ( .A(n2263), .B(n2264), .Z(n2262) );
  AND U5362 ( .A(n2265), .B(n2266), .Z(n2264) );
  NAND U5363 ( .A(n2267), .B(n852), .Z(n2266) );
  ANDN U5364 ( .B(n2268), .A(n2269), .Z(n852) );
  NAND U5365 ( .A(n2270), .B(n2271), .Z(n2267) );
  AND U5366 ( .A(n2272), .B(n2273), .Z(n2271) );
  AND U5367 ( .A(n2274), .B(n2275), .Z(n2272) );
  NANDN U5368 ( .A(n1456), .B(a_bus[4]), .Z(n2275) );
  AND U5369 ( .A(n2276), .B(n2277), .Z(n1456) );
  AND U5370 ( .A(n1945), .B(n2278), .Z(n2277) );
  NAND U5371 ( .A(n1168), .B(n1394), .Z(n2278) );
  NANDN U5372 ( .A(n2228), .B(n1606), .Z(n1945) );
  ANDN U5373 ( .B(\Shifter/N75 ), .A(n1174), .Z(n1606) );
  AND U5374 ( .A(n2279), .B(n2280), .Z(n2276) );
  NAND U5375 ( .A(n1405), .B(n1316), .Z(n2279) );
  NAND U5376 ( .A(n2281), .B(n2282), .Z(n1316) );
  ANDN U5377 ( .B(n2228), .A(n1174), .Z(n1405) );
  AND U5378 ( .A(n2283), .B(n2284), .Z(n2270) );
  NAND U5379 ( .A(n2285), .B(n863), .Z(n2284) );
  AND U5380 ( .A(n1394), .B(n1361), .Z(n863) );
  ANDN U5381 ( .B(n1174), .A(a_bus[2]), .Z(n1394) );
  NAND U5382 ( .A(n2286), .B(n865), .Z(n2265) );
  NOR U5383 ( .A(n2268), .B(n2269), .Z(n865) );
  NAND U5384 ( .A(n2287), .B(n2288), .Z(n2286) );
  AND U5385 ( .A(n2289), .B(n2273), .Z(n2288) );
  NAND U5386 ( .A(n870), .B(n1161), .Z(n2273) );
  NAND U5387 ( .A(n2290), .B(n2291), .Z(n1161) );
  AND U5388 ( .A(n2292), .B(n2293), .Z(n2291) );
  NANDN U5389 ( .A(n881), .B(b_bus[11]), .Z(n2293) );
  IV U5390 ( .A(n969), .Z(b_bus[11]) );
  NANDN U5391 ( .A(n882), .B(b_bus[12]), .Z(n2292) );
  IV U5392 ( .A(n965), .Z(b_bus[12]) );
  AND U5393 ( .A(n2294), .B(n2295), .Z(n2290) );
  NANDN U5394 ( .A(n885), .B(b_bus[14]), .Z(n2295) );
  IV U5395 ( .A(n960), .Z(b_bus[14]) );
  NANDN U5396 ( .A(n886), .B(b_bus[13]), .Z(n2294) );
  IV U5397 ( .A(n964), .Z(b_bus[13]) );
  AND U5398 ( .A(n2296), .B(n2228), .Z(n870) );
  AND U5399 ( .A(n2274), .B(n2297), .Z(n2289) );
  NANDN U5400 ( .A(n1458), .B(a_bus[4]), .Z(n2297) );
  AND U5401 ( .A(n2298), .B(n2299), .Z(n1458) );
  NAND U5402 ( .A(a_bus[3]), .B(n1172), .Z(n2299) );
  IV U5403 ( .A(n2300), .Z(n1172) );
  MUX U5404 ( .A(n1325), .B(n1324), .S(a_bus[2]), .Z(n2300) );
  NANDN U5405 ( .A(n881), .B(\Shifter/N75 ), .Z(n1324) );
  IV U5406 ( .A(n907), .Z(\Shifter/N75 ) );
  AND U5407 ( .A(n2281), .B(n2282), .Z(n1325) );
  AND U5408 ( .A(n2301), .B(n2302), .Z(n2282) );
  NANDN U5409 ( .A(n881), .B(b_bus[27]), .Z(n2302) );
  NANDN U5410 ( .A(n882), .B(b_bus[28]), .Z(n2301) );
  AND U5411 ( .A(n2303), .B(n2304), .Z(n2281) );
  NANDN U5412 ( .A(n885), .B(b_bus[30]), .Z(n2304) );
  NANDN U5413 ( .A(n886), .B(b_bus[29]), .Z(n2303) );
  AND U5414 ( .A(n2280), .B(n2305), .Z(n2298) );
  NAND U5415 ( .A(n1360), .B(n1168), .Z(n2305) );
  NAND U5416 ( .A(n2306), .B(n2307), .Z(n1168) );
  AND U5417 ( .A(n2308), .B(n2309), .Z(n2307) );
  NANDN U5418 ( .A(n881), .B(b_bus[19]), .Z(n2309) );
  NANDN U5419 ( .A(n882), .B(b_bus[20]), .Z(n2308) );
  AND U5420 ( .A(n2310), .B(n2311), .Z(n2306) );
  NANDN U5421 ( .A(n885), .B(b_bus[22]), .Z(n2311) );
  NANDN U5422 ( .A(n886), .B(b_bus[21]), .Z(n2310) );
  NAND U5423 ( .A(n1175), .B(n1403), .Z(n2280) );
  NAND U5424 ( .A(n2312), .B(n2313), .Z(n1175) );
  AND U5425 ( .A(n2314), .B(n2315), .Z(n2313) );
  NANDN U5426 ( .A(n881), .B(b_bus[23]), .Z(n2315) );
  NANDN U5427 ( .A(n882), .B(b_bus[24]), .Z(n2314) );
  AND U5428 ( .A(n2316), .B(n2317), .Z(n2312) );
  NANDN U5429 ( .A(n885), .B(b_bus[26]), .Z(n2317) );
  NANDN U5430 ( .A(n886), .B(b_bus[25]), .Z(n2316) );
  NANDN U5431 ( .A(n2072), .B(n874), .Z(n2274) );
  AND U5432 ( .A(n1403), .B(n1361), .Z(n874) );
  ANDN U5433 ( .B(n1174), .A(n2228), .Z(n1403) );
  AND U5434 ( .A(n2318), .B(n2319), .Z(n2072) );
  AND U5435 ( .A(n2320), .B(n2321), .Z(n2319) );
  NANDN U5436 ( .A(n881), .B(b_bus[7]), .Z(n2321) );
  IV U5437 ( .A(n984), .Z(b_bus[7]) );
  NANDN U5438 ( .A(n882), .B(b_bus[8]), .Z(n2320) );
  IV U5439 ( .A(n980), .Z(b_bus[8]) );
  AND U5440 ( .A(n2322), .B(n2323), .Z(n2318) );
  NANDN U5441 ( .A(n885), .B(b_bus[10]), .Z(n2323) );
  NANDN U5442 ( .A(n886), .B(b_bus[9]), .Z(n2322) );
  AND U5443 ( .A(n2283), .B(n2324), .Z(n2287) );
  NAND U5444 ( .A(n2285), .B(n876), .Z(n2324) );
  ANDN U5445 ( .B(n1360), .A(a_bus[4]), .Z(n876) );
  AND U5446 ( .A(n1174), .B(n2228), .Z(n1360) );
  NAND U5447 ( .A(n2325), .B(n2326), .Z(n2285) );
  AND U5448 ( .A(n2327), .B(n2328), .Z(n2326) );
  NANDN U5449 ( .A(n881), .B(b_bus[3]), .Z(n2328) );
  NANDN U5450 ( .A(n882), .B(b_bus[4]), .Z(n2327) );
  IV U5451 ( .A(n990), .Z(b_bus[4]) );
  AND U5452 ( .A(n2329), .B(n2330), .Z(n2325) );
  NANDN U5453 ( .A(n885), .B(b_bus[6]), .Z(n2330) );
  IV U5454 ( .A(n985), .Z(b_bus[6]) );
  NANDN U5455 ( .A(n886), .B(b_bus[5]), .Z(n2329) );
  IV U5456 ( .A(n989), .Z(b_bus[5]) );
  NAND U5457 ( .A(n888), .B(n1170), .Z(n2283) );
  NAND U5458 ( .A(n2331), .B(n2332), .Z(n1170) );
  AND U5459 ( .A(n2333), .B(n2334), .Z(n2332) );
  NANDN U5460 ( .A(n881), .B(b_bus[15]), .Z(n2334) );
  IV U5461 ( .A(n959), .Z(b_bus[15]) );
  NAND U5462 ( .A(n1003), .B(n1004), .Z(n881) );
  NANDN U5463 ( .A(n882), .B(b_bus[16]), .Z(n2333) );
  NAND U5464 ( .A(n1003), .B(a_bus[0]), .Z(n882) );
  IV U5465 ( .A(a_bus[1]), .Z(n1003) );
  AND U5466 ( .A(n2335), .B(n2336), .Z(n2331) );
  NANDN U5467 ( .A(n885), .B(b_bus[18]), .Z(n2336) );
  NAND U5468 ( .A(a_bus[1]), .B(a_bus[0]), .Z(n885) );
  NANDN U5469 ( .A(n886), .B(b_bus[17]), .Z(n2335) );
  IV U5470 ( .A(n954), .Z(b_bus[17]) );
  NAND U5471 ( .A(n1004), .B(a_bus[1]), .Z(n886) );
  MUX U5472 ( .A(reg_source[1]), .B(imm[7]), .S(n1015), .Z(a_bus[1]) );
  IV U5473 ( .A(a_bus[0]), .Z(n1004) );
  MUX U5474 ( .A(reg_source[0]), .B(imm[6]), .S(n1015), .Z(a_bus[0]) );
  ANDN U5475 ( .B(n2296), .A(n2228), .Z(n888) );
  IV U5476 ( .A(a_bus[2]), .Z(n2228) );
  ANDN U5477 ( .B(n1361), .A(n1174), .Z(n2296) );
  AND U5478 ( .A(n2337), .B(n2338), .Z(n2263) );
  NAND U5479 ( .A(n848), .B(\Shifter/sll_27/ML_int[4][3] ), .Z(n2338) );
  ANDN U5480 ( .B(\Shifter/sll_27/ML_int[3][3] ), .A(a_bus[3]), .Z(
        \Shifter/sll_27/ML_int[4][3] ) );
  ANDN U5481 ( .B(\Shifter/sll_27/ML_int[2][3] ), .A(a_bus[2]), .Z(
        \Shifter/sll_27/ML_int[3][3] ) );
  MUX U5482 ( .A(reg_source[2]), .B(imm[8]), .S(n1015), .Z(a_bus[2]) );
  ANDN U5483 ( .B(n1361), .A(n1408), .Z(n848) );
  NAND U5484 ( .A(n2269), .B(n2268), .Z(n1408) );
  AND U5485 ( .A(n2339), .B(n2340), .Z(n2268) );
  AND U5486 ( .A(n7), .B(n2341), .Z(n2339) );
  NANDN U5487 ( .A(n548), .B(n2342), .Z(n2341) );
  NAND U5488 ( .A(imm[1]), .B(imm[0]), .Z(n2342) );
  ANDN U5489 ( .B(n549), .A(imm[0]), .Z(n548) );
  NANDN U5490 ( .A(n2343), .B(n2340), .Z(n2269) );
  IV U5491 ( .A(a_bus[4]), .Z(n1361) );
  MUX U5492 ( .A(reg_source[4]), .B(imm[10]), .S(n1015), .Z(a_bus[4]) );
  NAND U5493 ( .A(\ALU/U2/U1/Z_0 ), .B(\ALU/N111 ), .Z(n2337) );
  AND U5494 ( .A(n2344), .B(n2345), .Z(n2261) );
  AND U5495 ( .A(n2346), .B(n2347), .Z(n2345) );
  NANDN U5496 ( .A(n891), .B(\ALU/N111 ), .Z(n2347) );
  NAND U5497 ( .A(n903), .B(n2348), .Z(n891) );
  NAND U5498 ( .A(n2349), .B(n1026), .Z(n2346) );
  ANDN U5499 ( .B(n901), .A(n903), .Z(n1026) );
  AND U5500 ( .A(n1019), .B(n2350), .Z(n901) );
  XOR U5501 ( .A(a_bus[3]), .B(b_bus[3]), .Z(n2349) );
  AND U5502 ( .A(n2351), .B(n2352), .Z(n2344) );
  NAND U5503 ( .A(n2353), .B(n897), .Z(n2352) );
  ANDN U5504 ( .B(n2354), .A(n903), .Z(n897) );
  AND U5505 ( .A(b_bus[3]), .B(a_bus[3]), .Z(n2353) );
  IV U5506 ( .A(n994), .Z(b_bus[3]) );
  MUX U5507 ( .A(n1022), .B(n1023), .S(n2355), .Z(n2351) );
  AND U5508 ( .A(n994), .B(n1174), .Z(n2355) );
  IV U5509 ( .A(a_bus[3]), .Z(n1174) );
  MUX U5510 ( .A(reg_source[3]), .B(imm[9]), .S(n1015), .Z(a_bus[3]) );
  AND U5511 ( .A(n2356), .B(n2340), .Z(n1015) );
  ANDN U5512 ( .B(n547), .A(n821), .Z(n2340) );
  AND U5513 ( .A(n2357), .B(n569), .Z(n547) );
  AND U5514 ( .A(n7), .B(n2358), .Z(n2356) );
  NANDN U5515 ( .A(n2359), .B(n2360), .Z(n2358) );
  NAND U5516 ( .A(n543), .B(n2361), .Z(n2360) );
  NAND U5517 ( .A(n2362), .B(n2363), .Z(n1023) );
  AND U5518 ( .A(n2364), .B(imm[0]), .Z(n2363) );
  AND U5519 ( .A(n10), .B(imm[2]), .Z(n2364) );
  NOR U5520 ( .A(n2343), .B(n444), .Z(n2362) );
  NAND U5521 ( .A(imm[1]), .B(n7), .Z(n2343) );
  NANDN U5522 ( .A(n903), .B(n2348), .Z(n1022) );
  AND U5523 ( .A(n1019), .B(n1017), .Z(n2348) );
  XOR U5524 ( .A(n974), .B(n2365), .Z(\ALU/r67/B_AS[9] ) );
  IV U5525 ( .A(b_bus[9]), .Z(n974) );
  NAND U5526 ( .A(n2366), .B(n2367), .Z(b_bus[9]) );
  NAND U5527 ( .A(n2368), .B(imm[9]), .Z(n2367) );
  NANDN U5528 ( .A(n2369), .B(reg_target[9]), .Z(n2366) );
  XOR U5529 ( .A(n980), .B(n2365), .Z(\ALU/r67/B_AS[8] ) );
  NOR U5530 ( .A(n2370), .B(n2371), .Z(n980) );
  ANDN U5531 ( .B(reg_target[8]), .A(n2369), .Z(n2371) );
  ANDN U5532 ( .B(imm[8]), .A(n2372), .Z(n2370) );
  XOR U5533 ( .A(n984), .B(n2365), .Z(\ALU/r67/B_AS[7] ) );
  NOR U5534 ( .A(n2373), .B(n2374), .Z(n984) );
  ANDN U5535 ( .B(imm[7]), .A(n2372), .Z(n2374) );
  ANDN U5536 ( .B(reg_target[7]), .A(n2369), .Z(n2373) );
  XOR U5537 ( .A(n985), .B(n2365), .Z(\ALU/r67/B_AS[6] ) );
  NOR U5538 ( .A(n2375), .B(n2376), .Z(n985) );
  ANDN U5539 ( .B(reg_target[6]), .A(n2369), .Z(n2376) );
  ANDN U5540 ( .B(imm[6]), .A(n2372), .Z(n2375) );
  XOR U5541 ( .A(n989), .B(n2365), .Z(\ALU/r67/B_AS[5] ) );
  NOR U5542 ( .A(n2377), .B(n2378), .Z(n989) );
  ANDN U5543 ( .B(imm[5]), .A(n2372), .Z(n2378) );
  ANDN U5544 ( .B(reg_target[5]), .A(n2369), .Z(n2377) );
  XOR U5545 ( .A(n990), .B(n2365), .Z(\ALU/r67/B_AS[4] ) );
  NOR U5546 ( .A(n2379), .B(n2380), .Z(n990) );
  ANDN U5547 ( .B(reg_target[4]), .A(n2369), .Z(n2380) );
  ANDN U5548 ( .B(imm[4]), .A(n2372), .Z(n2379) );
  XOR U5549 ( .A(n994), .B(n2365), .Z(\ALU/r67/B_AS[3] ) );
  NOR U5550 ( .A(n2381), .B(n2382), .Z(n994) );
  ANDN U5551 ( .B(imm[3]), .A(n2372), .Z(n2382) );
  ANDN U5552 ( .B(reg_target[3]), .A(n2369), .Z(n2381) );
  XOR U5553 ( .A(n907), .B(n2365), .Z(\ALU/r67/B_AS[31] ) );
  AND U5554 ( .A(n2383), .B(n918), .Z(n907) );
  NANDN U5555 ( .A(n2369), .B(reg_target[31]), .Z(n2383) );
  XOR U5556 ( .A(n1764), .B(n2365), .Z(\ALU/r67/B_AS[30] ) );
  IV U5557 ( .A(b_bus[30]), .Z(n1764) );
  NAND U5558 ( .A(n2384), .B(n918), .Z(b_bus[30]) );
  NANDN U5559 ( .A(n2369), .B(reg_target[30]), .Z(n2384) );
  XOR U5560 ( .A(n995), .B(n2365), .Z(\ALU/r67/B_AS[2] ) );
  NOR U5561 ( .A(n2385), .B(n2386), .Z(n995) );
  ANDN U5562 ( .B(reg_target[2]), .A(n2369), .Z(n2386) );
  ANDN U5563 ( .B(imm[2]), .A(n2372), .Z(n2385) );
  XOR U5564 ( .A(n1719), .B(n2365), .Z(\ALU/r67/B_AS[29] ) );
  IV U5565 ( .A(b_bus[29]), .Z(n1719) );
  NAND U5566 ( .A(n919), .B(n918), .Z(b_bus[29]) );
  NANDN U5567 ( .A(n2369), .B(reg_target[29]), .Z(n919) );
  XOR U5568 ( .A(n920), .B(n2365), .Z(\ALU/r67/B_AS[28] ) );
  NAND U5569 ( .A(n1014), .B(n918), .Z(b_bus[28]) );
  NANDN U5570 ( .A(n2369), .B(reg_target[28]), .Z(n1014) );
  XOR U5571 ( .A(n1667), .B(n2365), .Z(\ALU/r67/B_AS[27] ) );
  IV U5572 ( .A(b_bus[27]), .Z(n1667) );
  NAND U5573 ( .A(n925), .B(n918), .Z(b_bus[27]) );
  NANDN U5574 ( .A(n2369), .B(reg_target[27]), .Z(n925) );
  XOR U5575 ( .A(n926), .B(n2365), .Z(\ALU/r67/B_AS[26] ) );
  NAND U5576 ( .A(n1013), .B(n918), .Z(b_bus[26]) );
  NANDN U5577 ( .A(n2369), .B(reg_target[26]), .Z(n1013) );
  XOR U5578 ( .A(n1617), .B(n2365), .Z(\ALU/r67/B_AS[25] ) );
  IV U5579 ( .A(b_bus[25]), .Z(n1617) );
  NAND U5580 ( .A(n931), .B(n918), .Z(b_bus[25]) );
  NANDN U5581 ( .A(n2369), .B(reg_target[25]), .Z(n931) );
  XOR U5582 ( .A(n932), .B(n2365), .Z(\ALU/r67/B_AS[24] ) );
  NAND U5583 ( .A(n1012), .B(n918), .Z(b_bus[24]) );
  NANDN U5584 ( .A(n2369), .B(reg_target[24]), .Z(n1012) );
  XOR U5585 ( .A(n1562), .B(n2365), .Z(\ALU/r67/B_AS[23] ) );
  IV U5586 ( .A(b_bus[23]), .Z(n1562) );
  NAND U5587 ( .A(n937), .B(n918), .Z(b_bus[23]) );
  NANDN U5588 ( .A(n2369), .B(reg_target[23]), .Z(n937) );
  XOR U5589 ( .A(n938), .B(n2365), .Z(\ALU/r67/B_AS[22] ) );
  NAND U5590 ( .A(n1011), .B(n918), .Z(b_bus[22]) );
  NANDN U5591 ( .A(n2369), .B(reg_target[22]), .Z(n1011) );
  XOR U5592 ( .A(n1515), .B(n2365), .Z(\ALU/r67/B_AS[21] ) );
  IV U5593 ( .A(b_bus[21]), .Z(n1515) );
  NAND U5594 ( .A(n943), .B(n918), .Z(b_bus[21]) );
  NANDN U5595 ( .A(n2369), .B(reg_target[21]), .Z(n943) );
  XOR U5596 ( .A(n944), .B(n2365), .Z(\ALU/r67/B_AS[20] ) );
  NAND U5597 ( .A(n1010), .B(n918), .Z(b_bus[20]) );
  NANDN U5598 ( .A(n2369), .B(reg_target[20]), .Z(n1010) );
  XOR U5599 ( .A(n1001), .B(n2365), .Z(\ALU/r67/B_AS[1] ) );
  IV U5600 ( .A(b_bus[1]), .Z(n1001) );
  NAND U5601 ( .A(n2387), .B(n2388), .Z(b_bus[1]) );
  NAND U5602 ( .A(imm[1]), .B(n2368), .Z(n2388) );
  NANDN U5603 ( .A(n2369), .B(reg_target[1]), .Z(n2387) );
  XOR U5604 ( .A(n1466), .B(n2365), .Z(\ALU/r67/B_AS[19] ) );
  IV U5605 ( .A(b_bus[19]), .Z(n1466) );
  NAND U5606 ( .A(n949), .B(n918), .Z(b_bus[19]) );
  NANDN U5607 ( .A(n2369), .B(reg_target[19]), .Z(n949) );
  XOR U5608 ( .A(n950), .B(n2365), .Z(\ALU/r67/B_AS[18] ) );
  NAND U5609 ( .A(n1009), .B(n918), .Z(b_bus[18]) );
  NANDN U5610 ( .A(n2369), .B(reg_target[18]), .Z(n1009) );
  XOR U5611 ( .A(n954), .B(n2365), .Z(\ALU/r67/B_AS[17] ) );
  NOR U5612 ( .A(n2389), .B(n2390), .Z(n954) );
  ANDN U5613 ( .B(reg_target[17]), .A(n2369), .Z(n2390) );
  ANDN U5614 ( .B(imm[15]), .A(n2391), .Z(n2389) );
  XOR U5615 ( .A(n955), .B(n2365), .Z(\ALU/r67/B_AS[16] ) );
  NAND U5616 ( .A(n1008), .B(n918), .Z(b_bus[16]) );
  NANDN U5617 ( .A(n2391), .B(imm[15]), .Z(n918) );
  NANDN U5618 ( .A(n2369), .B(reg_target[16]), .Z(n1008) );
  XOR U5619 ( .A(n959), .B(n2365), .Z(\ALU/r67/B_AS[15] ) );
  NOR U5620 ( .A(n2392), .B(n2393), .Z(n959) );
  ANDN U5621 ( .B(reg_target[15]), .A(n2369), .Z(n2393) );
  ANDN U5622 ( .B(imm[15]), .A(n2372), .Z(n2392) );
  XOR U5623 ( .A(n960), .B(n2365), .Z(\ALU/r67/B_AS[14] ) );
  NOR U5624 ( .A(n2394), .B(n2395), .Z(n960) );
  ANDN U5625 ( .B(imm[14]), .A(n2372), .Z(n2395) );
  ANDN U5626 ( .B(reg_target[14]), .A(n2369), .Z(n2394) );
  XOR U5627 ( .A(n964), .B(n2365), .Z(\ALU/r67/B_AS[13] ) );
  NOR U5628 ( .A(n2396), .B(n2397), .Z(n964) );
  ANDN U5629 ( .B(reg_target[13]), .A(n2369), .Z(n2397) );
  ANDN U5630 ( .B(imm[13]), .A(n2372), .Z(n2396) );
  XOR U5631 ( .A(n965), .B(n2365), .Z(\ALU/r67/B_AS[12] ) );
  NOR U5632 ( .A(n2398), .B(n2399), .Z(n965) );
  ANDN U5633 ( .B(imm[12]), .A(n2372), .Z(n2399) );
  ANDN U5634 ( .B(reg_target[12]), .A(n2369), .Z(n2398) );
  XOR U5635 ( .A(n969), .B(n2365), .Z(\ALU/r67/B_AS[11] ) );
  NOR U5636 ( .A(n2400), .B(n2401), .Z(n969) );
  ANDN U5637 ( .B(reg_target[11]), .A(n2369), .Z(n2401) );
  ANDN U5638 ( .B(imm[11]), .A(n2372), .Z(n2400) );
  XOR U5639 ( .A(n977), .B(n2365), .Z(\ALU/r67/B_AS[10] ) );
  IV U5640 ( .A(\ALU/U2/U1/Z_0 ), .Z(n2365) );
  IV U5641 ( .A(b_bus[10]), .Z(n977) );
  NAND U5642 ( .A(n2402), .B(n2403), .Z(b_bus[10]) );
  NAND U5643 ( .A(n2368), .B(imm[10]), .Z(n2403) );
  NANDN U5644 ( .A(n2369), .B(reg_target[10]), .Z(n2402) );
  XNOR U5645 ( .A(n1005), .B(\ALU/U2/U1/Z_0 ), .Z(\ALU/r67/B_AS[0] ) );
  IV U5646 ( .A(b_bus[0]), .Z(n1005) );
  NAND U5647 ( .A(n2404), .B(n2405), .Z(b_bus[0]) );
  NAND U5648 ( .A(imm[0]), .B(n2368), .Z(n2405) );
  IV U5649 ( .A(n2372), .Z(n2368) );
  AND U5650 ( .A(n2391), .B(n2406), .Z(n2372) );
  NANDN U5651 ( .A(n2369), .B(reg_target[0]), .Z(n2404) );
  NAND U5652 ( .A(n2406), .B(n2391), .Z(n2369) );
  AND U5653 ( .A(n2407), .B(n2408), .Z(n2391) );
  ANDN U5654 ( .B(n2409), .A(n2410), .Z(n2407) );
  NANDN U5655 ( .A(n431), .B(n2411), .Z(n2409) );
  NANDN U5656 ( .A(n2412), .B(n125), .Z(n2411) );
  NANDN U5657 ( .A(n431), .B(n2413), .Z(n2406) );
  NAND U5658 ( .A(n2414), .B(n825), .Z(n2413) );
  AND U5659 ( .A(n2354), .B(n903), .Z(\ALU/U2/U1/Z_0 ) );
  IV U5660 ( .A(n1018), .Z(n903) );
  NAND U5661 ( .A(n2415), .B(n2416), .Z(n1018) );
  NAND U5662 ( .A(n2417), .B(n7), .Z(n2416) );
  NAND U5663 ( .A(n2418), .B(n2419), .Z(n2417) );
  AND U5664 ( .A(n1770), .B(n2420), .Z(n2419) );
  AND U5665 ( .A(n2421), .B(n2422), .Z(n2420) );
  NANDN U5666 ( .A(n444), .B(n2423), .Z(n2422) );
  NANDN U5667 ( .A(n110), .B(n2424), .Z(n2423) );
  ANDN U5668 ( .B(n549), .A(n2361), .Z(n110) );
  NAND U5669 ( .A(n448), .B(n540), .Z(n2421) );
  AND U5670 ( .A(n2425), .B(imm[1]), .Z(n540) );
  AND U5671 ( .A(n543), .B(n2361), .Z(n2425) );
  IV U5672 ( .A(imm[0]), .Z(n543) );
  AND U5673 ( .A(n793), .B(n794), .Z(n2418) );
  AND U5674 ( .A(n2426), .B(n2427), .Z(n2415) );
  NANDN U5675 ( .A(n431), .B(n2428), .Z(n2427) );
  NAND U5676 ( .A(n2414), .B(n2429), .Z(n2428) );
  ANDN U5677 ( .B(n125), .A(n2430), .Z(n2429) );
  NOR U5678 ( .A(n1017), .B(n1019), .Z(n2354) );
  NAND U5679 ( .A(n2431), .B(n2432), .Z(n1019) );
  AND U5680 ( .A(n2426), .B(n2433), .Z(n2432) );
  ANDN U5681 ( .B(n2408), .A(n2410), .Z(n2433) );
  AND U5682 ( .A(n2434), .B(n2054), .Z(n2410) );
  ANDN U5683 ( .B(n2435), .A(n2436), .Z(n2054) );
  OR U5684 ( .A(n2412), .B(n89), .Z(n2434) );
  NAND U5685 ( .A(n130), .B(n125), .Z(n89) );
  NAND U5686 ( .A(n458), .B(n241), .Z(n2408) );
  AND U5687 ( .A(n2435), .B(n2436), .Z(n241) );
  NOR U5688 ( .A(n132), .B(opcode[30]), .Z(n2435) );
  NAND U5689 ( .A(n2437), .B(n2438), .Z(n458) );
  ANDN U5690 ( .B(n125), .A(n818), .Z(n2438) );
  OR U5691 ( .A(n2439), .B(opcode[26]), .Z(n125) );
  ANDN U5692 ( .B(n825), .A(n2412), .Z(n2437) );
  NAND U5693 ( .A(n821), .B(n128), .Z(n2412) );
  NAND U5694 ( .A(n2440), .B(n2441), .Z(n2426) );
  AND U5695 ( .A(n122), .B(n10), .Z(n2441) );
  NOR U5696 ( .A(opcode[22]), .B(opcode[21]), .Z(n122) );
  ANDN U5697 ( .B(n24), .A(n121), .Z(n2440) );
  OR U5698 ( .A(opcode[24]), .B(opcode[25]), .Z(n121) );
  AND U5699 ( .A(n2442), .B(opcode[30]), .Z(n24) );
  AND U5700 ( .A(n132), .B(n2436), .Z(n2442) );
  IV U5701 ( .A(opcode[29]), .Z(n2436) );
  IV U5702 ( .A(opcode[31]), .Z(n132) );
  AND U5703 ( .A(n2443), .B(n2444), .Z(n2431) );
  NAND U5704 ( .A(n2445), .B(n7), .Z(n2444) );
  NAND U5705 ( .A(n2446), .B(n793), .Z(n2445) );
  ANDN U5706 ( .B(n2447), .A(n2448), .Z(n793) );
  IV U5707 ( .A(n2414), .Z(n2448) );
  ANDN U5708 ( .B(n127), .A(n2430), .Z(n2447) );
  NANDN U5709 ( .A(n2449), .B(n2450), .Z(n127) );
  AND U5710 ( .A(opcode[26]), .B(opcode[28]), .Z(n2450) );
  AND U5711 ( .A(n794), .B(n2451), .Z(n2446) );
  NAND U5712 ( .A(n10), .B(n2452), .Z(n2451) );
  NAND U5713 ( .A(n2453), .B(n2454), .Z(n2452) );
  NANDN U5714 ( .A(n444), .B(n2455), .Z(n2454) );
  NANDN U5715 ( .A(n2456), .B(n542), .Z(n2455) );
  NAND U5716 ( .A(n2361), .B(n549), .Z(n542) );
  MUX U5717 ( .A(n2457), .B(n549), .S(imm[0]), .Z(n2456) );
  AND U5718 ( .A(imm[1]), .B(imm[2]), .Z(n2457) );
  AND U5719 ( .A(n2458), .B(n1770), .Z(n2453) );
  NAND U5720 ( .A(n549), .B(n108), .Z(n1770) );
  ANDN U5721 ( .B(n2357), .A(n569), .Z(n108) );
  NOR U5722 ( .A(imm[4]), .B(imm[5]), .Z(n2357) );
  NAND U5723 ( .A(n557), .B(n21), .Z(n794) );
  NOR U5724 ( .A(opcode[17]), .B(opcode[18]), .Z(n21) );
  AND U5725 ( .A(n2459), .B(n17), .Z(n557) );
  IV U5726 ( .A(opcode[19]), .Z(n2459) );
  NANDN U5727 ( .A(n431), .B(n2460), .Z(n2443) );
  NAND U5728 ( .A(n2461), .B(n2462), .Z(n2460) );
  AND U5729 ( .A(n821), .B(n128), .Z(n2462) );
  IV U5730 ( .A(n17), .Z(n128) );
  AND U5731 ( .A(n2463), .B(opcode[26]), .Z(n17) );
  IV U5732 ( .A(n10), .Z(n821) );
  AND U5733 ( .A(n130), .B(n2414), .Z(n2461) );
  NOR U5734 ( .A(n817), .B(n818), .Z(n2414) );
  IV U5735 ( .A(n2464), .Z(n130) );
  IV U5736 ( .A(n2350), .Z(n1017) );
  NAND U5737 ( .A(n2465), .B(n2466), .Z(n2350) );
  NANDN U5738 ( .A(n431), .B(n2467), .Z(n2466) );
  NAND U5739 ( .A(n131), .B(n825), .Z(n2467) );
  NOR U5740 ( .A(n2464), .B(n2430), .Z(n825) );
  ANDN U5741 ( .B(opcode[26]), .A(n2439), .Z(n2464) );
  NAND U5742 ( .A(opcode[27]), .B(n2468), .Z(n2439) );
  IV U5743 ( .A(n817), .Z(n131) );
  AND U5744 ( .A(n2469), .B(opcode[27]), .Z(n817) );
  AND U5745 ( .A(n2470), .B(opcode[28]), .Z(n2469) );
  NAND U5746 ( .A(opcode[29]), .B(n2471), .Z(n431) );
  NAND U5747 ( .A(n2472), .B(n7), .Z(n2465) );
  ANDN U5748 ( .B(n2471), .A(opcode[29]), .Z(n7) );
  NOR U5749 ( .A(opcode[31]), .B(opcode[30]), .Z(n2471) );
  NAND U5750 ( .A(n2473), .B(n90), .Z(n2472) );
  NOR U5751 ( .A(n818), .B(n2430), .Z(n90) );
  NOR U5752 ( .A(opcode[26]), .B(n2474), .Z(n2430) );
  ANDN U5753 ( .B(opcode[26]), .A(n2474), .Z(n818) );
  NAND U5754 ( .A(opcode[28]), .B(n2449), .Z(n2474) );
  NAND U5755 ( .A(n10), .B(n2475), .Z(n2473) );
  NAND U5756 ( .A(n2476), .B(n2458), .Z(n2475) );
  NANDN U5757 ( .A(n572), .B(n553), .Z(n2458) );
  AND U5758 ( .A(n2477), .B(imm[0]), .Z(n553) );
  AND U5759 ( .A(n2361), .B(imm[1]), .Z(n2477) );
  IV U5760 ( .A(n448), .Z(n572) );
  AND U5761 ( .A(n2478), .B(imm[5]), .Z(n448) );
  AND U5762 ( .A(n571), .B(imm[3]), .Z(n2478) );
  NANDN U5763 ( .A(n444), .B(n2479), .Z(n2476) );
  NANDN U5764 ( .A(n2359), .B(n2424), .Z(n2479) );
  NANDN U5765 ( .A(imm[0]), .B(imm[2]), .Z(n2424) );
  ANDN U5766 ( .B(n2361), .A(n549), .Z(n2359) );
  IV U5767 ( .A(imm[1]), .Z(n549) );
  IV U5768 ( .A(imm[2]), .Z(n2361) );
  NAND U5769 ( .A(n2480), .B(imm[5]), .Z(n444) );
  AND U5770 ( .A(n569), .B(n571), .Z(n2480) );
  IV U5771 ( .A(imm[4]), .Z(n571) );
  IV U5772 ( .A(imm[3]), .Z(n569) );
  AND U5773 ( .A(n2463), .B(n2470), .Z(n10) );
  IV U5774 ( .A(opcode[26]), .Z(n2470) );
  AND U5775 ( .A(n2449), .B(n2468), .Z(n2463) );
  IV U5776 ( .A(opcode[28]), .Z(n2468) );
  IV U5777 ( .A(opcode[27]), .Z(n2449) );
endmodule

