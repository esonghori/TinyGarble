
module aes_seq ( clk, rst, g_init, e_init, o );
  input [127:0] g_init;
  input [127:0] e_init;
  output [127:0] o;
  input clk, rst;
  wire   N5, N6, N7, n7, \e/n118 , \e/n117 , \e/n116 , \e/n115 , \e/n114 ,
         \e/n113 , \e/n112 , \e/n111 , \e/n110 , \e/n109 , \e/n108 , \e/n107 ,
         \e/n106 , \e/n105 , \e/n104 , \e/n103 , \e/n102 , \e/n101 , \e/n100 ,
         \e/n99 , \e/n98 , \e/n97 , \e/n96 , \e/n95 , \e/n94 , \e/n93 ,
         \e/n92 , \e/n91 , \e/n90 , \e/n89 , \e/n88 , \e/n87 , \e/n85 ,
         \e/n84 , \e/n83 , \e/n82 , \e/n81 , \e/n80 , \e/n79 , \e/n78 ,
         \e/n77 , \e/n76 , \e/n75 , \e/n74 , \e/n73 , \e/n72 , \e/n71 ,
         \e/n70 , \e/n69 , \e/n68 , \e/n67 , \e/n66 , \e/n65 , \e/n64 ,
         \e/n63 , \e/n62 , \e/n61 , \e/n60 , \e/n59 , \e/n58 , \e/n57 ,
         \e/n56 , \e/n55 , \e/n54 , \e/Q[7] , \e/Q[6] , \e/Q[5] , \e/Q[4] ,
         \e/Q[3] , \e/Q[2] , \e/Q[1] , \e/Q[0] , \e/t[8] , \e/t[9] , \e/t[10] ,
         \e/t[11] , \e/t[12] , \e/t[13] , \e/t[14] , \e/t[15] , \e/t[16] ,
         \e/t[17] , \e/t[18] , \e/t[19] , \e/t[20] , \e/t[21] , \e/t[22] ,
         \e/t[23] , \e/t[24] , \e/t[25] , \e/t[26] , \e/t[27] , \e/t[28] ,
         \e/t[29] , \e/t[30] , \e/t[31] , \b/n6877 , \b/n6876 , \b/n6875 ,
         \b/n6874 , \b/n6872 , \b/n6871 , \b/n6870 , \b/n6869 , \b/n6868 ,
         \b/n6867 , \b/n6863 , \b/n6861 , \b/n6860 , \b/n6859 , \b/n6857 ,
         \b/n6854 , \b/n6853 , \b/n6852 , \b/n6851 , \b/n6850 , \b/n6849 ,
         \b/n6848 , \b/n6847 , \b/n6846 , \b/n6845 , \b/n6844 , \b/n6843 ,
         \b/n6842 , \b/n6841 , \b/n6840 , \b/n6839 , \b/n6838 , \b/n6837 ,
         \b/n6836 , \b/n6835 , \b/n6834 , \b/n6833 , \b/n6832 , \b/n6831 ,
         \b/n6830 , \b/n6829 , \b/n6828 , \b/n6827 , \b/n6826 , \b/n6825 ,
         \b/n6824 , \b/n6823 , \b/n6822 , \b/n6821 , \b/n6820 , \b/n6819 ,
         \b/n6818 , \b/n6817 , \b/n6816 , \b/n6815 , \b/n6814 , \b/n6813 ,
         \b/n6812 , \b/n6811 , \b/n6810 , \b/n6809 , \b/n6808 , \b/n6807 ,
         \b/n6806 , \b/n6805 , \b/n6804 , \b/n6803 , \b/n6802 , \b/n6801 ,
         \b/n6800 , \b/n6799 , \b/n6798 , \b/n6797 , \b/n6796 , \b/n6795 ,
         \b/n6794 , \b/n6793 , \b/n6792 , \b/n6791 , \b/n6790 , \b/n6789 ,
         \b/n6788 , \b/n6787 , \b/n6786 , \b/n6785 , \b/n6784 , \b/n6783 ,
         \b/n6782 , \b/n6781 , \b/n6780 , \b/n6779 , \b/n6778 , \b/n6777 ,
         \b/n6776 , \b/n6775 , \b/n6774 , \b/n6773 , \b/n6772 , \b/n6771 ,
         \b/n6770 , \b/n6769 , \b/n6768 , \b/n6767 , \b/n6766 , \b/n6765 ,
         \b/n6764 , \b/n6763 , \b/n6762 , \b/n6761 , \b/n6760 , \b/n6759 ,
         \b/n6758 , \b/n6757 , \b/n6756 , \b/n6755 , \b/n6754 , \b/n6753 ,
         \b/n6752 , \b/n6751 , \b/n6750 , \b/n6749 , \b/n6748 , \b/n6747 ,
         \b/n6746 , \b/n6745 , \b/n6744 , \b/n6743 , \b/n6742 , \b/n6741 ,
         \b/n6740 , \b/n6739 , \b/n6738 , \b/n6737 , \b/n6736 , \b/n6735 ,
         \b/n6734 , \b/n6733 , \b/n6732 , \b/n6731 , \b/n6730 , \b/n6729 ,
         \b/n6728 , \b/n6727 , \b/n6726 , \b/n6725 , \b/n6724 , \b/n6723 ,
         \b/n6722 , \b/n6721 , \b/n6720 , \b/n6719 , \b/n6718 , \b/n6717 ,
         \b/n6716 , \b/n6715 , \b/n6714 , \b/n6713 , \b/n6712 , \b/n6711 ,
         \b/n6710 , \b/n6709 , \b/n6708 , \b/n6707 , \b/n6706 , \b/n6705 ,
         \b/n6704 , \b/n6703 , \b/n6702 , \b/n6701 , \b/n6700 , \b/n6699 ,
         \b/n6698 , \b/n6697 , \b/n6696 , \b/n6695 , \b/n6694 , \b/n6693 ,
         \b/n6692 , \b/n6691 , \b/n6690 , \b/n6689 , \b/n6688 , \b/n6687 ,
         \b/n6686 , \b/n6685 , \b/n6684 , \b/n6683 , \b/n6682 , \b/n6681 ,
         \b/n6680 , \b/n6679 , \b/n6678 , \b/n6677 , \b/n6676 , \b/n6675 ,
         \b/n6674 , \b/n6673 , \b/n6672 , \b/n6671 , \b/n6670 , \b/n6669 ,
         \b/n6668 , \b/n6667 , \b/n6666 , \b/n6665 , \b/n6664 , \b/n6663 ,
         \b/n6662 , \b/n6661 , \b/n6660 , \b/n6659 , \b/n6658 , \b/n6657 ,
         \b/n6656 , \b/n6655 , \b/n6654 , \b/n6653 , \b/n6652 , \b/n6651 ,
         \b/n6650 , \b/n6649 , \b/n6648 , \b/n6647 , \b/n6646 , \b/n6645 ,
         \b/n6644 , \b/n6643 , \b/n6642 , \b/n6641 , \b/n6640 , \b/n6639 ,
         \b/n6638 , \b/n6637 , \b/n6636 , \b/n6635 , \b/n6634 , \b/n6633 ,
         \b/n6632 , \b/n6631 , \b/n6630 , \b/n6629 , \b/n6628 , \b/n6627 ,
         \b/n6626 , \b/n6625 , \b/n6624 , \b/n6623 , \b/n6622 , \b/n6621 ,
         \b/n6620 , \b/n6619 , \b/n6618 , \b/n6617 , \b/n6616 , \b/n6615 ,
         \b/n6614 , \b/n6613 , \b/n6612 , \b/n6611 , \b/n6610 , \b/n6609 ,
         \b/n6608 , \b/n6607 , \b/n6606 , \b/n6605 , \b/n6604 , \b/n6603 ,
         \b/n6602 , \b/n6601 , \b/n6600 , \b/n6599 , \b/n6598 , \b/n6597 ,
         \b/n6596 , \b/n6595 , \b/n6594 , \b/n6593 , \b/n6592 , \b/n6591 ,
         \b/n6590 , \b/n6589 , \b/n6588 , \b/n6587 , \b/n6586 , \b/n6585 ,
         \b/n6584 , \b/n6583 , \b/n6582 , \b/n6581 , \b/n6580 , \b/n6579 ,
         \b/n6578 , \b/n6577 , \b/n6576 , \b/n6575 , \b/n6574 , \b/n6573 ,
         \b/n6572 , \b/n6571 , \b/n6570 , \b/n6569 , \b/n6568 , \b/n6567 ,
         \b/n6566 , \b/n6565 , \b/n6564 , \b/n6563 , \b/n6562 , \b/n6561 ,
         \b/n6560 , \b/n6558 , \b/n6557 , \b/n6556 , \b/n6555 , \b/n6554 ,
         \b/n6552 , \b/n6551 , \b/n6550 , \b/n6549 , \b/n6548 , \b/n6547 ,
         \b/n6546 , \b/n6545 , \b/n6544 , \b/n6543 , \b/n6542 , \b/n6540 ,
         \b/n6539 , \b/n6538 , \b/n6536 , \b/n6535 , \b/n6534 , \b/n6533 ,
         \b/n6532 , \b/n6531 , \b/n6530 , \b/n6529 , \b/n6528 , \b/n6527 ,
         \b/n6526 , \b/n6525 , \b/n6524 , \b/n6523 , \b/n6522 , \b/n6521 ,
         \b/n6520 , \b/n6519 , \b/n6518 , \b/n6517 , \b/n6516 , \b/n6515 ,
         \b/n6513 , \b/n6512 , \b/n6511 , \b/n6510 , \b/n6509 , \b/n6508 ,
         \b/n6504 , \b/n6502 , \b/n6501 , \b/n6500 , \b/n6498 , \b/n6495 ,
         \b/n6494 , \b/n6493 , \b/n6492 , \b/n6491 , \b/n6490 , \b/n6489 ,
         \b/n6488 , \b/n6487 , \b/n6486 , \b/n6485 , \b/n6484 , \b/n6483 ,
         \b/n6482 , \b/n6481 , \b/n6480 , \b/n6479 , \b/n6478 , \b/n6477 ,
         \b/n6476 , \b/n6475 , \b/n6474 , \b/n6473 , \b/n6472 , \b/n6471 ,
         \b/n6470 , \b/n6469 , \b/n6468 , \b/n6467 , \b/n6466 , \b/n6465 ,
         \b/n6464 , \b/n6463 , \b/n6462 , \b/n6461 , \b/n6460 , \b/n6459 ,
         \b/n6458 , \b/n6457 , \b/n6456 , \b/n6455 , \b/n6454 , \b/n6453 ,
         \b/n6452 , \b/n6451 , \b/n6450 , \b/n6449 , \b/n6448 , \b/n6447 ,
         \b/n6446 , \b/n6445 , \b/n6444 , \b/n6443 , \b/n6442 , \b/n6441 ,
         \b/n6440 , \b/n6439 , \b/n6438 , \b/n6437 , \b/n6436 , \b/n6435 ,
         \b/n6434 , \b/n6433 , \b/n6432 , \b/n6431 , \b/n6430 , \b/n6429 ,
         \b/n6428 , \b/n6427 , \b/n6426 , \b/n6425 , \b/n6424 , \b/n6423 ,
         \b/n6422 , \b/n6421 , \b/n6420 , \b/n6419 , \b/n6418 , \b/n6417 ,
         \b/n6416 , \b/n6415 , \b/n6414 , \b/n6413 , \b/n6412 , \b/n6411 ,
         \b/n6410 , \b/n6409 , \b/n6408 , \b/n6407 , \b/n6406 , \b/n6405 ,
         \b/n6404 , \b/n6403 , \b/n6402 , \b/n6401 , \b/n6400 , \b/n6399 ,
         \b/n6398 , \b/n6397 , \b/n6396 , \b/n6395 , \b/n6394 , \b/n6393 ,
         \b/n6392 , \b/n6391 , \b/n6390 , \b/n6389 , \b/n6388 , \b/n6387 ,
         \b/n6386 , \b/n6385 , \b/n6384 , \b/n6383 , \b/n6382 , \b/n6381 ,
         \b/n6380 , \b/n6379 , \b/n6378 , \b/n6377 , \b/n6376 , \b/n6375 ,
         \b/n6374 , \b/n6373 , \b/n6372 , \b/n6371 , \b/n6370 , \b/n6369 ,
         \b/n6368 , \b/n6367 , \b/n6366 , \b/n6365 , \b/n6364 , \b/n6363 ,
         \b/n6362 , \b/n6361 , \b/n6360 , \b/n6359 , \b/n6358 , \b/n6357 ,
         \b/n6356 , \b/n6355 , \b/n6354 , \b/n6353 , \b/n6352 , \b/n6351 ,
         \b/n6350 , \b/n6349 , \b/n6348 , \b/n6347 , \b/n6346 , \b/n6345 ,
         \b/n6344 , \b/n6343 , \b/n6342 , \b/n6341 , \b/n6340 , \b/n6339 ,
         \b/n6338 , \b/n6337 , \b/n6336 , \b/n6335 , \b/n6334 , \b/n6333 ,
         \b/n6332 , \b/n6331 , \b/n6330 , \b/n6329 , \b/n6328 , \b/n6327 ,
         \b/n6326 , \b/n6325 , \b/n6324 , \b/n6323 , \b/n6322 , \b/n6321 ,
         \b/n6320 , \b/n6319 , \b/n6318 , \b/n6317 , \b/n6316 , \b/n6315 ,
         \b/n6314 , \b/n6313 , \b/n6312 , \b/n6311 , \b/n6310 , \b/n6309 ,
         \b/n6308 , \b/n6307 , \b/n6306 , \b/n6305 , \b/n6304 , \b/n6303 ,
         \b/n6302 , \b/n6301 , \b/n6300 , \b/n6299 , \b/n6298 , \b/n6297 ,
         \b/n6296 , \b/n6295 , \b/n6294 , \b/n6293 , \b/n6292 , \b/n6291 ,
         \b/n6290 , \b/n6289 , \b/n6288 , \b/n6287 , \b/n6286 , \b/n6285 ,
         \b/n6284 , \b/n6283 , \b/n6282 , \b/n6281 , \b/n6280 , \b/n6279 ,
         \b/n6278 , \b/n6277 , \b/n6276 , \b/n6275 , \b/n6274 , \b/n6273 ,
         \b/n6272 , \b/n6271 , \b/n6270 , \b/n6269 , \b/n6268 , \b/n6267 ,
         \b/n6266 , \b/n6265 , \b/n6264 , \b/n6263 , \b/n6262 , \b/n6261 ,
         \b/n6260 , \b/n6259 , \b/n6258 , \b/n6257 , \b/n6256 , \b/n6255 ,
         \b/n6254 , \b/n6253 , \b/n6252 , \b/n6251 , \b/n6250 , \b/n6249 ,
         \b/n6248 , \b/n6247 , \b/n6246 , \b/n6245 , \b/n6244 , \b/n6243 ,
         \b/n6242 , \b/n6241 , \b/n6240 , \b/n6239 , \b/n6238 , \b/n6237 ,
         \b/n6236 , \b/n6235 , \b/n6234 , \b/n6233 , \b/n6232 , \b/n6231 ,
         \b/n6230 , \b/n6229 , \b/n6228 , \b/n6227 , \b/n6226 , \b/n6225 ,
         \b/n6224 , \b/n6223 , \b/n6222 , \b/n6221 , \b/n6220 , \b/n6219 ,
         \b/n6218 , \b/n6217 , \b/n6216 , \b/n6215 , \b/n6214 , \b/n6213 ,
         \b/n6212 , \b/n6211 , \b/n6210 , \b/n6209 , \b/n6208 , \b/n6207 ,
         \b/n6206 , \b/n6205 , \b/n6204 , \b/n6203 , \b/n6202 , \b/n6201 ,
         \b/n6199 , \b/n6198 , \b/n6197 , \b/n6196 , \b/n6195 , \b/n6193 ,
         \b/n6192 , \b/n6191 , \b/n6190 , \b/n6189 , \b/n6188 , \b/n6187 ,
         \b/n6186 , \b/n6185 , \b/n6184 , \b/n6183 , \b/n6181 , \b/n6180 ,
         \b/n6179 , \b/n6177 , \b/n6176 , \b/n6175 , \b/n6174 , \b/n6173 ,
         \b/n6172 , \b/n6171 , \b/n6170 , \b/n6169 , \b/n6168 , \b/n6167 ,
         \b/n6166 , \b/n6165 , \b/n6164 , \b/n6163 , \b/n6162 , \b/n6161 ,
         \b/n6160 , \b/n6159 , \b/n6158 , \b/n6157 , \b/n6156 , \b/n6154 ,
         \b/n6153 , \b/n6152 , \b/n6151 , \b/n6150 , \b/n6149 , \b/n6145 ,
         \b/n6143 , \b/n6142 , \b/n6141 , \b/n6139 , \b/n6136 , \b/n6135 ,
         \b/n6134 , \b/n6133 , \b/n6132 , \b/n6131 , \b/n6130 , \b/n6129 ,
         \b/n6128 , \b/n6127 , \b/n6126 , \b/n6125 , \b/n6124 , \b/n6123 ,
         \b/n6122 , \b/n6121 , \b/n6120 , \b/n6119 , \b/n6118 , \b/n6117 ,
         \b/n6116 , \b/n6115 , \b/n6114 , \b/n6113 , \b/n6112 , \b/n6111 ,
         \b/n6110 , \b/n6109 , \b/n6108 , \b/n6107 , \b/n6106 , \b/n6105 ,
         \b/n6104 , \b/n6103 , \b/n6102 , \b/n6101 , \b/n6100 , \b/n6099 ,
         \b/n6098 , \b/n6097 , \b/n6096 , \b/n6095 , \b/n6094 , \b/n6093 ,
         \b/n6092 , \b/n6091 , \b/n6090 , \b/n6089 , \b/n6088 , \b/n6087 ,
         \b/n6086 , \b/n6085 , \b/n6084 , \b/n6083 , \b/n6082 , \b/n6081 ,
         \b/n6080 , \b/n6079 , \b/n6078 , \b/n6077 , \b/n6076 , \b/n6075 ,
         \b/n6074 , \b/n6073 , \b/n6072 , \b/n6071 , \b/n6070 , \b/n6069 ,
         \b/n6068 , \b/n6067 , \b/n6066 , \b/n6065 , \b/n6064 , \b/n6063 ,
         \b/n6062 , \b/n6061 , \b/n6060 , \b/n6059 , \b/n6058 , \b/n6057 ,
         \b/n6056 , \b/n6055 , \b/n6054 , \b/n6053 , \b/n6052 , \b/n6051 ,
         \b/n6050 , \b/n6049 , \b/n6048 , \b/n6047 , \b/n6046 , \b/n6045 ,
         \b/n6044 , \b/n6043 , \b/n6042 , \b/n6041 , \b/n6040 , \b/n6039 ,
         \b/n6038 , \b/n6037 , \b/n6036 , \b/n6035 , \b/n6034 , \b/n6033 ,
         \b/n6032 , \b/n6031 , \b/n6030 , \b/n6029 , \b/n6028 , \b/n6027 ,
         \b/n6026 , \b/n6025 , \b/n6024 , \b/n6023 , \b/n6022 , \b/n6021 ,
         \b/n6020 , \b/n6019 , \b/n6018 , \b/n6017 , \b/n6016 , \b/n6015 ,
         \b/n6014 , \b/n6013 , \b/n6012 , \b/n6011 , \b/n6010 , \b/n6009 ,
         \b/n6008 , \b/n6007 , \b/n6006 , \b/n6005 , \b/n6004 , \b/n6003 ,
         \b/n6002 , \b/n6001 , \b/n6000 , \b/n5999 , \b/n5998 , \b/n5997 ,
         \b/n5996 , \b/n5995 , \b/n5994 , \b/n5993 , \b/n5992 , \b/n5991 ,
         \b/n5990 , \b/n5989 , \b/n5988 , \b/n5987 , \b/n5986 , \b/n5985 ,
         \b/n5984 , \b/n5983 , \b/n5982 , \b/n5981 , \b/n5980 , \b/n5979 ,
         \b/n5978 , \b/n5977 , \b/n5976 , \b/n5975 , \b/n5974 , \b/n5973 ,
         \b/n5972 , \b/n5971 , \b/n5970 , \b/n5969 , \b/n5968 , \b/n5967 ,
         \b/n5966 , \b/n5965 , \b/n5964 , \b/n5963 , \b/n5962 , \b/n5961 ,
         \b/n5960 , \b/n5959 , \b/n5958 , \b/n5957 , \b/n5956 , \b/n5955 ,
         \b/n5954 , \b/n5953 , \b/n5952 , \b/n5951 , \b/n5950 , \b/n5949 ,
         \b/n5948 , \b/n5947 , \b/n5946 , \b/n5945 , \b/n5944 , \b/n5943 ,
         \b/n5942 , \b/n5941 , \b/n5940 , \b/n5939 , \b/n5938 , \b/n5937 ,
         \b/n5936 , \b/n5935 , \b/n5934 , \b/n5933 , \b/n5932 , \b/n5931 ,
         \b/n5930 , \b/n5929 , \b/n5928 , \b/n5927 , \b/n5926 , \b/n5925 ,
         \b/n5924 , \b/n5923 , \b/n5922 , \b/n5921 , \b/n5920 , \b/n5919 ,
         \b/n5918 , \b/n5917 , \b/n5916 , \b/n5915 , \b/n5914 , \b/n5913 ,
         \b/n5912 , \b/n5911 , \b/n5910 , \b/n5909 , \b/n5908 , \b/n5907 ,
         \b/n5906 , \b/n5905 , \b/n5904 , \b/n5903 , \b/n5902 , \b/n5901 ,
         \b/n5900 , \b/n5899 , \b/n5898 , \b/n5897 , \b/n5896 , \b/n5895 ,
         \b/n5894 , \b/n5893 , \b/n5892 , \b/n5891 , \b/n5890 , \b/n5889 ,
         \b/n5888 , \b/n5887 , \b/n5886 , \b/n5885 , \b/n5884 , \b/n5883 ,
         \b/n5882 , \b/n5881 , \b/n5880 , \b/n5879 , \b/n5878 , \b/n5877 ,
         \b/n5876 , \b/n5875 , \b/n5874 , \b/n5873 , \b/n5872 , \b/n5871 ,
         \b/n5870 , \b/n5869 , \b/n5868 , \b/n5867 , \b/n5866 , \b/n5865 ,
         \b/n5864 , \b/n5863 , \b/n5862 , \b/n5861 , \b/n5860 , \b/n5859 ,
         \b/n5858 , \b/n5857 , \b/n5856 , \b/n5855 , \b/n5854 , \b/n5853 ,
         \b/n5852 , \b/n5851 , \b/n5850 , \b/n5849 , \b/n5848 , \b/n5847 ,
         \b/n5846 , \b/n5845 , \b/n5844 , \b/n5843 , \b/n5842 , \b/n5840 ,
         \b/n5839 , \b/n5838 , \b/n5837 , \b/n5836 , \b/n5834 , \b/n5833 ,
         \b/n5832 , \b/n5831 , \b/n5830 , \b/n5829 , \b/n5828 , \b/n5827 ,
         \b/n5826 , \b/n5825 , \b/n5824 , \b/n5822 , \b/n5821 , \b/n5820 ,
         \b/n5818 , \b/n5817 , \b/n5816 , \b/n5815 , \b/n5814 , \b/n5813 ,
         \b/n5812 , \b/n5811 , \b/n5810 , \b/n5809 , \b/n5808 , \b/n5807 ,
         \b/n5806 , \b/n5805 , \b/n5804 , \b/n5803 , \b/n5802 , \b/n5801 ,
         \b/n5800 , \b/n5799 , \b/n5798 , \b/n5797 , \b/n5795 , \b/n5794 ,
         \b/n5793 , \b/n5792 , \b/n5791 , \b/n5790 , \b/n5786 , \b/n5785 ,
         \b/n5783 , \b/n5782 , \b/n5779 , \b/n5777 , \b/n5776 , \b/n5775 ,
         \b/n5774 , \b/n5773 , \b/n5772 , \b/n5771 , \b/n5770 , \b/n5769 ,
         \b/n5768 , \b/n5767 , \b/n5766 , \b/n5765 , \b/n5764 , \b/n5763 ,
         \b/n5762 , \b/n5761 , \b/n5760 , \b/n5759 , \b/n5758 , \b/n5757 ,
         \b/n5756 , \b/n5755 , \b/n5754 , \b/n5753 , \b/n5752 , \b/n5751 ,
         \b/n5750 , \b/n5749 , \b/n5748 , \b/n5747 , \b/n5746 , \b/n5745 ,
         \b/n5744 , \b/n5743 , \b/n5742 , \b/n5741 , \b/n5740 , \b/n5739 ,
         \b/n5738 , \b/n5737 , \b/n5736 , \b/n5735 , \b/n5734 , \b/n5733 ,
         \b/n5732 , \b/n5731 , \b/n5730 , \b/n5729 , \b/n5728 , \b/n5727 ,
         \b/n5726 , \b/n5725 , \b/n5724 , \b/n5723 , \b/n5722 , \b/n5721 ,
         \b/n5720 , \b/n5719 , \b/n5718 , \b/n5717 , \b/n5716 , \b/n5715 ,
         \b/n5714 , \b/n5713 , \b/n5712 , \b/n5711 , \b/n5710 , \b/n5709 ,
         \b/n5708 , \b/n5707 , \b/n5706 , \b/n5705 , \b/n5704 , \b/n5703 ,
         \b/n5702 , \b/n5701 , \b/n5700 , \b/n5699 , \b/n5698 , \b/n5697 ,
         \b/n5696 , \b/n5695 , \b/n5694 , \b/n5693 , \b/n5692 , \b/n5691 ,
         \b/n5690 , \b/n5689 , \b/n5688 , \b/n5687 , \b/n5686 , \b/n5685 ,
         \b/n5684 , \b/n5683 , \b/n5682 , \b/n5681 , \b/n5680 , \b/n5679 ,
         \b/n5678 , \b/n5677 , \b/n5676 , \b/n5675 , \b/n5674 , \b/n5673 ,
         \b/n5672 , \b/n5671 , \b/n5670 , \b/n5669 , \b/n5668 , \b/n5667 ,
         \b/n5666 , \b/n5665 , \b/n5664 , \b/n5663 , \b/n5662 , \b/n5661 ,
         \b/n5660 , \b/n5659 , \b/n5658 , \b/n5657 , \b/n5656 , \b/n5655 ,
         \b/n5654 , \b/n5653 , \b/n5652 , \b/n5651 , \b/n5650 , \b/n5649 ,
         \b/n5648 , \b/n5647 , \b/n5646 , \b/n5645 , \b/n5644 , \b/n5643 ,
         \b/n5642 , \b/n5641 , \b/n5640 , \b/n5639 , \b/n5638 , \b/n5637 ,
         \b/n5636 , \b/n5635 , \b/n5634 , \b/n5633 , \b/n5632 , \b/n5631 ,
         \b/n5630 , \b/n5629 , \b/n5628 , \b/n5627 , \b/n5626 , \b/n5625 ,
         \b/n5624 , \b/n5623 , \b/n5622 , \b/n5621 , \b/n5620 , \b/n5619 ,
         \b/n5618 , \b/n5617 , \b/n5616 , \b/n5615 , \b/n5614 , \b/n5613 ,
         \b/n5612 , \b/n5611 , \b/n5610 , \b/n5609 , \b/n5608 , \b/n5607 ,
         \b/n5606 , \b/n5605 , \b/n5604 , \b/n5603 , \b/n5602 , \b/n5601 ,
         \b/n5600 , \b/n5599 , \b/n5598 , \b/n5597 , \b/n5596 , \b/n5595 ,
         \b/n5594 , \b/n5593 , \b/n5592 , \b/n5591 , \b/n5590 , \b/n5589 ,
         \b/n5588 , \b/n5587 , \b/n5586 , \b/n5585 , \b/n5584 , \b/n5583 ,
         \b/n5582 , \b/n5581 , \b/n5580 , \b/n5579 , \b/n5578 , \b/n5577 ,
         \b/n5576 , \b/n5575 , \b/n5574 , \b/n5573 , \b/n5572 , \b/n5571 ,
         \b/n5570 , \b/n5569 , \b/n5568 , \b/n5567 , \b/n5566 , \b/n5565 ,
         \b/n5564 , \b/n5563 , \b/n5562 , \b/n5561 , \b/n5560 , \b/n5559 ,
         \b/n5558 , \b/n5557 , \b/n5556 , \b/n5555 , \b/n5554 , \b/n5553 ,
         \b/n5552 , \b/n5551 , \b/n5550 , \b/n5549 , \b/n5548 , \b/n5547 ,
         \b/n5546 , \b/n5545 , \b/n5544 , \b/n5543 , \b/n5542 , \b/n5541 ,
         \b/n5540 , \b/n5539 , \b/n5538 , \b/n5537 , \b/n5536 , \b/n5535 ,
         \b/n5534 , \b/n5533 , \b/n5532 , \b/n5531 , \b/n5530 , \b/n5529 ,
         \b/n5528 , \b/n5527 , \b/n5526 , \b/n5525 , \b/n5524 , \b/n5523 ,
         \b/n5522 , \b/n5521 , \b/n5520 , \b/n5519 , \b/n5518 , \b/n5517 ,
         \b/n5516 , \b/n5515 , \b/n5514 , \b/n5513 , \b/n5512 , \b/n5511 ,
         \b/n5510 , \b/n5509 , \b/n5508 , \b/n5507 , \b/n5506 , \b/n5505 ,
         \b/n5504 , \b/n5503 , \b/n5502 , \b/n5501 , \b/n5500 , \b/n5499 ,
         \b/n5498 , \b/n5497 , \b/n5496 , \b/n5495 , \b/n5494 , \b/n5493 ,
         \b/n5492 , \b/n5491 , \b/n5490 , \b/n5489 , \b/n5488 , \b/n5487 ,
         \b/n5486 , \b/n5485 , \b/n5483 , \b/n5482 , \b/n5481 , \b/n5480 ,
         \b/n5479 , \b/n5478 , \b/n5476 , \b/n5475 , \b/n5474 , \b/n5473 ,
         \b/n5472 , \b/n5471 , \b/n5470 , \b/n5469 , \b/n5468 , \b/n5467 ,
         \b/n5466 , \b/n5464 , \b/n5463 , \b/n5462 , \b/n5461 , \b/n5460 ,
         \b/n5459 , \b/n5458 , \b/n5457 , \b/n5456 , \b/n5454 , \b/n5453 ,
         \b/n5452 , \b/n5451 , \b/n5450 , \b/n5449 , \b/n5448 , \b/n5447 ,
         \b/n5446 , \b/n5445 , \b/n5444 , \b/n5443 , \b/n5442 , \b/n5441 ,
         \b/n5440 , \b/n5439 , \b/n5437 , \b/n5436 , \b/n5435 , \b/n5434 ,
         \b/n5433 , \b/n5432 , \b/n5428 , \b/n5426 , \b/n5425 , \b/n5424 ,
         \b/n5422 , \b/n5419 , \b/n5418 , \b/n5417 , \b/n5416 , \b/n5415 ,
         \b/n5414 , \b/n5413 , \b/n5412 , \b/n5411 , \b/n5410 , \b/n5409 ,
         \b/n5408 , \b/n5407 , \b/n5406 , \b/n5405 , \b/n5404 , \b/n5403 ,
         \b/n5402 , \b/n5401 , \b/n5400 , \b/n5399 , \b/n5398 , \b/n5397 ,
         \b/n5396 , \b/n5395 , \b/n5394 , \b/n5393 , \b/n5392 , \b/n5391 ,
         \b/n5390 , \b/n5389 , \b/n5388 , \b/n5387 , \b/n5386 , \b/n5385 ,
         \b/n5384 , \b/n5383 , \b/n5382 , \b/n5381 , \b/n5380 , \b/n5379 ,
         \b/n5378 , \b/n5377 , \b/n5376 , \b/n5375 , \b/n5374 , \b/n5373 ,
         \b/n5372 , \b/n5371 , \b/n5370 , \b/n5369 , \b/n5368 , \b/n5367 ,
         \b/n5366 , \b/n5365 , \b/n5364 , \b/n5363 , \b/n5362 , \b/n5361 ,
         \b/n5360 , \b/n5359 , \b/n5358 , \b/n5357 , \b/n5356 , \b/n5355 ,
         \b/n5354 , \b/n5353 , \b/n5352 , \b/n5351 , \b/n5350 , \b/n5349 ,
         \b/n5348 , \b/n5347 , \b/n5346 , \b/n5345 , \b/n5344 , \b/n5343 ,
         \b/n5342 , \b/n5341 , \b/n5340 , \b/n5339 , \b/n5338 , \b/n5337 ,
         \b/n5336 , \b/n5335 , \b/n5334 , \b/n5333 , \b/n5332 , \b/n5331 ,
         \b/n5330 , \b/n5329 , \b/n5328 , \b/n5327 , \b/n5326 , \b/n5325 ,
         \b/n5324 , \b/n5323 , \b/n5322 , \b/n5321 , \b/n5320 , \b/n5319 ,
         \b/n5318 , \b/n5317 , \b/n5316 , \b/n5315 , \b/n5314 , \b/n5313 ,
         \b/n5312 , \b/n5311 , \b/n5310 , \b/n5309 , \b/n5308 , \b/n5307 ,
         \b/n5306 , \b/n5305 , \b/n5304 , \b/n5303 , \b/n5302 , \b/n5301 ,
         \b/n5300 , \b/n5299 , \b/n5298 , \b/n5297 , \b/n5296 , \b/n5295 ,
         \b/n5294 , \b/n5293 , \b/n5292 , \b/n5291 , \b/n5290 , \b/n5289 ,
         \b/n5288 , \b/n5287 , \b/n5286 , \b/n5285 , \b/n5284 , \b/n5283 ,
         \b/n5282 , \b/n5281 , \b/n5280 , \b/n5279 , \b/n5278 , \b/n5277 ,
         \b/n5276 , \b/n5275 , \b/n5274 , \b/n5273 , \b/n5272 , \b/n5271 ,
         \b/n5270 , \b/n5269 , \b/n5268 , \b/n5267 , \b/n5266 , \b/n5265 ,
         \b/n5264 , \b/n5263 , \b/n5262 , \b/n5261 , \b/n5260 , \b/n5259 ,
         \b/n5258 , \b/n5257 , \b/n5256 , \b/n5255 , \b/n5254 , \b/n5253 ,
         \b/n5252 , \b/n5251 , \b/n5250 , \b/n5249 , \b/n5248 , \b/n5247 ,
         \b/n5246 , \b/n5245 , \b/n5244 , \b/n5243 , \b/n5242 , \b/n5241 ,
         \b/n5240 , \b/n5239 , \b/n5238 , \b/n5237 , \b/n5236 , \b/n5235 ,
         \b/n5234 , \b/n5233 , \b/n5232 , \b/n5231 , \b/n5230 , \b/n5229 ,
         \b/n5228 , \b/n5227 , \b/n5226 , \b/n5225 , \b/n5224 , \b/n5223 ,
         \b/n5222 , \b/n5221 , \b/n5220 , \b/n5219 , \b/n5218 , \b/n5217 ,
         \b/n5216 , \b/n5215 , \b/n5214 , \b/n5213 , \b/n5212 , \b/n5211 ,
         \b/n5210 , \b/n5209 , \b/n5208 , \b/n5207 , \b/n5206 , \b/n5205 ,
         \b/n5204 , \b/n5203 , \b/n5202 , \b/n5201 , \b/n5200 , \b/n5199 ,
         \b/n5198 , \b/n5197 , \b/n5196 , \b/n5195 , \b/n5194 , \b/n5193 ,
         \b/n5192 , \b/n5191 , \b/n5190 , \b/n5189 , \b/n5188 , \b/n5187 ,
         \b/n5186 , \b/n5185 , \b/n5184 , \b/n5183 , \b/n5182 , \b/n5181 ,
         \b/n5180 , \b/n5179 , \b/n5178 , \b/n5177 , \b/n5176 , \b/n5175 ,
         \b/n5174 , \b/n5173 , \b/n5172 , \b/n5171 , \b/n5170 , \b/n5169 ,
         \b/n5168 , \b/n5167 , \b/n5166 , \b/n5165 , \b/n5164 , \b/n5163 ,
         \b/n5162 , \b/n5161 , \b/n5160 , \b/n5159 , \b/n5158 , \b/n5157 ,
         \b/n5156 , \b/n5155 , \b/n5154 , \b/n5153 , \b/n5152 , \b/n5151 ,
         \b/n5150 , \b/n5149 , \b/n5148 , \b/n5147 , \b/n5146 , \b/n5145 ,
         \b/n5144 , \b/n5143 , \b/n5142 , \b/n5141 , \b/n5140 , \b/n5139 ,
         \b/n5138 , \b/n5137 , \b/n5136 , \b/n5135 , \b/n5134 , \b/n5133 ,
         \b/n5132 , \b/n5131 , \b/n5130 , \b/n5129 , \b/n5128 , \b/n5127 ,
         \b/n5126 , \b/n5125 , \b/n5123 , \b/n5122 , \b/n5121 , \b/n5120 ,
         \b/n5119 , \b/n5117 , \b/n5116 , \b/n5115 , \b/n5114 , \b/n5113 ,
         \b/n5112 , \b/n5111 , \b/n5110 , \b/n5109 , \b/n5108 , \b/n5107 ,
         \b/n5105 , \b/n5104 , \b/n5103 , \b/n5101 , \b/n5100 , \b/n5099 ,
         \b/n5098 , \b/n5097 , \b/n5096 , \b/n5095 , \b/n5094 , \b/n5093 ,
         \b/n5092 , \b/n5091 , \b/n5090 , \b/n5089 , \b/n5088 , \b/n5087 ,
         \b/n5086 , \b/n5085 , \b/n5084 , \b/n5083 , \b/n5082 , \b/n5081 ,
         \b/n5080 , \b/n5078 , \b/n5077 , \b/n5076 , \b/n5075 , \b/n5074 ,
         \b/n5073 , \b/n5069 , \b/n5067 , \b/n5066 , \b/n5065 , \b/n5063 ,
         \b/n5060 , \b/n5059 , \b/n5058 , \b/n5057 , \b/n5056 , \b/n5055 ,
         \b/n5054 , \b/n5053 , \b/n5052 , \b/n5051 , \b/n5050 , \b/n5049 ,
         \b/n5048 , \b/n5047 , \b/n5046 , \b/n5045 , \b/n5044 , \b/n5043 ,
         \b/n5042 , \b/n5041 , \b/n5040 , \b/n5039 , \b/n5038 , \b/n5037 ,
         \b/n5036 , \b/n5035 , \b/n5034 , \b/n5033 , \b/n5032 , \b/n5031 ,
         \b/n5030 , \b/n5029 , \b/n5028 , \b/n5027 , \b/n5026 , \b/n5025 ,
         \b/n5024 , \b/n5023 , \b/n5022 , \b/n5021 , \b/n5020 , \b/n5019 ,
         \b/n5018 , \b/n5017 , \b/n5016 , \b/n5015 , \b/n5014 , \b/n5013 ,
         \b/n5012 , \b/n5011 , \b/n5010 , \b/n5009 , \b/n5008 , \b/n5007 ,
         \b/n5006 , \b/n5005 , \b/n5004 , \b/n5003 , \b/n5002 , \b/n5001 ,
         \b/n5000 , \b/n4999 , \b/n4998 , \b/n4997 , \b/n4996 , \b/n4995 ,
         \b/n4994 , \b/n4993 , \b/n4992 , \b/n4991 , \b/n4990 , \b/n4989 ,
         \b/n4988 , \b/n4987 , \b/n4986 , \b/n4985 , \b/n4984 , \b/n4983 ,
         \b/n4982 , \b/n4981 , \b/n4980 , \b/n4979 , \b/n4978 , \b/n4977 ,
         \b/n4976 , \b/n4975 , \b/n4974 , \b/n4973 , \b/n4972 , \b/n4971 ,
         \b/n4970 , \b/n4969 , \b/n4968 , \b/n4967 , \b/n4966 , \b/n4965 ,
         \b/n4964 , \b/n4963 , \b/n4962 , \b/n4961 , \b/n4960 , \b/n4959 ,
         \b/n4958 , \b/n4957 , \b/n4956 , \b/n4955 , \b/n4954 , \b/n4953 ,
         \b/n4952 , \b/n4951 , \b/n4950 , \b/n4949 , \b/n4948 , \b/n4947 ,
         \b/n4946 , \b/n4945 , \b/n4944 , \b/n4943 , \b/n4942 , \b/n4941 ,
         \b/n4940 , \b/n4939 , \b/n4938 , \b/n4937 , \b/n4936 , \b/n4935 ,
         \b/n4934 , \b/n4933 , \b/n4932 , \b/n4931 , \b/n4930 , \b/n4929 ,
         \b/n4928 , \b/n4927 , \b/n4926 , \b/n4925 , \b/n4924 , \b/n4923 ,
         \b/n4922 , \b/n4921 , \b/n4920 , \b/n4919 , \b/n4918 , \b/n4917 ,
         \b/n4916 , \b/n4915 , \b/n4914 , \b/n4913 , \b/n4912 , \b/n4911 ,
         \b/n4910 , \b/n4909 , \b/n4908 , \b/n4907 , \b/n4906 , \b/n4905 ,
         \b/n4904 , \b/n4903 , \b/n4902 , \b/n4901 , \b/n4900 , \b/n4899 ,
         \b/n4898 , \b/n4897 , \b/n4896 , \b/n4895 , \b/n4894 , \b/n4893 ,
         \b/n4892 , \b/n4891 , \b/n4890 , \b/n4889 , \b/n4888 , \b/n4887 ,
         \b/n4886 , \b/n4885 , \b/n4884 , \b/n4883 , \b/n4882 , \b/n4881 ,
         \b/n4880 , \b/n4879 , \b/n4878 , \b/n4877 , \b/n4876 , \b/n4875 ,
         \b/n4874 , \b/n4873 , \b/n4872 , \b/n4871 , \b/n4870 , \b/n4869 ,
         \b/n4868 , \b/n4867 , \b/n4866 , \b/n4865 , \b/n4864 , \b/n4863 ,
         \b/n4862 , \b/n4861 , \b/n4860 , \b/n4859 , \b/n4858 , \b/n4857 ,
         \b/n4856 , \b/n4855 , \b/n4854 , \b/n4853 , \b/n4852 , \b/n4851 ,
         \b/n4850 , \b/n4849 , \b/n4848 , \b/n4847 , \b/n4846 , \b/n4845 ,
         \b/n4844 , \b/n4843 , \b/n4842 , \b/n4841 , \b/n4840 , \b/n4839 ,
         \b/n4838 , \b/n4837 , \b/n4836 , \b/n4835 , \b/n4834 , \b/n4833 ,
         \b/n4832 , \b/n4831 , \b/n4830 , \b/n4829 , \b/n4828 , \b/n4827 ,
         \b/n4826 , \b/n4825 , \b/n4824 , \b/n4823 , \b/n4822 , \b/n4821 ,
         \b/n4820 , \b/n4819 , \b/n4818 , \b/n4817 , \b/n4816 , \b/n4815 ,
         \b/n4814 , \b/n4813 , \b/n4812 , \b/n4811 , \b/n4810 , \b/n4809 ,
         \b/n4808 , \b/n4807 , \b/n4806 , \b/n4805 , \b/n4804 , \b/n4803 ,
         \b/n4802 , \b/n4801 , \b/n4800 , \b/n4799 , \b/n4798 , \b/n4797 ,
         \b/n4796 , \b/n4795 , \b/n4794 , \b/n4793 , \b/n4792 , \b/n4791 ,
         \b/n4790 , \b/n4789 , \b/n4788 , \b/n4787 , \b/n4786 , \b/n4785 ,
         \b/n4784 , \b/n4783 , \b/n4782 , \b/n4781 , \b/n4780 , \b/n4779 ,
         \b/n4778 , \b/n4777 , \b/n4776 , \b/n4775 , \b/n4774 , \b/n4773 ,
         \b/n4772 , \b/n4771 , \b/n4770 , \b/n4769 , \b/n4768 , \b/n4767 ,
         \b/n4766 , \b/n4764 , \b/n4763 , \b/n4762 , \b/n4761 , \b/n4760 ,
         \b/n4758 , \b/n4757 , \b/n4756 , \b/n4755 , \b/n4754 , \b/n4753 ,
         \b/n4752 , \b/n4751 , \b/n4750 , \b/n4749 , \b/n4748 , \b/n4746 ,
         \b/n4745 , \b/n4744 , \b/n4742 , \b/n4741 , \b/n4740 , \b/n4739 ,
         \b/n4738 , \b/n4737 , \b/n4736 , \b/n4735 , \b/n4734 , \b/n4733 ,
         \b/n4732 , \b/n4731 , \b/n4730 , \b/n4729 , \b/n4728 , \b/n4727 ,
         \b/n4726 , \b/n4725 , \b/n4724 , \b/n4723 , \b/n4722 , \b/n4721 ,
         \b/n4719 , \b/n4718 , \b/n4717 , \b/n4716 , \b/n4715 , \b/n4714 ,
         \b/n4710 , \b/n4708 , \b/n4707 , \b/n4706 , \b/n4704 , \b/n4701 ,
         \b/n4700 , \b/n4699 , \b/n4698 , \b/n4697 , \b/n4696 , \b/n4695 ,
         \b/n4694 , \b/n4693 , \b/n4692 , \b/n4691 , \b/n4690 , \b/n4689 ,
         \b/n4688 , \b/n4687 , \b/n4686 , \b/n4685 , \b/n4684 , \b/n4683 ,
         \b/n4682 , \b/n4681 , \b/n4680 , \b/n4679 , \b/n4678 , \b/n4677 ,
         \b/n4676 , \b/n4675 , \b/n4674 , \b/n4673 , \b/n4672 , \b/n4671 ,
         \b/n4670 , \b/n4669 , \b/n4668 , \b/n4667 , \b/n4666 , \b/n4665 ,
         \b/n4664 , \b/n4663 , \b/n4662 , \b/n4661 , \b/n4660 , \b/n4659 ,
         \b/n4658 , \b/n4657 , \b/n4656 , \b/n4655 , \b/n4654 , \b/n4653 ,
         \b/n4652 , \b/n4651 , \b/n4650 , \b/n4649 , \b/n4648 , \b/n4647 ,
         \b/n4646 , \b/n4645 , \b/n4644 , \b/n4643 , \b/n4642 , \b/n4641 ,
         \b/n4640 , \b/n4639 , \b/n4638 , \b/n4637 , \b/n4636 , \b/n4635 ,
         \b/n4634 , \b/n4633 , \b/n4632 , \b/n4631 , \b/n4630 , \b/n4629 ,
         \b/n4628 , \b/n4627 , \b/n4626 , \b/n4625 , \b/n4624 , \b/n4623 ,
         \b/n4622 , \b/n4621 , \b/n4620 , \b/n4619 , \b/n4618 , \b/n4617 ,
         \b/n4616 , \b/n4615 , \b/n4614 , \b/n4613 , \b/n4612 , \b/n4611 ,
         \b/n4610 , \b/n4609 , \b/n4608 , \b/n4607 , \b/n4606 , \b/n4605 ,
         \b/n4604 , \b/n4603 , \b/n4602 , \b/n4601 , \b/n4600 , \b/n4599 ,
         \b/n4598 , \b/n4597 , \b/n4596 , \b/n4595 , \b/n4594 , \b/n4593 ,
         \b/n4592 , \b/n4591 , \b/n4590 , \b/n4589 , \b/n4588 , \b/n4587 ,
         \b/n4586 , \b/n4585 , \b/n4584 , \b/n4583 , \b/n4582 , \b/n4581 ,
         \b/n4580 , \b/n4579 , \b/n4578 , \b/n4577 , \b/n4576 , \b/n4575 ,
         \b/n4574 , \b/n4573 , \b/n4572 , \b/n4571 , \b/n4570 , \b/n4569 ,
         \b/n4568 , \b/n4567 , \b/n4566 , \b/n4565 , \b/n4564 , \b/n4563 ,
         \b/n4562 , \b/n4561 , \b/n4560 , \b/n4559 , \b/n4558 , \b/n4557 ,
         \b/n4556 , \b/n4555 , \b/n4554 , \b/n4553 , \b/n4552 , \b/n4551 ,
         \b/n4550 , \b/n4549 , \b/n4548 , \b/n4547 , \b/n4546 , \b/n4545 ,
         \b/n4544 , \b/n4543 , \b/n4542 , \b/n4541 , \b/n4540 , \b/n4539 ,
         \b/n4538 , \b/n4537 , \b/n4536 , \b/n4535 , \b/n4534 , \b/n4533 ,
         \b/n4532 , \b/n4531 , \b/n4530 , \b/n4529 , \b/n4528 , \b/n4527 ,
         \b/n4526 , \b/n4525 , \b/n4524 , \b/n4523 , \b/n4522 , \b/n4521 ,
         \b/n4520 , \b/n4519 , \b/n4518 , \b/n4517 , \b/n4516 , \b/n4515 ,
         \b/n4514 , \b/n4513 , \b/n4512 , \b/n4511 , \b/n4510 , \b/n4509 ,
         \b/n4508 , \b/n4507 , \b/n4506 , \b/n4505 , \b/n4504 , \b/n4503 ,
         \b/n4502 , \b/n4501 , \b/n4500 , \b/n4499 , \b/n4498 , \b/n4497 ,
         \b/n4496 , \b/n4495 , \b/n4494 , \b/n4493 , \b/n4492 , \b/n4491 ,
         \b/n4490 , \b/n4489 , \b/n4488 , \b/n4487 , \b/n4486 , \b/n4485 ,
         \b/n4484 , \b/n4483 , \b/n4482 , \b/n4481 , \b/n4480 , \b/n4479 ,
         \b/n4478 , \b/n4477 , \b/n4476 , \b/n4475 , \b/n4474 , \b/n4473 ,
         \b/n4472 , \b/n4471 , \b/n4470 , \b/n4469 , \b/n4468 , \b/n4467 ,
         \b/n4466 , \b/n4465 , \b/n4464 , \b/n4463 , \b/n4462 , \b/n4461 ,
         \b/n4460 , \b/n4459 , \b/n4458 , \b/n4457 , \b/n4456 , \b/n4455 ,
         \b/n4454 , \b/n4453 , \b/n4452 , \b/n4451 , \b/n4450 , \b/n4449 ,
         \b/n4448 , \b/n4447 , \b/n4446 , \b/n4445 , \b/n4444 , \b/n4443 ,
         \b/n4442 , \b/n4441 , \b/n4440 , \b/n4439 , \b/n4438 , \b/n4437 ,
         \b/n4436 , \b/n4435 , \b/n4434 , \b/n4433 , \b/n4432 , \b/n4431 ,
         \b/n4430 , \b/n4429 , \b/n4428 , \b/n4427 , \b/n4426 , \b/n4425 ,
         \b/n4424 , \b/n4423 , \b/n4422 , \b/n4421 , \b/n4420 , \b/n4419 ,
         \b/n4418 , \b/n4417 , \b/n4416 , \b/n4415 , \b/n4414 , \b/n4413 ,
         \b/n4412 , \b/n4411 , \b/n4410 , \b/n4409 , \b/n4408 , \b/n4407 ,
         \b/n4405 , \b/n4404 , \b/n4403 , \b/n4402 , \b/n4401 , \b/n4399 ,
         \b/n4398 , \b/n4397 , \b/n4396 , \b/n4395 , \b/n4394 , \b/n4393 ,
         \b/n4392 , \b/n4391 , \b/n4390 , \b/n4389 , \b/n4387 , \b/n4386 ,
         \b/n4385 , \b/n4383 , \b/n4382 , \b/n4381 , \b/n4380 , \b/n4379 ,
         \b/n4378 , \b/n4377 , \b/n4376 , \b/n4375 , \b/n4374 , \b/n4373 ,
         \b/n4372 , \b/n4371 , \b/n4370 , \b/n4369 , \b/n4368 , \b/n4367 ,
         \b/n4366 , \b/n4365 , \b/n4364 , \b/n4363 , \b/n4362 , \b/n4360 ,
         \b/n4359 , \b/n4358 , \b/n4357 , \b/n4356 , \b/n4355 , \b/n4351 ,
         \b/n4349 , \b/n4348 , \b/n4347 , \b/n4345 , \b/n4342 , \b/n4341 ,
         \b/n4340 , \b/n4339 , \b/n4338 , \b/n4337 , \b/n4336 , \b/n4335 ,
         \b/n4334 , \b/n4333 , \b/n4332 , \b/n4331 , \b/n4330 , \b/n4329 ,
         \b/n4328 , \b/n4327 , \b/n4326 , \b/n4325 , \b/n4324 , \b/n4323 ,
         \b/n4322 , \b/n4321 , \b/n4320 , \b/n4319 , \b/n4318 , \b/n4317 ,
         \b/n4316 , \b/n4315 , \b/n4314 , \b/n4313 , \b/n4312 , \b/n4311 ,
         \b/n4310 , \b/n4309 , \b/n4308 , \b/n4307 , \b/n4306 , \b/n4305 ,
         \b/n4304 , \b/n4303 , \b/n4302 , \b/n4301 , \b/n4300 , \b/n4299 ,
         \b/n4298 , \b/n4297 , \b/n4296 , \b/n4295 , \b/n4294 , \b/n4293 ,
         \b/n4292 , \b/n4291 , \b/n4290 , \b/n4289 , \b/n4288 , \b/n4287 ,
         \b/n4286 , \b/n4285 , \b/n4284 , \b/n4283 , \b/n4282 , \b/n4281 ,
         \b/n4280 , \b/n4279 , \b/n4278 , \b/n4277 , \b/n4276 , \b/n4275 ,
         \b/n4274 , \b/n4273 , \b/n4272 , \b/n4271 , \b/n4270 , \b/n4269 ,
         \b/n4268 , \b/n4267 , \b/n4266 , \b/n4265 , \b/n4264 , \b/n4263 ,
         \b/n4262 , \b/n4261 , \b/n4260 , \b/n4259 , \b/n4258 , \b/n4257 ,
         \b/n4256 , \b/n4255 , \b/n4254 , \b/n4253 , \b/n4252 , \b/n4251 ,
         \b/n4250 , \b/n4249 , \b/n4248 , \b/n4247 , \b/n4246 , \b/n4245 ,
         \b/n4244 , \b/n4243 , \b/n4242 , \b/n4241 , \b/n4240 , \b/n4239 ,
         \b/n4238 , \b/n4237 , \b/n4236 , \b/n4235 , \b/n4234 , \b/n4233 ,
         \b/n4232 , \b/n4231 , \b/n4230 , \b/n4229 , \b/n4228 , \b/n4227 ,
         \b/n4226 , \b/n4225 , \b/n4224 , \b/n4223 , \b/n4222 , \b/n4221 ,
         \b/n4220 , \b/n4219 , \b/n4218 , \b/n4217 , \b/n4216 , \b/n4215 ,
         \b/n4214 , \b/n4213 , \b/n4212 , \b/n4211 , \b/n4210 , \b/n4209 ,
         \b/n4208 , \b/n4207 , \b/n4206 , \b/n4205 , \b/n4204 , \b/n4203 ,
         \b/n4202 , \b/n4201 , \b/n4200 , \b/n4199 , \b/n4198 , \b/n4197 ,
         \b/n4196 , \b/n4195 , \b/n4194 , \b/n4193 , \b/n4192 , \b/n4191 ,
         \b/n4190 , \b/n4189 , \b/n4188 , \b/n4187 , \b/n4186 , \b/n4185 ,
         \b/n4184 , \b/n4183 , \b/n4182 , \b/n4181 , \b/n4180 , \b/n4179 ,
         \b/n4178 , \b/n4177 , \b/n4176 , \b/n4175 , \b/n4174 , \b/n4173 ,
         \b/n4172 , \b/n4171 , \b/n4170 , \b/n4169 , \b/n4168 , \b/n4167 ,
         \b/n4166 , \b/n4165 , \b/n4164 , \b/n4163 , \b/n4162 , \b/n4161 ,
         \b/n4160 , \b/n4159 , \b/n4158 , \b/n4157 , \b/n4156 , \b/n4155 ,
         \b/n4154 , \b/n4153 , \b/n4152 , \b/n4151 , \b/n4150 , \b/n4149 ,
         \b/n4148 , \b/n4147 , \b/n4146 , \b/n4145 , \b/n4144 , \b/n4143 ,
         \b/n4142 , \b/n4141 , \b/n4140 , \b/n4139 , \b/n4138 , \b/n4137 ,
         \b/n4136 , \b/n4135 , \b/n4134 , \b/n4133 , \b/n4132 , \b/n4131 ,
         \b/n4130 , \b/n4129 , \b/n4128 , \b/n4127 , \b/n4126 , \b/n4125 ,
         \b/n4124 , \b/n4123 , \b/n4122 , \b/n4121 , \b/n4120 , \b/n4119 ,
         \b/n4118 , \b/n4117 , \b/n4116 , \b/n4115 , \b/n4114 , \b/n4113 ,
         \b/n4112 , \b/n4111 , \b/n4110 , \b/n4109 , \b/n4108 , \b/n4107 ,
         \b/n4106 , \b/n4105 , \b/n4104 , \b/n4103 , \b/n4102 , \b/n4101 ,
         \b/n4100 , \b/n4099 , \b/n4098 , \b/n4097 , \b/n4096 , \b/n4095 ,
         \b/n4094 , \b/n4093 , \b/n4092 , \b/n4091 , \b/n4090 , \b/n4089 ,
         \b/n4088 , \b/n4087 , \b/n4086 , \b/n4085 , \b/n4084 , \b/n4083 ,
         \b/n4082 , \b/n4081 , \b/n4080 , \b/n4079 , \b/n4078 , \b/n4077 ,
         \b/n4076 , \b/n4075 , \b/n4074 , \b/n4073 , \b/n4072 , \b/n4071 ,
         \b/n4070 , \b/n4069 , \b/n4068 , \b/n4067 , \b/n4066 , \b/n4065 ,
         \b/n4064 , \b/n4063 , \b/n4062 , \b/n4061 , \b/n4060 , \b/n4059 ,
         \b/n4058 , \b/n4057 , \b/n4056 , \b/n4055 , \b/n4054 , \b/n4053 ,
         \b/n4052 , \b/n4051 , \b/n4050 , \b/n4049 , \b/n4048 , \b/n4046 ,
         \b/n4045 , \b/n4044 , \b/n4043 , \b/n4042 , \b/n4040 , \b/n4039 ,
         \b/n4038 , \b/n4037 , \b/n4036 , \b/n4035 , \b/n4034 , \b/n4033 ,
         \b/n4032 , \b/n4031 , \b/n4030 , \b/n4028 , \b/n4027 , \b/n4026 ,
         \b/n4024 , \b/n4023 , \b/n4022 , \b/n4021 , \b/n4020 , \b/n4019 ,
         \b/n4018 , \b/n4017 , \b/n4016 , \b/n4015 , \b/n4014 , \b/n4013 ,
         \b/n4012 , \b/n4011 , \b/n4010 , \b/n4009 , \b/n4008 , \b/n4007 ,
         \b/n4006 , \b/n4005 , \b/n4004 , \b/n4003 , \b/n4001 , \b/n4000 ,
         \b/n3999 , \b/n3998 , \b/n3997 , \b/n3996 , \b/n3992 , \b/n3990 ,
         \b/n3989 , \b/n3988 , \b/n3986 , \b/n3983 , \b/n3982 , \b/n3981 ,
         \b/n3980 , \b/n3979 , \b/n3978 , \b/n3977 , \b/n3976 , \b/n3975 ,
         \b/n3974 , \b/n3973 , \b/n3972 , \b/n3971 , \b/n3970 , \b/n3969 ,
         \b/n3968 , \b/n3967 , \b/n3966 , \b/n3965 , \b/n3964 , \b/n3963 ,
         \b/n3962 , \b/n3961 , \b/n3960 , \b/n3959 , \b/n3958 , \b/n3957 ,
         \b/n3956 , \b/n3955 , \b/n3954 , \b/n3953 , \b/n3952 , \b/n3951 ,
         \b/n3950 , \b/n3949 , \b/n3948 , \b/n3947 , \b/n3946 , \b/n3945 ,
         \b/n3944 , \b/n3943 , \b/n3942 , \b/n3941 , \b/n3940 , \b/n3939 ,
         \b/n3938 , \b/n3937 , \b/n3936 , \b/n3935 , \b/n3934 , \b/n3933 ,
         \b/n3932 , \b/n3931 , \b/n3930 , \b/n3929 , \b/n3928 , \b/n3927 ,
         \b/n3926 , \b/n3925 , \b/n3924 , \b/n3923 , \b/n3922 , \b/n3921 ,
         \b/n3920 , \b/n3919 , \b/n3918 , \b/n3917 , \b/n3916 , \b/n3915 ,
         \b/n3914 , \b/n3913 , \b/n3912 , \b/n3911 , \b/n3910 , \b/n3909 ,
         \b/n3908 , \b/n3907 , \b/n3906 , \b/n3905 , \b/n3904 , \b/n3903 ,
         \b/n3902 , \b/n3901 , \b/n3900 , \b/n3899 , \b/n3898 , \b/n3897 ,
         \b/n3896 , \b/n3895 , \b/n3894 , \b/n3893 , \b/n3892 , \b/n3891 ,
         \b/n3890 , \b/n3889 , \b/n3888 , \b/n3887 , \b/n3886 , \b/n3885 ,
         \b/n3884 , \b/n3883 , \b/n3882 , \b/n3881 , \b/n3880 , \b/n3879 ,
         \b/n3878 , \b/n3877 , \b/n3876 , \b/n3875 , \b/n3874 , \b/n3873 ,
         \b/n3872 , \b/n3871 , \b/n3870 , \b/n3869 , \b/n3868 , \b/n3867 ,
         \b/n3866 , \b/n3865 , \b/n3864 , \b/n3863 , \b/n3862 , \b/n3861 ,
         \b/n3860 , \b/n3859 , \b/n3858 , \b/n3857 , \b/n3856 , \b/n3855 ,
         \b/n3854 , \b/n3853 , \b/n3852 , \b/n3851 , \b/n3850 , \b/n3849 ,
         \b/n3848 , \b/n3847 , \b/n3846 , \b/n3845 , \b/n3844 , \b/n3843 ,
         \b/n3842 , \b/n3841 , \b/n3840 , \b/n3839 , \b/n3838 , \b/n3837 ,
         \b/n3836 , \b/n3835 , \b/n3834 , \b/n3833 , \b/n3832 , \b/n3831 ,
         \b/n3830 , \b/n3829 , \b/n3828 , \b/n3827 , \b/n3826 , \b/n3825 ,
         \b/n3824 , \b/n3823 , \b/n3822 , \b/n3821 , \b/n3820 , \b/n3819 ,
         \b/n3818 , \b/n3817 , \b/n3816 , \b/n3815 , \b/n3814 , \b/n3813 ,
         \b/n3812 , \b/n3811 , \b/n3810 , \b/n3809 , \b/n3808 , \b/n3807 ,
         \b/n3806 , \b/n3805 , \b/n3804 , \b/n3803 , \b/n3802 , \b/n3801 ,
         \b/n3800 , \b/n3799 , \b/n3798 , \b/n3797 , \b/n3796 , \b/n3795 ,
         \b/n3794 , \b/n3793 , \b/n3792 , \b/n3791 , \b/n3790 , \b/n3789 ,
         \b/n3788 , \b/n3787 , \b/n3786 , \b/n3785 , \b/n3784 , \b/n3783 ,
         \b/n3782 , \b/n3781 , \b/n3780 , \b/n3779 , \b/n3778 , \b/n3777 ,
         \b/n3776 , \b/n3775 , \b/n3774 , \b/n3773 , \b/n3772 , \b/n3771 ,
         \b/n3770 , \b/n3769 , \b/n3768 , \b/n3767 , \b/n3766 , \b/n3765 ,
         \b/n3764 , \b/n3763 , \b/n3762 , \b/n3761 , \b/n3760 , \b/n3759 ,
         \b/n3758 , \b/n3757 , \b/n3756 , \b/n3755 , \b/n3754 , \b/n3753 ,
         \b/n3752 , \b/n3751 , \b/n3750 , \b/n3749 , \b/n3748 , \b/n3747 ,
         \b/n3746 , \b/n3745 , \b/n3744 , \b/n3743 , \b/n3742 , \b/n3741 ,
         \b/n3740 , \b/n3739 , \b/n3738 , \b/n3737 , \b/n3736 , \b/n3735 ,
         \b/n3734 , \b/n3733 , \b/n3732 , \b/n3731 , \b/n3730 , \b/n3729 ,
         \b/n3728 , \b/n3727 , \b/n3726 , \b/n3725 , \b/n3724 , \b/n3723 ,
         \b/n3722 , \b/n3721 , \b/n3720 , \b/n3719 , \b/n3718 , \b/n3717 ,
         \b/n3716 , \b/n3715 , \b/n3714 , \b/n3713 , \b/n3712 , \b/n3711 ,
         \b/n3710 , \b/n3709 , \b/n3708 , \b/n3707 , \b/n3706 , \b/n3705 ,
         \b/n3704 , \b/n3703 , \b/n3702 , \b/n3701 , \b/n3700 , \b/n3699 ,
         \b/n3698 , \b/n3697 , \b/n3696 , \b/n3695 , \b/n3694 , \b/n3693 ,
         \b/n3692 , \b/n3691 , \b/n3690 , \b/n3689 , \b/n3687 , \b/n3686 ,
         \b/n3685 , \b/n3684 , \b/n3683 , \b/n3681 , \b/n3680 , \b/n3679 ,
         \b/n3678 , \b/n3677 , \b/n3676 , \b/n3675 , \b/n3674 , \b/n3673 ,
         \b/n3672 , \b/n3671 , \b/n3669 , \b/n3668 , \b/n3667 , \b/n3665 ,
         \b/n3664 , \b/n3663 , \b/n3662 , \b/n3661 , \b/n3660 , \b/n3659 ,
         \b/n3658 , \b/n3657 , \b/n3656 , \b/n3655 , \b/n3654 , \b/n3653 ,
         \b/n3652 , \b/n3651 , \b/n3650 , \b/n3649 , \b/n3648 , \b/n3647 ,
         \b/n3646 , \b/n3645 , \b/n3644 , \b/n3642 , \b/n3641 , \b/n3640 ,
         \b/n3639 , \b/n3638 , \b/n3637 , \b/n3633 , \b/n3631 , \b/n3630 ,
         \b/n3629 , \b/n3627 , \b/n3624 , \b/n3623 , \b/n3622 , \b/n3621 ,
         \b/n3620 , \b/n3619 , \b/n3618 , \b/n3617 , \b/n3616 , \b/n3615 ,
         \b/n3614 , \b/n3613 , \b/n3612 , \b/n3611 , \b/n3610 , \b/n3609 ,
         \b/n3608 , \b/n3607 , \b/n3606 , \b/n3605 , \b/n3604 , \b/n3603 ,
         \b/n3602 , \b/n3601 , \b/n3600 , \b/n3599 , \b/n3598 , \b/n3597 ,
         \b/n3596 , \b/n3595 , \b/n3594 , \b/n3593 , \b/n3592 , \b/n3591 ,
         \b/n3590 , \b/n3589 , \b/n3588 , \b/n3587 , \b/n3586 , \b/n3585 ,
         \b/n3584 , \b/n3583 , \b/n3582 , \b/n3581 , \b/n3580 , \b/n3579 ,
         \b/n3578 , \b/n3577 , \b/n3576 , \b/n3575 , \b/n3574 , \b/n3573 ,
         \b/n3572 , \b/n3571 , \b/n3570 , \b/n3569 , \b/n3568 , \b/n3567 ,
         \b/n3566 , \b/n3565 , \b/n3564 , \b/n3563 , \b/n3562 , \b/n3561 ,
         \b/n3560 , \b/n3559 , \b/n3558 , \b/n3557 , \b/n3556 , \b/n3555 ,
         \b/n3554 , \b/n3553 , \b/n3552 , \b/n3551 , \b/n3550 , \b/n3549 ,
         \b/n3548 , \b/n3547 , \b/n3546 , \b/n3545 , \b/n3544 , \b/n3543 ,
         \b/n3542 , \b/n3541 , \b/n3540 , \b/n3539 , \b/n3538 , \b/n3537 ,
         \b/n3536 , \b/n3535 , \b/n3534 , \b/n3533 , \b/n3532 , \b/n3531 ,
         \b/n3530 , \b/n3529 , \b/n3528 , \b/n3527 , \b/n3526 , \b/n3525 ,
         \b/n3524 , \b/n3523 , \b/n3522 , \b/n3521 , \b/n3520 , \b/n3519 ,
         \b/n3518 , \b/n3517 , \b/n3516 , \b/n3515 , \b/n3514 , \b/n3513 ,
         \b/n3512 , \b/n3511 , \b/n3510 , \b/n3509 , \b/n3508 , \b/n3507 ,
         \b/n3506 , \b/n3505 , \b/n3504 , \b/n3503 , \b/n3502 , \b/n3501 ,
         \b/n3500 , \b/n3499 , \b/n3498 , \b/n3497 , \b/n3496 , \b/n3495 ,
         \b/n3494 , \b/n3493 , \b/n3492 , \b/n3491 , \b/n3490 , \b/n3489 ,
         \b/n3488 , \b/n3487 , \b/n3486 , \b/n3485 , \b/n3484 , \b/n3483 ,
         \b/n3482 , \b/n3481 , \b/n3480 , \b/n3479 , \b/n3478 , \b/n3477 ,
         \b/n3476 , \b/n3475 , \b/n3474 , \b/n3473 , \b/n3472 , \b/n3471 ,
         \b/n3470 , \b/n3469 , \b/n3468 , \b/n3467 , \b/n3466 , \b/n3465 ,
         \b/n3464 , \b/n3463 , \b/n3462 , \b/n3461 , \b/n3460 , \b/n3459 ,
         \b/n3458 , \b/n3457 , \b/n3456 , \b/n3455 , \b/n3454 , \b/n3453 ,
         \b/n3452 , \b/n3451 , \b/n3450 , \b/n3449 , \b/n3448 , \b/n3447 ,
         \b/n3446 , \b/n3445 , \b/n3444 , \b/n3443 , \b/n3442 , \b/n3441 ,
         \b/n3440 , \b/n3439 , \b/n3438 , \b/n3437 , \b/n3436 , \b/n3435 ,
         \b/n3434 , \b/n3433 , \b/n3432 , \b/n3431 , \b/n3430 , \b/n3429 ,
         \b/n3428 , \b/n3427 , \b/n3426 , \b/n3425 , \b/n3424 , \b/n3423 ,
         \b/n3422 , \b/n3421 , \b/n3420 , \b/n3419 , \b/n3418 , \b/n3417 ,
         \b/n3416 , \b/n3415 , \b/n3414 , \b/n3413 , \b/n3412 , \b/n3411 ,
         \b/n3410 , \b/n3409 , \b/n3408 , \b/n3407 , \b/n3406 , \b/n3405 ,
         \b/n3404 , \b/n3403 , \b/n3402 , \b/n3401 , \b/n3400 , \b/n3399 ,
         \b/n3398 , \b/n3397 , \b/n3396 , \b/n3395 , \b/n3394 , \b/n3393 ,
         \b/n3392 , \b/n3391 , \b/n3390 , \b/n3389 , \b/n3388 , \b/n3387 ,
         \b/n3386 , \b/n3385 , \b/n3384 , \b/n3383 , \b/n3382 , \b/n3381 ,
         \b/n3380 , \b/n3379 , \b/n3378 , \b/n3377 , \b/n3376 , \b/n3375 ,
         \b/n3374 , \b/n3373 , \b/n3372 , \b/n3371 , \b/n3370 , \b/n3369 ,
         \b/n3368 , \b/n3367 , \b/n3366 , \b/n3365 , \b/n3364 , \b/n3363 ,
         \b/n3362 , \b/n3361 , \b/n3360 , \b/n3359 , \b/n3358 , \b/n3357 ,
         \b/n3356 , \b/n3355 , \b/n3354 , \b/n3353 , \b/n3352 , \b/n3351 ,
         \b/n3350 , \b/n3349 , \b/n3348 , \b/n3347 , \b/n3346 , \b/n3345 ,
         \b/n3344 , \b/n3343 , \b/n3342 , \b/n3341 , \b/n3340 , \b/n3339 ,
         \b/n3338 , \b/n3337 , \b/n3336 , \b/n3335 , \b/n3334 , \b/n3333 ,
         \b/n3332 , \b/n3331 , \b/n3330 , \b/n3328 , \b/n3327 , \b/n3326 ,
         \b/n3325 , \b/n3324 , \b/n3322 , \b/n3321 , \b/n3320 , \b/n3319 ,
         \b/n3318 , \b/n3317 , \b/n3316 , \b/n3315 , \b/n3314 , \b/n3313 ,
         \b/n3312 , \b/n3310 , \b/n3309 , \b/n3308 , \b/n3306 , \b/n3305 ,
         \b/n3304 , \b/n3303 , \b/n3302 , \b/n3301 , \b/n3300 , \b/n3299 ,
         \b/n3298 , \b/n3297 , \b/n3296 , \b/n3295 , \b/n3294 , \b/n3293 ,
         \b/n3292 , \b/n3291 , \b/n3290 , \b/n3289 , \b/n3288 , \b/n3287 ,
         \b/n3286 , \b/n3285 , \b/n3283 , \b/n3282 , \b/n3281 , \b/n3280 ,
         \b/n3279 , \b/n3278 , \b/n3274 , \b/n3272 , \b/n3271 , \b/n3270 ,
         \b/n3268 , \b/n3265 , \b/n3264 , \b/n3263 , \b/n3262 , \b/n3261 ,
         \b/n3260 , \b/n3259 , \b/n3258 , \b/n3257 , \b/n3256 , \b/n3255 ,
         \b/n3254 , \b/n3253 , \b/n3252 , \b/n3251 , \b/n3250 , \b/n3249 ,
         \b/n3248 , \b/n3247 , \b/n3246 , \b/n3245 , \b/n3244 , \b/n3243 ,
         \b/n3242 , \b/n3241 , \b/n3240 , \b/n3239 , \b/n3238 , \b/n3237 ,
         \b/n3236 , \b/n3235 , \b/n3234 , \b/n3233 , \b/n3232 , \b/n3231 ,
         \b/n3230 , \b/n3229 , \b/n3228 , \b/n3227 , \b/n3226 , \b/n3225 ,
         \b/n3224 , \b/n3223 , \b/n3222 , \b/n3221 , \b/n3220 , \b/n3219 ,
         \b/n3218 , \b/n3217 , \b/n3216 , \b/n3215 , \b/n3214 , \b/n3213 ,
         \b/n3212 , \b/n3211 , \b/n3210 , \b/n3209 , \b/n3208 , \b/n3207 ,
         \b/n3206 , \b/n3205 , \b/n3204 , \b/n3203 , \b/n3202 , \b/n3201 ,
         \b/n3200 , \b/n3199 , \b/n3198 , \b/n3197 , \b/n3196 , \b/n3195 ,
         \b/n3194 , \b/n3193 , \b/n3192 , \b/n3191 , \b/n3190 , \b/n3189 ,
         \b/n3188 , \b/n3187 , \b/n3186 , \b/n3185 , \b/n3184 , \b/n3183 ,
         \b/n3182 , \b/n3181 , \b/n3180 , \b/n3179 , \b/n3178 , \b/n3177 ,
         \b/n3176 , \b/n3175 , \b/n3174 , \b/n3173 , \b/n3172 , \b/n3171 ,
         \b/n3170 , \b/n3169 , \b/n3168 , \b/n3167 , \b/n3166 , \b/n3165 ,
         \b/n3164 , \b/n3163 , \b/n3162 , \b/n3161 , \b/n3160 , \b/n3159 ,
         \b/n3158 , \b/n3157 , \b/n3156 , \b/n3155 , \b/n3154 , \b/n3153 ,
         \b/n3152 , \b/n3151 , \b/n3150 , \b/n3149 , \b/n3148 , \b/n3147 ,
         \b/n3146 , \b/n3145 , \b/n3144 , \b/n3143 , \b/n3142 , \b/n3141 ,
         \b/n3140 , \b/n3139 , \b/n3138 , \b/n3137 , \b/n3136 , \b/n3135 ,
         \b/n3134 , \b/n3133 , \b/n3132 , \b/n3131 , \b/n3130 , \b/n3129 ,
         \b/n3128 , \b/n3127 , \b/n3126 , \b/n3125 , \b/n3124 , \b/n3123 ,
         \b/n3122 , \b/n3121 , \b/n3120 , \b/n3119 , \b/n3118 , \b/n3117 ,
         \b/n3116 , \b/n3115 , \b/n3114 , \b/n3113 , \b/n3112 , \b/n3111 ,
         \b/n3110 , \b/n3109 , \b/n3108 , \b/n3107 , \b/n3106 , \b/n3105 ,
         \b/n3104 , \b/n3103 , \b/n3102 , \b/n3101 , \b/n3100 , \b/n3099 ,
         \b/n3098 , \b/n3097 , \b/n3096 , \b/n3095 , \b/n3094 , \b/n3093 ,
         \b/n3092 , \b/n3091 , \b/n3090 , \b/n3089 , \b/n3088 , \b/n3087 ,
         \b/n3086 , \b/n3085 , \b/n3084 , \b/n3083 , \b/n3082 , \b/n3081 ,
         \b/n3080 , \b/n3079 , \b/n3078 , \b/n3077 , \b/n3076 , \b/n3075 ,
         \b/n3074 , \b/n3073 , \b/n3072 , \b/n3071 , \b/n3070 , \b/n3069 ,
         \b/n3068 , \b/n3067 , \b/n3066 , \b/n3065 , \b/n3064 , \b/n3063 ,
         \b/n3062 , \b/n3061 , \b/n3060 , \b/n3059 , \b/n3058 , \b/n3057 ,
         \b/n3056 , \b/n3055 , \b/n3054 , \b/n3053 , \b/n3052 , \b/n3051 ,
         \b/n3050 , \b/n3049 , \b/n3048 , \b/n3047 , \b/n3046 , \b/n3045 ,
         \b/n3044 , \b/n3043 , \b/n3042 , \b/n3041 , \b/n3040 , \b/n3039 ,
         \b/n3038 , \b/n3037 , \b/n3036 , \b/n3035 , \b/n3034 , \b/n3033 ,
         \b/n3032 , \b/n3031 , \b/n3030 , \b/n3029 , \b/n3028 , \b/n3027 ,
         \b/n3026 , \b/n3025 , \b/n3024 , \b/n3023 , \b/n3022 , \b/n3021 ,
         \b/n3020 , \b/n3019 , \b/n3018 , \b/n3017 , \b/n3016 , \b/n3015 ,
         \b/n3014 , \b/n3013 , \b/n3012 , \b/n3011 , \b/n3010 , \b/n3009 ,
         \b/n3008 , \b/n3007 , \b/n3006 , \b/n3005 , \b/n3004 , \b/n3003 ,
         \b/n3002 , \b/n3001 , \b/n3000 , \b/n2999 , \b/n2998 , \b/n2997 ,
         \b/n2996 , \b/n2995 , \b/n2994 , \b/n2993 , \b/n2992 , \b/n2991 ,
         \b/n2990 , \b/n2989 , \b/n2988 , \b/n2987 , \b/n2986 , \b/n2985 ,
         \b/n2984 , \b/n2983 , \b/n2982 , \b/n2981 , \b/n2980 , \b/n2979 ,
         \b/n2978 , \b/n2977 , \b/n2976 , \b/n2975 , \b/n2974 , \b/n2973 ,
         \b/n2972 , \b/n2971 , \b/n2969 , \b/n2968 , \b/n2967 , \b/n2966 ,
         \b/n2965 , \b/n2963 , \b/n2962 , \b/n2961 , \b/n2960 , \b/n2959 ,
         \b/n2958 , \b/n2957 , \b/n2956 , \b/n2955 , \b/n2954 , \b/n2953 ,
         \b/n2951 , \b/n2950 , \b/n2949 , \b/n2947 , \b/n2946 , \b/n2945 ,
         \b/n2944 , \b/n2943 , \b/n2942 , \b/n2941 , \b/n2940 , \b/n2939 ,
         \b/n2938 , \b/n2937 , \b/n2936 , \b/n2935 , \b/n2934 , \b/n2933 ,
         \b/n2932 , \b/n2931 , \b/n2930 , \b/n2929 , \b/n2928 , \b/n2927 ,
         \b/n2926 , \b/n2924 , \b/n2923 , \b/n2922 , \b/n2921 , \b/n2920 ,
         \b/n2919 , \b/n2915 , \b/n2913 , \b/n2912 , \b/n2911 , \b/n2909 ,
         \b/n2906 , \b/n2905 , \b/n2904 , \b/n2903 , \b/n2902 , \b/n2901 ,
         \b/n2900 , \b/n2899 , \b/n2898 , \b/n2897 , \b/n2896 , \b/n2895 ,
         \b/n2894 , \b/n2893 , \b/n2892 , \b/n2891 , \b/n2890 , \b/n2889 ,
         \b/n2888 , \b/n2887 , \b/n2886 , \b/n2885 , \b/n2884 , \b/n2883 ,
         \b/n2882 , \b/n2881 , \b/n2880 , \b/n2879 , \b/n2878 , \b/n2877 ,
         \b/n2876 , \b/n2875 , \b/n2874 , \b/n2873 , \b/n2872 , \b/n2871 ,
         \b/n2870 , \b/n2869 , \b/n2868 , \b/n2867 , \b/n2866 , \b/n2865 ,
         \b/n2864 , \b/n2863 , \b/n2862 , \b/n2861 , \b/n2860 , \b/n2859 ,
         \b/n2858 , \b/n2857 , \b/n2856 , \b/n2855 , \b/n2854 , \b/n2853 ,
         \b/n2852 , \b/n2851 , \b/n2850 , \b/n2849 , \b/n2848 , \b/n2847 ,
         \b/n2846 , \b/n2845 , \b/n2844 , \b/n2843 , \b/n2842 , \b/n2841 ,
         \b/n2840 , \b/n2839 , \b/n2838 , \b/n2837 , \b/n2836 , \b/n2835 ,
         \b/n2834 , \b/n2833 , \b/n2832 , \b/n2831 , \b/n2830 , \b/n2829 ,
         \b/n2828 , \b/n2827 , \b/n2826 , \b/n2825 , \b/n2824 , \b/n2823 ,
         \b/n2822 , \b/n2821 , \b/n2820 , \b/n2819 , \b/n2818 , \b/n2817 ,
         \b/n2816 , \b/n2815 , \b/n2814 , \b/n2813 , \b/n2812 , \b/n2811 ,
         \b/n2810 , \b/n2809 , \b/n2808 , \b/n2807 , \b/n2806 , \b/n2805 ,
         \b/n2804 , \b/n2803 , \b/n2802 , \b/n2801 , \b/n2800 , \b/n2799 ,
         \b/n2798 , \b/n2797 , \b/n2796 , \b/n2795 , \b/n2794 , \b/n2793 ,
         \b/n2792 , \b/n2791 , \b/n2790 , \b/n2789 , \b/n2788 , \b/n2787 ,
         \b/n2786 , \b/n2785 , \b/n2784 , \b/n2783 , \b/n2782 , \b/n2781 ,
         \b/n2780 , \b/n2779 , \b/n2778 , \b/n2777 , \b/n2776 , \b/n2775 ,
         \b/n2774 , \b/n2773 , \b/n2772 , \b/n2771 , \b/n2770 , \b/n2769 ,
         \b/n2768 , \b/n2767 , \b/n2766 , \b/n2765 , \b/n2764 , \b/n2763 ,
         \b/n2762 , \b/n2761 , \b/n2760 , \b/n2759 , \b/n2758 , \b/n2757 ,
         \b/n2756 , \b/n2755 , \b/n2754 , \b/n2753 , \b/n2752 , \b/n2751 ,
         \b/n2750 , \b/n2749 , \b/n2748 , \b/n2747 , \b/n2746 , \b/n2745 ,
         \b/n2744 , \b/n2743 , \b/n2742 , \b/n2741 , \b/n2740 , \b/n2739 ,
         \b/n2738 , \b/n2737 , \b/n2736 , \b/n2735 , \b/n2734 , \b/n2733 ,
         \b/n2732 , \b/n2731 , \b/n2730 , \b/n2729 , \b/n2728 , \b/n2727 ,
         \b/n2726 , \b/n2725 , \b/n2724 , \b/n2723 , \b/n2722 , \b/n2721 ,
         \b/n2720 , \b/n2719 , \b/n2718 , \b/n2717 , \b/n2716 , \b/n2715 ,
         \b/n2714 , \b/n2713 , \b/n2712 , \b/n2711 , \b/n2710 , \b/n2709 ,
         \b/n2708 , \b/n2707 , \b/n2706 , \b/n2705 , \b/n2704 , \b/n2703 ,
         \b/n2702 , \b/n2701 , \b/n2700 , \b/n2699 , \b/n2698 , \b/n2697 ,
         \b/n2696 , \b/n2695 , \b/n2694 , \b/n2693 , \b/n2692 , \b/n2691 ,
         \b/n2690 , \b/n2689 , \b/n2688 , \b/n2687 , \b/n2686 , \b/n2685 ,
         \b/n2684 , \b/n2683 , \b/n2682 , \b/n2681 , \b/n2680 , \b/n2679 ,
         \b/n2678 , \b/n2677 , \b/n2676 , \b/n2675 , \b/n2674 , \b/n2673 ,
         \b/n2672 , \b/n2671 , \b/n2670 , \b/n2669 , \b/n2668 , \b/n2667 ,
         \b/n2666 , \b/n2665 , \b/n2664 , \b/n2663 , \b/n2662 , \b/n2661 ,
         \b/n2660 , \b/n2659 , \b/n2658 , \b/n2657 , \b/n2656 , \b/n2655 ,
         \b/n2654 , \b/n2653 , \b/n2652 , \b/n2651 , \b/n2650 , \b/n2649 ,
         \b/n2648 , \b/n2647 , \b/n2646 , \b/n2645 , \b/n2644 , \b/n2643 ,
         \b/n2642 , \b/n2641 , \b/n2640 , \b/n2639 , \b/n2638 , \b/n2637 ,
         \b/n2636 , \b/n2635 , \b/n2634 , \b/n2633 , \b/n2632 , \b/n2631 ,
         \b/n2630 , \b/n2629 , \b/n2628 , \b/n2627 , \b/n2626 , \b/n2625 ,
         \b/n2624 , \b/n2623 , \b/n2622 , \b/n2621 , \b/n2620 , \b/n2619 ,
         \b/n2618 , \b/n2617 , \b/n2616 , \b/n2615 , \b/n2614 , \b/n2613 ,
         \b/n2612 , \b/n2610 , \b/n2609 , \b/n2608 , \b/n2607 , \b/n2606 ,
         \b/n2604 , \b/n2603 , \b/n2602 , \b/n2601 , \b/n2600 , \b/n2599 ,
         \b/n2598 , \b/n2597 , \b/n2596 , \b/n2595 , \b/n2594 , \b/n2592 ,
         \b/n2591 , \b/n2590 , \b/n2588 , \b/n2587 , \b/n2586 , \b/n2585 ,
         \b/n2584 , \b/n2583 , \b/n2582 , \b/n2581 , \b/n2580 , \b/n2579 ,
         \b/n2578 , \b/n2577 , \b/n2576 , \b/n2575 , \b/n2574 , \b/n2573 ,
         \b/n2572 , \b/n2571 , \b/n2570 , \b/n2569 , \b/n2568 , \b/n2567 ,
         \b/n2565 , \b/n2564 , \b/n2563 , \b/n2562 , \b/n2561 , \b/n2560 ,
         \b/n2556 , \b/n2554 , \b/n2553 , \b/n2552 , \b/n2550 , \b/n2547 ,
         \b/n2546 , \b/n2545 , \b/n2544 , \b/n2543 , \b/n2542 , \b/n2541 ,
         \b/n2540 , \b/n2539 , \b/n2538 , \b/n2537 , \b/n2536 , \b/n2535 ,
         \b/n2534 , \b/n2533 , \b/n2532 , \b/n2531 , \b/n2530 , \b/n2529 ,
         \b/n2528 , \b/n2527 , \b/n2526 , \b/n2525 , \b/n2524 , \b/n2523 ,
         \b/n2522 , \b/n2521 , \b/n2520 , \b/n2519 , \b/n2518 , \b/n2517 ,
         \b/n2516 , \b/n2515 , \b/n2514 , \b/n2513 , \b/n2512 , \b/n2511 ,
         \b/n2510 , \b/n2509 , \b/n2508 , \b/n2507 , \b/n2506 , \b/n2505 ,
         \b/n2504 , \b/n2503 , \b/n2502 , \b/n2501 , \b/n2500 , \b/n2499 ,
         \b/n2498 , \b/n2497 , \b/n2496 , \b/n2495 , \b/n2494 , \b/n2493 ,
         \b/n2492 , \b/n2491 , \b/n2490 , \b/n2489 , \b/n2488 , \b/n2487 ,
         \b/n2486 , \b/n2485 , \b/n2484 , \b/n2483 , \b/n2482 , \b/n2481 ,
         \b/n2480 , \b/n2479 , \b/n2478 , \b/n2477 , \b/n2476 , \b/n2475 ,
         \b/n2474 , \b/n2473 , \b/n2472 , \b/n2471 , \b/n2470 , \b/n2469 ,
         \b/n2468 , \b/n2467 , \b/n2466 , \b/n2465 , \b/n2464 , \b/n2463 ,
         \b/n2462 , \b/n2461 , \b/n2460 , \b/n2459 , \b/n2458 , \b/n2457 ,
         \b/n2456 , \b/n2455 , \b/n2454 , \b/n2453 , \b/n2452 , \b/n2451 ,
         \b/n2450 , \b/n2449 , \b/n2448 , \b/n2447 , \b/n2446 , \b/n2445 ,
         \b/n2444 , \b/n2443 , \b/n2442 , \b/n2441 , \b/n2440 , \b/n2439 ,
         \b/n2438 , \b/n2437 , \b/n2436 , \b/n2435 , \b/n2434 , \b/n2433 ,
         \b/n2432 , \b/n2431 , \b/n2430 , \b/n2429 , \b/n2428 , \b/n2427 ,
         \b/n2426 , \b/n2425 , \b/n2424 , \b/n2423 , \b/n2422 , \b/n2421 ,
         \b/n2420 , \b/n2419 , \b/n2418 , \b/n2417 , \b/n2416 , \b/n2415 ,
         \b/n2414 , \b/n2413 , \b/n2412 , \b/n2411 , \b/n2410 , \b/n2409 ,
         \b/n2408 , \b/n2407 , \b/n2406 , \b/n2405 , \b/n2404 , \b/n2403 ,
         \b/n2402 , \b/n2401 , \b/n2400 , \b/n2399 , \b/n2398 , \b/n2397 ,
         \b/n2396 , \b/n2395 , \b/n2394 , \b/n2393 , \b/n2392 , \b/n2391 ,
         \b/n2390 , \b/n2389 , \b/n2388 , \b/n2387 , \b/n2386 , \b/n2385 ,
         \b/n2384 , \b/n2383 , \b/n2382 , \b/n2381 , \b/n2380 , \b/n2379 ,
         \b/n2378 , \b/n2377 , \b/n2376 , \b/n2375 , \b/n2374 , \b/n2373 ,
         \b/n2372 , \b/n2371 , \b/n2370 , \b/n2369 , \b/n2368 , \b/n2367 ,
         \b/n2366 , \b/n2365 , \b/n2364 , \b/n2363 , \b/n2362 , \b/n2361 ,
         \b/n2360 , \b/n2359 , \b/n2358 , \b/n2357 , \b/n2356 , \b/n2355 ,
         \b/n2354 , \b/n2353 , \b/n2352 , \b/n2351 , \b/n2350 , \b/n2349 ,
         \b/n2348 , \b/n2347 , \b/n2346 , \b/n2345 , \b/n2344 , \b/n2343 ,
         \b/n2342 , \b/n2341 , \b/n2340 , \b/n2339 , \b/n2338 , \b/n2337 ,
         \b/n2336 , \b/n2335 , \b/n2334 , \b/n2333 , \b/n2332 , \b/n2331 ,
         \b/n2330 , \b/n2329 , \b/n2328 , \b/n2327 , \b/n2326 , \b/n2325 ,
         \b/n2324 , \b/n2323 , \b/n2322 , \b/n2321 , \b/n2320 , \b/n2319 ,
         \b/n2318 , \b/n2317 , \b/n2316 , \b/n2315 , \b/n2314 , \b/n2313 ,
         \b/n2312 , \b/n2311 , \b/n2310 , \b/n2309 , \b/n2308 , \b/n2307 ,
         \b/n2306 , \b/n2305 , \b/n2304 , \b/n2303 , \b/n2302 , \b/n2301 ,
         \b/n2300 , \b/n2299 , \b/n2298 , \b/n2297 , \b/n2296 , \b/n2295 ,
         \b/n2294 , \b/n2293 , \b/n2292 , \b/n2291 , \b/n2290 , \b/n2289 ,
         \b/n2288 , \b/n2287 , \b/n2286 , \b/n2285 , \b/n2284 , \b/n2283 ,
         \b/n2282 , \b/n2281 , \b/n2280 , \b/n2279 , \b/n2278 , \b/n2277 ,
         \b/n2276 , \b/n2275 , \b/n2274 , \b/n2273 , \b/n2272 , \b/n2271 ,
         \b/n2270 , \b/n2269 , \b/n2268 , \b/n2267 , \b/n2266 , \b/n2265 ,
         \b/n2264 , \b/n2263 , \b/n2262 , \b/n2261 , \b/n2260 , \b/n2259 ,
         \b/n2258 , \b/n2257 , \b/n2256 , \b/n2255 , \b/n2254 , \b/n2253 ,
         \b/n2251 , \b/n2250 , \b/n2249 , \b/n2248 , \b/n2247 , \b/n2245 ,
         \b/n2244 , \b/n2243 , \b/n2242 , \b/n2241 , \b/n2240 , \b/n2239 ,
         \b/n2238 , \b/n2237 , \b/n2236 , \b/n2235 , \b/n2233 , \b/n2232 ,
         \b/n2231 , \b/n2229 , \b/n2228 , \b/n2227 , \b/n2226 , \b/n2225 ,
         \b/n2224 , \b/n2223 , \b/n2222 , \b/n2221 , \b/n2220 , \b/n2219 ,
         \b/n2218 , \b/n2217 , \b/n2216 , \b/n2215 , \b/n2214 , \b/n2213 ,
         \b/n2212 , \b/n2211 , \b/n2210 , \b/n2209 , \b/n2208 , \b/n2206 ,
         \b/n2205 , \b/n2204 , \b/n2203 , \b/n2202 , \b/n2201 , \b/n2197 ,
         \b/n2195 , \b/n2194 , \b/n2193 , \b/n2191 , \b/n2188 , \b/n2187 ,
         \b/n2186 , \b/n2185 , \b/n2184 , \b/n2183 , \b/n2182 , \b/n2181 ,
         \b/n2180 , \b/n2179 , \b/n2178 , \b/n2177 , \b/n2176 , \b/n2175 ,
         \b/n2174 , \b/n2173 , \b/n2172 , \b/n2171 , \b/n2170 , \b/n2169 ,
         \b/n2168 , \b/n2167 , \b/n2166 , \b/n2165 , \b/n2164 , \b/n2163 ,
         \b/n2162 , \b/n2161 , \b/n2160 , \b/n2159 , \b/n2158 , \b/n2157 ,
         \b/n2156 , \b/n2155 , \b/n2154 , \b/n2153 , \b/n2152 , \b/n2151 ,
         \b/n2150 , \b/n2149 , \b/n2148 , \b/n2147 , \b/n2146 , \b/n2145 ,
         \b/n2144 , \b/n2143 , \b/n2142 , \b/n2141 , \b/n2140 , \b/n2139 ,
         \b/n2138 , \b/n2137 , \b/n2136 , \b/n2135 , \b/n2134 , \b/n2133 ,
         \b/n2132 , \b/n2131 , \b/n2130 , \b/n2129 , \b/n2128 , \b/n2127 ,
         \b/n2126 , \b/n2125 , \b/n2124 , \b/n2123 , \b/n2122 , \b/n2121 ,
         \b/n2120 , \b/n2119 , \b/n2118 , \b/n2117 , \b/n2116 , \b/n2115 ,
         \b/n2114 , \b/n2113 , \b/n2112 , \b/n2111 , \b/n2110 , \b/n2109 ,
         \b/n2108 , \b/n2107 , \b/n2106 , \b/n2105 , \b/n2104 , \b/n2103 ,
         \b/n2102 , \b/n2101 , \b/n2100 , \b/n2099 , \b/n2098 , \b/n2097 ,
         \b/n2096 , \b/n2095 , \b/n2094 , \b/n2093 , \b/n2092 , \b/n2091 ,
         \b/n2090 , \b/n2089 , \b/n2088 , \b/n2087 , \b/n2086 , \b/n2085 ,
         \b/n2084 , \b/n2083 , \b/n2082 , \b/n2081 , \b/n2080 , \b/n2079 ,
         \b/n2078 , \b/n2077 , \b/n2076 , \b/n2075 , \b/n2074 , \b/n2073 ,
         \b/n2072 , \b/n2071 , \b/n2070 , \b/n2069 , \b/n2068 , \b/n2067 ,
         \b/n2066 , \b/n2065 , \b/n2064 , \b/n2063 , \b/n2062 , \b/n2061 ,
         \b/n2060 , \b/n2059 , \b/n2058 , \b/n2057 , \b/n2056 , \b/n2055 ,
         \b/n2054 , \b/n2053 , \b/n2052 , \b/n2051 , \b/n2050 , \b/n2049 ,
         \b/n2048 , \b/n2047 , \b/n2046 , \b/n2045 , \b/n2044 , \b/n2043 ,
         \b/n2042 , \b/n2041 , \b/n2040 , \b/n2039 , \b/n2038 , \b/n2037 ,
         \b/n2036 , \b/n2035 , \b/n2034 , \b/n2033 , \b/n2032 , \b/n2031 ,
         \b/n2030 , \b/n2029 , \b/n2028 , \b/n2027 , \b/n2026 , \b/n2025 ,
         \b/n2024 , \b/n2023 , \b/n2022 , \b/n2021 , \b/n2020 , \b/n2019 ,
         \b/n2018 , \b/n2017 , \b/n2016 , \b/n2015 , \b/n2014 , \b/n2013 ,
         \b/n2012 , \b/n2011 , \b/n2010 , \b/n2009 , \b/n2008 , \b/n2007 ,
         \b/n2006 , \b/n2005 , \b/n2004 , \b/n2003 , \b/n2002 , \b/n2001 ,
         \b/n2000 , \b/n1999 , \b/n1998 , \b/n1997 , \b/n1996 , \b/n1995 ,
         \b/n1994 , \b/n1993 , \b/n1992 , \b/n1991 , \b/n1990 , \b/n1989 ,
         \b/n1988 , \b/n1987 , \b/n1986 , \b/n1985 , \b/n1984 , \b/n1983 ,
         \b/n1982 , \b/n1981 , \b/n1980 , \b/n1979 , \b/n1978 , \b/n1977 ,
         \b/n1976 , \b/n1975 , \b/n1974 , \b/n1973 , \b/n1972 , \b/n1971 ,
         \b/n1970 , \b/n1969 , \b/n1968 , \b/n1967 , \b/n1966 , \b/n1965 ,
         \b/n1964 , \b/n1963 , \b/n1962 , \b/n1961 , \b/n1960 , \b/n1959 ,
         \b/n1958 , \b/n1957 , \b/n1956 , \b/n1955 , \b/n1954 , \b/n1953 ,
         \b/n1952 , \b/n1951 , \b/n1950 , \b/n1949 , \b/n1948 , \b/n1947 ,
         \b/n1946 , \b/n1945 , \b/n1944 , \b/n1943 , \b/n1942 , \b/n1941 ,
         \b/n1940 , \b/n1939 , \b/n1938 , \b/n1937 , \b/n1936 , \b/n1935 ,
         \b/n1934 , \b/n1933 , \b/n1932 , \b/n1931 , \b/n1930 , \b/n1929 ,
         \b/n1928 , \b/n1927 , \b/n1926 , \b/n1925 , \b/n1924 , \b/n1923 ,
         \b/n1922 , \b/n1921 , \b/n1920 , \b/n1919 , \b/n1918 , \b/n1917 ,
         \b/n1916 , \b/n1915 , \b/n1914 , \b/n1913 , \b/n1912 , \b/n1911 ,
         \b/n1910 , \b/n1909 , \b/n1908 , \b/n1907 , \b/n1906 , \b/n1905 ,
         \b/n1904 , \b/n1903 , \b/n1902 , \b/n1901 , \b/n1900 , \b/n1899 ,
         \b/n1898 , \b/n1897 , \b/n1896 , \b/n1895 , \b/n1894 , \b/n1892 ,
         \b/n1891 , \b/n1890 , \b/n1889 , \b/n1888 , \b/n1886 , \b/n1885 ,
         \b/n1884 , \b/n1883 , \b/n1882 , \b/n1881 , \b/n1880 , \b/n1879 ,
         \b/n1878 , \b/n1877 , \b/n1876 , \b/n1874 , \b/n1873 , \b/n1872 ,
         \b/n1870 , \b/n1869 , \b/n1868 , \b/n1867 , \b/n1866 , \b/n1865 ,
         \b/n1864 , \b/n1863 , \b/n1862 , \b/n1861 , \b/n1860 , \b/n1859 ,
         \b/n1858 , \b/n1857 , \b/n1856 , \b/n1855 , \b/n1854 , \b/n1853 ,
         \b/n1852 , \b/n1851 , \b/n1850 , \b/n1849 , \b/n1847 , \b/n1846 ,
         \b/n1845 , \b/n1844 , \b/n1843 , \b/n1842 , \b/n1838 , \b/n1837 ,
         \b/n1835 , \b/n1834 , \b/n1831 , \b/n1829 , \b/n1828 , \b/n1827 ,
         \b/n1826 , \b/n1825 , \b/n1824 , \b/n1823 , \b/n1822 , \b/n1821 ,
         \b/n1820 , \b/n1819 , \b/n1818 , \b/n1817 , \b/n1816 , \b/n1815 ,
         \b/n1814 , \b/n1813 , \b/n1812 , \b/n1811 , \b/n1810 , \b/n1809 ,
         \b/n1808 , \b/n1807 , \b/n1806 , \b/n1805 , \b/n1804 , \b/n1803 ,
         \b/n1802 , \b/n1801 , \b/n1800 , \b/n1799 , \b/n1798 , \b/n1797 ,
         \b/n1796 , \b/n1795 , \b/n1794 , \b/n1793 , \b/n1792 , \b/n1791 ,
         \b/n1790 , \b/n1789 , \b/n1788 , \b/n1787 , \b/n1786 , \b/n1785 ,
         \b/n1784 , \b/n1783 , \b/n1782 , \b/n1781 , \b/n1780 , \b/n1779 ,
         \b/n1778 , \b/n1777 , \b/n1776 , \b/n1775 , \b/n1774 , \b/n1773 ,
         \b/n1772 , \b/n1771 , \b/n1770 , \b/n1769 , \b/n1768 , \b/n1767 ,
         \b/n1766 , \b/n1765 , \b/n1764 , \b/n1763 , \b/n1762 , \b/n1761 ,
         \b/n1760 , \b/n1759 , \b/n1758 , \b/n1757 , \b/n1756 , \b/n1755 ,
         \b/n1754 , \b/n1753 , \b/n1752 , \b/n1751 , \b/n1750 , \b/n1749 ,
         \b/n1748 , \b/n1747 , \b/n1746 , \b/n1745 , \b/n1744 , \b/n1743 ,
         \b/n1742 , \b/n1741 , \b/n1740 , \b/n1739 , \b/n1738 , \b/n1737 ,
         \b/n1736 , \b/n1735 , \b/n1734 , \b/n1733 , \b/n1732 , \b/n1731 ,
         \b/n1730 , \b/n1729 , \b/n1728 , \b/n1727 , \b/n1726 , \b/n1725 ,
         \b/n1724 , \b/n1723 , \b/n1722 , \b/n1721 , \b/n1720 , \b/n1719 ,
         \b/n1718 , \b/n1717 , \b/n1716 , \b/n1715 , \b/n1714 , \b/n1713 ,
         \b/n1712 , \b/n1711 , \b/n1710 , \b/n1709 , \b/n1708 , \b/n1707 ,
         \b/n1706 , \b/n1705 , \b/n1704 , \b/n1703 , \b/n1702 , \b/n1701 ,
         \b/n1700 , \b/n1699 , \b/n1698 , \b/n1697 , \b/n1696 , \b/n1695 ,
         \b/n1694 , \b/n1693 , \b/n1692 , \b/n1691 , \b/n1690 , \b/n1689 ,
         \b/n1688 , \b/n1687 , \b/n1686 , \b/n1685 , \b/n1684 , \b/n1683 ,
         \b/n1682 , \b/n1681 , \b/n1680 , \b/n1679 , \b/n1678 , \b/n1677 ,
         \b/n1676 , \b/n1675 , \b/n1674 , \b/n1673 , \b/n1672 , \b/n1671 ,
         \b/n1670 , \b/n1669 , \b/n1668 , \b/n1667 , \b/n1666 , \b/n1665 ,
         \b/n1664 , \b/n1663 , \b/n1662 , \b/n1661 , \b/n1660 , \b/n1659 ,
         \b/n1658 , \b/n1657 , \b/n1656 , \b/n1655 , \b/n1654 , \b/n1653 ,
         \b/n1652 , \b/n1651 , \b/n1650 , \b/n1649 , \b/n1648 , \b/n1647 ,
         \b/n1646 , \b/n1645 , \b/n1644 , \b/n1643 , \b/n1642 , \b/n1641 ,
         \b/n1640 , \b/n1639 , \b/n1638 , \b/n1637 , \b/n1636 , \b/n1635 ,
         \b/n1634 , \b/n1633 , \b/n1632 , \b/n1631 , \b/n1630 , \b/n1629 ,
         \b/n1628 , \b/n1627 , \b/n1626 , \b/n1625 , \b/n1624 , \b/n1623 ,
         \b/n1622 , \b/n1621 , \b/n1620 , \b/n1619 , \b/n1618 , \b/n1617 ,
         \b/n1616 , \b/n1615 , \b/n1614 , \b/n1613 , \b/n1612 , \b/n1611 ,
         \b/n1610 , \b/n1609 , \b/n1608 , \b/n1607 , \b/n1606 , \b/n1605 ,
         \b/n1604 , \b/n1603 , \b/n1602 , \b/n1601 , \b/n1600 , \b/n1599 ,
         \b/n1598 , \b/n1597 , \b/n1596 , \b/n1595 , \b/n1594 , \b/n1593 ,
         \b/n1592 , \b/n1591 , \b/n1590 , \b/n1589 , \b/n1588 , \b/n1587 ,
         \b/n1586 , \b/n1585 , \b/n1584 , \b/n1583 , \b/n1582 , \b/n1581 ,
         \b/n1580 , \b/n1579 , \b/n1578 , \b/n1577 , \b/n1576 , \b/n1575 ,
         \b/n1574 , \b/n1573 , \b/n1572 , \b/n1571 , \b/n1570 , \b/n1569 ,
         \b/n1568 , \b/n1567 , \b/n1566 , \b/n1565 , \b/n1564 , \b/n1563 ,
         \b/n1562 , \b/n1561 , \b/n1560 , \b/n1559 , \b/n1558 , \b/n1557 ,
         \b/n1556 , \b/n1555 , \b/n1554 , \b/n1553 , \b/n1552 , \b/n1551 ,
         \b/n1550 , \b/n1549 , \b/n1548 , \b/n1547 , \b/n1546 , \b/n1545 ,
         \b/n1544 , \b/n1543 , \b/n1542 , \b/n1541 , \b/n1540 , \b/n1539 ,
         \b/n1538 , \b/n1537 , \b/n1536 , \b/n1535 , \b/n1533 , \b/n1532 ,
         \b/n1531 , \b/n1530 , \b/n1529 , \b/n1528 , \b/n1526 , \b/n1525 ,
         \b/n1524 , \b/n1523 , \b/n1522 , \b/n1521 , \b/n1520 , \b/n1519 ,
         \b/n1518 , \b/n1517 , \b/n1515 , \b/n1514 , \b/n1513 , \b/n1512 ,
         \b/n1511 , \b/n1510 , \b/n1509 , \b/n1508 , \b/n1507 , \b/n1505 ,
         \b/n1504 , \b/n1503 , \b/n1502 , \b/n1501 , \b/n1500 , \b/n1499 ,
         \b/n1498 , \b/n1497 , \b/n1496 , \b/n1495 , \b/n1494 , \b/n1493 ,
         \b/n1492 , \b/n1491 , \b/n1490 , \b/n1488 , \b/n1487 , \b/n1486 ,
         \b/n1485 , \b/n1484 , \b/n1483 , \b/n1479 , \b/n1477 , \b/n1476 ,
         \b/n1475 , \b/n1473 , \b/n1470 , \b/n1469 , \b/n1468 , \b/n1467 ,
         \b/n1466 , \b/n1465 , \b/n1464 , \b/n1463 , \b/n1462 , \b/n1461 ,
         \b/n1460 , \b/n1459 , \b/n1458 , \b/n1457 , \b/n1456 , \b/n1455 ,
         \b/n1454 , \b/n1453 , \b/n1452 , \b/n1451 , \b/n1450 , \b/n1449 ,
         \b/n1448 , \b/n1447 , \b/n1446 , \b/n1445 , \b/n1444 , \b/n1443 ,
         \b/n1442 , \b/n1441 , \b/n1440 , \b/n1439 , \b/n1438 , \b/n1437 ,
         \b/n1436 , \b/n1435 , \b/n1434 , \b/n1433 , \b/n1432 , \b/n1431 ,
         \b/n1430 , \b/n1429 , \b/n1428 , \b/n1427 , \b/n1426 , \b/n1425 ,
         \b/n1424 , \b/n1423 , \b/n1422 , \b/n1421 , \b/n1420 , \b/n1419 ,
         \b/n1418 , \b/n1417 , \b/n1416 , \b/n1415 , \b/n1414 , \b/n1413 ,
         \b/n1412 , \b/n1411 , \b/n1410 , \b/n1409 , \b/n1408 , \b/n1407 ,
         \b/n1406 , \b/n1405 , \b/n1404 , \b/n1403 , \b/n1402 , \b/n1401 ,
         \b/n1400 , \b/n1399 , \b/n1398 , \b/n1397 , \b/n1396 , \b/n1395 ,
         \b/n1394 , \b/n1393 , \b/n1392 , \b/n1391 , \b/n1390 , \b/n1389 ,
         \b/n1388 , \b/n1387 , \b/n1386 , \b/n1385 , \b/n1384 , \b/n1383 ,
         \b/n1382 , \b/n1381 , \b/n1380 , \b/n1379 , \b/n1378 , \b/n1377 ,
         \b/n1376 , \b/n1375 , \b/n1374 , \b/n1373 , \b/n1372 , \b/n1371 ,
         \b/n1370 , \b/n1369 , \b/n1368 , \b/n1367 , \b/n1366 , \b/n1365 ,
         \b/n1364 , \b/n1363 , \b/n1362 , \b/n1361 , \b/n1360 , \b/n1359 ,
         \b/n1358 , \b/n1357 , \b/n1356 , \b/n1355 , \b/n1354 , \b/n1353 ,
         \b/n1352 , \b/n1351 , \b/n1350 , \b/n1349 , \b/n1348 , \b/n1347 ,
         \b/n1346 , \b/n1345 , \b/n1344 , \b/n1343 , \b/n1342 , \b/n1341 ,
         \b/n1340 , \b/n1339 , \b/n1338 , \b/n1337 , \b/n1336 , \b/n1335 ,
         \b/n1334 , \b/n1333 , \b/n1332 , \b/n1331 , \b/n1330 , \b/n1329 ,
         \b/n1328 , \b/n1327 , \b/n1326 , \b/n1325 , \b/n1324 , \b/n1323 ,
         \b/n1322 , \b/n1321 , \b/n1320 , \b/n1319 , \b/n1318 , \b/n1317 ,
         \b/n1316 , \b/n1315 , \b/n1314 , \b/n1313 , \b/n1312 , \b/n1311 ,
         \b/n1310 , \b/n1309 , \b/n1308 , \b/n1307 , \b/n1306 , \b/n1305 ,
         \b/n1304 , \b/n1303 , \b/n1302 , \b/n1301 , \b/n1300 , \b/n1299 ,
         \b/n1298 , \b/n1297 , \b/n1296 , \b/n1295 , \b/n1294 , \b/n1293 ,
         \b/n1292 , \b/n1291 , \b/n1290 , \b/n1289 , \b/n1288 , \b/n1287 ,
         \b/n1286 , \b/n1285 , \b/n1284 , \b/n1283 , \b/n1282 , \b/n1281 ,
         \b/n1280 , \b/n1279 , \b/n1278 , \b/n1277 , \b/n1276 , \b/n1275 ,
         \b/n1274 , \b/n1273 , \b/n1272 , \b/n1271 , \b/n1270 , \b/n1269 ,
         \b/n1268 , \b/n1267 , \b/n1266 , \b/n1265 , \b/n1264 , \b/n1263 ,
         \b/n1262 , \b/n1261 , \b/n1260 , \b/n1259 , \b/n1258 , \b/n1257 ,
         \b/n1256 , \b/n1255 , \b/n1254 , \b/n1253 , \b/n1252 , \b/n1251 ,
         \b/n1250 , \b/n1249 , \b/n1248 , \b/n1247 , \b/n1246 , \b/n1245 ,
         \b/n1244 , \b/n1243 , \b/n1242 , \b/n1241 , \b/n1240 , \b/n1239 ,
         \b/n1238 , \b/n1237 , \b/n1236 , \b/n1235 , \b/n1234 , \b/n1233 ,
         \b/n1232 , \b/n1231 , \b/n1230 , \b/n1229 , \b/n1228 , \b/n1227 ,
         \b/n1226 , \b/n1225 , \b/n1224 , \b/n1223 , \b/n1222 , \b/n1221 ,
         \b/n1220 , \b/n1219 , \b/n1218 , \b/n1217 , \b/n1216 , \b/n1215 ,
         \b/n1214 , \b/n1213 , \b/n1212 , \b/n1211 , \b/n1210 , \b/n1209 ,
         \b/n1208 , \b/n1207 , \b/n1206 , \b/n1205 , \b/n1204 , \b/n1203 ,
         \b/n1202 , \b/n1201 , \b/n1200 , \b/n1199 , \b/n1198 , \b/n1197 ,
         \b/n1196 , \b/n1195 , \b/n1194 , \b/n1193 , \b/n1192 , \b/n1191 ,
         \b/n1190 , \b/n1189 , \b/n1188 , \b/n1187 , \b/n1186 , \b/n1185 ,
         \b/n1184 , \b/n1183 , \b/n1182 , \b/n1181 , \b/n1180 , \b/n1179 ,
         \b/n1178 , \b/n1177 , \b/n1176 , \b/n1174 , \b/n1173 , \b/n1172 ,
         \b/n1171 , \b/n1170 , \b/n1168 , \b/n1167 , \b/n1166 , \b/n1165 ,
         \b/n1164 , \b/n1163 , \b/n1162 , \b/n1161 , \b/n1160 , \b/n1159 ,
         \b/n1158 , \b/n1156 , \b/n1155 , \b/n1154 , \b/n1152 , \b/n1151 ,
         \b/n1150 , \b/n1149 , \b/n1148 , \b/n1147 , \b/n1146 , \b/n1145 ,
         \b/n1144 , \b/n1143 , \b/n1142 , \b/n1141 , \b/n1140 , \b/n1139 ,
         \b/n1138 , \b/n1137 , \b/n1136 , \b/n1135 , \b/n1134 , \b/n1132 ,
         \b/n1131 , \b/n1130 , \b/n1129 , \b/n1128 , \b/n1127 , \b/n1126 ,
         \b/n1125 , \b/n1124 , \b/n1123 , \b/n1122 , \b/n1121 , \b/n1120 ,
         \b/n1119 , \b/n1118 , \b/n1117 , \b/n1116 , \b/n1114 , \b/n1113 ,
         \b/n1112 , \b/n1111 , \b/n1110 , \b/n1109 , \b/n1108 , \b/n1106 ,
         \b/n1105 , \b/n1104 , \b/n1102 , \b/n1101 , \b/n1099 , \b/n1098 ,
         \b/n1095 , \b/n1094 , \b/n1093 , \b/n1092 , \b/n1091 , \b/n1090 ,
         \b/n1087 , \b/n1086 , \b/n1085 , \b/n1084 , \b/n1082 , \b/n1080 ,
         \b/n1079 , \b/n1078 , \b/n1077 , \b/n1076 , \b/n1074 , \b/n1073 ,
         \b/n1072 , \b/n1070 , \b/n1069 , \b/n1067 , \b/n1066 , \b/n1065 ,
         \b/n1063 , \b/n1061 , \b/n1060 , \b/n1059 , \b/n1058 , \b/n1056 ,
         \b/n1055 , \b/n1054 , \b/n1053 , \b/n1052 , \b/n1050 , \b/n1049 ,
         \b/n1048 , \b/n1047 , \b/n1046 , \b/n1045 , \b/n1043 , \b/n1042 ,
         \b/n1041 , \b/n1040 , \b/n1039 , \b/n1038 , \b/n1036 , \b/n1035 ,
         \b/n1034 , \b/n1033 , \b/n1032 , \b/n1031 , \b/n1030 , \b/n1029 ,
         \b/n1027 , \b/n1026 , \b/n1023 , \b/n1022 , \b/n1021 , \b/n1020 ,
         \b/n1019 , \b/n1018 , \b/n1015 , \b/n1014 , \b/n1013 , \b/n1012 ,
         \b/n1010 , \b/n1009 , \b/n1008 , \b/n1007 , \b/n1006 , \b/n1004 ,
         \b/n1003 , \b/n1002 , \b/n1000 , \b/n999 , \b/n997 , \b/n996 ,
         \b/n995 , \b/n993 , \b/n991 , \b/n990 , \b/n989 , \b/n988 , \b/n987 ,
         \b/n986 , \b/n985 , \b/n984 , \b/n983 , \b/n982 , \b/n981 , \b/n980 ,
         \b/n979 , \b/n978 , \b/n977 , \b/n976 , \b/n975 , \b/n973 , \b/n972 ,
         \b/n971 , \b/n970 , \b/n969 , \b/n968 , \b/n967 , \b/n965 , \b/n964 ,
         \b/n963 , \b/n961 , \b/n960 , \b/n958 , \b/n957 , \b/n954 , \b/n953 ,
         \b/n952 , \b/n951 , \b/n950 , \b/n949 , \b/n946 , \b/n945 , \b/n944 ,
         \b/n943 , \b/n941 , \b/n939 , \b/n938 , \b/n937 , \b/n936 , \b/n935 ,
         \b/n933 , \b/n932 , \b/n931 , \b/n929 , \b/n928 , \b/n926 , \b/n925 ,
         \b/n924 , \b/n922 , \b/n920 , \b/n919 , \b/n918 , \b/n917 , \b/n916 ,
         \b/n915 , \b/n914 , \b/n913 , \b/n912 , \b/n911 , \b/n910 , \b/n909 ,
         \b/n908 , \b/n907 , \b/n906 , \b/n905 , \b/n904 , \b/n902 , \b/n901 ,
         \b/n900 , \b/n899 , \b/n898 , \b/n897 , \b/n896 , \b/n894 , \b/n893 ,
         \b/n892 , \b/n890 , \b/n889 , \b/n887 , \b/n886 , \b/n883 , \b/n882 ,
         \b/n881 , \b/n880 , \b/n879 , \b/n878 , \b/n875 , \b/n874 , \b/n873 ,
         \b/n872 , \b/n870 , \b/n868 , \b/n867 , \b/n866 , \b/n865 , \b/n864 ,
         \b/n862 , \b/n861 , \b/n860 , \b/n858 , \b/n857 , \b/n855 , \b/n854 ,
         \b/n853 , \b/n851 , \b/n849 , \b/n848 , \b/n847 , \b/n846 , \b/n845 ,
         \b/n844 , \b/n843 , \b/n842 , \b/n841 , \b/n840 , \b/n839 , \b/n838 ,
         \b/n837 , \b/n836 , \b/n835 , \b/n834 , \b/n833 , \b/n831 , \b/n830 ,
         \b/n829 , \b/n828 , \b/n827 , \b/n826 , \b/n825 , \b/n823 , \b/n822 ,
         \b/n821 , \b/n819 , \b/n818 , \b/n816 , \b/n815 , \b/n812 , \b/n811 ,
         \b/n810 , \b/n809 , \b/n808 , \b/n807 , \b/n804 , \b/n803 , \b/n802 ,
         \b/n801 , \b/n799 , \b/n797 , \b/n796 , \b/n795 , \b/n794 , \b/n793 ,
         \b/n791 , \b/n790 , \b/n789 , \b/n787 , \b/n786 , \b/n784 , \b/n783 ,
         \b/n782 , \b/n780 , \b/n778 , \b/n777 , \b/n776 , \b/n775 , \b/n774 ,
         \b/n773 , \b/n772 , \b/n771 , \b/n770 , \b/n769 , \b/n768 , \b/n767 ,
         \b/n766 , \b/n765 , \b/n764 , \b/n763 , \b/n762 , \b/n760 , \b/n759 ,
         \b/n758 , \b/n757 , \b/n756 , \b/n755 , \b/n754 , \b/n752 , \b/n751 ,
         \b/n750 , \b/n748 , \b/n747 , \b/n745 , \b/n744 , \b/n741 , \b/n740 ,
         \b/n739 , \b/n738 , \b/n737 , \b/n736 , \b/n733 , \b/n732 , \b/n731 ,
         \b/n730 , \b/n728 , \b/n726 , \b/n725 , \b/n724 , \b/n723 , \b/n722 ,
         \b/n720 , \b/n719 , \b/n718 , \b/n716 , \b/n715 , \b/n713 , \b/n712 ,
         \b/n711 , \b/n709 , \b/n707 , \b/n706 , \b/n705 , \b/n704 , \b/n703 ,
         \b/n702 , \b/n701 , \b/n700 , \b/n699 , \b/n698 , \b/n697 , \b/n696 ,
         \b/n695 , \b/n694 , \b/n693 , \b/n692 , \b/n691 , \b/n689 , \b/n688 ,
         \b/n687 , \b/n686 , \b/n685 , \b/n684 , \b/n683 , \b/n681 , \b/n680 ,
         \b/n679 , \b/n677 , \b/n676 , \b/n674 , \b/n673 , \b/n670 , \b/n669 ,
         \b/n668 , \b/n667 , \b/n666 , \b/n665 , \b/n662 , \b/n661 , \b/n660 ,
         \b/n659 , \b/n657 , \b/n655 , \b/n654 , \b/n653 , \b/n652 , \b/n651 ,
         \b/n649 , \b/n648 , \b/n647 , \b/n645 , \b/n644 , \b/n642 , \b/n641 ,
         \b/n640 , \b/n638 , \b/n636 , \b/n635 , \b/n634 , \b/n633 , \b/n632 ,
         \b/n631 , \b/n630 , \b/n629 , \b/n628 , \b/n627 , \b/n626 , \b/n625 ,
         \b/n624 , \b/n623 , \b/n622 , \b/n621 , \b/n620 , \b/n618 , \b/n617 ,
         \b/n616 , \b/n615 , \b/n614 , \b/n613 , \b/n612 , \b/n610 , \b/n609 ,
         \b/n608 , \b/n606 , \b/n605 , \b/n603 , \b/n602 , \b/n599 , \b/n598 ,
         \b/n597 , \b/n596 , \b/n595 , \b/n594 , \b/n591 , \b/n590 , \b/n589 ,
         \b/n588 , \b/n586 , \b/n584 , \b/n583 , \b/n582 , \b/n581 , \b/n580 ,
         \b/n578 , \b/n577 , \b/n576 , \b/n574 , \b/n573 , \b/n571 , \b/n570 ,
         \b/n569 , \b/n567 , \b/n565 , \b/n564 , \b/n563 , \b/n562 , \b/n561 ,
         \b/n560 , \b/n559 , \b/n558 , \b/n557 , \b/n556 , \b/n555 , \b/n554 ,
         \b/n553 , \b/n552 , \b/n551 , \b/n550 , \b/n549 , \b/n547 , \b/n546 ,
         \b/n545 , \b/n544 , \b/n543 , \b/n542 , \b/n541 , \b/n539 , \b/n538 ,
         \b/n537 , \b/n535 , \b/n534 , \b/n532 , \b/n531 , \b/n528 , \b/n527 ,
         \b/n526 , \b/n525 , \b/n524 , \b/n523 , \b/n520 , \b/n519 , \b/n518 ,
         \b/n517 , \b/n515 , \b/n513 , \b/n512 , \b/n511 , \b/n510 , \b/n509 ,
         \b/n507 , \b/n506 , \b/n505 , \b/n503 , \b/n502 , \b/n500 , \b/n499 ,
         \b/n498 , \b/n496 , \b/n494 , \b/n493 , \b/n492 , \b/n491 , \b/n490 ,
         \b/n489 , \b/n488 , \b/n487 , \b/n486 , \b/n485 , \b/n484 , \b/n483 ,
         \b/n482 , \b/n481 , \b/n480 , \b/n479 , \b/n478 , \b/n476 , \b/n475 ,
         \b/n474 , \b/n473 , \b/n472 , \b/n471 , \b/n470 , \b/n468 , \b/n467 ,
         \b/n466 , \b/n464 , \b/n463 , \b/n461 , \b/n460 , \b/n457 , \b/n456 ,
         \b/n455 , \b/n454 , \b/n453 , \b/n452 , \b/n449 , \b/n448 , \b/n447 ,
         \b/n446 , \b/n444 , \b/n442 , \b/n441 , \b/n440 , \b/n439 , \b/n438 ,
         \b/n436 , \b/n435 , \b/n434 , \b/n432 , \b/n431 , \b/n429 , \b/n428 ,
         \b/n427 , \b/n425 , \b/n423 , \b/n422 , \b/n421 , \b/n420 , \b/n419 ,
         \b/n418 , \b/n417 , \b/n416 , \b/n415 , \b/n414 , \b/n413 , \b/n412 ,
         \b/n411 , \b/n410 , \b/n409 , \b/n408 , \b/n407 , \b/n405 , \b/n404 ,
         \b/n403 , \b/n402 , \b/n401 , \b/n400 , \b/n399 , \b/n397 , \b/n396 ,
         \b/n395 , \b/n393 , \b/n392 , \b/n390 , \b/n389 , \b/n386 , \b/n385 ,
         \b/n384 , \b/n383 , \b/n382 , \b/n381 , \b/n378 , \b/n377 , \b/n376 ,
         \b/n375 , \b/n373 , \b/n371 , \b/n370 , \b/n369 , \b/n368 , \b/n367 ,
         \b/n365 , \b/n364 , \b/n363 , \b/n361 , \b/n360 , \b/n358 , \b/n357 ,
         \b/n356 , \b/n354 , \b/n352 , \b/n351 , \b/n350 , \b/n349 , \b/n348 ,
         \b/n347 , \b/n346 , \b/n345 , \b/n344 , \b/n343 , \b/n342 , \b/n341 ,
         \b/n340 , \b/n339 , \b/n338 , \b/n337 , \b/n336 , \b/n334 , \b/n333 ,
         \b/n332 , \b/n331 , \b/n330 , \b/n329 , \b/n328 , \b/n326 , \b/n325 ,
         \b/n324 , \b/n322 , \b/n321 , \b/n319 , \b/n318 , \b/n315 , \b/n314 ,
         \b/n313 , \b/n312 , \b/n311 , \b/n310 , \b/n307 , \b/n306 , \b/n305 ,
         \b/n304 , \b/n302 , \b/n300 , \b/n299 , \b/n298 , \b/n297 , \b/n296 ,
         \b/n294 , \b/n293 , \b/n292 , \b/n290 , \b/n289 , \b/n287 , \b/n286 ,
         \b/n285 , \b/n283 , \b/n281 , \b/n280 , \b/n279 , \b/n278 , \b/n277 ,
         \b/n276 , \b/n275 , \b/n274 , \b/n273 , \b/n272 , \b/n271 , \b/n270 ,
         \b/n269 , \b/n266 , \b/n265 , \b/n264 , \b/n262 , \b/n260 , \b/n259 ,
         \b/n258 , \b/n257 , \b/n256 , \b/n255 , \b/n253 , \b/n251 , \b/n250 ,
         \b/n249 , \b/n248 , \b/n247 , \b/n244 , \b/n243 , \b/n242 , \b/n241 ,
         \b/n240 , \b/n239 , \b/n238 , \b/n237 , \b/n236 , \b/n235 , \b/n233 ,
         \b/n232 , \b/n229 , \b/n228 , \b/n227 , \b/n226 , \b/n225 , \b/n224 ,
         \b/n221 , \b/n220 , \b/n219 , \b/n218 , \b/n217 , \b/n216 , \b/n215 ,
         \b/n213 , \b/n211 , \b/n210 , \b/n209 , \b/n208 , \b/n207 , \b/n206 ,
         \b/n205 , \b/n204 , \b/n203 , \b/n202 , \b/n201 , \b/n200 , \b/n199 ,
         \b/n198 , \b/n197 , \b/n196 , \b/n195 , \b/n193 , \b/n192 , \b/n191 ,
         \b/n190 , \b/n189 , \b/n188 , \b/n187 , \b/n185 , \b/n184 , \b/n183 ,
         \b/n181 , \b/n180 , \b/n178 , \b/n177 , \b/n174 , \b/n173 , \b/n172 ,
         \b/n171 , \b/n170 , \b/n169 , \b/n166 , \b/n165 , \b/n164 , \b/n163 ,
         \b/n161 , \b/n159 , \b/n158 , \b/n157 , \b/n156 , \b/n155 , \b/n153 ,
         \b/n152 , \b/n151 , \b/n149 , \b/n148 , \b/n146 , \b/n145 , \b/n144 ,
         \b/n142 , \b/n140 , \b/n139 , \b/n138 , \b/n137 , \b/n136 , \b/n135 ,
         \b/n134 , \b/n133 , \b/n132 , \b/n131 , \b/n130 , \b/n129 , \b/n128 ,
         \b/n127 , \b/n126 , \b/n125 , \b/n124 , \b/n122 , \b/n121 , \b/n120 ,
         \b/n119 , \b/n118 , \b/n117 , \b/n116 , \b/n114 , \b/n113 , \b/n112 ,
         \b/n110 , \b/n109 , \b/n107 , \b/n106 , \b/n103 , \b/n102 , \b/n101 ,
         \b/n100 , \b/n99 , \b/n98 , \b/n95 , \b/n94 , \b/n93 , \b/n92 ,
         \b/n90 , \b/n88 , \b/n87 , \b/n86 , \b/n85 , \b/n84 , \b/n82 ,
         \b/n81 , \b/n80 , \b/n78 , \b/n77 , \b/n75 , \b/n74 , \b/n73 ,
         \b/n71 , \b/n69 , \b/n68 , \b/n67 , \b/n66 , \b/n65 , \b/n64 ,
         \b/n63 , \b/n62 , \b/n61 , \b/n60 , \b/n59 , \b/n58 , \b/n57 ,
         \b/n56 , \b/n55 , \b/n54 , \b/n53 , \b/n51 , \b/n50 , \b/n49 ,
         \b/n48 , \b/n47 , \b/n46 , \b/n45 , \b/n43 , \b/n42 , \b/n41 ,
         \b/n39 , \b/n38 , \b/n36 , \b/n35 , \b/n32 , \b/n31 , \b/n30 ,
         \b/n29 , \b/n28 , \b/n27 , \b/n24 , \b/n23 , \b/n22 , \b/n21 ,
         \b/n19 , \b/n17 , \b/n16 , \b/n15 , \b/n14 , \b/n13 , \b/n11 ,
         \b/n10 , \b/n9 , \b/n7 , \b/n6 , \b/n4 , \b/n3 , \b/n2 , \d/n468 ,
         \d/n467 , \d/n466 , \d/n465 , \d/n464 , \d/n463 , \d/n462 , \d/n461 ,
         \d/n460 , \d/n459 , \d/n458 , \d/n457 , \d/n456 , \d/n455 , \d/n454 ,
         \d/n453 , \d/n452 , \d/n451 , \d/n450 , \d/n449 , \d/n448 , \d/n447 ,
         \d/n446 , \d/n445 , \d/n444 , \d/n443 , \d/n442 , \d/n441 , \d/n440 ,
         \d/n439 , \d/n438 , \d/n437 , \d/n436 , \d/n435 , \d/n434 , \d/n433 ,
         \d/n432 , \d/n431 , \d/n430 , \d/n429 , \d/n428 , \d/n427 , \d/n426 ,
         \d/n425 , \d/n424 , \d/n423 , \d/n422 , \d/n421 , \d/n420 , \d/n419 ,
         \d/n418 , \d/n417 , \d/n416 , \d/n415 , \d/n414 , \d/n413 , \d/n412 ,
         \d/n411 , \d/n410 , \d/n409 , \d/n408 , \d/n407 , \d/n406 , \d/n405 ,
         \d/n404 , \d/n403 , \d/n402 , \d/n401 , \d/n400 , \d/n399 , \d/n398 ,
         \d/n397 , \d/n396 , \d/n395 , \d/n394 , \d/n393 , \d/n392 , \d/n391 ,
         \d/n390 , \d/n389 , \d/n388 , \d/n387 , \d/n386 , \d/n385 , \d/n384 ,
         \d/n383 , \d/n382 , \d/n381 , \d/n380 , \d/n379 , \d/n378 , \d/n377 ,
         \d/n376 , \d/n375 , \d/n374 , \d/n373 , \d/n372 , \d/n371 , \d/n370 ,
         \d/n369 , \d/n368 , \d/n367 , \d/n366 , \d/n365 , \d/n364 , \d/n363 ,
         \d/n362 , \d/n361 , \d/n360 , \d/n359 , \d/n358 , \d/n357 , \d/n356 ,
         \d/n355 , \d/n354 , \d/n353 , \d/n352 , \d/n351 , \d/n350 , \d/n349 ,
         \d/n348 , \d/n347 , \d/n346 , \d/n345 , \d/n344 , \d/n343 , \d/n342 ,
         \d/n341 , \d/n340 , \d/n339 , \d/n338 , \d/n337 , \d/n336 , \d/n335 ,
         \d/n334 , \d/n333 , \d/n332 , \d/n331 , \d/n330 , \d/n329 , \d/n328 ,
         \d/n327 , \d/n326 , \d/n325 , \d/n324 , \d/n323 , \d/n322 , \d/n321 ,
         \d/n320 , \d/n319 , \d/n318 , \d/n317 , \d/n316 , \d/n315 , \d/n314 ,
         \d/n313 , \d/n312 , \d/n311 , \d/n310 , \d/n309 , \d/n308 , \d/n307 ,
         \d/n306 , \d/n305 , \d/n304 , \d/n303 , \d/n302 , \d/n301 , \d/n300 ,
         \d/n299 , \d/n298 , \d/n297 , \d/n296 , \d/n295 , \d/n294 , \d/n293 ,
         \d/n292 , \d/n291 , \d/n290 , \d/n289 , \d/n288 , \d/n287 , \d/n286 ,
         \d/n285 , \d/n284 , \d/n283 , \d/n282 , \d/n281 , \d/n280 , \d/n279 ,
         \d/n278 , \d/n277 , \d/n276 , \d/n275 , \d/n274 , \d/n273 , \d/n272 ,
         \d/n271 , \d/n270 , \d/n269 , \d/n268 , \d/n267 , \d/n266 , \d/n265 ,
         \d/n264 , \d/n263 , \d/n262 , \d/n261 , \d/n260 , \d/n259 , \d/n258 ,
         \d/n257 , \d/n256 , \d/n255 , \d/n254 , \d/n253 , \d/n252 , \d/n251 ,
         \d/n250 , \d/n249 , \d/n248 , \d/n247 , \d/n246 , \d/n245 , \d/n244 ,
         \d/n243 , \d/n242 , \d/n241 , \d/n240 , \d/n239 , \d/n238 , \d/n237 ,
         \d/n236 , \d/n235 , \d/n234 , \d/n233 , \d/n232 , \d/n231 , \d/n230 ,
         \d/n229 , \d/n228 , \d/n227 , \d/n226 , \d/n225 , \d/n224 , \d/n223 ,
         \d/n222 , \d/n221 , \d/n220 , \d/n219 , \d/n218 , \d/n217 , \d/n216 ,
         \d/n215 , \d/n214 , \d/n213 , \d/n212 , \d/n211 , \d/n210 , \d/n209 ,
         \d/n208 , \d/n207 , \d/n206 , \d/n205 , \d/n204 , \d/n203 , \d/n202 ,
         \d/n201 , \d/n200 , \d/n199 , \d/n198 , \d/n197 , \d/n196 , \d/n195 ,
         \d/n194 , \d/n193 , \d/n192 , \d/n191 , \d/n190 , \d/n189 , \d/n188 ,
         \d/n187 , \d/n186 , \d/n185 , \d/n184 , \d/n183 , \d/n182 , \d/n181 ,
         \d/n180 , \d/n179 , \d/n178 , \d/n177 , \d/n176 , \d/n175 , \d/n174 ,
         \d/n173 , \d/n172 , \d/n171 , \d/n170 , \d/n169 , \d/n168 , \d/n167 ,
         \d/n166 , \d/n165 , \d/n164 , \d/n163 , \d/n162 , \d/n161 , \d/n160 ,
         \d/n159 , \d/n158 , \d/n157 , \d/n156 , \d/n155 , \d/n154 , \d/n153 ,
         \d/n152 , \d/n151 , \d/n150 , \d/n149 , \d/n148 , \d/n147 , \d/n146 ,
         \d/n145 , \d/n144 , \d/n143 , \d/n142 , \d/n141 , \d/n140 , \d/n139 ,
         \d/n138 , \d/n137 , \d/n136 , \d/n135 , \d/n134 , \d/n133 , \d/n132 ,
         \d/n131 , \d/n130 , \d/n129 , \d/n128 , \d/n127 , \d/n126 , \d/n125 ,
         \d/n124 , \d/n123 , \d/n122 , \d/n121 , \d/n120 , \d/n119 , \d/n118 ,
         \d/n117 , n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082;
  wire   [127:0] key;
  wire   [3:0] counter;
  wire   [127:0] nextKey;
  wire   [127:0] msg;
  wire   [127:0] mix_col_out;
  wire   [127:0] shift_row_out;

  DFF \counter_reg[0]  ( .D(n7), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[0]) );
  DFF \counter_reg[1]  ( .D(N5), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[1]) );
  DFF \counter_reg[2]  ( .D(N6), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[2]) );
  DFF \counter_reg[3]  ( .D(N7), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[3]) );
  DFF \key_reg[0]  ( .D(nextKey[0]), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(
        key[0]) );
  DFF \key_reg[1]  ( .D(nextKey[1]), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(
        key[1]) );
  DFF \key_reg[2]  ( .D(nextKey[2]), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(
        key[2]) );
  DFF \key_reg[3]  ( .D(nextKey[3]), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(
        key[3]) );
  DFF \key_reg[4]  ( .D(nextKey[4]), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(
        key[4]) );
  DFF \key_reg[5]  ( .D(nextKey[5]), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(
        key[5]) );
  DFF \key_reg[6]  ( .D(nextKey[6]), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(
        key[6]) );
  DFF \key_reg[7]  ( .D(nextKey[7]), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(
        key[7]) );
  DFF \key_reg[8]  ( .D(nextKey[8]), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(
        key[8]) );
  DFF \key_reg[9]  ( .D(nextKey[9]), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(
        key[9]) );
  DFF \key_reg[10]  ( .D(nextKey[10]), .CLK(clk), .RST(rst), .I(g_init[10]), 
        .Q(key[10]) );
  DFF \key_reg[11]  ( .D(nextKey[11]), .CLK(clk), .RST(rst), .I(g_init[11]), 
        .Q(key[11]) );
  DFF \key_reg[12]  ( .D(nextKey[12]), .CLK(clk), .RST(rst), .I(g_init[12]), 
        .Q(key[12]) );
  DFF \key_reg[13]  ( .D(nextKey[13]), .CLK(clk), .RST(rst), .I(g_init[13]), 
        .Q(key[13]) );
  DFF \key_reg[14]  ( .D(nextKey[14]), .CLK(clk), .RST(rst), .I(g_init[14]), 
        .Q(key[14]) );
  DFF \key_reg[15]  ( .D(nextKey[15]), .CLK(clk), .RST(rst), .I(g_init[15]), 
        .Q(key[15]) );
  DFF \key_reg[16]  ( .D(nextKey[16]), .CLK(clk), .RST(rst), .I(g_init[16]), 
        .Q(key[16]) );
  DFF \key_reg[17]  ( .D(nextKey[17]), .CLK(clk), .RST(rst), .I(g_init[17]), 
        .Q(key[17]) );
  DFF \key_reg[18]  ( .D(nextKey[18]), .CLK(clk), .RST(rst), .I(g_init[18]), 
        .Q(key[18]) );
  DFF \key_reg[19]  ( .D(nextKey[19]), .CLK(clk), .RST(rst), .I(g_init[19]), 
        .Q(key[19]) );
  DFF \key_reg[20]  ( .D(nextKey[20]), .CLK(clk), .RST(rst), .I(g_init[20]), 
        .Q(key[20]) );
  DFF \key_reg[21]  ( .D(nextKey[21]), .CLK(clk), .RST(rst), .I(g_init[21]), 
        .Q(key[21]) );
  DFF \key_reg[22]  ( .D(nextKey[22]), .CLK(clk), .RST(rst), .I(g_init[22]), 
        .Q(key[22]) );
  DFF \key_reg[23]  ( .D(nextKey[23]), .CLK(clk), .RST(rst), .I(g_init[23]), 
        .Q(key[23]) );
  DFF \key_reg[24]  ( .D(nextKey[24]), .CLK(clk), .RST(rst), .I(g_init[24]), 
        .Q(key[24]) );
  DFF \key_reg[25]  ( .D(nextKey[25]), .CLK(clk), .RST(rst), .I(g_init[25]), 
        .Q(key[25]) );
  DFF \key_reg[26]  ( .D(nextKey[26]), .CLK(clk), .RST(rst), .I(g_init[26]), 
        .Q(key[26]) );
  DFF \key_reg[27]  ( .D(nextKey[27]), .CLK(clk), .RST(rst), .I(g_init[27]), 
        .Q(key[27]) );
  DFF \key_reg[28]  ( .D(nextKey[28]), .CLK(clk), .RST(rst), .I(g_init[28]), 
        .Q(key[28]) );
  DFF \key_reg[29]  ( .D(nextKey[29]), .CLK(clk), .RST(rst), .I(g_init[29]), 
        .Q(key[29]) );
  DFF \key_reg[30]  ( .D(nextKey[30]), .CLK(clk), .RST(rst), .I(g_init[30]), 
        .Q(key[30]) );
  DFF \key_reg[31]  ( .D(nextKey[31]), .CLK(clk), .RST(rst), .I(g_init[31]), 
        .Q(key[31]) );
  DFF \key_reg[32]  ( .D(nextKey[32]), .CLK(clk), .RST(rst), .I(g_init[32]), 
        .Q(key[32]) );
  DFF \key_reg[33]  ( .D(nextKey[33]), .CLK(clk), .RST(rst), .I(g_init[33]), 
        .Q(key[33]) );
  DFF \key_reg[34]  ( .D(nextKey[34]), .CLK(clk), .RST(rst), .I(g_init[34]), 
        .Q(key[34]) );
  DFF \key_reg[35]  ( .D(nextKey[35]), .CLK(clk), .RST(rst), .I(g_init[35]), 
        .Q(key[35]) );
  DFF \key_reg[36]  ( .D(nextKey[36]), .CLK(clk), .RST(rst), .I(g_init[36]), 
        .Q(key[36]) );
  DFF \key_reg[37]  ( .D(nextKey[37]), .CLK(clk), .RST(rst), .I(g_init[37]), 
        .Q(key[37]) );
  DFF \key_reg[38]  ( .D(nextKey[38]), .CLK(clk), .RST(rst), .I(g_init[38]), 
        .Q(key[38]) );
  DFF \key_reg[39]  ( .D(nextKey[39]), .CLK(clk), .RST(rst), .I(g_init[39]), 
        .Q(key[39]) );
  DFF \key_reg[40]  ( .D(nextKey[40]), .CLK(clk), .RST(rst), .I(g_init[40]), 
        .Q(key[40]) );
  DFF \key_reg[41]  ( .D(nextKey[41]), .CLK(clk), .RST(rst), .I(g_init[41]), 
        .Q(key[41]) );
  DFF \key_reg[42]  ( .D(nextKey[42]), .CLK(clk), .RST(rst), .I(g_init[42]), 
        .Q(key[42]) );
  DFF \key_reg[43]  ( .D(nextKey[43]), .CLK(clk), .RST(rst), .I(g_init[43]), 
        .Q(key[43]) );
  DFF \key_reg[44]  ( .D(nextKey[44]), .CLK(clk), .RST(rst), .I(g_init[44]), 
        .Q(key[44]) );
  DFF \key_reg[45]  ( .D(nextKey[45]), .CLK(clk), .RST(rst), .I(g_init[45]), 
        .Q(key[45]) );
  DFF \key_reg[46]  ( .D(nextKey[46]), .CLK(clk), .RST(rst), .I(g_init[46]), 
        .Q(key[46]) );
  DFF \key_reg[47]  ( .D(nextKey[47]), .CLK(clk), .RST(rst), .I(g_init[47]), 
        .Q(key[47]) );
  DFF \key_reg[48]  ( .D(nextKey[48]), .CLK(clk), .RST(rst), .I(g_init[48]), 
        .Q(key[48]) );
  DFF \key_reg[49]  ( .D(nextKey[49]), .CLK(clk), .RST(rst), .I(g_init[49]), 
        .Q(key[49]) );
  DFF \key_reg[50]  ( .D(nextKey[50]), .CLK(clk), .RST(rst), .I(g_init[50]), 
        .Q(key[50]) );
  DFF \key_reg[51]  ( .D(nextKey[51]), .CLK(clk), .RST(rst), .I(g_init[51]), 
        .Q(key[51]) );
  DFF \key_reg[52]  ( .D(nextKey[52]), .CLK(clk), .RST(rst), .I(g_init[52]), 
        .Q(key[52]) );
  DFF \key_reg[53]  ( .D(nextKey[53]), .CLK(clk), .RST(rst), .I(g_init[53]), 
        .Q(key[53]) );
  DFF \key_reg[54]  ( .D(nextKey[54]), .CLK(clk), .RST(rst), .I(g_init[54]), 
        .Q(key[54]) );
  DFF \key_reg[55]  ( .D(nextKey[55]), .CLK(clk), .RST(rst), .I(g_init[55]), 
        .Q(key[55]) );
  DFF \key_reg[56]  ( .D(nextKey[56]), .CLK(clk), .RST(rst), .I(g_init[56]), 
        .Q(key[56]) );
  DFF \key_reg[57]  ( .D(nextKey[57]), .CLK(clk), .RST(rst), .I(g_init[57]), 
        .Q(key[57]) );
  DFF \key_reg[58]  ( .D(nextKey[58]), .CLK(clk), .RST(rst), .I(g_init[58]), 
        .Q(key[58]) );
  DFF \key_reg[59]  ( .D(nextKey[59]), .CLK(clk), .RST(rst), .I(g_init[59]), 
        .Q(key[59]) );
  DFF \key_reg[60]  ( .D(nextKey[60]), .CLK(clk), .RST(rst), .I(g_init[60]), 
        .Q(key[60]) );
  DFF \key_reg[61]  ( .D(nextKey[61]), .CLK(clk), .RST(rst), .I(g_init[61]), 
        .Q(key[61]) );
  DFF \key_reg[62]  ( .D(nextKey[62]), .CLK(clk), .RST(rst), .I(g_init[62]), 
        .Q(key[62]) );
  DFF \key_reg[63]  ( .D(nextKey[63]), .CLK(clk), .RST(rst), .I(g_init[63]), 
        .Q(key[63]) );
  DFF \key_reg[64]  ( .D(nextKey[64]), .CLK(clk), .RST(rst), .I(g_init[64]), 
        .Q(key[64]) );
  DFF \key_reg[65]  ( .D(nextKey[65]), .CLK(clk), .RST(rst), .I(g_init[65]), 
        .Q(key[65]) );
  DFF \key_reg[66]  ( .D(nextKey[66]), .CLK(clk), .RST(rst), .I(g_init[66]), 
        .Q(key[66]) );
  DFF \key_reg[67]  ( .D(nextKey[67]), .CLK(clk), .RST(rst), .I(g_init[67]), 
        .Q(key[67]) );
  DFF \key_reg[68]  ( .D(nextKey[68]), .CLK(clk), .RST(rst), .I(g_init[68]), 
        .Q(key[68]) );
  DFF \key_reg[69]  ( .D(nextKey[69]), .CLK(clk), .RST(rst), .I(g_init[69]), 
        .Q(key[69]) );
  DFF \key_reg[70]  ( .D(nextKey[70]), .CLK(clk), .RST(rst), .I(g_init[70]), 
        .Q(key[70]) );
  DFF \key_reg[71]  ( .D(nextKey[71]), .CLK(clk), .RST(rst), .I(g_init[71]), 
        .Q(key[71]) );
  DFF \key_reg[72]  ( .D(nextKey[72]), .CLK(clk), .RST(rst), .I(g_init[72]), 
        .Q(key[72]) );
  DFF \key_reg[73]  ( .D(nextKey[73]), .CLK(clk), .RST(rst), .I(g_init[73]), 
        .Q(key[73]) );
  DFF \key_reg[74]  ( .D(nextKey[74]), .CLK(clk), .RST(rst), .I(g_init[74]), 
        .Q(key[74]) );
  DFF \key_reg[75]  ( .D(nextKey[75]), .CLK(clk), .RST(rst), .I(g_init[75]), 
        .Q(key[75]) );
  DFF \key_reg[76]  ( .D(nextKey[76]), .CLK(clk), .RST(rst), .I(g_init[76]), 
        .Q(key[76]) );
  DFF \key_reg[77]  ( .D(nextKey[77]), .CLK(clk), .RST(rst), .I(g_init[77]), 
        .Q(key[77]) );
  DFF \key_reg[78]  ( .D(nextKey[78]), .CLK(clk), .RST(rst), .I(g_init[78]), 
        .Q(key[78]) );
  DFF \key_reg[79]  ( .D(nextKey[79]), .CLK(clk), .RST(rst), .I(g_init[79]), 
        .Q(key[79]) );
  DFF \key_reg[80]  ( .D(nextKey[80]), .CLK(clk), .RST(rst), .I(g_init[80]), 
        .Q(key[80]) );
  DFF \key_reg[81]  ( .D(nextKey[81]), .CLK(clk), .RST(rst), .I(g_init[81]), 
        .Q(key[81]) );
  DFF \key_reg[82]  ( .D(nextKey[82]), .CLK(clk), .RST(rst), .I(g_init[82]), 
        .Q(key[82]) );
  DFF \key_reg[83]  ( .D(nextKey[83]), .CLK(clk), .RST(rst), .I(g_init[83]), 
        .Q(key[83]) );
  DFF \key_reg[84]  ( .D(nextKey[84]), .CLK(clk), .RST(rst), .I(g_init[84]), 
        .Q(key[84]) );
  DFF \key_reg[85]  ( .D(nextKey[85]), .CLK(clk), .RST(rst), .I(g_init[85]), 
        .Q(key[85]) );
  DFF \key_reg[86]  ( .D(nextKey[86]), .CLK(clk), .RST(rst), .I(g_init[86]), 
        .Q(key[86]) );
  DFF \key_reg[87]  ( .D(nextKey[87]), .CLK(clk), .RST(rst), .I(g_init[87]), 
        .Q(key[87]) );
  DFF \key_reg[88]  ( .D(nextKey[88]), .CLK(clk), .RST(rst), .I(g_init[88]), 
        .Q(key[88]) );
  DFF \key_reg[89]  ( .D(nextKey[89]), .CLK(clk), .RST(rst), .I(g_init[89]), 
        .Q(key[89]) );
  DFF \key_reg[90]  ( .D(nextKey[90]), .CLK(clk), .RST(rst), .I(g_init[90]), 
        .Q(key[90]) );
  DFF \key_reg[91]  ( .D(nextKey[91]), .CLK(clk), .RST(rst), .I(g_init[91]), 
        .Q(key[91]) );
  DFF \key_reg[92]  ( .D(nextKey[92]), .CLK(clk), .RST(rst), .I(g_init[92]), 
        .Q(key[92]) );
  DFF \key_reg[93]  ( .D(nextKey[93]), .CLK(clk), .RST(rst), .I(g_init[93]), 
        .Q(key[93]) );
  DFF \key_reg[94]  ( .D(nextKey[94]), .CLK(clk), .RST(rst), .I(g_init[94]), 
        .Q(key[94]) );
  DFF \key_reg[95]  ( .D(nextKey[95]), .CLK(clk), .RST(rst), .I(g_init[95]), 
        .Q(key[95]) );
  DFF \key_reg[96]  ( .D(n736), .CLK(clk), .RST(rst), .I(g_init[96]), .Q(
        key[96]) );
  DFF \key_reg[97]  ( .D(n735), .CLK(clk), .RST(rst), .I(g_init[97]), .Q(
        key[97]) );
  DFF \key_reg[98]  ( .D(n734), .CLK(clk), .RST(rst), .I(g_init[98]), .Q(
        key[98]) );
  DFF \key_reg[99]  ( .D(n733), .CLK(clk), .RST(rst), .I(g_init[99]), .Q(
        key[99]) );
  DFF \key_reg[100]  ( .D(n732), .CLK(clk), .RST(rst), .I(g_init[100]), .Q(
        key[100]) );
  DFF \key_reg[101]  ( .D(n731), .CLK(clk), .RST(rst), .I(g_init[101]), .Q(
        key[101]) );
  DFF \key_reg[102]  ( .D(n730), .CLK(clk), .RST(rst), .I(g_init[102]), .Q(
        key[102]) );
  DFF \key_reg[103]  ( .D(n729), .CLK(clk), .RST(rst), .I(g_init[103]), .Q(
        key[103]) );
  DFF \key_reg[104]  ( .D(nextKey[104]), .CLK(clk), .RST(rst), .I(g_init[104]), 
        .Q(key[104]) );
  DFF \key_reg[105]  ( .D(nextKey[105]), .CLK(clk), .RST(rst), .I(g_init[105]), 
        .Q(key[105]) );
  DFF \key_reg[106]  ( .D(nextKey[106]), .CLK(clk), .RST(rst), .I(g_init[106]), 
        .Q(key[106]) );
  DFF \key_reg[107]  ( .D(nextKey[107]), .CLK(clk), .RST(rst), .I(g_init[107]), 
        .Q(key[107]) );
  DFF \key_reg[108]  ( .D(nextKey[108]), .CLK(clk), .RST(rst), .I(g_init[108]), 
        .Q(key[108]) );
  DFF \key_reg[109]  ( .D(nextKey[109]), .CLK(clk), .RST(rst), .I(g_init[109]), 
        .Q(key[109]) );
  DFF \key_reg[110]  ( .D(nextKey[110]), .CLK(clk), .RST(rst), .I(g_init[110]), 
        .Q(key[110]) );
  DFF \key_reg[111]  ( .D(nextKey[111]), .CLK(clk), .RST(rst), .I(g_init[111]), 
        .Q(key[111]) );
  DFF \key_reg[112]  ( .D(nextKey[112]), .CLK(clk), .RST(rst), .I(g_init[112]), 
        .Q(key[112]) );
  DFF \key_reg[113]  ( .D(nextKey[113]), .CLK(clk), .RST(rst), .I(g_init[113]), 
        .Q(key[113]) );
  DFF \key_reg[114]  ( .D(nextKey[114]), .CLK(clk), .RST(rst), .I(g_init[114]), 
        .Q(key[114]) );
  DFF \key_reg[115]  ( .D(nextKey[115]), .CLK(clk), .RST(rst), .I(g_init[115]), 
        .Q(key[115]) );
  DFF \key_reg[116]  ( .D(nextKey[116]), .CLK(clk), .RST(rst), .I(g_init[116]), 
        .Q(key[116]) );
  DFF \key_reg[117]  ( .D(nextKey[117]), .CLK(clk), .RST(rst), .I(g_init[117]), 
        .Q(key[117]) );
  DFF \key_reg[118]  ( .D(nextKey[118]), .CLK(clk), .RST(rst), .I(g_init[118]), 
        .Q(key[118]) );
  DFF \key_reg[119]  ( .D(nextKey[119]), .CLK(clk), .RST(rst), .I(g_init[119]), 
        .Q(key[119]) );
  DFF \key_reg[120]  ( .D(nextKey[120]), .CLK(clk), .RST(rst), .I(g_init[120]), 
        .Q(key[120]) );
  DFF \key_reg[121]  ( .D(nextKey[121]), .CLK(clk), .RST(rst), .I(g_init[121]), 
        .Q(key[121]) );
  DFF \key_reg[122]  ( .D(nextKey[122]), .CLK(clk), .RST(rst), .I(g_init[122]), 
        .Q(key[122]) );
  DFF \key_reg[123]  ( .D(nextKey[123]), .CLK(clk), .RST(rst), .I(g_init[123]), 
        .Q(key[123]) );
  DFF \key_reg[124]  ( .D(nextKey[124]), .CLK(clk), .RST(rst), .I(g_init[124]), 
        .Q(key[124]) );
  DFF \key_reg[125]  ( .D(nextKey[125]), .CLK(clk), .RST(rst), .I(g_init[125]), 
        .Q(key[125]) );
  DFF \key_reg[126]  ( .D(nextKey[126]), .CLK(clk), .RST(rst), .I(g_init[126]), 
        .Q(key[126]) );
  DFF \key_reg[127]  ( .D(nextKey[127]), .CLK(clk), .RST(rst), .I(g_init[127]), 
        .Q(key[127]) );
  DFF \msg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(e_init[0]), .Q(msg[0])
         );
  DFF \msg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(e_init[1]), .Q(msg[1])
         );
  DFF \msg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(e_init[2]), .Q(msg[2])
         );
  DFF \msg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(e_init[3]), .Q(msg[3])
         );
  DFF \msg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(e_init[4]), .Q(msg[4])
         );
  DFF \msg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(e_init[5]), .Q(msg[5])
         );
  DFF \msg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(e_init[6]), .Q(msg[6])
         );
  DFF \msg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(e_init[7]), .Q(msg[7])
         );
  DFF \msg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(e_init[8]), .Q(msg[8])
         );
  DFF \msg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(e_init[9]), .Q(msg[9])
         );
  DFF \msg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(e_init[10]), .Q(
        msg[10]) );
  DFF \msg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(e_init[11]), .Q(
        msg[11]) );
  DFF \msg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(e_init[12]), .Q(
        msg[12]) );
  DFF \msg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(e_init[13]), .Q(
        msg[13]) );
  DFF \msg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(e_init[14]), .Q(
        msg[14]) );
  DFF \msg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(e_init[15]), .Q(
        msg[15]) );
  DFF \msg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(e_init[16]), .Q(
        msg[16]) );
  DFF \msg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(e_init[17]), .Q(
        msg[17]) );
  DFF \msg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(e_init[18]), .Q(
        msg[18]) );
  DFF \msg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(e_init[19]), .Q(
        msg[19]) );
  DFF \msg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(e_init[20]), .Q(
        msg[20]) );
  DFF \msg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(e_init[21]), .Q(
        msg[21]) );
  DFF \msg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(e_init[22]), .Q(
        msg[22]) );
  DFF \msg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(e_init[23]), .Q(
        msg[23]) );
  DFF \msg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(e_init[24]), .Q(
        msg[24]) );
  DFF \msg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(e_init[25]), .Q(
        msg[25]) );
  DFF \msg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(e_init[26]), .Q(
        msg[26]) );
  DFF \msg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(e_init[27]), .Q(
        msg[27]) );
  DFF \msg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(e_init[28]), .Q(
        msg[28]) );
  DFF \msg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(e_init[29]), .Q(
        msg[29]) );
  DFF \msg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(e_init[30]), .Q(
        msg[30]) );
  DFF \msg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(e_init[31]), .Q(
        msg[31]) );
  DFF \msg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(e_init[32]), .Q(
        msg[32]) );
  DFF \msg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(e_init[33]), .Q(
        msg[33]) );
  DFF \msg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(e_init[34]), .Q(
        msg[34]) );
  DFF \msg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(e_init[35]), .Q(
        msg[35]) );
  DFF \msg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(e_init[36]), .Q(
        msg[36]) );
  DFF \msg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(e_init[37]), .Q(
        msg[37]) );
  DFF \msg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(e_init[38]), .Q(
        msg[38]) );
  DFF \msg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(e_init[39]), .Q(
        msg[39]) );
  DFF \msg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(e_init[40]), .Q(
        msg[40]) );
  DFF \msg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(e_init[41]), .Q(
        msg[41]) );
  DFF \msg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(e_init[42]), .Q(
        msg[42]) );
  DFF \msg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(e_init[43]), .Q(
        msg[43]) );
  DFF \msg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(e_init[44]), .Q(
        msg[44]) );
  DFF \msg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(e_init[45]), .Q(
        msg[45]) );
  DFF \msg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(e_init[46]), .Q(
        msg[46]) );
  DFF \msg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(e_init[47]), .Q(
        msg[47]) );
  DFF \msg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(e_init[48]), .Q(
        msg[48]) );
  DFF \msg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(e_init[49]), .Q(
        msg[49]) );
  DFF \msg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(e_init[50]), .Q(
        msg[50]) );
  DFF \msg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(e_init[51]), .Q(
        msg[51]) );
  DFF \msg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(e_init[52]), .Q(
        msg[52]) );
  DFF \msg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(e_init[53]), .Q(
        msg[53]) );
  DFF \msg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(e_init[54]), .Q(
        msg[54]) );
  DFF \msg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(e_init[55]), .Q(
        msg[55]) );
  DFF \msg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(e_init[56]), .Q(
        msg[56]) );
  DFF \msg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(e_init[57]), .Q(
        msg[57]) );
  DFF \msg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(e_init[58]), .Q(
        msg[58]) );
  DFF \msg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(e_init[59]), .Q(
        msg[59]) );
  DFF \msg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(e_init[60]), .Q(
        msg[60]) );
  DFF \msg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(e_init[61]), .Q(
        msg[61]) );
  DFF \msg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(e_init[62]), .Q(
        msg[62]) );
  DFF \msg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(e_init[63]), .Q(
        msg[63]) );
  DFF \msg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(e_init[64]), .Q(
        msg[64]) );
  DFF \msg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(e_init[65]), .Q(
        msg[65]) );
  DFF \msg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(e_init[66]), .Q(
        msg[66]) );
  DFF \msg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(e_init[67]), .Q(
        msg[67]) );
  DFF \msg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(e_init[68]), .Q(
        msg[68]) );
  DFF \msg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(e_init[69]), .Q(
        msg[69]) );
  DFF \msg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(e_init[70]), .Q(
        msg[70]) );
  DFF \msg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(e_init[71]), .Q(
        msg[71]) );
  DFF \msg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(e_init[72]), .Q(
        msg[72]) );
  DFF \msg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(e_init[73]), .Q(
        msg[73]) );
  DFF \msg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(e_init[74]), .Q(
        msg[74]) );
  DFF \msg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(e_init[75]), .Q(
        msg[75]) );
  DFF \msg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(e_init[76]), .Q(
        msg[76]) );
  DFF \msg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(e_init[77]), .Q(
        msg[77]) );
  DFF \msg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(e_init[78]), .Q(
        msg[78]) );
  DFF \msg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(e_init[79]), .Q(
        msg[79]) );
  DFF \msg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(e_init[80]), .Q(
        msg[80]) );
  DFF \msg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(e_init[81]), .Q(
        msg[81]) );
  DFF \msg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(e_init[82]), .Q(
        msg[82]) );
  DFF \msg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(e_init[83]), .Q(
        msg[83]) );
  DFF \msg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(e_init[84]), .Q(
        msg[84]) );
  DFF \msg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(e_init[85]), .Q(
        msg[85]) );
  DFF \msg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(e_init[86]), .Q(
        msg[86]) );
  DFF \msg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(e_init[87]), .Q(
        msg[87]) );
  DFF \msg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(e_init[88]), .Q(
        msg[88]) );
  DFF \msg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(e_init[89]), .Q(
        msg[89]) );
  DFF \msg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(e_init[90]), .Q(
        msg[90]) );
  DFF \msg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(e_init[91]), .Q(
        msg[91]) );
  DFF \msg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(e_init[92]), .Q(
        msg[92]) );
  DFF \msg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(e_init[93]), .Q(
        msg[93]) );
  DFF \msg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(e_init[94]), .Q(
        msg[94]) );
  DFF \msg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(e_init[95]), .Q(
        msg[95]) );
  DFF \msg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(e_init[96]), .Q(
        msg[96]) );
  DFF \msg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(e_init[97]), .Q(
        msg[97]) );
  DFF \msg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(e_init[98]), .Q(
        msg[98]) );
  DFF \msg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(e_init[99]), .Q(
        msg[99]) );
  DFF \msg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(e_init[100]), .Q(
        msg[100]) );
  DFF \msg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(e_init[101]), .Q(
        msg[101]) );
  DFF \msg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(e_init[102]), .Q(
        msg[102]) );
  DFF \msg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(e_init[103]), .Q(
        msg[103]) );
  DFF \msg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(e_init[104]), .Q(
        msg[104]) );
  DFF \msg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(e_init[105]), .Q(
        msg[105]) );
  DFF \msg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(e_init[106]), .Q(
        msg[106]) );
  DFF \msg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(e_init[107]), .Q(
        msg[107]) );
  DFF \msg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(e_init[108]), .Q(
        msg[108]) );
  DFF \msg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(e_init[109]), .Q(
        msg[109]) );
  DFF \msg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(e_init[110]), .Q(
        msg[110]) );
  DFF \msg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(e_init[111]), .Q(
        msg[111]) );
  DFF \msg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(e_init[112]), .Q(
        msg[112]) );
  DFF \msg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(e_init[113]), .Q(
        msg[113]) );
  DFF \msg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(e_init[114]), .Q(
        msg[114]) );
  DFF \msg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(e_init[115]), .Q(
        msg[115]) );
  DFF \msg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(e_init[116]), .Q(
        msg[116]) );
  DFF \msg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(e_init[117]), .Q(
        msg[117]) );
  DFF \msg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(e_init[118]), .Q(
        msg[118]) );
  DFF \msg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(e_init[119]), .Q(
        msg[119]) );
  DFF \msg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(e_init[120]), .Q(
        msg[120]) );
  DFF \msg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(e_init[121]), .Q(
        msg[121]) );
  DFF \msg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(e_init[122]), .Q(
        msg[122]) );
  DFF \msg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(e_init[123]), .Q(
        msg[123]) );
  DFF \msg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .I(e_init[124]), .Q(
        msg[124]) );
  DFF \msg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .I(e_init[125]), .Q(
        msg[125]) );
  DFF \msg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .I(e_init[126]), .Q(
        msg[126]) );
  DFF \msg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(e_init[127]), .Q(
        msg[127]) );
  XOR \e/U223  ( .A(\e/n87 ), .B(\e/n54 ), .Z(\e/n95 ) );
  XOR \e/U222  ( .A(\e/Q[0] ), .B(key[0]), .Z(\e/n54 ) );
  XOR \e/U221  ( .A(\e/n88 ), .B(\e/n55 ), .Z(\e/n96 ) );
  XOR \e/U220  ( .A(\e/Q[1] ), .B(key[1]), .Z(\e/n55 ) );
  XOR \e/U219  ( .A(\e/n89 ), .B(\e/n56 ), .Z(\e/n97 ) );
  XOR \e/U218  ( .A(\e/Q[2] ), .B(key[2]), .Z(\e/n56 ) );
  XOR \e/U217  ( .A(\e/n90 ), .B(\e/n57 ), .Z(\e/n98 ) );
  XOR \e/U216  ( .A(\e/Q[3] ), .B(key[3]), .Z(\e/n57 ) );
  XOR \e/U215  ( .A(\e/n91 ), .B(\e/n58 ), .Z(\e/n99 ) );
  XOR \e/U214  ( .A(\e/Q[4] ), .B(key[4]), .Z(\e/n58 ) );
  XOR \e/U213  ( .A(\e/n92 ), .B(\e/n59 ), .Z(\e/n100 ) );
  XOR \e/U212  ( .A(\e/Q[5] ), .B(key[5]), .Z(\e/n59 ) );
  XOR \e/U211  ( .A(\e/n93 ), .B(\e/n60 ), .Z(\e/n101 ) );
  XOR \e/U210  ( .A(\e/Q[6] ), .B(key[6]), .Z(\e/n60 ) );
  XOR \e/U209  ( .A(\e/n94 ), .B(\e/n61 ), .Z(\e/n102 ) );
  XOR \e/U208  ( .A(\e/Q[7] ), .B(key[7]), .Z(\e/n61 ) );
  XOR \e/U207  ( .A(key[32]), .B(\e/n95 ), .Z(\e/n103 ) );
  XOR \e/U206  ( .A(key[33]), .B(\e/n96 ), .Z(\e/n104 ) );
  XOR \e/U205  ( .A(key[34]), .B(\e/n97 ), .Z(\e/n105 ) );
  XOR \e/U204  ( .A(key[35]), .B(\e/n98 ), .Z(\e/n106 ) );
  XOR \e/U203  ( .A(key[36]), .B(\e/n99 ), .Z(\e/n107 ) );
  XOR \e/U202  ( .A(key[37]), .B(\e/n100 ), .Z(\e/n108 ) );
  XOR \e/U201  ( .A(key[38]), .B(\e/n101 ), .Z(\e/n109 ) );
  XOR \e/U200  ( .A(key[39]), .B(\e/n102 ), .Z(\e/n110 ) );
  XOR \e/U199  ( .A(key[64]), .B(\e/n103 ), .Z(\e/n111 ) );
  XOR \e/U198  ( .A(key[65]), .B(\e/n104 ), .Z(\e/n112 ) );
  XOR \e/U197  ( .A(key[66]), .B(\e/n105 ), .Z(\e/n113 ) );
  XOR \e/U196  ( .A(key[67]), .B(\e/n106 ), .Z(\e/n114 ) );
  XOR \e/U195  ( .A(key[68]), .B(\e/n107 ), .Z(\e/n115 ) );
  XOR \e/U194  ( .A(key[69]), .B(\e/n108 ), .Z(\e/n116 ) );
  XOR \e/U193  ( .A(key[70]), .B(\e/n109 ), .Z(\e/n117 ) );
  XOR \e/U192  ( .A(key[71]), .B(\e/n110 ), .Z(\e/n118 ) );
  XOR \e/U183  ( .A(key[8]), .B(\e/n62 ), .Z(nextKey[40]) );
  XOR \e/U182  ( .A(\e/t[8] ), .B(key[40]), .Z(\e/n62 ) );
  XOR \e/U181  ( .A(key[9]), .B(\e/n63 ), .Z(nextKey[41]) );
  XOR \e/U180  ( .A(\e/t[9] ), .B(key[41]), .Z(\e/n63 ) );
  XOR \e/U179  ( .A(key[10]), .B(\e/n64 ), .Z(nextKey[42]) );
  XOR \e/U178  ( .A(\e/t[10] ), .B(key[42]), .Z(\e/n64 ) );
  XOR \e/U177  ( .A(key[11]), .B(\e/n65 ), .Z(nextKey[43]) );
  XOR \e/U176  ( .A(\e/t[11] ), .B(key[43]), .Z(\e/n65 ) );
  XOR \e/U175  ( .A(key[12]), .B(\e/n66 ), .Z(nextKey[44]) );
  XOR \e/U174  ( .A(\e/t[12] ), .B(key[44]), .Z(\e/n66 ) );
  XOR \e/U173  ( .A(key[13]), .B(\e/n67 ), .Z(nextKey[45]) );
  XOR \e/U172  ( .A(\e/t[13] ), .B(key[45]), .Z(\e/n67 ) );
  XOR \e/U171  ( .A(key[14]), .B(\e/n68 ), .Z(nextKey[46]) );
  XOR \e/U170  ( .A(\e/t[14] ), .B(key[46]), .Z(\e/n68 ) );
  XOR \e/U169  ( .A(key[15]), .B(\e/n69 ), .Z(nextKey[47]) );
  XOR \e/U168  ( .A(\e/t[15] ), .B(key[47]), .Z(\e/n69 ) );
  XOR \e/U167  ( .A(key[16]), .B(\e/n70 ), .Z(nextKey[48]) );
  XOR \e/U166  ( .A(\e/t[16] ), .B(key[48]), .Z(\e/n70 ) );
  XOR \e/U165  ( .A(key[17]), .B(\e/n71 ), .Z(nextKey[49]) );
  XOR \e/U164  ( .A(\e/t[17] ), .B(key[49]), .Z(\e/n71 ) );
  XOR \e/U163  ( .A(key[18]), .B(\e/n72 ), .Z(nextKey[50]) );
  XOR \e/U162  ( .A(\e/t[18] ), .B(key[50]), .Z(\e/n72 ) );
  XOR \e/U161  ( .A(key[19]), .B(\e/n73 ), .Z(nextKey[51]) );
  XOR \e/U160  ( .A(\e/t[19] ), .B(key[51]), .Z(\e/n73 ) );
  XOR \e/U159  ( .A(key[20]), .B(\e/n74 ), .Z(nextKey[52]) );
  XOR \e/U158  ( .A(\e/t[20] ), .B(key[52]), .Z(\e/n74 ) );
  XOR \e/U157  ( .A(key[21]), .B(\e/n75 ), .Z(nextKey[53]) );
  XOR \e/U156  ( .A(\e/t[21] ), .B(key[53]), .Z(\e/n75 ) );
  XOR \e/U155  ( .A(key[22]), .B(\e/n76 ), .Z(nextKey[54]) );
  XOR \e/U154  ( .A(\e/t[22] ), .B(key[54]), .Z(\e/n76 ) );
  XOR \e/U153  ( .A(key[23]), .B(\e/n77 ), .Z(nextKey[55]) );
  XOR \e/U152  ( .A(\e/t[23] ), .B(key[55]), .Z(\e/n77 ) );
  XOR \e/U151  ( .A(key[24]), .B(\e/n78 ), .Z(nextKey[56]) );
  XOR \e/U150  ( .A(\e/t[24] ), .B(key[56]), .Z(\e/n78 ) );
  XOR \e/U149  ( .A(key[25]), .B(\e/n79 ), .Z(nextKey[57]) );
  XOR \e/U148  ( .A(\e/t[25] ), .B(key[57]), .Z(\e/n79 ) );
  XOR \e/U147  ( .A(key[26]), .B(\e/n80 ), .Z(nextKey[58]) );
  XOR \e/U146  ( .A(\e/t[26] ), .B(key[58]), .Z(\e/n80 ) );
  XOR \e/U145  ( .A(key[27]), .B(\e/n81 ), .Z(nextKey[59]) );
  XOR \e/U144  ( .A(\e/t[27] ), .B(key[59]), .Z(\e/n81 ) );
  XOR \e/U143  ( .A(key[28]), .B(\e/n82 ), .Z(nextKey[60]) );
  XOR \e/U142  ( .A(\e/t[28] ), .B(key[60]), .Z(\e/n82 ) );
  XOR \e/U141  ( .A(key[29]), .B(\e/n83 ), .Z(nextKey[61]) );
  XOR \e/U140  ( .A(\e/t[29] ), .B(key[61]), .Z(\e/n83 ) );
  XOR \e/U139  ( .A(key[30]), .B(\e/n84 ), .Z(nextKey[62]) );
  XOR \e/U138  ( .A(\e/t[30] ), .B(key[62]), .Z(\e/n84 ) );
  XOR \e/U137  ( .A(key[31]), .B(\e/n85 ), .Z(nextKey[63]) );
  XOR \e/U136  ( .A(\e/t[31] ), .B(key[63]), .Z(\e/n85 ) );
  XOR \e/U135  ( .A(key[72]), .B(nextKey[40]), .Z(nextKey[72]) );
  XOR \e/U134  ( .A(key[73]), .B(nextKey[41]), .Z(nextKey[73]) );
  XOR \e/U133  ( .A(key[74]), .B(nextKey[42]), .Z(nextKey[74]) );
  XOR \e/U132  ( .A(key[75]), .B(nextKey[43]), .Z(nextKey[75]) );
  XOR \e/U131  ( .A(key[76]), .B(nextKey[44]), .Z(nextKey[76]) );
  XOR \e/U130  ( .A(key[77]), .B(nextKey[45]), .Z(nextKey[77]) );
  XOR \e/U129  ( .A(key[78]), .B(nextKey[46]), .Z(nextKey[78]) );
  XOR \e/U128  ( .A(key[79]), .B(nextKey[47]), .Z(nextKey[79]) );
  XOR \e/U127  ( .A(key[80]), .B(nextKey[48]), .Z(nextKey[80]) );
  XOR \e/U126  ( .A(key[81]), .B(nextKey[49]), .Z(nextKey[81]) );
  XOR \e/U125  ( .A(key[82]), .B(nextKey[50]), .Z(nextKey[82]) );
  XOR \e/U124  ( .A(key[83]), .B(nextKey[51]), .Z(nextKey[83]) );
  XOR \e/U123  ( .A(key[84]), .B(nextKey[52]), .Z(nextKey[84]) );
  XOR \e/U122  ( .A(key[85]), .B(nextKey[53]), .Z(nextKey[85]) );
  XOR \e/U121  ( .A(key[86]), .B(nextKey[54]), .Z(nextKey[86]) );
  XOR \e/U120  ( .A(key[87]), .B(nextKey[55]), .Z(nextKey[87]) );
  XOR \e/U119  ( .A(key[88]), .B(nextKey[56]), .Z(nextKey[88]) );
  XOR \e/U118  ( .A(key[89]), .B(nextKey[57]), .Z(nextKey[89]) );
  XOR \e/U117  ( .A(key[90]), .B(nextKey[58]), .Z(nextKey[90]) );
  XOR \e/U116  ( .A(key[91]), .B(nextKey[59]), .Z(nextKey[91]) );
  XOR \e/U115  ( .A(key[92]), .B(nextKey[60]), .Z(nextKey[92]) );
  XOR \e/U114  ( .A(key[93]), .B(nextKey[61]), .Z(nextKey[93]) );
  XOR \e/U113  ( .A(key[94]), .B(nextKey[62]), .Z(nextKey[94]) );
  XOR \e/U112  ( .A(key[95]), .B(nextKey[63]), .Z(nextKey[95]) );
  XOR \e/U111  ( .A(key[104]), .B(nextKey[72]), .Z(nextKey[104]) );
  XOR \e/U110  ( .A(key[105]), .B(nextKey[73]), .Z(nextKey[105]) );
  XOR \e/U109  ( .A(key[106]), .B(nextKey[74]), .Z(nextKey[106]) );
  XOR \e/U108  ( .A(key[107]), .B(nextKey[75]), .Z(nextKey[107]) );
  XOR \e/U107  ( .A(key[108]), .B(nextKey[76]), .Z(nextKey[108]) );
  XOR \e/U106  ( .A(key[109]), .B(nextKey[77]), .Z(nextKey[109]) );
  XOR \e/U105  ( .A(key[110]), .B(nextKey[78]), .Z(nextKey[110]) );
  XOR \e/U104  ( .A(key[111]), .B(nextKey[79]), .Z(nextKey[111]) );
  XOR \e/U103  ( .A(key[112]), .B(nextKey[80]), .Z(nextKey[112]) );
  XOR \e/U102  ( .A(key[113]), .B(nextKey[81]), .Z(nextKey[113]) );
  XOR \e/U101  ( .A(key[114]), .B(nextKey[82]), .Z(nextKey[114]) );
  XOR \e/U100  ( .A(key[115]), .B(nextKey[83]), .Z(nextKey[115]) );
  XOR \e/U99  ( .A(key[116]), .B(nextKey[84]), .Z(nextKey[116]) );
  XOR \e/U98  ( .A(key[117]), .B(nextKey[85]), .Z(nextKey[117]) );
  XOR \e/U97  ( .A(key[118]), .B(nextKey[86]), .Z(nextKey[118]) );
  XOR \e/U96  ( .A(key[119]), .B(nextKey[87]), .Z(nextKey[119]) );
  XOR \e/U95  ( .A(key[120]), .B(nextKey[88]), .Z(nextKey[120]) );
  XOR \e/U94  ( .A(key[121]), .B(nextKey[89]), .Z(nextKey[121]) );
  XOR \e/U93  ( .A(key[122]), .B(nextKey[90]), .Z(nextKey[122]) );
  XOR \e/U92  ( .A(key[123]), .B(nextKey[91]), .Z(nextKey[123]) );
  XOR \e/U91  ( .A(key[124]), .B(nextKey[92]), .Z(nextKey[124]) );
  XOR \e/U90  ( .A(key[125]), .B(nextKey[93]), .Z(nextKey[125]) );
  XOR \e/U89  ( .A(key[126]), .B(nextKey[94]), .Z(nextKey[126]) );
  XOR \e/U88  ( .A(key[127]), .B(nextKey[95]), .Z(nextKey[127]) );
  MUX \b/U7005  ( .IN0(msg[124]), .IN1(\b/n6519 ), .SEL(msg[121]), .F(
        \b/n6877 ) );
  MUX \b/U7004  ( .IN0(msg[124]), .IN1(\b/n6528 ), .SEL(msg[121]), .F(
        \b/n6876 ) );
  MUX \b/U7003  ( .IN0(\b/n6520 ), .IN1(\b/n6523 ), .SEL(msg[121]), .F(
        \b/n6875 ) );
  MUX \b/U7002  ( .IN0(\b/n6525 ), .IN1(\b/n60 ), .SEL(msg[121]), .F(\b/n6874 ) );
  MUX \b/U7000  ( .IN0(\b/n6528 ), .IN1(\b/n6519 ), .SEL(msg[122]), .F(
        \b/n6701 ) );
  MUX \b/U6999  ( .IN0(\b/n6521 ), .IN1(\b/n71 ), .SEL(msg[122]), .F(\b/n6702 ) );
  MUX \b/U6998  ( .IN0(\b/n14 ), .IN1(\b/n24 ), .SEL(msg[121]), .F(\b/n6665 )
         );
  MUX \b/U6997  ( .IN0(\b/n6549 ), .IN1(\b/n6860 ), .SEL(msg[127]), .F(
        \b/n6872 ) );
  MUX \b/U6996  ( .IN0(\b/n6523 ), .IN1(\b/n6519 ), .SEL(msg[121]), .F(
        \b/n6863 ) );
  MUX \b/U6995  ( .IN0(\b/n66 ), .IN1(\b/n6525 ), .SEL(msg[121]), .F(\b/n6871 ) );
  MUX \b/U6994  ( .IN0(msg[123]), .IN1(\b/n60 ), .SEL(msg[121]), .F(\b/n6870 )
         );
  MUX \b/U6993  ( .IN0(\b/n6528 ), .IN1(\b/n66 ), .SEL(msg[121]), .F(\b/n6869 ) );
  MUX \b/U6992  ( .IN0(msg[124]), .IN1(\b/n6525 ), .SEL(msg[121]), .F(
        \b/n6868 ) );
  MUX \b/U6991  ( .IN0(\b/n51 ), .IN1(\b/n30 ), .SEL(msg[125]), .F(\b/n6575 )
         );
  MUX \b/U6990  ( .IN0(\b/n6520 ), .IN1(\b/n24 ), .SEL(msg[121]), .F(\b/n6867 ) );
  NANDN \b/U6987  ( .B(\b/n6526 ), .A(msg[127]), .Z(\b/n6840 ) );
  NAND \b/U6986  ( .A(msg[127]), .B(\b/n27 ), .Z(\b/n6808 ) );
  NAND \b/U6985  ( .A(msg[127]), .B(\b/n39 ), .Z(\b/n6749 ) );
  NAND \b/U6984  ( .A(msg[127]), .B(\b/n6857 ), .Z(\b/n6782 ) );
  NAND \b/U6983  ( .A(msg[127]), .B(\b/n6777 ), .Z(\b/n6740 ) );
  NAND \b/U6981  ( .A(\b/n71 ), .B(\b/n60 ), .Z(\b/n6861 ) );
  NAND \b/U6980  ( .A(msg[127]), .B(\b/n6859 ), .Z(\b/n6854 ) );
  NAND \b/U6979  ( .A(n728), .B(msg[127]), .Z(\b/n6834 ) );
  NAND \b/U6977  ( .A(msg[122]), .B(\b/n6528 ), .Z(\b/n6694 ) );
  NAND \b/U6976  ( .A(\b/n60 ), .B(msg[121]), .Z(\b/n6649 ) );
  NAND \b/U6975  ( .A(msg[127]), .B(\b/n6863 ), .Z(\b/n6648 ) );
  NAND \b/U6973  ( .A(\b/n6861 ), .B(msg[127]), .Z(\b/n6664 ) );
  NAND \b/U6972  ( .A(\b/n6682 ), .B(\b/n6528 ), .Z(\b/n6860 ) );
  NANDN \b/U6971  ( .B(\b/n14 ), .A(\b/n71 ), .Z(\b/n6859 ) );
  NAND \b/U6969  ( .A(msg[121]), .B(\b/n6528 ), .Z(\b/n6580 ) );
  NAND \b/U6968  ( .A(\b/n14 ), .B(\b/n71 ), .Z(\b/n6857 ) );
  NAND \b/U6965  ( .A(msg[121]), .B(\b/n6523 ), .Z(\b/n6682 ) );
  ANDN \b/U6963  ( .A(msg[122]), .B(msg[121]), .Z(\b/n6710 ) );
  AND \b/U6962  ( .A(\b/n6520 ), .B(\b/n6854 ), .Z(\b/n6625 ) );
  MUX \b/U6961  ( .IN0(\b/n6853 ), .IN1(\b/n6837 ), .SEL(msg[126]), .F(
        shift_row_out[31]) );
  MUX \b/U6960  ( .IN0(\b/n6852 ), .IN1(\b/n6845 ), .SEL(msg[120]), .F(
        \b/n6853 ) );
  MUX \b/U6959  ( .IN0(\b/n6851 ), .IN1(\b/n6848 ), .SEL(msg[125]), .F(
        \b/n6852 ) );
  MUX \b/U6958  ( .IN0(\b/n6850 ), .IN1(\b/n6849 ), .SEL(msg[122]), .F(
        \b/n6851 ) );
  MUX \b/U6957  ( .IN0(msg[124]), .IN1(\b/n31 ), .SEL(msg[127]), .F(\b/n6850 )
         );
  MUX \b/U6956  ( .IN0(\b/n6521 ), .IN1(\b/n35 ), .SEL(msg[127]), .F(\b/n6849 ) );
  MUX \b/U6955  ( .IN0(\b/n6847 ), .IN1(\b/n6846 ), .SEL(msg[122]), .F(
        \b/n6848 ) );
  MUX \b/U6954  ( .IN0(\b/n6579 ), .IN1(\b/n27 ), .SEL(msg[127]), .F(\b/n6847 ) );
  MUX \b/U6953  ( .IN0(\b/n6531 ), .IN1(\b/n6542 ), .SEL(msg[127]), .F(
        \b/n6846 ) );
  MUX \b/U6952  ( .IN0(\b/n6844 ), .IN1(\b/n6841 ), .SEL(msg[125]), .F(
        \b/n6845 ) );
  MUX \b/U6951  ( .IN0(\b/n6843 ), .IN1(\b/n6842 ), .SEL(msg[122]), .F(
        \b/n6844 ) );
  MUX \b/U6950  ( .IN0(\b/n6555 ), .IN1(\b/n6530 ), .SEL(msg[127]), .F(
        \b/n6843 ) );
  MUX \b/U6949  ( .IN0(\b/n39 ), .IN1(\b/n6551 ), .SEL(msg[127]), .F(\b/n6842 ) );
  MUX \b/U6948  ( .IN0(\b/n6839 ), .IN1(\b/n6838 ), .SEL(msg[122]), .F(
        \b/n6841 ) );
  AND \b/U6947  ( .A(\b/n29 ), .B(\b/n6840 ), .Z(\b/n6839 ) );
  MUX \b/U6946  ( .IN0(\b/n6535 ), .IN1(n727), .SEL(msg[127]), .F(\b/n6838 )
         );
  MUX \b/U6945  ( .IN0(\b/n6836 ), .IN1(\b/n6828 ), .SEL(msg[120]), .F(
        \b/n6837 ) );
  MUX \b/U6944  ( .IN0(\b/n6835 ), .IN1(\b/n6831 ), .SEL(msg[125]), .F(
        \b/n6836 ) );
  MUX \b/U6943  ( .IN0(\b/n6832 ), .IN1(\b/n6833 ), .SEL(msg[122]), .F(
        \b/n6835 ) );
  NAND \b/U6942  ( .A(\b/n6649 ), .B(\b/n6834 ), .Z(\b/n6833 ) );
  MUX \b/U6941  ( .IN0(\b/n69 ), .IN1(\b/n61 ), .SEL(msg[127]), .F(\b/n6832 )
         );
  MUX \b/U6940  ( .IN0(\b/n6830 ), .IN1(\b/n6829 ), .SEL(msg[122]), .F(
        \b/n6831 ) );
  MUX \b/U6939  ( .IN0(\b/n6525 ), .IN1(\b/n6519 ), .SEL(msg[127]), .F(
        \b/n6830 ) );
  MUX \b/U6938  ( .IN0(\b/n62 ), .IN1(\b/n6556 ), .SEL(msg[127]), .F(\b/n6829 ) );
  MUX \b/U6937  ( .IN0(\b/n6827 ), .IN1(\b/n6824 ), .SEL(msg[125]), .F(
        \b/n6828 ) );
  MUX \b/U6936  ( .IN0(\b/n6826 ), .IN1(\b/n6825 ), .SEL(msg[122]), .F(
        \b/n6827 ) );
  MUX \b/U6935  ( .IN0(\b/n6560 ), .IN1(\b/n6546 ), .SEL(msg[127]), .F(
        \b/n6826 ) );
  MUX \b/U6934  ( .IN0(\b/n15 ), .IN1(\b/n6528 ), .SEL(msg[127]), .F(\b/n6825 ) );
  MUX \b/U6933  ( .IN0(\b/n6823 ), .IN1(\b/n6822 ), .SEL(msg[122]), .F(
        \b/n6824 ) );
  MUX \b/U6932  ( .IN0(\b/n6561 ), .IN1(\b/n6569 ), .SEL(msg[127]), .F(
        \b/n6823 ) );
  MUX \b/U6931  ( .IN0(\b/n6554 ), .IN1(\b/n6821 ), .SEL(msg[127]), .F(
        \b/n6822 ) );
  MUX \b/U6930  ( .IN0(\b/n66 ), .IN1(\b/n24 ), .SEL(msg[121]), .F(\b/n6821 )
         );
  MUX \b/U6929  ( .IN0(\b/n6820 ), .IN1(\b/n6802 ), .SEL(msg[126]), .F(
        shift_row_out[30]) );
  MUX \b/U6928  ( .IN0(\b/n6819 ), .IN1(\b/n6810 ), .SEL(msg[120]), .F(
        \b/n6820 ) );
  MUX \b/U6927  ( .IN0(\b/n6818 ), .IN1(\b/n6813 ), .SEL(msg[125]), .F(
        \b/n6819 ) );
  MUX \b/U6926  ( .IN0(\b/n6817 ), .IN1(\b/n6815 ), .SEL(msg[122]), .F(
        \b/n6818 ) );
  MUX \b/U6925  ( .IN0(\b/n6816 ), .IN1(\b/n6532 ), .SEL(msg[127]), .F(
        \b/n6817 ) );
  MUX \b/U6924  ( .IN0(\b/n66 ), .IN1(\b/n6519 ), .SEL(msg[121]), .F(\b/n6816 ) );
  MUX \b/U6923  ( .IN0(\b/n6814 ), .IN1(\b/n54 ), .SEL(msg[127]), .F(\b/n6815 ) );
  MUX \b/U6922  ( .IN0(\b/n6519 ), .IN1(\b/n6520 ), .SEL(msg[121]), .F(
        \b/n6814 ) );
  MUX \b/U6921  ( .IN0(\b/n6812 ), .IN1(\b/n6811 ), .SEL(msg[122]), .F(
        \b/n6813 ) );
  MUX \b/U6920  ( .IN0(n726), .IN1(\b/n6600 ), .SEL(msg[127]), .F(\b/n6812 )
         );
  MUX \b/U6919  ( .IN0(\b/n6558 ), .IN1(\b/n6565 ), .SEL(msg[127]), .F(
        \b/n6811 ) );
  MUX \b/U6918  ( .IN0(\b/n6809 ), .IN1(\b/n6805 ), .SEL(msg[125]), .F(
        \b/n6810 ) );
  MUX \b/U6917  ( .IN0(\b/n6807 ), .IN1(\b/n6806 ), .SEL(msg[122]), .F(
        \b/n6809 ) );
  AND \b/U6916  ( .A(\b/n7 ), .B(\b/n6808 ), .Z(\b/n6807 ) );
  MUX \b/U6915  ( .IN0(\b/n6635 ), .IN1(msg[123]), .SEL(msg[127]), .F(
        \b/n6806 ) );
  MUX \b/U6914  ( .IN0(\b/n6804 ), .IN1(\b/n6803 ), .SEL(msg[122]), .F(
        \b/n6805 ) );
  MUX \b/U6913  ( .IN0(\b/n50 ), .IN1(\b/n6523 ), .SEL(msg[127]), .F(\b/n6804 ) );
  MUX \b/U6911  ( .IN0(\b/n6801 ), .IN1(\b/n6794 ), .SEL(msg[120]), .F(
        \b/n6802 ) );
  MUX \b/U6910  ( .IN0(\b/n6800 ), .IN1(\b/n6797 ), .SEL(msg[125]), .F(
        \b/n6801 ) );
  MUX \b/U6909  ( .IN0(\b/n6799 ), .IN1(\b/n6798 ), .SEL(msg[122]), .F(
        \b/n6800 ) );
  MUX \b/U6908  ( .IN0(\b/n46 ), .IN1(\b/n6527 ), .SEL(msg[127]), .F(\b/n6799 ) );
  MUX \b/U6907  ( .IN0(\b/n6531 ), .IN1(n727), .SEL(msg[127]), .F(\b/n6798 )
         );
  MUX \b/U6906  ( .IN0(\b/n6796 ), .IN1(\b/n6795 ), .SEL(msg[122]), .F(
        \b/n6797 ) );
  MUX \b/U6905  ( .IN0(\b/n6547 ), .IN1(\b/n11 ), .SEL(msg[127]), .F(\b/n6796 ) );
  MUX \b/U6904  ( .IN0(\b/n31 ), .IN1(\b/n61 ), .SEL(msg[127]), .F(\b/n6795 )
         );
  MUX \b/U6903  ( .IN0(\b/n6793 ), .IN1(\b/n6789 ), .SEL(msg[125]), .F(
        \b/n6794 ) );
  MUX \b/U6902  ( .IN0(\b/n6792 ), .IN1(\b/n6791 ), .SEL(msg[122]), .F(
        \b/n6793 ) );
  MUX \b/U6901  ( .IN0(\b/n6536 ), .IN1(\b/n61 ), .SEL(msg[127]), .F(\b/n6792 ) );
  MUX \b/U6900  ( .IN0(\b/n6790 ), .IN1(\b/n6557 ), .SEL(msg[127]), .F(
        \b/n6791 ) );
  NANDN \b/U6899  ( .B(msg[124]), .A(msg[121]), .Z(\b/n6790 ) );
  MUX \b/U6898  ( .IN0(\b/n6788 ), .IN1(\b/n6786 ), .SEL(msg[122]), .F(
        \b/n6789 ) );
  MUX \b/U6897  ( .IN0(\b/n24 ), .IN1(\b/n6787 ), .SEL(msg[127]), .F(\b/n6788 ) );
  MUX \b/U6896  ( .IN0(\b/n51 ), .IN1(\b/n41 ), .SEL(msg[121]), .F(\b/n6787 )
         );
  MUX \b/U6895  ( .IN0(\b/n13 ), .IN1(\b/n6532 ), .SEL(msg[127]), .F(\b/n6786 ) );
  NANDN \b/U6894  ( .B(\b/n14 ), .A(msg[121]), .Z(\b/n6532 ) );
  MUX \b/U6893  ( .IN0(\b/n6785 ), .IN1(\b/n6764 ), .SEL(msg[126]), .F(
        shift_row_out[29]) );
  MUX \b/U6892  ( .IN0(\b/n6784 ), .IN1(\b/n6774 ), .SEL(msg[120]), .F(
        \b/n6785 ) );
  MUX \b/U6891  ( .IN0(\b/n6783 ), .IN1(\b/n6779 ), .SEL(msg[125]), .F(
        \b/n6784 ) );
  MUX \b/U6890  ( .IN0(\b/n6780 ), .IN1(\b/n6781 ), .SEL(msg[122]), .F(
        \b/n6783 ) );
  AND \b/U6889  ( .A(\b/n6550 ), .B(\b/n6782 ), .Z(\b/n6781 ) );
  MUX \b/U6888  ( .IN0(\b/n6528 ), .IN1(\b/n62 ), .SEL(msg[127]), .F(\b/n6780 ) );
  MUX \b/U6887  ( .IN0(\b/n6778 ), .IN1(\b/n6776 ), .SEL(msg[122]), .F(
        \b/n6779 ) );
  MUX \b/U6886  ( .IN0(\b/n17 ), .IN1(\b/n6777 ), .SEL(msg[127]), .F(\b/n6778 ) );
  NAND \b/U6885  ( .A(\b/n41 ), .B(\b/n71 ), .Z(\b/n6777 ) );
  MUX \b/U6884  ( .IN0(\b/n6528 ), .IN1(\b/n6775 ), .SEL(msg[127]), .F(
        \b/n6776 ) );
  NAND \b/U6883  ( .A(\b/n6519 ), .B(\b/n6580 ), .Z(\b/n6775 ) );
  MUX \b/U6882  ( .IN0(\b/n6773 ), .IN1(\b/n6769 ), .SEL(msg[125]), .F(
        \b/n6774 ) );
  MUX \b/U6881  ( .IN0(\b/n6772 ), .IN1(\b/n6771 ), .SEL(msg[122]), .F(
        \b/n6773 ) );
  MUX \b/U6880  ( .IN0(\b/n6540 ), .IN1(\b/n64 ), .SEL(msg[127]), .F(\b/n6772 ) );
  MUX \b/U6879  ( .IN0(\b/n6565 ), .IN1(\b/n6770 ), .SEL(msg[127]), .F(
        \b/n6771 ) );
  MUX \b/U6878  ( .IN0(\b/n60 ), .IN1(\b/n41 ), .SEL(msg[121]), .F(\b/n6770 )
         );
  MUX \b/U6877  ( .IN0(\b/n6768 ), .IN1(\b/n6767 ), .SEL(msg[122]), .F(
        \b/n6769 ) );
  MUX \b/U6876  ( .IN0(\b/n58 ), .IN1(n725), .SEL(msg[127]), .F(\b/n6768 ) );
  MUX \b/U6875  ( .IN0(\b/n6766 ), .IN1(\b/n6765 ), .SEL(msg[127]), .F(
        \b/n6767 ) );
  AND \b/U6874  ( .A(\b/n6525 ), .B(\b/n6600 ), .Z(\b/n6766 ) );
  MUX \b/U6873  ( .IN0(\b/n30 ), .IN1(\b/n14 ), .SEL(msg[121]), .F(\b/n6765 )
         );
  MUX \b/U6872  ( .IN0(\b/n6763 ), .IN1(\b/n6754 ), .SEL(msg[120]), .F(
        \b/n6764 ) );
  MUX \b/U6871  ( .IN0(\b/n6762 ), .IN1(\b/n6758 ), .SEL(msg[125]), .F(
        \b/n6763 ) );
  MUX \b/U6870  ( .IN0(\b/n6761 ), .IN1(\b/n6759 ), .SEL(msg[122]), .F(
        \b/n6762 ) );
  MUX \b/U6869  ( .IN0(\b/n6531 ), .IN1(\b/n6760 ), .SEL(msg[127]), .F(
        \b/n6761 ) );
  NAND \b/U6868  ( .A(msg[121]), .B(\b/n30 ), .Z(\b/n6760 ) );
  MUX \b/U6867  ( .IN0(\b/n14 ), .IN1(\b/n67 ), .SEL(msg[127]), .F(\b/n6759 )
         );
  MUX \b/U6866  ( .IN0(\b/n6757 ), .IN1(\b/n6756 ), .SEL(msg[122]), .F(
        \b/n6758 ) );
  MUX \b/U6865  ( .IN0(\b/n6557 ), .IN1(\b/n32 ), .SEL(msg[127]), .F(\b/n6757 ) );
  MUX \b/U6864  ( .IN0(\b/n6755 ), .IN1(\b/n6520 ), .SEL(n724), .F(\b/n6756 )
         );
  AND \b/U6863  ( .A(msg[127]), .B(msg[123]), .Z(\b/n6755 ) );
  MUX \b/U6862  ( .IN0(\b/n6753 ), .IN1(\b/n6750 ), .SEL(msg[125]), .F(
        \b/n6754 ) );
  MUX \b/U6861  ( .IN0(\b/n6752 ), .IN1(\b/n6751 ), .SEL(msg[122]), .F(
        \b/n6753 ) );
  MUX \b/U6860  ( .IN0(\b/n6681 ), .IN1(\b/n6520 ), .SEL(msg[127]), .F(
        \b/n6752 ) );
  MUX \b/U6859  ( .IN0(n723), .IN1(\b/n65 ), .SEL(msg[127]), .F(\b/n6751 ) );
  MUX \b/U6858  ( .IN0(\b/n6748 ), .IN1(\b/n6747 ), .SEL(msg[122]), .F(
        \b/n6750 ) );
  AND \b/U6857  ( .A(\b/n6749 ), .B(\b/n6649 ), .Z(\b/n6748 ) );
  MUX \b/U6856  ( .IN0(\b/n16 ), .IN1(\b/n60 ), .SEL(msg[127]), .F(\b/n6747 )
         );
  MUX \b/U6855  ( .IN0(\b/n6746 ), .IN1(\b/n6729 ), .SEL(msg[126]), .F(
        shift_row_out[28]) );
  MUX \b/U6854  ( .IN0(\b/n6745 ), .IN1(\b/n6737 ), .SEL(msg[120]), .F(
        \b/n6746 ) );
  MUX \b/U6853  ( .IN0(\b/n6744 ), .IN1(\b/n6741 ), .SEL(msg[125]), .F(
        \b/n6745 ) );
  MUX \b/U6852  ( .IN0(\b/n6743 ), .IN1(\b/n6742 ), .SEL(msg[122]), .F(
        \b/n6744 ) );
  MUX \b/U6851  ( .IN0(\b/n42 ), .IN1(\b/n63 ), .SEL(msg[127]), .F(\b/n6743 )
         );
  MUX \b/U6850  ( .IN0(\b/n6600 ), .IN1(\b/n6565 ), .SEL(msg[127]), .F(
        \b/n6742 ) );
  NAND \b/U6849  ( .A(msg[121]), .B(\b/n6519 ), .Z(\b/n6600 ) );
  MUX \b/U6848  ( .IN0(\b/n6738 ), .IN1(\b/n6739 ), .SEL(msg[122]), .F(
        \b/n6741 ) );
  AND \b/U6847  ( .A(\b/n6550 ), .B(\b/n6740 ), .Z(\b/n6739 ) );
  MUX \b/U6846  ( .IN0(\b/n6548 ), .IN1(\b/n45 ), .SEL(msg[127]), .F(\b/n6738 ) );
  MUX \b/U6845  ( .IN0(\b/n6736 ), .IN1(\b/n6733 ), .SEL(msg[125]), .F(
        \b/n6737 ) );
  MUX \b/U6844  ( .IN0(\b/n6735 ), .IN1(\b/n6734 ), .SEL(msg[122]), .F(
        \b/n6736 ) );
  MUX \b/U6843  ( .IN0(\b/n7 ), .IN1(\b/n53 ), .SEL(msg[127]), .F(\b/n6735 )
         );
  MUX \b/U6842  ( .IN0(\b/n14 ), .IN1(\b/n6528 ), .SEL(msg[127]), .F(\b/n6734 ) );
  MUX \b/U6841  ( .IN0(\b/n6732 ), .IN1(\b/n6730 ), .SEL(msg[122]), .F(
        \b/n6733 ) );
  MUX \b/U6840  ( .IN0(\b/n6544 ), .IN1(\b/n6731 ), .SEL(msg[127]), .F(
        \b/n6732 ) );
  AND \b/U6839  ( .A(\b/n6528 ), .B(\b/n71 ), .Z(\b/n6731 ) );
  MUX \b/U6838  ( .IN0(\b/n29 ), .IN1(\b/n48 ), .SEL(msg[127]), .F(\b/n6730 )
         );
  MUX \b/U6837  ( .IN0(\b/n6728 ), .IN1(\b/n6722 ), .SEL(msg[120]), .F(
        \b/n6729 ) );
  MUX \b/U6836  ( .IN0(\b/n6727 ), .IN1(\b/n6725 ), .SEL(msg[125]), .F(
        \b/n6728 ) );
  MUX \b/U6835  ( .IN0(\b/n6726 ), .IN1(\b/n6522 ), .SEL(msg[122]), .F(
        \b/n6727 ) );
  MUX \b/U6834  ( .IN0(\b/n6542 ), .IN1(\b/n50 ), .SEL(msg[127]), .F(\b/n6726 ) );
  MUX \b/U6833  ( .IN0(\b/n6724 ), .IN1(\b/n6723 ), .SEL(msg[122]), .F(
        \b/n6725 ) );
  MUX \b/U6832  ( .IN0(n722), .IN1(\b/n42 ), .SEL(msg[127]), .F(\b/n6724 ) );
  MUX \b/U6831  ( .IN0(\b/n6552 ), .IN1(\b/n6555 ), .SEL(msg[127]), .F(
        \b/n6723 ) );
  MUX \b/U6830  ( .IN0(\b/n6721 ), .IN1(\b/n6718 ), .SEL(msg[125]), .F(
        \b/n6722 ) );
  MUX \b/U6829  ( .IN0(\b/n6720 ), .IN1(\b/n6719 ), .SEL(msg[122]), .F(
        \b/n6721 ) );
  MUX \b/U6828  ( .IN0(\b/n15 ), .IN1(\b/n6524 ), .SEL(msg[127]), .F(\b/n6720 ) );
  MUX \b/U6827  ( .IN0(\b/n60 ), .IN1(\b/n6546 ), .SEL(msg[127]), .F(\b/n6719 ) );
  MUX \b/U6826  ( .IN0(\b/n3 ), .IN1(\b/n6717 ), .SEL(msg[122]), .F(\b/n6718 )
         );
  MUX \b/U6825  ( .IN0(\b/n23 ), .IN1(\b/n6528 ), .SEL(msg[127]), .F(\b/n6717 ) );
  MUX \b/U6824  ( .IN0(\b/n6716 ), .IN1(\b/n6697 ), .SEL(msg[126]), .F(
        shift_row_out[27]) );
  MUX \b/U6823  ( .IN0(\b/n6715 ), .IN1(\b/n6707 ), .SEL(msg[120]), .F(
        \b/n6716 ) );
  MUX \b/U6822  ( .IN0(\b/n6714 ), .IN1(\b/n6711 ), .SEL(msg[125]), .F(
        \b/n6715 ) );
  MUX \b/U6821  ( .IN0(\b/n6713 ), .IN1(\b/n6712 ), .SEL(msg[127]), .F(
        \b/n6714 ) );
  MUX \b/U6820  ( .IN0(\b/n6536 ), .IN1(\b/n48 ), .SEL(msg[122]), .F(\b/n6713 ) );
  MUX \b/U6819  ( .IN0(n725), .IN1(\b/n6 ), .SEL(msg[122]), .F(\b/n6712 ) );
  MUX \b/U6818  ( .IN0(\b/n6709 ), .IN1(\b/n6708 ), .SEL(msg[127]), .F(
        \b/n6711 ) );
  AND \b/U6817  ( .A(\b/n6710 ), .B(msg[124]), .Z(\b/n6709 ) );
  MUX \b/U6816  ( .IN0(\b/n36 ), .IN1(\b/n6549 ), .SEL(msg[122]), .F(\b/n6708 ) );
  MUX \b/U6815  ( .IN0(\b/n6706 ), .IN1(\b/n6703 ), .SEL(msg[125]), .F(
        \b/n6707 ) );
  MUX \b/U6814  ( .IN0(\b/n6705 ), .IN1(\b/n6704 ), .SEL(msg[127]), .F(
        \b/n6706 ) );
  MUX \b/U6813  ( .IN0(\b/n6540 ), .IN1(n721), .SEL(msg[122]), .F(\b/n6705 )
         );
  MUX \b/U6812  ( .IN0(\b/n4 ), .IN1(\b/n23 ), .SEL(msg[122]), .F(\b/n6704 )
         );
  MUX \b/U6811  ( .IN0(\b/n6699 ), .IN1(\b/n6700 ), .SEL(msg[127]), .F(
        \b/n6703 ) );
  NAND \b/U6810  ( .A(\b/n6701 ), .B(\b/n6702 ), .Z(\b/n6700 ) );
  MUX \b/U6809  ( .IN0(\b/n49 ), .IN1(\b/n6698 ), .SEL(msg[122]), .F(\b/n6699 ) );
  MUX \b/U6808  ( .IN0(\b/n24 ), .IN1(\b/n66 ), .SEL(msg[121]), .F(\b/n6698 )
         );
  MUX \b/U6807  ( .IN0(\b/n6696 ), .IN1(\b/n6687 ), .SEL(msg[120]), .F(
        \b/n6697 ) );
  MUX \b/U6806  ( .IN0(\b/n6695 ), .IN1(\b/n6691 ), .SEL(msg[125]), .F(
        \b/n6696 ) );
  MUX \b/U6805  ( .IN0(\b/n6693 ), .IN1(\b/n6692 ), .SEL(msg[127]), .F(
        \b/n6695 ) );
  NAND \b/U6804  ( .A(\b/n14 ), .B(\b/n6694 ), .Z(\b/n6693 ) );
  MUX \b/U6803  ( .IN0(\b/n65 ), .IN1(\b/n27 ), .SEL(msg[122]), .F(\b/n6692 )
         );
  MUX \b/U6802  ( .IN0(\b/n6690 ), .IN1(\b/n6688 ), .SEL(msg[127]), .F(
        \b/n6691 ) );
  MUX \b/U6801  ( .IN0(\b/n6531 ), .IN1(\b/n6689 ), .SEL(msg[122]), .F(
        \b/n6690 ) );
  AND \b/U6800  ( .A(msg[121]), .B(\b/n14 ), .Z(\b/n6689 ) );
  MUX \b/U6799  ( .IN0(\b/n19 ), .IN1(\b/n6550 ), .SEL(msg[122]), .F(\b/n6688 ) );
  MUX \b/U6798  ( .IN0(\b/n6686 ), .IN1(\b/n6680 ), .SEL(msg[125]), .F(
        \b/n6687 ) );
  MUX \b/U6797  ( .IN0(\b/n6685 ), .IN1(\b/n6683 ), .SEL(msg[127]), .F(
        \b/n6686 ) );
  MUX \b/U6796  ( .IN0(\b/n6684 ), .IN1(\b/n6520 ), .SEL(\b/n6568 ), .F(
        \b/n6685 ) );
  MUX \b/U6795  ( .IN0(msg[123]), .IN1(msg[124]), .SEL(msg[122]), .F(\b/n6684 ) );
  MUX \b/U6794  ( .IN0(\b/n6550 ), .IN1(\b/n6681 ), .SEL(msg[122]), .F(
        \b/n6683 ) );
  NAND \b/U6793  ( .A(\b/n6520 ), .B(\b/n6682 ), .Z(\b/n6681 ) );
  MUX \b/U6792  ( .IN0(\b/n6677 ), .IN1(\b/n6678 ), .SEL(msg[127]), .F(
        \b/n6680 ) );
  AND \b/U6791  ( .A(\b/n47 ), .B(\b/n6679 ), .Z(\b/n6678 ) );
  MUX \b/U6790  ( .IN0(\b/n28 ), .IN1(\b/n6521 ), .SEL(msg[122]), .F(\b/n6677 ) );
  MUX \b/U6789  ( .IN0(\b/n6676 ), .IN1(\b/n6660 ), .SEL(msg[126]), .F(
        shift_row_out[26]) );
  MUX \b/U6788  ( .IN0(\b/n6675 ), .IN1(\b/n6667 ), .SEL(msg[120]), .F(
        \b/n6676 ) );
  MUX \b/U6787  ( .IN0(\b/n6674 ), .IN1(\b/n6670 ), .SEL(msg[125]), .F(
        \b/n6675 ) );
  MUX \b/U6786  ( .IN0(\b/n6673 ), .IN1(\b/n6671 ), .SEL(msg[122]), .F(
        \b/n6674 ) );
  MUX \b/U6785  ( .IN0(\b/n36 ), .IN1(\b/n6672 ), .SEL(msg[127]), .F(\b/n6673 ) );
  MUX \b/U6784  ( .IN0(\b/n6528 ), .IN1(\b/n14 ), .SEL(msg[121]), .F(\b/n6672 ) );
  MUX \b/U6783  ( .IN0(\b/n6567 ), .IN1(\b/n54 ), .SEL(msg[127]), .F(\b/n6671 ) );
  MUX \b/U6782  ( .IN0(\b/n6669 ), .IN1(\b/n6668 ), .SEL(msg[122]), .F(
        \b/n6670 ) );
  MUX \b/U6781  ( .IN0(\b/n6521 ), .IN1(\b/n21 ), .SEL(msg[127]), .F(\b/n6669 ) );
  MUX \b/U6780  ( .IN0(\b/n57 ), .IN1(\b/n6554 ), .SEL(msg[127]), .F(\b/n6668 ) );
  MUX \b/U6779  ( .IN0(\b/n6666 ), .IN1(\b/n6662 ), .SEL(msg[125]), .F(
        \b/n6667 ) );
  MUX \b/U6778  ( .IN0(\b/n6663 ), .IN1(\b/n3 ), .SEL(msg[122]), .F(\b/n6666 )
         );
  NAND \b/U6777  ( .A(\b/n6664 ), .B(\b/n6665 ), .Z(\b/n6663 ) );
  MUX \b/U6776  ( .IN0(n723), .IN1(\b/n6661 ), .SEL(\b/n6566 ), .F(\b/n6662 )
         );
  MUX \b/U6775  ( .IN0(\b/n35 ), .IN1(\b/n6533 ), .SEL(msg[122]), .F(\b/n6661 ) );
  MUX \b/U6774  ( .IN0(\b/n6659 ), .IN1(\b/n6651 ), .SEL(msg[120]), .F(
        \b/n6660 ) );
  MUX \b/U6773  ( .IN0(\b/n6658 ), .IN1(\b/n6655 ), .SEL(msg[125]), .F(
        \b/n6659 ) );
  MUX \b/U6772  ( .IN0(\b/n6657 ), .IN1(\b/n6656 ), .SEL(msg[122]), .F(
        \b/n6658 ) );
  MUX \b/U6771  ( .IN0(\b/n63 ), .IN1(msg[121]), .SEL(msg[127]), .F(\b/n6657 )
         );
  MUX \b/U6770  ( .IN0(n726), .IN1(\b/n6534 ), .SEL(msg[127]), .F(\b/n6656 )
         );
  MUX \b/U6769  ( .IN0(\b/n6654 ), .IN1(\b/n6653 ), .SEL(msg[122]), .F(
        \b/n6655 ) );
  MUX \b/U6768  ( .IN0(\b/n68 ), .IN1(\b/n62 ), .SEL(msg[127]), .F(\b/n6654 )
         );
  MUX \b/U6767  ( .IN0(n726), .IN1(\b/n6652 ), .SEL(msg[127]), .F(\b/n6653 )
         );
  MUX \b/U6766  ( .IN0(\b/n14 ), .IN1(\b/n51 ), .SEL(msg[121]), .F(\b/n6652 )
         );
  MUX \b/U6765  ( .IN0(\b/n6650 ), .IN1(\b/n6644 ), .SEL(msg[125]), .F(
        \b/n6651 ) );
  MUX \b/U6764  ( .IN0(\b/n6647 ), .IN1(\b/n6646 ), .SEL(msg[122]), .F(
        \b/n6650 ) );
  NAND \b/U6763  ( .A(\b/n6648 ), .B(\b/n6649 ), .Z(\b/n6647 ) );
  MUX \b/U6762  ( .IN0(\b/n6520 ), .IN1(\b/n6645 ), .SEL(n724), .F(\b/n6646 )
         );
  MUX \b/U6761  ( .IN0(msg[123]), .IN1(\b/n24 ), .SEL(msg[127]), .F(\b/n6645 )
         );
  MUX \b/U6760  ( .IN0(\b/n6643 ), .IN1(\b/n6642 ), .SEL(msg[122]), .F(
        \b/n6644 ) );
  MUX \b/U6759  ( .IN0(\b/n6565 ), .IN1(\b/n22 ), .SEL(msg[127]), .F(\b/n6643 ) );
  MUX \b/U6758  ( .IN0(\b/n6561 ), .IN1(\b/n6641 ), .SEL(msg[127]), .F(
        \b/n6642 ) );
  MUX \b/U6757  ( .IN0(\b/n6523 ), .IN1(\b/n6528 ), .SEL(msg[121]), .F(
        \b/n6641 ) );
  MUX \b/U6756  ( .IN0(\b/n6640 ), .IN1(\b/n6622 ), .SEL(msg[126]), .F(
        shift_row_out[25]) );
  MUX \b/U6755  ( .IN0(\b/n6639 ), .IN1(\b/n6630 ), .SEL(msg[120]), .F(
        \b/n6640 ) );
  MUX \b/U6754  ( .IN0(\b/n6638 ), .IN1(\b/n6634 ), .SEL(msg[125]), .F(
        \b/n6639 ) );
  MUX \b/U6753  ( .IN0(\b/n6637 ), .IN1(\b/n6636 ), .SEL(msg[122]), .F(
        \b/n6638 ) );
  MUX \b/U6752  ( .IN0(\b/n59 ), .IN1(n728), .SEL(msg[127]), .F(\b/n6637 ) );
  MUX \b/U6751  ( .IN0(\b/n6635 ), .IN1(n722), .SEL(msg[127]), .F(\b/n6636 )
         );
  NAND \b/U6750  ( .A(\b/n71 ), .B(\b/n30 ), .Z(\b/n6635 ) );
  MUX \b/U6749  ( .IN0(\b/n6633 ), .IN1(\b/n6632 ), .SEL(msg[122]), .F(
        \b/n6634 ) );
  MUX \b/U6748  ( .IN0(\b/n7 ), .IN1(\b/n6535 ), .SEL(msg[127]), .F(\b/n6633 )
         );
  MUX \b/U6747  ( .IN0(\b/n6525 ), .IN1(\b/n6631 ), .SEL(msg[127]), .F(
        \b/n6632 ) );
  AND \b/U6746  ( .A(msg[121]), .B(msg[124]), .Z(\b/n6631 ) );
  MUX \b/U6745  ( .IN0(\b/n6629 ), .IN1(\b/n6626 ), .SEL(msg[125]), .F(
        \b/n6630 ) );
  MUX \b/U6744  ( .IN0(\b/n6628 ), .IN1(\b/n6627 ), .SEL(msg[122]), .F(
        \b/n6629 ) );
  MUX \b/U6743  ( .IN0(\b/n6564 ), .IN1(\b/n68 ), .SEL(msg[127]), .F(\b/n6628 ) );
  MUX \b/U6742  ( .IN0(\b/n43 ), .IN1(\b/n6533 ), .SEL(msg[127]), .F(\b/n6627 ) );
  MUX \b/U6741  ( .IN0(\b/n6623 ), .IN1(\b/n6624 ), .SEL(msg[122]), .F(
        \b/n6626 ) );
  AND \b/U6740  ( .A(\b/n6625 ), .B(\b/n6580 ), .Z(\b/n6624 ) );
  MUX \b/U6739  ( .IN0(\b/n6539 ), .IN1(\b/n6528 ), .SEL(msg[127]), .F(
        \b/n6623 ) );
  MUX \b/U6738  ( .IN0(\b/n6621 ), .IN1(\b/n6613 ), .SEL(msg[120]), .F(
        \b/n6622 ) );
  MUX \b/U6737  ( .IN0(\b/n6620 ), .IN1(\b/n6616 ), .SEL(msg[125]), .F(
        \b/n6621 ) );
  MUX \b/U6736  ( .IN0(\b/n6619 ), .IN1(\b/n6618 ), .SEL(msg[122]), .F(
        \b/n6620 ) );
  MUX \b/U6735  ( .IN0(\b/n6527 ), .IN1(\b/n32 ), .SEL(msg[127]), .F(\b/n6619 ) );
  MUX \b/U6734  ( .IN0(\b/n6617 ), .IN1(\b/n16 ), .SEL(msg[127]), .F(\b/n6618 ) );
  MUX \b/U6733  ( .IN0(\b/n6525 ), .IN1(\b/n24 ), .SEL(msg[121]), .F(\b/n6617 ) );
  MUX \b/U6732  ( .IN0(\b/n6615 ), .IN1(\b/n6614 ), .SEL(msg[122]), .F(
        \b/n6616 ) );
  MUX \b/U6731  ( .IN0(\b/n63 ), .IN1(\b/n41 ), .SEL(msg[127]), .F(\b/n6615 )
         );
  MUX \b/U6730  ( .IN0(\b/n59 ), .IN1(\b/n19 ), .SEL(msg[127]), .F(\b/n6614 )
         );
  MUX \b/U6729  ( .IN0(\b/n6612 ), .IN1(\b/n6607 ), .SEL(msg[125]), .F(
        \b/n6613 ) );
  MUX \b/U6728  ( .IN0(\b/n6611 ), .IN1(\b/n6608 ), .SEL(msg[122]), .F(
        \b/n6612 ) );
  MUX \b/U6727  ( .IN0(\b/n6609 ), .IN1(\b/n6610 ), .SEL(msg[127]), .F(
        \b/n6611 ) );
  NAND \b/U6726  ( .A(\b/n6528 ), .B(\b/n6600 ), .Z(\b/n6610 ) );
  MUX \b/U6725  ( .IN0(\b/n6528 ), .IN1(\b/n24 ), .SEL(msg[121]), .F(\b/n6609 ) );
  MUX \b/U6724  ( .IN0(\b/n6545 ), .IN1(\b/n6543 ), .SEL(msg[127]), .F(
        \b/n6608 ) );
  MUX \b/U6723  ( .IN0(\b/n6563 ), .IN1(\b/n6606 ), .SEL(msg[122]), .F(
        \b/n6607 ) );
  MUX \b/U6722  ( .IN0(\b/n30 ), .IN1(\b/n62 ), .SEL(msg[127]), .F(\b/n6606 )
         );
  MUX \b/U6721  ( .IN0(\b/n6605 ), .IN1(\b/n6588 ), .SEL(msg[126]), .F(
        shift_row_out[24]) );
  MUX \b/U6720  ( .IN0(\b/n6604 ), .IN1(\b/n6596 ), .SEL(msg[120]), .F(
        \b/n6605 ) );
  MUX \b/U6719  ( .IN0(\b/n6603 ), .IN1(\b/n6601 ), .SEL(msg[122]), .F(
        \b/n6604 ) );
  MUX \b/U6718  ( .IN0(\b/n4 ), .IN1(\b/n6602 ), .SEL(msg[127]), .F(\b/n6603 )
         );
  MUX \b/U6717  ( .IN0(\b/n57 ), .IN1(\b/n60 ), .SEL(msg[125]), .F(\b/n6602 )
         );
  MUX \b/U6716  ( .IN0(\b/n6598 ), .IN1(\b/n6597 ), .SEL(msg[127]), .F(
        \b/n6601 ) );
  NAND \b/U6715  ( .A(\b/n6599 ), .B(\b/n6600 ), .Z(\b/n6598 ) );
  MUX \b/U6714  ( .IN0(\b/n56 ), .IN1(\b/n71 ), .SEL(msg[125]), .F(\b/n6597 )
         );
  MUX \b/U6713  ( .IN0(\b/n6595 ), .IN1(\b/n6591 ), .SEL(msg[122]), .F(
        \b/n6596 ) );
  MUX \b/U6712  ( .IN0(\b/n6594 ), .IN1(\b/n6592 ), .SEL(msg[127]), .F(
        \b/n6595 ) );
  MUX \b/U6711  ( .IN0(\b/n6593 ), .IN1(\b/n9 ), .SEL(msg[125]), .F(\b/n6594 )
         );
  NAND \b/U6710  ( .A(\b/n71 ), .B(\b/n6520 ), .Z(\b/n6593 ) );
  MUX \b/U6708  ( .IN0(\b/n6590 ), .IN1(\b/n6589 ), .SEL(msg[127]), .F(
        \b/n6591 ) );
  MUX \b/U6707  ( .IN0(n723), .IN1(\b/n6 ), .SEL(msg[125]), .F(\b/n6590 ) );
  MUX \b/U6706  ( .IN0(\b/n58 ), .IN1(\b/n14 ), .SEL(msg[125]), .F(\b/n6589 )
         );
  MUX \b/U6705  ( .IN0(\b/n6587 ), .IN1(\b/n6577 ), .SEL(msg[120]), .F(
        \b/n6588 ) );
  MUX \b/U6704  ( .IN0(\b/n6586 ), .IN1(\b/n6582 ), .SEL(msg[122]), .F(
        \b/n6587 ) );
  MUX \b/U6703  ( .IN0(\b/n6585 ), .IN1(\b/n6584 ), .SEL(msg[127]), .F(
        \b/n6586 ) );
  MUX \b/U6702  ( .IN0(n721), .IN1(\b/n10 ), .SEL(msg[125]), .F(\b/n6585 ) );
  MUX \b/U6701  ( .IN0(\b/n6583 ), .IN1(\b/n47 ), .SEL(msg[125]), .F(\b/n6584 ) );
  NAND \b/U6700  ( .A(\b/n6519 ), .B(\b/n6521 ), .Z(\b/n6583 ) );
  MUX \b/U6699  ( .IN0(\b/n6581 ), .IN1(\b/n6578 ), .SEL(msg[127]), .F(
        \b/n6582 ) );
  MUX \b/U6698  ( .IN0(\b/n17 ), .IN1(\b/n6579 ), .SEL(msg[125]), .F(\b/n6581 ) );
  NAND \b/U6697  ( .A(\b/n6523 ), .B(\b/n6580 ), .Z(\b/n6579 ) );
  MUX \b/U6696  ( .IN0(\b/n6538 ), .IN1(\b/n6529 ), .SEL(msg[125]), .F(
        \b/n6578 ) );
  MUX \b/U6695  ( .IN0(\b/n6576 ), .IN1(\b/n6572 ), .SEL(msg[122]), .F(
        \b/n6577 ) );
  MUX \b/U6694  ( .IN0(\b/n6574 ), .IN1(\b/n6573 ), .SEL(msg[127]), .F(
        \b/n6576 ) );
  NAND \b/U6693  ( .A(\b/n6575 ), .B(\b/n6562 ), .Z(\b/n6574 ) );
  MUX \b/U6692  ( .IN0(msg[123]), .IN1(\b/n6554 ), .SEL(msg[125]), .F(
        \b/n6573 ) );
  MUX \b/U6691  ( .IN0(\b/n6571 ), .IN1(\b/n6570 ), .SEL(msg[127]), .F(
        \b/n6572 ) );
  MUX \b/U6690  ( .IN0(\b/n22 ), .IN1(\b/n38 ), .SEL(msg[125]), .F(\b/n6571 )
         );
  MUX \b/U6689  ( .IN0(\b/n55 ), .IN1(\b/n43 ), .SEL(msg[125]), .F(\b/n6570 )
         );
  XOR \b/U6688  ( .A(\b/n6520 ), .B(msg[121]), .Z(\b/n6569 ) );
  XOR \b/U6687  ( .A(msg[121]), .B(msg[122]), .Z(\b/n6568 ) );
  XOR \b/U6686  ( .A(msg[121]), .B(msg[123]), .Z(\b/n6567 ) );
  XOR \b/U6685  ( .A(msg[122]), .B(msg[127]), .Z(\b/n6566 ) );
  XOR \b/U6684  ( .A(\b/n71 ), .B(\b/n14 ), .Z(\b/n6565 ) );
  XOR \b/U6683  ( .A(msg[121]), .B(\b/n60 ), .Z(\b/n6564 ) );
  XOR \b/U6681  ( .A(msg[121]), .B(msg[125]), .Z(\b/n6562 ) );
  NAND \b/U6680  ( .A(msg[121]), .B(msg[123]), .Z(\b/n6561 ) );
  MUX \b/U6679  ( .IN0(\b/n6520 ), .IN1(\b/n14 ), .SEL(msg[121]), .F(\b/n6560 ) );
  MUX \b/U6677  ( .IN0(msg[123]), .IN1(\b/n51 ), .SEL(msg[121]), .F(\b/n6558 )
         );
  MUX \b/U6676  ( .IN0(\b/n30 ), .IN1(\b/n51 ), .SEL(msg[121]), .F(\b/n6557 )
         );
  MUX \b/U6675  ( .IN0(\b/n6523 ), .IN1(\b/n6525 ), .SEL(msg[121]), .F(
        \b/n6556 ) );
  MUX \b/U6674  ( .IN0(msg[124]), .IN1(\b/n30 ), .SEL(msg[121]), .F(\b/n6555 )
         );
  OR \b/U6673  ( .A(msg[121]), .B(msg[124]), .Z(\b/n6554 ) );
  NAND \b/U6671  ( .A(\b/n51 ), .B(\b/n71 ), .Z(\b/n6552 ) );
  MUX \b/U6670  ( .IN0(\b/n51 ), .IN1(msg[124]), .SEL(msg[121]), .F(\b/n6551 )
         );
  MUX \b/U6669  ( .IN0(\b/n6519 ), .IN1(\b/n6528 ), .SEL(msg[121]), .F(
        \b/n6550 ) );
  MUX \b/U6668  ( .IN0(\b/n66 ), .IN1(msg[124]), .SEL(msg[121]), .F(\b/n6549 )
         );
  MUX \b/U6667  ( .IN0(\b/n24 ), .IN1(\b/n51 ), .SEL(msg[121]), .F(\b/n6548 )
         );
  MUX \b/U6666  ( .IN0(\b/n6519 ), .IN1(msg[124]), .SEL(msg[121]), .F(
        \b/n6547 ) );
  MUX \b/U6665  ( .IN0(\b/n41 ), .IN1(\b/n30 ), .SEL(msg[121]), .F(\b/n6546 )
         );
  XOR \b/U6664  ( .A(\b/n24 ), .B(msg[121]), .Z(\b/n6545 ) );
  MUX \b/U6663  ( .IN0(\b/n6525 ), .IN1(\b/n41 ), .SEL(msg[121]), .F(\b/n6544 ) );
  NANDN \b/U6662  ( .B(msg[121]), .A(msg[123]), .Z(\b/n6543 ) );
  MUX \b/U6661  ( .IN0(\b/n14 ), .IN1(msg[123]), .SEL(msg[121]), .F(\b/n6542 )
         );
  NAND \b/U6659  ( .A(\b/n6523 ), .B(\b/n71 ), .Z(\b/n6540 ) );
  MUX \b/U6658  ( .IN0(msg[124]), .IN1(\b/n6520 ), .SEL(msg[121]), .F(
        \b/n6539 ) );
  MUX \b/U6657  ( .IN0(\b/n41 ), .IN1(msg[123]), .SEL(msg[121]), .F(\b/n6538 )
         );
  MUX \b/U6655  ( .IN0(msg[124]), .IN1(\b/n60 ), .SEL(msg[121]), .F(\b/n6536 )
         );
  MUX \b/U6654  ( .IN0(\b/n14 ), .IN1(\b/n66 ), .SEL(msg[121]), .F(\b/n6535 )
         );
  NAND \b/U6653  ( .A(\b/n6521 ), .B(\b/n14 ), .Z(\b/n6534 ) );
  MUX \b/U6652  ( .IN0(\b/n6520 ), .IN1(\b/n6528 ), .SEL(msg[121]), .F(
        \b/n6533 ) );
  NAND \b/U6651  ( .A(\b/n6532 ), .B(\b/n6519 ), .Z(\b/n6531 ) );
  MUX \b/U6650  ( .IN0(\b/n6523 ), .IN1(\b/n66 ), .SEL(msg[121]), .F(\b/n6530 ) );
  MUX \b/U6649  ( .IN0(\b/n66 ), .IN1(\b/n30 ), .SEL(msg[121]), .F(\b/n6529 )
         );
  NANDN \b/U6648  ( .B(msg[123]), .A(msg[124]), .Z(\b/n6528 ) );
  MUX \b/U6647  ( .IN0(\b/n6523 ), .IN1(msg[123]), .SEL(msg[121]), .F(
        \b/n6527 ) );
  OR \b/U6646  ( .A(msg[123]), .B(msg[124]), .Z(\b/n6523 ) );
  MUX \b/U6645  ( .IN0(\b/n14 ), .IN1(\b/n30 ), .SEL(msg[121]), .F(\b/n6526 )
         );
  XOR \b/U6644  ( .A(\b/n24 ), .B(msg[123]), .Z(\b/n6525 ) );
  NANDN \b/U6643  ( .B(msg[123]), .A(msg[121]), .Z(\b/n6524 ) );
  NAND \b/U6642  ( .A(\b/n6523 ), .B(\b/n6521 ), .Z(\b/n6522 ) );
  NAND \b/U6641  ( .A(msg[121]), .B(\b/n6520 ), .Z(\b/n6521 ) );
  NANDN \b/U6640  ( .B(msg[124]), .A(msg[123]), .Z(\b/n6520 ) );
  NAND \b/U6639  ( .A(msg[123]), .B(msg[124]), .Z(\b/n6519 ) );
  MUX \b/U6638  ( .IN0(msg[116]), .IN1(\b/n6160 ), .SEL(msg[113]), .F(
        \b/n6518 ) );
  MUX \b/U6637  ( .IN0(msg[116]), .IN1(\b/n6169 ), .SEL(msg[113]), .F(
        \b/n6517 ) );
  MUX \b/U6636  ( .IN0(\b/n6161 ), .IN1(\b/n6164 ), .SEL(msg[113]), .F(
        \b/n6516 ) );
  MUX \b/U6635  ( .IN0(\b/n6166 ), .IN1(\b/n131 ), .SEL(msg[113]), .F(
        \b/n6515 ) );
  MUX \b/U6633  ( .IN0(\b/n6169 ), .IN1(\b/n6160 ), .SEL(msg[114]), .F(
        \b/n6342 ) );
  MUX \b/U6632  ( .IN0(\b/n6162 ), .IN1(\b/n142 ), .SEL(msg[114]), .F(
        \b/n6343 ) );
  MUX \b/U6631  ( .IN0(\b/n85 ), .IN1(\b/n95 ), .SEL(msg[113]), .F(\b/n6306 )
         );
  MUX \b/U6630  ( .IN0(\b/n6190 ), .IN1(\b/n6501 ), .SEL(msg[119]), .F(
        \b/n6513 ) );
  MUX \b/U6629  ( .IN0(\b/n6164 ), .IN1(\b/n6160 ), .SEL(msg[113]), .F(
        \b/n6504 ) );
  MUX \b/U6628  ( .IN0(\b/n137 ), .IN1(\b/n6166 ), .SEL(msg[113]), .F(
        \b/n6512 ) );
  MUX \b/U6627  ( .IN0(msg[115]), .IN1(\b/n131 ), .SEL(msg[113]), .F(\b/n6511 ) );
  MUX \b/U6626  ( .IN0(\b/n6169 ), .IN1(\b/n137 ), .SEL(msg[113]), .F(
        \b/n6510 ) );
  MUX \b/U6625  ( .IN0(msg[116]), .IN1(\b/n6166 ), .SEL(msg[113]), .F(
        \b/n6509 ) );
  MUX \b/U6624  ( .IN0(\b/n122 ), .IN1(\b/n101 ), .SEL(msg[117]), .F(\b/n6216 ) );
  MUX \b/U6623  ( .IN0(\b/n6161 ), .IN1(\b/n95 ), .SEL(msg[113]), .F(\b/n6508 ) );
  NANDN \b/U6620  ( .B(\b/n6167 ), .A(msg[119]), .Z(\b/n6481 ) );
  NAND \b/U6619  ( .A(msg[119]), .B(\b/n98 ), .Z(\b/n6449 ) );
  NAND \b/U6618  ( .A(msg[119]), .B(\b/n110 ), .Z(\b/n6390 ) );
  NAND \b/U6617  ( .A(msg[119]), .B(\b/n6498 ), .Z(\b/n6423 ) );
  NAND \b/U6616  ( .A(msg[119]), .B(\b/n6418 ), .Z(\b/n6381 ) );
  NAND \b/U6614  ( .A(\b/n142 ), .B(\b/n131 ), .Z(\b/n6502 ) );
  NAND \b/U6613  ( .A(msg[119]), .B(\b/n6500 ), .Z(\b/n6495 ) );
  NAND \b/U6612  ( .A(n720), .B(msg[119]), .Z(\b/n6475 ) );
  NAND \b/U6610  ( .A(msg[114]), .B(\b/n6169 ), .Z(\b/n6335 ) );
  NAND \b/U6609  ( .A(\b/n131 ), .B(msg[113]), .Z(\b/n6290 ) );
  NAND \b/U6608  ( .A(msg[119]), .B(\b/n6504 ), .Z(\b/n6289 ) );
  NAND \b/U6606  ( .A(\b/n6502 ), .B(msg[119]), .Z(\b/n6305 ) );
  NAND \b/U6605  ( .A(\b/n6323 ), .B(\b/n6169 ), .Z(\b/n6501 ) );
  NANDN \b/U6604  ( .B(\b/n85 ), .A(\b/n142 ), .Z(\b/n6500 ) );
  NAND \b/U6602  ( .A(msg[113]), .B(\b/n6169 ), .Z(\b/n6221 ) );
  NAND \b/U6601  ( .A(\b/n85 ), .B(\b/n142 ), .Z(\b/n6498 ) );
  NAND \b/U6598  ( .A(msg[113]), .B(\b/n6164 ), .Z(\b/n6323 ) );
  ANDN \b/U6596  ( .A(msg[114]), .B(msg[113]), .Z(\b/n6351 ) );
  AND \b/U6595  ( .A(\b/n6161 ), .B(\b/n6495 ), .Z(\b/n6266 ) );
  MUX \b/U6594  ( .IN0(\b/n6494 ), .IN1(\b/n6478 ), .SEL(msg[118]), .F(
        shift_row_out[55]) );
  MUX \b/U6593  ( .IN0(\b/n6493 ), .IN1(\b/n6486 ), .SEL(msg[112]), .F(
        \b/n6494 ) );
  MUX \b/U6592  ( .IN0(\b/n6492 ), .IN1(\b/n6489 ), .SEL(msg[117]), .F(
        \b/n6493 ) );
  MUX \b/U6591  ( .IN0(\b/n6491 ), .IN1(\b/n6490 ), .SEL(msg[114]), .F(
        \b/n6492 ) );
  MUX \b/U6590  ( .IN0(msg[116]), .IN1(\b/n102 ), .SEL(msg[119]), .F(\b/n6491 ) );
  MUX \b/U6589  ( .IN0(\b/n6162 ), .IN1(\b/n106 ), .SEL(msg[119]), .F(
        \b/n6490 ) );
  MUX \b/U6588  ( .IN0(\b/n6488 ), .IN1(\b/n6487 ), .SEL(msg[114]), .F(
        \b/n6489 ) );
  MUX \b/U6587  ( .IN0(\b/n6220 ), .IN1(\b/n98 ), .SEL(msg[119]), .F(\b/n6488 ) );
  MUX \b/U6586  ( .IN0(\b/n6172 ), .IN1(\b/n6183 ), .SEL(msg[119]), .F(
        \b/n6487 ) );
  MUX \b/U6585  ( .IN0(\b/n6485 ), .IN1(\b/n6482 ), .SEL(msg[117]), .F(
        \b/n6486 ) );
  MUX \b/U6584  ( .IN0(\b/n6484 ), .IN1(\b/n6483 ), .SEL(msg[114]), .F(
        \b/n6485 ) );
  MUX \b/U6583  ( .IN0(\b/n6196 ), .IN1(\b/n6171 ), .SEL(msg[119]), .F(
        \b/n6484 ) );
  MUX \b/U6582  ( .IN0(\b/n110 ), .IN1(\b/n6192 ), .SEL(msg[119]), .F(
        \b/n6483 ) );
  MUX \b/U6581  ( .IN0(\b/n6480 ), .IN1(\b/n6479 ), .SEL(msg[114]), .F(
        \b/n6482 ) );
  AND \b/U6580  ( .A(\b/n100 ), .B(\b/n6481 ), .Z(\b/n6480 ) );
  MUX \b/U6579  ( .IN0(\b/n6176 ), .IN1(n719), .SEL(msg[119]), .F(\b/n6479 )
         );
  MUX \b/U6578  ( .IN0(\b/n6477 ), .IN1(\b/n6469 ), .SEL(msg[112]), .F(
        \b/n6478 ) );
  MUX \b/U6577  ( .IN0(\b/n6476 ), .IN1(\b/n6472 ), .SEL(msg[117]), .F(
        \b/n6477 ) );
  MUX \b/U6576  ( .IN0(\b/n6473 ), .IN1(\b/n6474 ), .SEL(msg[114]), .F(
        \b/n6476 ) );
  NAND \b/U6575  ( .A(\b/n6290 ), .B(\b/n6475 ), .Z(\b/n6474 ) );
  MUX \b/U6574  ( .IN0(\b/n140 ), .IN1(\b/n132 ), .SEL(msg[119]), .F(\b/n6473 ) );
  MUX \b/U6573  ( .IN0(\b/n6471 ), .IN1(\b/n6470 ), .SEL(msg[114]), .F(
        \b/n6472 ) );
  MUX \b/U6572  ( .IN0(\b/n6166 ), .IN1(\b/n6160 ), .SEL(msg[119]), .F(
        \b/n6471 ) );
  MUX \b/U6571  ( .IN0(\b/n133 ), .IN1(\b/n6197 ), .SEL(msg[119]), .F(
        \b/n6470 ) );
  MUX \b/U6570  ( .IN0(\b/n6468 ), .IN1(\b/n6465 ), .SEL(msg[117]), .F(
        \b/n6469 ) );
  MUX \b/U6569  ( .IN0(\b/n6467 ), .IN1(\b/n6466 ), .SEL(msg[114]), .F(
        \b/n6468 ) );
  MUX \b/U6568  ( .IN0(\b/n6201 ), .IN1(\b/n6187 ), .SEL(msg[119]), .F(
        \b/n6467 ) );
  MUX \b/U6567  ( .IN0(\b/n86 ), .IN1(\b/n6169 ), .SEL(msg[119]), .F(\b/n6466 ) );
  MUX \b/U6566  ( .IN0(\b/n6464 ), .IN1(\b/n6463 ), .SEL(msg[114]), .F(
        \b/n6465 ) );
  MUX \b/U6565  ( .IN0(\b/n6202 ), .IN1(\b/n6210 ), .SEL(msg[119]), .F(
        \b/n6464 ) );
  MUX \b/U6564  ( .IN0(\b/n6195 ), .IN1(\b/n6462 ), .SEL(msg[119]), .F(
        \b/n6463 ) );
  MUX \b/U6563  ( .IN0(\b/n137 ), .IN1(\b/n95 ), .SEL(msg[113]), .F(\b/n6462 )
         );
  MUX \b/U6562  ( .IN0(\b/n6461 ), .IN1(\b/n6443 ), .SEL(msg[118]), .F(
        shift_row_out[54]) );
  MUX \b/U6561  ( .IN0(\b/n6460 ), .IN1(\b/n6451 ), .SEL(msg[112]), .F(
        \b/n6461 ) );
  MUX \b/U6560  ( .IN0(\b/n6459 ), .IN1(\b/n6454 ), .SEL(msg[117]), .F(
        \b/n6460 ) );
  MUX \b/U6559  ( .IN0(\b/n6458 ), .IN1(\b/n6456 ), .SEL(msg[114]), .F(
        \b/n6459 ) );
  MUX \b/U6558  ( .IN0(\b/n6457 ), .IN1(\b/n6173 ), .SEL(msg[119]), .F(
        \b/n6458 ) );
  MUX \b/U6557  ( .IN0(\b/n137 ), .IN1(\b/n6160 ), .SEL(msg[113]), .F(
        \b/n6457 ) );
  MUX \b/U6556  ( .IN0(\b/n6455 ), .IN1(\b/n125 ), .SEL(msg[119]), .F(
        \b/n6456 ) );
  MUX \b/U6555  ( .IN0(\b/n6160 ), .IN1(\b/n6161 ), .SEL(msg[113]), .F(
        \b/n6455 ) );
  MUX \b/U6554  ( .IN0(\b/n6453 ), .IN1(\b/n6452 ), .SEL(msg[114]), .F(
        \b/n6454 ) );
  MUX \b/U6553  ( .IN0(n718), .IN1(\b/n6241 ), .SEL(msg[119]), .F(\b/n6453 )
         );
  MUX \b/U6552  ( .IN0(\b/n6199 ), .IN1(\b/n6206 ), .SEL(msg[119]), .F(
        \b/n6452 ) );
  MUX \b/U6551  ( .IN0(\b/n6450 ), .IN1(\b/n6446 ), .SEL(msg[117]), .F(
        \b/n6451 ) );
  MUX \b/U6550  ( .IN0(\b/n6448 ), .IN1(\b/n6447 ), .SEL(msg[114]), .F(
        \b/n6450 ) );
  AND \b/U6549  ( .A(\b/n78 ), .B(\b/n6449 ), .Z(\b/n6448 ) );
  MUX \b/U6548  ( .IN0(\b/n6276 ), .IN1(msg[115]), .SEL(msg[119]), .F(
        \b/n6447 ) );
  MUX \b/U6547  ( .IN0(\b/n6445 ), .IN1(\b/n6444 ), .SEL(msg[114]), .F(
        \b/n6446 ) );
  MUX \b/U6546  ( .IN0(\b/n121 ), .IN1(\b/n6164 ), .SEL(msg[119]), .F(
        \b/n6445 ) );
  MUX \b/U6544  ( .IN0(\b/n6442 ), .IN1(\b/n6435 ), .SEL(msg[112]), .F(
        \b/n6443 ) );
  MUX \b/U6543  ( .IN0(\b/n6441 ), .IN1(\b/n6438 ), .SEL(msg[117]), .F(
        \b/n6442 ) );
  MUX \b/U6542  ( .IN0(\b/n6440 ), .IN1(\b/n6439 ), .SEL(msg[114]), .F(
        \b/n6441 ) );
  MUX \b/U6541  ( .IN0(\b/n117 ), .IN1(\b/n6168 ), .SEL(msg[119]), .F(
        \b/n6440 ) );
  MUX \b/U6540  ( .IN0(\b/n6172 ), .IN1(n719), .SEL(msg[119]), .F(\b/n6439 )
         );
  MUX \b/U6539  ( .IN0(\b/n6437 ), .IN1(\b/n6436 ), .SEL(msg[114]), .F(
        \b/n6438 ) );
  MUX \b/U6538  ( .IN0(\b/n6188 ), .IN1(\b/n82 ), .SEL(msg[119]), .F(\b/n6437 ) );
  MUX \b/U6537  ( .IN0(\b/n102 ), .IN1(\b/n132 ), .SEL(msg[119]), .F(\b/n6436 ) );
  MUX \b/U6536  ( .IN0(\b/n6434 ), .IN1(\b/n6430 ), .SEL(msg[117]), .F(
        \b/n6435 ) );
  MUX \b/U6535  ( .IN0(\b/n6433 ), .IN1(\b/n6432 ), .SEL(msg[114]), .F(
        \b/n6434 ) );
  MUX \b/U6534  ( .IN0(\b/n6177 ), .IN1(\b/n132 ), .SEL(msg[119]), .F(
        \b/n6433 ) );
  MUX \b/U6533  ( .IN0(\b/n6431 ), .IN1(\b/n6198 ), .SEL(msg[119]), .F(
        \b/n6432 ) );
  NANDN \b/U6532  ( .B(msg[116]), .A(msg[113]), .Z(\b/n6431 ) );
  MUX \b/U6531  ( .IN0(\b/n6429 ), .IN1(\b/n6427 ), .SEL(msg[114]), .F(
        \b/n6430 ) );
  MUX \b/U6530  ( .IN0(\b/n95 ), .IN1(\b/n6428 ), .SEL(msg[119]), .F(\b/n6429 ) );
  MUX \b/U6529  ( .IN0(\b/n122 ), .IN1(\b/n112 ), .SEL(msg[113]), .F(\b/n6428 ) );
  MUX \b/U6528  ( .IN0(\b/n84 ), .IN1(\b/n6173 ), .SEL(msg[119]), .F(\b/n6427 ) );
  NANDN \b/U6527  ( .B(\b/n85 ), .A(msg[113]), .Z(\b/n6173 ) );
  MUX \b/U6526  ( .IN0(\b/n6426 ), .IN1(\b/n6405 ), .SEL(msg[118]), .F(
        shift_row_out[53]) );
  MUX \b/U6525  ( .IN0(\b/n6425 ), .IN1(\b/n6415 ), .SEL(msg[112]), .F(
        \b/n6426 ) );
  MUX \b/U6524  ( .IN0(\b/n6424 ), .IN1(\b/n6420 ), .SEL(msg[117]), .F(
        \b/n6425 ) );
  MUX \b/U6523  ( .IN0(\b/n6421 ), .IN1(\b/n6422 ), .SEL(msg[114]), .F(
        \b/n6424 ) );
  AND \b/U6522  ( .A(\b/n6191 ), .B(\b/n6423 ), .Z(\b/n6422 ) );
  MUX \b/U6521  ( .IN0(\b/n6169 ), .IN1(\b/n133 ), .SEL(msg[119]), .F(
        \b/n6421 ) );
  MUX \b/U6520  ( .IN0(\b/n6419 ), .IN1(\b/n6417 ), .SEL(msg[114]), .F(
        \b/n6420 ) );
  MUX \b/U6519  ( .IN0(\b/n88 ), .IN1(\b/n6418 ), .SEL(msg[119]), .F(\b/n6419 ) );
  NAND \b/U6518  ( .A(\b/n112 ), .B(\b/n142 ), .Z(\b/n6418 ) );
  MUX \b/U6517  ( .IN0(\b/n6169 ), .IN1(\b/n6416 ), .SEL(msg[119]), .F(
        \b/n6417 ) );
  NAND \b/U6516  ( .A(\b/n6160 ), .B(\b/n6221 ), .Z(\b/n6416 ) );
  MUX \b/U6515  ( .IN0(\b/n6414 ), .IN1(\b/n6410 ), .SEL(msg[117]), .F(
        \b/n6415 ) );
  MUX \b/U6514  ( .IN0(\b/n6413 ), .IN1(\b/n6412 ), .SEL(msg[114]), .F(
        \b/n6414 ) );
  MUX \b/U6513  ( .IN0(\b/n6181 ), .IN1(\b/n135 ), .SEL(msg[119]), .F(
        \b/n6413 ) );
  MUX \b/U6512  ( .IN0(\b/n6206 ), .IN1(\b/n6411 ), .SEL(msg[119]), .F(
        \b/n6412 ) );
  MUX \b/U6511  ( .IN0(\b/n131 ), .IN1(\b/n112 ), .SEL(msg[113]), .F(\b/n6411 ) );
  MUX \b/U6510  ( .IN0(\b/n6409 ), .IN1(\b/n6408 ), .SEL(msg[114]), .F(
        \b/n6410 ) );
  MUX \b/U6509  ( .IN0(\b/n129 ), .IN1(n717), .SEL(msg[119]), .F(\b/n6409 ) );
  MUX \b/U6508  ( .IN0(\b/n6407 ), .IN1(\b/n6406 ), .SEL(msg[119]), .F(
        \b/n6408 ) );
  AND \b/U6507  ( .A(\b/n6166 ), .B(\b/n6241 ), .Z(\b/n6407 ) );
  MUX \b/U6506  ( .IN0(\b/n101 ), .IN1(\b/n85 ), .SEL(msg[113]), .F(\b/n6406 )
         );
  MUX \b/U6505  ( .IN0(\b/n6404 ), .IN1(\b/n6395 ), .SEL(msg[112]), .F(
        \b/n6405 ) );
  MUX \b/U6504  ( .IN0(\b/n6403 ), .IN1(\b/n6399 ), .SEL(msg[117]), .F(
        \b/n6404 ) );
  MUX \b/U6503  ( .IN0(\b/n6402 ), .IN1(\b/n6400 ), .SEL(msg[114]), .F(
        \b/n6403 ) );
  MUX \b/U6502  ( .IN0(\b/n6172 ), .IN1(\b/n6401 ), .SEL(msg[119]), .F(
        \b/n6402 ) );
  NAND \b/U6501  ( .A(msg[113]), .B(\b/n101 ), .Z(\b/n6401 ) );
  MUX \b/U6500  ( .IN0(\b/n85 ), .IN1(\b/n138 ), .SEL(msg[119]), .F(\b/n6400 )
         );
  MUX \b/U6499  ( .IN0(\b/n6398 ), .IN1(\b/n6397 ), .SEL(msg[114]), .F(
        \b/n6399 ) );
  MUX \b/U6498  ( .IN0(\b/n6198 ), .IN1(\b/n103 ), .SEL(msg[119]), .F(
        \b/n6398 ) );
  MUX \b/U6497  ( .IN0(\b/n6396 ), .IN1(\b/n6161 ), .SEL(n716), .F(\b/n6397 )
         );
  AND \b/U6496  ( .A(msg[119]), .B(msg[115]), .Z(\b/n6396 ) );
  MUX \b/U6495  ( .IN0(\b/n6394 ), .IN1(\b/n6391 ), .SEL(msg[117]), .F(
        \b/n6395 ) );
  MUX \b/U6494  ( .IN0(\b/n6393 ), .IN1(\b/n6392 ), .SEL(msg[114]), .F(
        \b/n6394 ) );
  MUX \b/U6493  ( .IN0(\b/n6322 ), .IN1(\b/n6161 ), .SEL(msg[119]), .F(
        \b/n6393 ) );
  MUX \b/U6492  ( .IN0(n715), .IN1(\b/n136 ), .SEL(msg[119]), .F(\b/n6392 ) );
  MUX \b/U6491  ( .IN0(\b/n6389 ), .IN1(\b/n6388 ), .SEL(msg[114]), .F(
        \b/n6391 ) );
  AND \b/U6490  ( .A(\b/n6390 ), .B(\b/n6290 ), .Z(\b/n6389 ) );
  MUX \b/U6489  ( .IN0(\b/n87 ), .IN1(\b/n131 ), .SEL(msg[119]), .F(\b/n6388 )
         );
  MUX \b/U6488  ( .IN0(\b/n6387 ), .IN1(\b/n6370 ), .SEL(msg[118]), .F(
        shift_row_out[52]) );
  MUX \b/U6487  ( .IN0(\b/n6386 ), .IN1(\b/n6378 ), .SEL(msg[112]), .F(
        \b/n6387 ) );
  MUX \b/U6486  ( .IN0(\b/n6385 ), .IN1(\b/n6382 ), .SEL(msg[117]), .F(
        \b/n6386 ) );
  MUX \b/U6485  ( .IN0(\b/n6384 ), .IN1(\b/n6383 ), .SEL(msg[114]), .F(
        \b/n6385 ) );
  MUX \b/U6484  ( .IN0(\b/n113 ), .IN1(\b/n134 ), .SEL(msg[119]), .F(\b/n6384 ) );
  MUX \b/U6483  ( .IN0(\b/n6241 ), .IN1(\b/n6206 ), .SEL(msg[119]), .F(
        \b/n6383 ) );
  NAND \b/U6482  ( .A(msg[113]), .B(\b/n6160 ), .Z(\b/n6241 ) );
  MUX \b/U6481  ( .IN0(\b/n6379 ), .IN1(\b/n6380 ), .SEL(msg[114]), .F(
        \b/n6382 ) );
  AND \b/U6480  ( .A(\b/n6191 ), .B(\b/n6381 ), .Z(\b/n6380 ) );
  MUX \b/U6479  ( .IN0(\b/n6189 ), .IN1(\b/n116 ), .SEL(msg[119]), .F(
        \b/n6379 ) );
  MUX \b/U6478  ( .IN0(\b/n6377 ), .IN1(\b/n6374 ), .SEL(msg[117]), .F(
        \b/n6378 ) );
  MUX \b/U6477  ( .IN0(\b/n6376 ), .IN1(\b/n6375 ), .SEL(msg[114]), .F(
        \b/n6377 ) );
  MUX \b/U6476  ( .IN0(\b/n78 ), .IN1(\b/n124 ), .SEL(msg[119]), .F(\b/n6376 )
         );
  MUX \b/U6475  ( .IN0(\b/n85 ), .IN1(\b/n6169 ), .SEL(msg[119]), .F(\b/n6375 ) );
  MUX \b/U6474  ( .IN0(\b/n6373 ), .IN1(\b/n6371 ), .SEL(msg[114]), .F(
        \b/n6374 ) );
  MUX \b/U6473  ( .IN0(\b/n6185 ), .IN1(\b/n6372 ), .SEL(msg[119]), .F(
        \b/n6373 ) );
  AND \b/U6472  ( .A(\b/n6169 ), .B(\b/n142 ), .Z(\b/n6372 ) );
  MUX \b/U6471  ( .IN0(\b/n100 ), .IN1(\b/n119 ), .SEL(msg[119]), .F(\b/n6371 ) );
  MUX \b/U6470  ( .IN0(\b/n6369 ), .IN1(\b/n6363 ), .SEL(msg[112]), .F(
        \b/n6370 ) );
  MUX \b/U6469  ( .IN0(\b/n6368 ), .IN1(\b/n6366 ), .SEL(msg[117]), .F(
        \b/n6369 ) );
  MUX \b/U6468  ( .IN0(\b/n6367 ), .IN1(\b/n6163 ), .SEL(msg[114]), .F(
        \b/n6368 ) );
  MUX \b/U6467  ( .IN0(\b/n6183 ), .IN1(\b/n121 ), .SEL(msg[119]), .F(
        \b/n6367 ) );
  MUX \b/U6466  ( .IN0(\b/n6365 ), .IN1(\b/n6364 ), .SEL(msg[114]), .F(
        \b/n6366 ) );
  MUX \b/U6465  ( .IN0(n714), .IN1(\b/n113 ), .SEL(msg[119]), .F(\b/n6365 ) );
  MUX \b/U6464  ( .IN0(\b/n6193 ), .IN1(\b/n6196 ), .SEL(msg[119]), .F(
        \b/n6364 ) );
  MUX \b/U6463  ( .IN0(\b/n6362 ), .IN1(\b/n6359 ), .SEL(msg[117]), .F(
        \b/n6363 ) );
  MUX \b/U6462  ( .IN0(\b/n6361 ), .IN1(\b/n6360 ), .SEL(msg[114]), .F(
        \b/n6362 ) );
  MUX \b/U6461  ( .IN0(\b/n86 ), .IN1(\b/n6165 ), .SEL(msg[119]), .F(\b/n6361 ) );
  MUX \b/U6460  ( .IN0(\b/n131 ), .IN1(\b/n6187 ), .SEL(msg[119]), .F(
        \b/n6360 ) );
  MUX \b/U6459  ( .IN0(\b/n74 ), .IN1(\b/n6358 ), .SEL(msg[114]), .F(\b/n6359 ) );
  MUX \b/U6458  ( .IN0(\b/n94 ), .IN1(\b/n6169 ), .SEL(msg[119]), .F(\b/n6358 ) );
  MUX \b/U6457  ( .IN0(\b/n6357 ), .IN1(\b/n6338 ), .SEL(msg[118]), .F(
        shift_row_out[51]) );
  MUX \b/U6456  ( .IN0(\b/n6356 ), .IN1(\b/n6348 ), .SEL(msg[112]), .F(
        \b/n6357 ) );
  MUX \b/U6455  ( .IN0(\b/n6355 ), .IN1(\b/n6352 ), .SEL(msg[117]), .F(
        \b/n6356 ) );
  MUX \b/U6454  ( .IN0(\b/n6354 ), .IN1(\b/n6353 ), .SEL(msg[119]), .F(
        \b/n6355 ) );
  MUX \b/U6453  ( .IN0(\b/n6177 ), .IN1(\b/n119 ), .SEL(msg[114]), .F(
        \b/n6354 ) );
  MUX \b/U6452  ( .IN0(n717), .IN1(\b/n77 ), .SEL(msg[114]), .F(\b/n6353 ) );
  MUX \b/U6451  ( .IN0(\b/n6350 ), .IN1(\b/n6349 ), .SEL(msg[119]), .F(
        \b/n6352 ) );
  AND \b/U6450  ( .A(\b/n6351 ), .B(msg[116]), .Z(\b/n6350 ) );
  MUX \b/U6449  ( .IN0(\b/n107 ), .IN1(\b/n6190 ), .SEL(msg[114]), .F(
        \b/n6349 ) );
  MUX \b/U6448  ( .IN0(\b/n6347 ), .IN1(\b/n6344 ), .SEL(msg[117]), .F(
        \b/n6348 ) );
  MUX \b/U6447  ( .IN0(\b/n6346 ), .IN1(\b/n6345 ), .SEL(msg[119]), .F(
        \b/n6347 ) );
  MUX \b/U6446  ( .IN0(\b/n6181 ), .IN1(n713), .SEL(msg[114]), .F(\b/n6346 )
         );
  MUX \b/U6445  ( .IN0(\b/n75 ), .IN1(\b/n94 ), .SEL(msg[114]), .F(\b/n6345 )
         );
  MUX \b/U6444  ( .IN0(\b/n6340 ), .IN1(\b/n6341 ), .SEL(msg[119]), .F(
        \b/n6344 ) );
  NAND \b/U6443  ( .A(\b/n6342 ), .B(\b/n6343 ), .Z(\b/n6341 ) );
  MUX \b/U6442  ( .IN0(\b/n120 ), .IN1(\b/n6339 ), .SEL(msg[114]), .F(
        \b/n6340 ) );
  MUX \b/U6441  ( .IN0(\b/n95 ), .IN1(\b/n137 ), .SEL(msg[113]), .F(\b/n6339 )
         );
  MUX \b/U6440  ( .IN0(\b/n6337 ), .IN1(\b/n6328 ), .SEL(msg[112]), .F(
        \b/n6338 ) );
  MUX \b/U6439  ( .IN0(\b/n6336 ), .IN1(\b/n6332 ), .SEL(msg[117]), .F(
        \b/n6337 ) );
  MUX \b/U6438  ( .IN0(\b/n6334 ), .IN1(\b/n6333 ), .SEL(msg[119]), .F(
        \b/n6336 ) );
  NAND \b/U6437  ( .A(\b/n85 ), .B(\b/n6335 ), .Z(\b/n6334 ) );
  MUX \b/U6436  ( .IN0(\b/n136 ), .IN1(\b/n98 ), .SEL(msg[114]), .F(\b/n6333 )
         );
  MUX \b/U6435  ( .IN0(\b/n6331 ), .IN1(\b/n6329 ), .SEL(msg[119]), .F(
        \b/n6332 ) );
  MUX \b/U6434  ( .IN0(\b/n6172 ), .IN1(\b/n6330 ), .SEL(msg[114]), .F(
        \b/n6331 ) );
  AND \b/U6433  ( .A(msg[113]), .B(\b/n85 ), .Z(\b/n6330 ) );
  MUX \b/U6432  ( .IN0(\b/n90 ), .IN1(\b/n6191 ), .SEL(msg[114]), .F(\b/n6329 ) );
  MUX \b/U6431  ( .IN0(\b/n6327 ), .IN1(\b/n6321 ), .SEL(msg[117]), .F(
        \b/n6328 ) );
  MUX \b/U6430  ( .IN0(\b/n6326 ), .IN1(\b/n6324 ), .SEL(msg[119]), .F(
        \b/n6327 ) );
  MUX \b/U6429  ( .IN0(\b/n6325 ), .IN1(\b/n6161 ), .SEL(\b/n6209 ), .F(
        \b/n6326 ) );
  MUX \b/U6428  ( .IN0(msg[115]), .IN1(msg[116]), .SEL(msg[114]), .F(\b/n6325 ) );
  MUX \b/U6427  ( .IN0(\b/n6191 ), .IN1(\b/n6322 ), .SEL(msg[114]), .F(
        \b/n6324 ) );
  NAND \b/U6426  ( .A(\b/n6161 ), .B(\b/n6323 ), .Z(\b/n6322 ) );
  MUX \b/U6425  ( .IN0(\b/n6318 ), .IN1(\b/n6319 ), .SEL(msg[119]), .F(
        \b/n6321 ) );
  AND \b/U6424  ( .A(\b/n118 ), .B(\b/n6320 ), .Z(\b/n6319 ) );
  MUX \b/U6423  ( .IN0(\b/n99 ), .IN1(\b/n6162 ), .SEL(msg[114]), .F(\b/n6318 ) );
  MUX \b/U6422  ( .IN0(\b/n6317 ), .IN1(\b/n6301 ), .SEL(msg[118]), .F(
        shift_row_out[50]) );
  MUX \b/U6421  ( .IN0(\b/n6316 ), .IN1(\b/n6308 ), .SEL(msg[112]), .F(
        \b/n6317 ) );
  MUX \b/U6420  ( .IN0(\b/n6315 ), .IN1(\b/n6311 ), .SEL(msg[117]), .F(
        \b/n6316 ) );
  MUX \b/U6419  ( .IN0(\b/n6314 ), .IN1(\b/n6312 ), .SEL(msg[114]), .F(
        \b/n6315 ) );
  MUX \b/U6418  ( .IN0(\b/n107 ), .IN1(\b/n6313 ), .SEL(msg[119]), .F(
        \b/n6314 ) );
  MUX \b/U6417  ( .IN0(\b/n6169 ), .IN1(\b/n85 ), .SEL(msg[113]), .F(\b/n6313 ) );
  MUX \b/U6416  ( .IN0(\b/n6208 ), .IN1(\b/n125 ), .SEL(msg[119]), .F(
        \b/n6312 ) );
  MUX \b/U6415  ( .IN0(\b/n6310 ), .IN1(\b/n6309 ), .SEL(msg[114]), .F(
        \b/n6311 ) );
  MUX \b/U6414  ( .IN0(\b/n6162 ), .IN1(\b/n92 ), .SEL(msg[119]), .F(\b/n6310 ) );
  MUX \b/U6413  ( .IN0(\b/n128 ), .IN1(\b/n6195 ), .SEL(msg[119]), .F(
        \b/n6309 ) );
  MUX \b/U6412  ( .IN0(\b/n6307 ), .IN1(\b/n6303 ), .SEL(msg[117]), .F(
        \b/n6308 ) );
  MUX \b/U6411  ( .IN0(\b/n6304 ), .IN1(\b/n74 ), .SEL(msg[114]), .F(\b/n6307 ) );
  NAND \b/U6410  ( .A(\b/n6305 ), .B(\b/n6306 ), .Z(\b/n6304 ) );
  MUX \b/U6409  ( .IN0(n715), .IN1(\b/n6302 ), .SEL(\b/n6207 ), .F(\b/n6303 )
         );
  MUX \b/U6408  ( .IN0(\b/n106 ), .IN1(\b/n6174 ), .SEL(msg[114]), .F(
        \b/n6302 ) );
  MUX \b/U6407  ( .IN0(\b/n6300 ), .IN1(\b/n6292 ), .SEL(msg[112]), .F(
        \b/n6301 ) );
  MUX \b/U6406  ( .IN0(\b/n6299 ), .IN1(\b/n6296 ), .SEL(msg[117]), .F(
        \b/n6300 ) );
  MUX \b/U6405  ( .IN0(\b/n6298 ), .IN1(\b/n6297 ), .SEL(msg[114]), .F(
        \b/n6299 ) );
  MUX \b/U6404  ( .IN0(\b/n134 ), .IN1(msg[113]), .SEL(msg[119]), .F(\b/n6298 ) );
  MUX \b/U6403  ( .IN0(n718), .IN1(\b/n6175 ), .SEL(msg[119]), .F(\b/n6297 )
         );
  MUX \b/U6402  ( .IN0(\b/n6295 ), .IN1(\b/n6294 ), .SEL(msg[114]), .F(
        \b/n6296 ) );
  MUX \b/U6401  ( .IN0(\b/n139 ), .IN1(\b/n133 ), .SEL(msg[119]), .F(\b/n6295 ) );
  MUX \b/U6400  ( .IN0(n718), .IN1(\b/n6293 ), .SEL(msg[119]), .F(\b/n6294 )
         );
  MUX \b/U6399  ( .IN0(\b/n85 ), .IN1(\b/n122 ), .SEL(msg[113]), .F(\b/n6293 )
         );
  MUX \b/U6398  ( .IN0(\b/n6291 ), .IN1(\b/n6285 ), .SEL(msg[117]), .F(
        \b/n6292 ) );
  MUX \b/U6397  ( .IN0(\b/n6288 ), .IN1(\b/n6287 ), .SEL(msg[114]), .F(
        \b/n6291 ) );
  NAND \b/U6396  ( .A(\b/n6289 ), .B(\b/n6290 ), .Z(\b/n6288 ) );
  MUX \b/U6395  ( .IN0(\b/n6161 ), .IN1(\b/n6286 ), .SEL(n716), .F(\b/n6287 )
         );
  MUX \b/U6394  ( .IN0(msg[115]), .IN1(\b/n95 ), .SEL(msg[119]), .F(\b/n6286 )
         );
  MUX \b/U6393  ( .IN0(\b/n6284 ), .IN1(\b/n6283 ), .SEL(msg[114]), .F(
        \b/n6285 ) );
  MUX \b/U6392  ( .IN0(\b/n6206 ), .IN1(\b/n93 ), .SEL(msg[119]), .F(\b/n6284 ) );
  MUX \b/U6391  ( .IN0(\b/n6202 ), .IN1(\b/n6282 ), .SEL(msg[119]), .F(
        \b/n6283 ) );
  MUX \b/U6390  ( .IN0(\b/n6164 ), .IN1(\b/n6169 ), .SEL(msg[113]), .F(
        \b/n6282 ) );
  MUX \b/U6389  ( .IN0(\b/n6281 ), .IN1(\b/n6263 ), .SEL(msg[118]), .F(
        shift_row_out[49]) );
  MUX \b/U6388  ( .IN0(\b/n6280 ), .IN1(\b/n6271 ), .SEL(msg[112]), .F(
        \b/n6281 ) );
  MUX \b/U6387  ( .IN0(\b/n6279 ), .IN1(\b/n6275 ), .SEL(msg[117]), .F(
        \b/n6280 ) );
  MUX \b/U6386  ( .IN0(\b/n6278 ), .IN1(\b/n6277 ), .SEL(msg[114]), .F(
        \b/n6279 ) );
  MUX \b/U6385  ( .IN0(\b/n130 ), .IN1(n720), .SEL(msg[119]), .F(\b/n6278 ) );
  MUX \b/U6384  ( .IN0(\b/n6276 ), .IN1(n714), .SEL(msg[119]), .F(\b/n6277 )
         );
  NAND \b/U6383  ( .A(\b/n142 ), .B(\b/n101 ), .Z(\b/n6276 ) );
  MUX \b/U6382  ( .IN0(\b/n6274 ), .IN1(\b/n6273 ), .SEL(msg[114]), .F(
        \b/n6275 ) );
  MUX \b/U6381  ( .IN0(\b/n78 ), .IN1(\b/n6176 ), .SEL(msg[119]), .F(\b/n6274 ) );
  MUX \b/U6380  ( .IN0(\b/n6166 ), .IN1(\b/n6272 ), .SEL(msg[119]), .F(
        \b/n6273 ) );
  AND \b/U6379  ( .A(msg[113]), .B(msg[116]), .Z(\b/n6272 ) );
  MUX \b/U6378  ( .IN0(\b/n6270 ), .IN1(\b/n6267 ), .SEL(msg[117]), .F(
        \b/n6271 ) );
  MUX \b/U6377  ( .IN0(\b/n6269 ), .IN1(\b/n6268 ), .SEL(msg[114]), .F(
        \b/n6270 ) );
  MUX \b/U6376  ( .IN0(\b/n6205 ), .IN1(\b/n139 ), .SEL(msg[119]), .F(
        \b/n6269 ) );
  MUX \b/U6375  ( .IN0(\b/n114 ), .IN1(\b/n6174 ), .SEL(msg[119]), .F(
        \b/n6268 ) );
  MUX \b/U6374  ( .IN0(\b/n6264 ), .IN1(\b/n6265 ), .SEL(msg[114]), .F(
        \b/n6267 ) );
  AND \b/U6373  ( .A(\b/n6266 ), .B(\b/n6221 ), .Z(\b/n6265 ) );
  MUX \b/U6372  ( .IN0(\b/n6180 ), .IN1(\b/n6169 ), .SEL(msg[119]), .F(
        \b/n6264 ) );
  MUX \b/U6371  ( .IN0(\b/n6262 ), .IN1(\b/n6254 ), .SEL(msg[112]), .F(
        \b/n6263 ) );
  MUX \b/U6370  ( .IN0(\b/n6261 ), .IN1(\b/n6257 ), .SEL(msg[117]), .F(
        \b/n6262 ) );
  MUX \b/U6369  ( .IN0(\b/n6260 ), .IN1(\b/n6259 ), .SEL(msg[114]), .F(
        \b/n6261 ) );
  MUX \b/U6368  ( .IN0(\b/n6168 ), .IN1(\b/n103 ), .SEL(msg[119]), .F(
        \b/n6260 ) );
  MUX \b/U6367  ( .IN0(\b/n6258 ), .IN1(\b/n87 ), .SEL(msg[119]), .F(\b/n6259 ) );
  MUX \b/U6366  ( .IN0(\b/n6166 ), .IN1(\b/n95 ), .SEL(msg[113]), .F(\b/n6258 ) );
  MUX \b/U6365  ( .IN0(\b/n6256 ), .IN1(\b/n6255 ), .SEL(msg[114]), .F(
        \b/n6257 ) );
  MUX \b/U6364  ( .IN0(\b/n134 ), .IN1(\b/n112 ), .SEL(msg[119]), .F(\b/n6256 ) );
  MUX \b/U6363  ( .IN0(\b/n130 ), .IN1(\b/n90 ), .SEL(msg[119]), .F(\b/n6255 )
         );
  MUX \b/U6362  ( .IN0(\b/n6253 ), .IN1(\b/n6248 ), .SEL(msg[117]), .F(
        \b/n6254 ) );
  MUX \b/U6361  ( .IN0(\b/n6252 ), .IN1(\b/n6249 ), .SEL(msg[114]), .F(
        \b/n6253 ) );
  MUX \b/U6360  ( .IN0(\b/n6250 ), .IN1(\b/n6251 ), .SEL(msg[119]), .F(
        \b/n6252 ) );
  NAND \b/U6359  ( .A(\b/n6169 ), .B(\b/n6241 ), .Z(\b/n6251 ) );
  MUX \b/U6358  ( .IN0(\b/n6169 ), .IN1(\b/n95 ), .SEL(msg[113]), .F(\b/n6250 ) );
  MUX \b/U6357  ( .IN0(\b/n6186 ), .IN1(\b/n6184 ), .SEL(msg[119]), .F(
        \b/n6249 ) );
  MUX \b/U6356  ( .IN0(\b/n6204 ), .IN1(\b/n6247 ), .SEL(msg[114]), .F(
        \b/n6248 ) );
  MUX \b/U6355  ( .IN0(\b/n101 ), .IN1(\b/n133 ), .SEL(msg[119]), .F(\b/n6247 ) );
  MUX \b/U6354  ( .IN0(\b/n6246 ), .IN1(\b/n6229 ), .SEL(msg[118]), .F(
        shift_row_out[48]) );
  MUX \b/U6353  ( .IN0(\b/n6245 ), .IN1(\b/n6237 ), .SEL(msg[112]), .F(
        \b/n6246 ) );
  MUX \b/U6352  ( .IN0(\b/n6244 ), .IN1(\b/n6242 ), .SEL(msg[114]), .F(
        \b/n6245 ) );
  MUX \b/U6351  ( .IN0(\b/n75 ), .IN1(\b/n6243 ), .SEL(msg[119]), .F(\b/n6244 ) );
  MUX \b/U6350  ( .IN0(\b/n128 ), .IN1(\b/n131 ), .SEL(msg[117]), .F(\b/n6243 ) );
  MUX \b/U6349  ( .IN0(\b/n6239 ), .IN1(\b/n6238 ), .SEL(msg[119]), .F(
        \b/n6242 ) );
  NAND \b/U6348  ( .A(\b/n6240 ), .B(\b/n6241 ), .Z(\b/n6239 ) );
  MUX \b/U6347  ( .IN0(\b/n127 ), .IN1(\b/n142 ), .SEL(msg[117]), .F(\b/n6238 ) );
  MUX \b/U6346  ( .IN0(\b/n6236 ), .IN1(\b/n6232 ), .SEL(msg[114]), .F(
        \b/n6237 ) );
  MUX \b/U6345  ( .IN0(\b/n6235 ), .IN1(\b/n6233 ), .SEL(msg[119]), .F(
        \b/n6236 ) );
  MUX \b/U6344  ( .IN0(\b/n6234 ), .IN1(\b/n80 ), .SEL(msg[117]), .F(\b/n6235 ) );
  NAND \b/U6343  ( .A(\b/n142 ), .B(\b/n6161 ), .Z(\b/n6234 ) );
  MUX \b/U6341  ( .IN0(\b/n6231 ), .IN1(\b/n6230 ), .SEL(msg[119]), .F(
        \b/n6232 ) );
  MUX \b/U6340  ( .IN0(n715), .IN1(\b/n77 ), .SEL(msg[117]), .F(\b/n6231 ) );
  MUX \b/U6339  ( .IN0(\b/n129 ), .IN1(\b/n85 ), .SEL(msg[117]), .F(\b/n6230 )
         );
  MUX \b/U6338  ( .IN0(\b/n6228 ), .IN1(\b/n6218 ), .SEL(msg[112]), .F(
        \b/n6229 ) );
  MUX \b/U6337  ( .IN0(\b/n6227 ), .IN1(\b/n6223 ), .SEL(msg[114]), .F(
        \b/n6228 ) );
  MUX \b/U6336  ( .IN0(\b/n6226 ), .IN1(\b/n6225 ), .SEL(msg[119]), .F(
        \b/n6227 ) );
  MUX \b/U6335  ( .IN0(n713), .IN1(\b/n81 ), .SEL(msg[117]), .F(\b/n6226 ) );
  MUX \b/U6334  ( .IN0(\b/n6224 ), .IN1(\b/n118 ), .SEL(msg[117]), .F(
        \b/n6225 ) );
  NAND \b/U6333  ( .A(\b/n6160 ), .B(\b/n6162 ), .Z(\b/n6224 ) );
  MUX \b/U6332  ( .IN0(\b/n6222 ), .IN1(\b/n6219 ), .SEL(msg[119]), .F(
        \b/n6223 ) );
  MUX \b/U6331  ( .IN0(\b/n88 ), .IN1(\b/n6220 ), .SEL(msg[117]), .F(\b/n6222 ) );
  NAND \b/U6330  ( .A(\b/n6164 ), .B(\b/n6221 ), .Z(\b/n6220 ) );
  MUX \b/U6329  ( .IN0(\b/n6179 ), .IN1(\b/n6170 ), .SEL(msg[117]), .F(
        \b/n6219 ) );
  MUX \b/U6328  ( .IN0(\b/n6217 ), .IN1(\b/n6213 ), .SEL(msg[114]), .F(
        \b/n6218 ) );
  MUX \b/U6327  ( .IN0(\b/n6215 ), .IN1(\b/n6214 ), .SEL(msg[119]), .F(
        \b/n6217 ) );
  NAND \b/U6326  ( .A(\b/n6216 ), .B(\b/n6203 ), .Z(\b/n6215 ) );
  MUX \b/U6325  ( .IN0(msg[115]), .IN1(\b/n6195 ), .SEL(msg[117]), .F(
        \b/n6214 ) );
  MUX \b/U6324  ( .IN0(\b/n6212 ), .IN1(\b/n6211 ), .SEL(msg[119]), .F(
        \b/n6213 ) );
  MUX \b/U6323  ( .IN0(\b/n93 ), .IN1(\b/n109 ), .SEL(msg[117]), .F(\b/n6212 )
         );
  MUX \b/U6322  ( .IN0(\b/n126 ), .IN1(\b/n114 ), .SEL(msg[117]), .F(\b/n6211 ) );
  XOR \b/U6321  ( .A(\b/n6161 ), .B(msg[113]), .Z(\b/n6210 ) );
  XOR \b/U6320  ( .A(msg[113]), .B(msg[114]), .Z(\b/n6209 ) );
  XOR \b/U6319  ( .A(msg[113]), .B(msg[115]), .Z(\b/n6208 ) );
  XOR \b/U6318  ( .A(msg[114]), .B(msg[119]), .Z(\b/n6207 ) );
  XOR \b/U6317  ( .A(\b/n142 ), .B(\b/n85 ), .Z(\b/n6206 ) );
  XOR \b/U6316  ( .A(msg[113]), .B(\b/n131 ), .Z(\b/n6205 ) );
  XOR \b/U6314  ( .A(msg[113]), .B(msg[117]), .Z(\b/n6203 ) );
  NAND \b/U6313  ( .A(msg[113]), .B(msg[115]), .Z(\b/n6202 ) );
  MUX \b/U6312  ( .IN0(\b/n6161 ), .IN1(\b/n85 ), .SEL(msg[113]), .F(\b/n6201 ) );
  MUX \b/U6310  ( .IN0(msg[115]), .IN1(\b/n122 ), .SEL(msg[113]), .F(\b/n6199 ) );
  MUX \b/U6309  ( .IN0(\b/n101 ), .IN1(\b/n122 ), .SEL(msg[113]), .F(\b/n6198 ) );
  MUX \b/U6308  ( .IN0(\b/n6164 ), .IN1(\b/n6166 ), .SEL(msg[113]), .F(
        \b/n6197 ) );
  MUX \b/U6307  ( .IN0(msg[116]), .IN1(\b/n101 ), .SEL(msg[113]), .F(\b/n6196 ) );
  OR \b/U6306  ( .A(msg[113]), .B(msg[116]), .Z(\b/n6195 ) );
  NAND \b/U6304  ( .A(\b/n122 ), .B(\b/n142 ), .Z(\b/n6193 ) );
  MUX \b/U6303  ( .IN0(\b/n122 ), .IN1(msg[116]), .SEL(msg[113]), .F(\b/n6192 ) );
  MUX \b/U6302  ( .IN0(\b/n6160 ), .IN1(\b/n6169 ), .SEL(msg[113]), .F(
        \b/n6191 ) );
  MUX \b/U6301  ( .IN0(\b/n137 ), .IN1(msg[116]), .SEL(msg[113]), .F(\b/n6190 ) );
  MUX \b/U6300  ( .IN0(\b/n95 ), .IN1(\b/n122 ), .SEL(msg[113]), .F(\b/n6189 )
         );
  MUX \b/U6299  ( .IN0(\b/n6160 ), .IN1(msg[116]), .SEL(msg[113]), .F(
        \b/n6188 ) );
  MUX \b/U6298  ( .IN0(\b/n112 ), .IN1(\b/n101 ), .SEL(msg[113]), .F(\b/n6187 ) );
  XOR \b/U6297  ( .A(\b/n95 ), .B(msg[113]), .Z(\b/n6186 ) );
  MUX \b/U6296  ( .IN0(\b/n6166 ), .IN1(\b/n112 ), .SEL(msg[113]), .F(
        \b/n6185 ) );
  NANDN \b/U6295  ( .B(msg[113]), .A(msg[115]), .Z(\b/n6184 ) );
  MUX \b/U6294  ( .IN0(\b/n85 ), .IN1(msg[115]), .SEL(msg[113]), .F(\b/n6183 )
         );
  NAND \b/U6292  ( .A(\b/n6164 ), .B(\b/n142 ), .Z(\b/n6181 ) );
  MUX \b/U6291  ( .IN0(msg[116]), .IN1(\b/n6161 ), .SEL(msg[113]), .F(
        \b/n6180 ) );
  MUX \b/U6290  ( .IN0(\b/n112 ), .IN1(msg[115]), .SEL(msg[113]), .F(\b/n6179 ) );
  MUX \b/U6288  ( .IN0(msg[116]), .IN1(\b/n131 ), .SEL(msg[113]), .F(\b/n6177 ) );
  MUX \b/U6287  ( .IN0(\b/n85 ), .IN1(\b/n137 ), .SEL(msg[113]), .F(\b/n6176 )
         );
  NAND \b/U6286  ( .A(\b/n6162 ), .B(\b/n85 ), .Z(\b/n6175 ) );
  MUX \b/U6285  ( .IN0(\b/n6161 ), .IN1(\b/n6169 ), .SEL(msg[113]), .F(
        \b/n6174 ) );
  NAND \b/U6284  ( .A(\b/n6173 ), .B(\b/n6160 ), .Z(\b/n6172 ) );
  MUX \b/U6283  ( .IN0(\b/n6164 ), .IN1(\b/n137 ), .SEL(msg[113]), .F(
        \b/n6171 ) );
  MUX \b/U6282  ( .IN0(\b/n137 ), .IN1(\b/n101 ), .SEL(msg[113]), .F(\b/n6170 ) );
  NANDN \b/U6281  ( .B(msg[115]), .A(msg[116]), .Z(\b/n6169 ) );
  MUX \b/U6280  ( .IN0(\b/n6164 ), .IN1(msg[115]), .SEL(msg[113]), .F(
        \b/n6168 ) );
  OR \b/U6279  ( .A(msg[115]), .B(msg[116]), .Z(\b/n6164 ) );
  MUX \b/U6278  ( .IN0(\b/n85 ), .IN1(\b/n101 ), .SEL(msg[113]), .F(\b/n6167 )
         );
  XOR \b/U6277  ( .A(\b/n95 ), .B(msg[115]), .Z(\b/n6166 ) );
  NANDN \b/U6276  ( .B(msg[115]), .A(msg[113]), .Z(\b/n6165 ) );
  NAND \b/U6275  ( .A(\b/n6164 ), .B(\b/n6162 ), .Z(\b/n6163 ) );
  NAND \b/U6274  ( .A(msg[113]), .B(\b/n6161 ), .Z(\b/n6162 ) );
  NANDN \b/U6273  ( .B(msg[116]), .A(msg[115]), .Z(\b/n6161 ) );
  NAND \b/U6272  ( .A(msg[115]), .B(msg[116]), .Z(\b/n6160 ) );
  MUX \b/U6271  ( .IN0(msg[108]), .IN1(\b/n5801 ), .SEL(msg[105]), .F(
        \b/n6159 ) );
  MUX \b/U6270  ( .IN0(msg[108]), .IN1(\b/n5810 ), .SEL(msg[105]), .F(
        \b/n6158 ) );
  MUX \b/U6269  ( .IN0(\b/n5802 ), .IN1(\b/n5805 ), .SEL(msg[105]), .F(
        \b/n6157 ) );
  MUX \b/U6268  ( .IN0(\b/n5807 ), .IN1(\b/n202 ), .SEL(msg[105]), .F(
        \b/n6156 ) );
  MUX \b/U6266  ( .IN0(\b/n5810 ), .IN1(\b/n5801 ), .SEL(msg[106]), .F(
        \b/n5983 ) );
  MUX \b/U6265  ( .IN0(\b/n5803 ), .IN1(\b/n213 ), .SEL(msg[106]), .F(
        \b/n5984 ) );
  MUX \b/U6264  ( .IN0(\b/n156 ), .IN1(\b/n166 ), .SEL(msg[105]), .F(\b/n5947 ) );
  MUX \b/U6263  ( .IN0(\b/n5831 ), .IN1(\b/n6142 ), .SEL(msg[111]), .F(
        \b/n6154 ) );
  MUX \b/U6262  ( .IN0(\b/n5805 ), .IN1(\b/n5801 ), .SEL(msg[105]), .F(
        \b/n6145 ) );
  MUX \b/U6261  ( .IN0(\b/n208 ), .IN1(\b/n5807 ), .SEL(msg[105]), .F(
        \b/n6153 ) );
  MUX \b/U6260  ( .IN0(msg[107]), .IN1(\b/n202 ), .SEL(msg[105]), .F(\b/n6152 ) );
  MUX \b/U6259  ( .IN0(\b/n5810 ), .IN1(\b/n208 ), .SEL(msg[105]), .F(
        \b/n6151 ) );
  MUX \b/U6258  ( .IN0(msg[108]), .IN1(\b/n5807 ), .SEL(msg[105]), .F(
        \b/n6150 ) );
  MUX \b/U6257  ( .IN0(\b/n193 ), .IN1(\b/n172 ), .SEL(msg[109]), .F(\b/n5857 ) );
  MUX \b/U6256  ( .IN0(\b/n5802 ), .IN1(\b/n166 ), .SEL(msg[105]), .F(
        \b/n6149 ) );
  NANDN \b/U6253  ( .B(\b/n5808 ), .A(msg[111]), .Z(\b/n6122 ) );
  NAND \b/U6252  ( .A(msg[111]), .B(\b/n169 ), .Z(\b/n6090 ) );
  NAND \b/U6251  ( .A(msg[111]), .B(\b/n181 ), .Z(\b/n6031 ) );
  NAND \b/U6250  ( .A(msg[111]), .B(\b/n6139 ), .Z(\b/n6064 ) );
  NAND \b/U6249  ( .A(msg[111]), .B(\b/n6059 ), .Z(\b/n6022 ) );
  NAND \b/U6247  ( .A(\b/n213 ), .B(\b/n202 ), .Z(\b/n6143 ) );
  NAND \b/U6246  ( .A(msg[111]), .B(\b/n6141 ), .Z(\b/n6136 ) );
  NAND \b/U6245  ( .A(n712), .B(msg[111]), .Z(\b/n6116 ) );
  NAND \b/U6243  ( .A(msg[106]), .B(\b/n5810 ), .Z(\b/n5976 ) );
  NAND \b/U6242  ( .A(\b/n202 ), .B(msg[105]), .Z(\b/n5931 ) );
  NAND \b/U6241  ( .A(msg[111]), .B(\b/n6145 ), .Z(\b/n5930 ) );
  NAND \b/U6239  ( .A(\b/n6143 ), .B(msg[111]), .Z(\b/n5946 ) );
  NAND \b/U6238  ( .A(\b/n5964 ), .B(\b/n5810 ), .Z(\b/n6142 ) );
  NANDN \b/U6237  ( .B(\b/n156 ), .A(\b/n213 ), .Z(\b/n6141 ) );
  NAND \b/U6235  ( .A(msg[105]), .B(\b/n5810 ), .Z(\b/n5862 ) );
  NAND \b/U6234  ( .A(\b/n156 ), .B(\b/n213 ), .Z(\b/n6139 ) );
  NAND \b/U6231  ( .A(msg[105]), .B(\b/n5805 ), .Z(\b/n5964 ) );
  ANDN \b/U6229  ( .A(msg[106]), .B(msg[105]), .Z(\b/n5992 ) );
  AND \b/U6228  ( .A(\b/n5802 ), .B(\b/n6136 ), .Z(\b/n5907 ) );
  MUX \b/U6227  ( .IN0(\b/n6135 ), .IN1(\b/n6119 ), .SEL(msg[110]), .F(
        shift_row_out[79]) );
  MUX \b/U6226  ( .IN0(\b/n6134 ), .IN1(\b/n6127 ), .SEL(msg[104]), .F(
        \b/n6135 ) );
  MUX \b/U6225  ( .IN0(\b/n6133 ), .IN1(\b/n6130 ), .SEL(msg[109]), .F(
        \b/n6134 ) );
  MUX \b/U6224  ( .IN0(\b/n6132 ), .IN1(\b/n6131 ), .SEL(msg[106]), .F(
        \b/n6133 ) );
  MUX \b/U6223  ( .IN0(msg[108]), .IN1(\b/n173 ), .SEL(msg[111]), .F(\b/n6132 ) );
  MUX \b/U6222  ( .IN0(\b/n5803 ), .IN1(\b/n177 ), .SEL(msg[111]), .F(
        \b/n6131 ) );
  MUX \b/U6221  ( .IN0(\b/n6129 ), .IN1(\b/n6128 ), .SEL(msg[106]), .F(
        \b/n6130 ) );
  MUX \b/U6220  ( .IN0(\b/n5861 ), .IN1(\b/n169 ), .SEL(msg[111]), .F(
        \b/n6129 ) );
  MUX \b/U6219  ( .IN0(\b/n5813 ), .IN1(\b/n5824 ), .SEL(msg[111]), .F(
        \b/n6128 ) );
  MUX \b/U6218  ( .IN0(\b/n6126 ), .IN1(\b/n6123 ), .SEL(msg[109]), .F(
        \b/n6127 ) );
  MUX \b/U6217  ( .IN0(\b/n6125 ), .IN1(\b/n6124 ), .SEL(msg[106]), .F(
        \b/n6126 ) );
  MUX \b/U6216  ( .IN0(\b/n5837 ), .IN1(\b/n5812 ), .SEL(msg[111]), .F(
        \b/n6125 ) );
  MUX \b/U6215  ( .IN0(\b/n181 ), .IN1(\b/n5833 ), .SEL(msg[111]), .F(
        \b/n6124 ) );
  MUX \b/U6214  ( .IN0(\b/n6121 ), .IN1(\b/n6120 ), .SEL(msg[106]), .F(
        \b/n6123 ) );
  AND \b/U6213  ( .A(\b/n171 ), .B(\b/n6122 ), .Z(\b/n6121 ) );
  MUX \b/U6212  ( .IN0(\b/n5817 ), .IN1(n711), .SEL(msg[111]), .F(\b/n6120 )
         );
  MUX \b/U6211  ( .IN0(\b/n6118 ), .IN1(\b/n6110 ), .SEL(msg[104]), .F(
        \b/n6119 ) );
  MUX \b/U6210  ( .IN0(\b/n6117 ), .IN1(\b/n6113 ), .SEL(msg[109]), .F(
        \b/n6118 ) );
  MUX \b/U6209  ( .IN0(\b/n6114 ), .IN1(\b/n6115 ), .SEL(msg[106]), .F(
        \b/n6117 ) );
  NAND \b/U6208  ( .A(\b/n5931 ), .B(\b/n6116 ), .Z(\b/n6115 ) );
  MUX \b/U6207  ( .IN0(\b/n211 ), .IN1(\b/n203 ), .SEL(msg[111]), .F(\b/n6114 ) );
  MUX \b/U6206  ( .IN0(\b/n6112 ), .IN1(\b/n6111 ), .SEL(msg[106]), .F(
        \b/n6113 ) );
  MUX \b/U6205  ( .IN0(\b/n5807 ), .IN1(\b/n5801 ), .SEL(msg[111]), .F(
        \b/n6112 ) );
  MUX \b/U6204  ( .IN0(\b/n204 ), .IN1(\b/n5838 ), .SEL(msg[111]), .F(
        \b/n6111 ) );
  MUX \b/U6203  ( .IN0(\b/n6109 ), .IN1(\b/n6106 ), .SEL(msg[109]), .F(
        \b/n6110 ) );
  MUX \b/U6202  ( .IN0(\b/n6108 ), .IN1(\b/n6107 ), .SEL(msg[106]), .F(
        \b/n6109 ) );
  MUX \b/U6201  ( .IN0(\b/n5842 ), .IN1(\b/n5828 ), .SEL(msg[111]), .F(
        \b/n6108 ) );
  MUX \b/U6200  ( .IN0(\b/n157 ), .IN1(\b/n5810 ), .SEL(msg[111]), .F(
        \b/n6107 ) );
  MUX \b/U6199  ( .IN0(\b/n6105 ), .IN1(\b/n6104 ), .SEL(msg[106]), .F(
        \b/n6106 ) );
  MUX \b/U6198  ( .IN0(\b/n5843 ), .IN1(\b/n5851 ), .SEL(msg[111]), .F(
        \b/n6105 ) );
  MUX \b/U6197  ( .IN0(\b/n5836 ), .IN1(\b/n6103 ), .SEL(msg[111]), .F(
        \b/n6104 ) );
  MUX \b/U6196  ( .IN0(\b/n208 ), .IN1(\b/n166 ), .SEL(msg[105]), .F(\b/n6103 ) );
  MUX \b/U6195  ( .IN0(\b/n6102 ), .IN1(\b/n6084 ), .SEL(msg[110]), .F(
        shift_row_out[78]) );
  MUX \b/U6194  ( .IN0(\b/n6101 ), .IN1(\b/n6092 ), .SEL(msg[104]), .F(
        \b/n6102 ) );
  MUX \b/U6193  ( .IN0(\b/n6100 ), .IN1(\b/n6095 ), .SEL(msg[109]), .F(
        \b/n6101 ) );
  MUX \b/U6192  ( .IN0(\b/n6099 ), .IN1(\b/n6097 ), .SEL(msg[106]), .F(
        \b/n6100 ) );
  MUX \b/U6191  ( .IN0(\b/n6098 ), .IN1(\b/n5814 ), .SEL(msg[111]), .F(
        \b/n6099 ) );
  MUX \b/U6190  ( .IN0(\b/n208 ), .IN1(\b/n5801 ), .SEL(msg[105]), .F(
        \b/n6098 ) );
  MUX \b/U6189  ( .IN0(\b/n6096 ), .IN1(\b/n196 ), .SEL(msg[111]), .F(
        \b/n6097 ) );
  MUX \b/U6188  ( .IN0(\b/n5801 ), .IN1(\b/n5802 ), .SEL(msg[105]), .F(
        \b/n6096 ) );
  MUX \b/U6187  ( .IN0(\b/n6094 ), .IN1(\b/n6093 ), .SEL(msg[106]), .F(
        \b/n6095 ) );
  MUX \b/U6186  ( .IN0(n710), .IN1(\b/n5882 ), .SEL(msg[111]), .F(\b/n6094 )
         );
  MUX \b/U6185  ( .IN0(\b/n5840 ), .IN1(\b/n5847 ), .SEL(msg[111]), .F(
        \b/n6093 ) );
  MUX \b/U6184  ( .IN0(\b/n6091 ), .IN1(\b/n6087 ), .SEL(msg[109]), .F(
        \b/n6092 ) );
  MUX \b/U6183  ( .IN0(\b/n6089 ), .IN1(\b/n6088 ), .SEL(msg[106]), .F(
        \b/n6091 ) );
  AND \b/U6182  ( .A(\b/n149 ), .B(\b/n6090 ), .Z(\b/n6089 ) );
  MUX \b/U6181  ( .IN0(\b/n5917 ), .IN1(msg[107]), .SEL(msg[111]), .F(
        \b/n6088 ) );
  MUX \b/U6180  ( .IN0(\b/n6086 ), .IN1(\b/n6085 ), .SEL(msg[106]), .F(
        \b/n6087 ) );
  MUX \b/U6179  ( .IN0(\b/n192 ), .IN1(\b/n5805 ), .SEL(msg[111]), .F(
        \b/n6086 ) );
  MUX \b/U6177  ( .IN0(\b/n6083 ), .IN1(\b/n6076 ), .SEL(msg[104]), .F(
        \b/n6084 ) );
  MUX \b/U6176  ( .IN0(\b/n6082 ), .IN1(\b/n6079 ), .SEL(msg[109]), .F(
        \b/n6083 ) );
  MUX \b/U6175  ( .IN0(\b/n6081 ), .IN1(\b/n6080 ), .SEL(msg[106]), .F(
        \b/n6082 ) );
  MUX \b/U6174  ( .IN0(\b/n188 ), .IN1(\b/n5809 ), .SEL(msg[111]), .F(
        \b/n6081 ) );
  MUX \b/U6173  ( .IN0(\b/n5813 ), .IN1(n711), .SEL(msg[111]), .F(\b/n6080 )
         );
  MUX \b/U6172  ( .IN0(\b/n6078 ), .IN1(\b/n6077 ), .SEL(msg[106]), .F(
        \b/n6079 ) );
  MUX \b/U6171  ( .IN0(\b/n5829 ), .IN1(\b/n153 ), .SEL(msg[111]), .F(
        \b/n6078 ) );
  MUX \b/U6170  ( .IN0(\b/n173 ), .IN1(\b/n203 ), .SEL(msg[111]), .F(\b/n6077 ) );
  MUX \b/U6169  ( .IN0(\b/n6075 ), .IN1(\b/n6071 ), .SEL(msg[109]), .F(
        \b/n6076 ) );
  MUX \b/U6168  ( .IN0(\b/n6074 ), .IN1(\b/n6073 ), .SEL(msg[106]), .F(
        \b/n6075 ) );
  MUX \b/U6167  ( .IN0(\b/n5818 ), .IN1(\b/n203 ), .SEL(msg[111]), .F(
        \b/n6074 ) );
  MUX \b/U6166  ( .IN0(\b/n6072 ), .IN1(\b/n5839 ), .SEL(msg[111]), .F(
        \b/n6073 ) );
  NANDN \b/U6165  ( .B(msg[108]), .A(msg[105]), .Z(\b/n6072 ) );
  MUX \b/U6164  ( .IN0(\b/n6070 ), .IN1(\b/n6068 ), .SEL(msg[106]), .F(
        \b/n6071 ) );
  MUX \b/U6163  ( .IN0(\b/n166 ), .IN1(\b/n6069 ), .SEL(msg[111]), .F(
        \b/n6070 ) );
  MUX \b/U6162  ( .IN0(\b/n193 ), .IN1(\b/n183 ), .SEL(msg[105]), .F(\b/n6069 ) );
  MUX \b/U6161  ( .IN0(\b/n155 ), .IN1(\b/n5814 ), .SEL(msg[111]), .F(
        \b/n6068 ) );
  NANDN \b/U6160  ( .B(\b/n156 ), .A(msg[105]), .Z(\b/n5814 ) );
  MUX \b/U6159  ( .IN0(\b/n6067 ), .IN1(\b/n6046 ), .SEL(msg[110]), .F(
        shift_row_out[77]) );
  MUX \b/U6158  ( .IN0(\b/n6066 ), .IN1(\b/n6056 ), .SEL(msg[104]), .F(
        \b/n6067 ) );
  MUX \b/U6157  ( .IN0(\b/n6065 ), .IN1(\b/n6061 ), .SEL(msg[109]), .F(
        \b/n6066 ) );
  MUX \b/U6156  ( .IN0(\b/n6062 ), .IN1(\b/n6063 ), .SEL(msg[106]), .F(
        \b/n6065 ) );
  AND \b/U6155  ( .A(\b/n5832 ), .B(\b/n6064 ), .Z(\b/n6063 ) );
  MUX \b/U6154  ( .IN0(\b/n5810 ), .IN1(\b/n204 ), .SEL(msg[111]), .F(
        \b/n6062 ) );
  MUX \b/U6153  ( .IN0(\b/n6060 ), .IN1(\b/n6058 ), .SEL(msg[106]), .F(
        \b/n6061 ) );
  MUX \b/U6152  ( .IN0(\b/n159 ), .IN1(\b/n6059 ), .SEL(msg[111]), .F(
        \b/n6060 ) );
  NAND \b/U6151  ( .A(\b/n183 ), .B(\b/n213 ), .Z(\b/n6059 ) );
  MUX \b/U6150  ( .IN0(\b/n5810 ), .IN1(\b/n6057 ), .SEL(msg[111]), .F(
        \b/n6058 ) );
  NAND \b/U6149  ( .A(\b/n5801 ), .B(\b/n5862 ), .Z(\b/n6057 ) );
  MUX \b/U6148  ( .IN0(\b/n6055 ), .IN1(\b/n6051 ), .SEL(msg[109]), .F(
        \b/n6056 ) );
  MUX \b/U6147  ( .IN0(\b/n6054 ), .IN1(\b/n6053 ), .SEL(msg[106]), .F(
        \b/n6055 ) );
  MUX \b/U6146  ( .IN0(\b/n5822 ), .IN1(\b/n206 ), .SEL(msg[111]), .F(
        \b/n6054 ) );
  MUX \b/U6145  ( .IN0(\b/n5847 ), .IN1(\b/n6052 ), .SEL(msg[111]), .F(
        \b/n6053 ) );
  MUX \b/U6144  ( .IN0(\b/n202 ), .IN1(\b/n183 ), .SEL(msg[105]), .F(\b/n6052 ) );
  MUX \b/U6143  ( .IN0(\b/n6050 ), .IN1(\b/n6049 ), .SEL(msg[106]), .F(
        \b/n6051 ) );
  MUX \b/U6142  ( .IN0(\b/n200 ), .IN1(n709), .SEL(msg[111]), .F(\b/n6050 ) );
  MUX \b/U6141  ( .IN0(\b/n6048 ), .IN1(\b/n6047 ), .SEL(msg[111]), .F(
        \b/n6049 ) );
  AND \b/U6140  ( .A(\b/n5807 ), .B(\b/n5882 ), .Z(\b/n6048 ) );
  MUX \b/U6139  ( .IN0(\b/n172 ), .IN1(\b/n156 ), .SEL(msg[105]), .F(\b/n6047 ) );
  MUX \b/U6138  ( .IN0(\b/n6045 ), .IN1(\b/n6036 ), .SEL(msg[104]), .F(
        \b/n6046 ) );
  MUX \b/U6137  ( .IN0(\b/n6044 ), .IN1(\b/n6040 ), .SEL(msg[109]), .F(
        \b/n6045 ) );
  MUX \b/U6136  ( .IN0(\b/n6043 ), .IN1(\b/n6041 ), .SEL(msg[106]), .F(
        \b/n6044 ) );
  MUX \b/U6135  ( .IN0(\b/n5813 ), .IN1(\b/n6042 ), .SEL(msg[111]), .F(
        \b/n6043 ) );
  NAND \b/U6134  ( .A(msg[105]), .B(\b/n172 ), .Z(\b/n6042 ) );
  MUX \b/U6133  ( .IN0(\b/n156 ), .IN1(\b/n209 ), .SEL(msg[111]), .F(\b/n6041 ) );
  MUX \b/U6132  ( .IN0(\b/n6039 ), .IN1(\b/n6038 ), .SEL(msg[106]), .F(
        \b/n6040 ) );
  MUX \b/U6131  ( .IN0(\b/n5839 ), .IN1(\b/n174 ), .SEL(msg[111]), .F(
        \b/n6039 ) );
  MUX \b/U6130  ( .IN0(\b/n6037 ), .IN1(\b/n5802 ), .SEL(n708), .F(\b/n6038 )
         );
  AND \b/U6129  ( .A(msg[111]), .B(msg[107]), .Z(\b/n6037 ) );
  MUX \b/U6128  ( .IN0(\b/n6035 ), .IN1(\b/n6032 ), .SEL(msg[109]), .F(
        \b/n6036 ) );
  MUX \b/U6127  ( .IN0(\b/n6034 ), .IN1(\b/n6033 ), .SEL(msg[106]), .F(
        \b/n6035 ) );
  MUX \b/U6126  ( .IN0(\b/n5963 ), .IN1(\b/n5802 ), .SEL(msg[111]), .F(
        \b/n6034 ) );
  MUX \b/U6125  ( .IN0(n707), .IN1(\b/n207 ), .SEL(msg[111]), .F(\b/n6033 ) );
  MUX \b/U6124  ( .IN0(\b/n6030 ), .IN1(\b/n6029 ), .SEL(msg[106]), .F(
        \b/n6032 ) );
  AND \b/U6123  ( .A(\b/n6031 ), .B(\b/n5931 ), .Z(\b/n6030 ) );
  MUX \b/U6122  ( .IN0(\b/n158 ), .IN1(\b/n202 ), .SEL(msg[111]), .F(\b/n6029 ) );
  MUX \b/U6121  ( .IN0(\b/n6028 ), .IN1(\b/n6011 ), .SEL(msg[110]), .F(
        shift_row_out[76]) );
  MUX \b/U6120  ( .IN0(\b/n6027 ), .IN1(\b/n6019 ), .SEL(msg[104]), .F(
        \b/n6028 ) );
  MUX \b/U6119  ( .IN0(\b/n6026 ), .IN1(\b/n6023 ), .SEL(msg[109]), .F(
        \b/n6027 ) );
  MUX \b/U6118  ( .IN0(\b/n6025 ), .IN1(\b/n6024 ), .SEL(msg[106]), .F(
        \b/n6026 ) );
  MUX \b/U6117  ( .IN0(\b/n184 ), .IN1(\b/n205 ), .SEL(msg[111]), .F(\b/n6025 ) );
  MUX \b/U6116  ( .IN0(\b/n5882 ), .IN1(\b/n5847 ), .SEL(msg[111]), .F(
        \b/n6024 ) );
  NAND \b/U6115  ( .A(msg[105]), .B(\b/n5801 ), .Z(\b/n5882 ) );
  MUX \b/U6114  ( .IN0(\b/n6020 ), .IN1(\b/n6021 ), .SEL(msg[106]), .F(
        \b/n6023 ) );
  AND \b/U6113  ( .A(\b/n5832 ), .B(\b/n6022 ), .Z(\b/n6021 ) );
  MUX \b/U6112  ( .IN0(\b/n5830 ), .IN1(\b/n187 ), .SEL(msg[111]), .F(
        \b/n6020 ) );
  MUX \b/U6111  ( .IN0(\b/n6018 ), .IN1(\b/n6015 ), .SEL(msg[109]), .F(
        \b/n6019 ) );
  MUX \b/U6110  ( .IN0(\b/n6017 ), .IN1(\b/n6016 ), .SEL(msg[106]), .F(
        \b/n6018 ) );
  MUX \b/U6109  ( .IN0(\b/n149 ), .IN1(\b/n195 ), .SEL(msg[111]), .F(\b/n6017 ) );
  MUX \b/U6108  ( .IN0(\b/n156 ), .IN1(\b/n5810 ), .SEL(msg[111]), .F(
        \b/n6016 ) );
  MUX \b/U6107  ( .IN0(\b/n6014 ), .IN1(\b/n6012 ), .SEL(msg[106]), .F(
        \b/n6015 ) );
  MUX \b/U6106  ( .IN0(\b/n5826 ), .IN1(\b/n6013 ), .SEL(msg[111]), .F(
        \b/n6014 ) );
  AND \b/U6105  ( .A(\b/n5810 ), .B(\b/n213 ), .Z(\b/n6013 ) );
  MUX \b/U6104  ( .IN0(\b/n171 ), .IN1(\b/n190 ), .SEL(msg[111]), .F(\b/n6012 ) );
  MUX \b/U6103  ( .IN0(\b/n6010 ), .IN1(\b/n6004 ), .SEL(msg[104]), .F(
        \b/n6011 ) );
  MUX \b/U6102  ( .IN0(\b/n6009 ), .IN1(\b/n6007 ), .SEL(msg[109]), .F(
        \b/n6010 ) );
  MUX \b/U6101  ( .IN0(\b/n6008 ), .IN1(\b/n5804 ), .SEL(msg[106]), .F(
        \b/n6009 ) );
  MUX \b/U6100  ( .IN0(\b/n5824 ), .IN1(\b/n192 ), .SEL(msg[111]), .F(
        \b/n6008 ) );
  MUX \b/U6099  ( .IN0(\b/n6006 ), .IN1(\b/n6005 ), .SEL(msg[106]), .F(
        \b/n6007 ) );
  MUX \b/U6098  ( .IN0(n706), .IN1(\b/n184 ), .SEL(msg[111]), .F(\b/n6006 ) );
  MUX \b/U6097  ( .IN0(\b/n5834 ), .IN1(\b/n5837 ), .SEL(msg[111]), .F(
        \b/n6005 ) );
  MUX \b/U6096  ( .IN0(\b/n6003 ), .IN1(\b/n6000 ), .SEL(msg[109]), .F(
        \b/n6004 ) );
  MUX \b/U6095  ( .IN0(\b/n6002 ), .IN1(\b/n6001 ), .SEL(msg[106]), .F(
        \b/n6003 ) );
  MUX \b/U6094  ( .IN0(\b/n157 ), .IN1(\b/n5806 ), .SEL(msg[111]), .F(
        \b/n6002 ) );
  MUX \b/U6093  ( .IN0(\b/n202 ), .IN1(\b/n5828 ), .SEL(msg[111]), .F(
        \b/n6001 ) );
  MUX \b/U6092  ( .IN0(\b/n145 ), .IN1(\b/n5999 ), .SEL(msg[106]), .F(
        \b/n6000 ) );
  MUX \b/U6091  ( .IN0(\b/n165 ), .IN1(\b/n5810 ), .SEL(msg[111]), .F(
        \b/n5999 ) );
  MUX \b/U6090  ( .IN0(\b/n5998 ), .IN1(\b/n5979 ), .SEL(msg[110]), .F(
        shift_row_out[75]) );
  MUX \b/U6089  ( .IN0(\b/n5997 ), .IN1(\b/n5989 ), .SEL(msg[104]), .F(
        \b/n5998 ) );
  MUX \b/U6088  ( .IN0(\b/n5996 ), .IN1(\b/n5993 ), .SEL(msg[109]), .F(
        \b/n5997 ) );
  MUX \b/U6087  ( .IN0(\b/n5995 ), .IN1(\b/n5994 ), .SEL(msg[111]), .F(
        \b/n5996 ) );
  MUX \b/U6086  ( .IN0(\b/n5818 ), .IN1(\b/n190 ), .SEL(msg[106]), .F(
        \b/n5995 ) );
  MUX \b/U6085  ( .IN0(n709), .IN1(\b/n148 ), .SEL(msg[106]), .F(\b/n5994 ) );
  MUX \b/U6084  ( .IN0(\b/n5991 ), .IN1(\b/n5990 ), .SEL(msg[111]), .F(
        \b/n5993 ) );
  AND \b/U6083  ( .A(\b/n5992 ), .B(msg[108]), .Z(\b/n5991 ) );
  MUX \b/U6082  ( .IN0(\b/n178 ), .IN1(\b/n5831 ), .SEL(msg[106]), .F(
        \b/n5990 ) );
  MUX \b/U6081  ( .IN0(\b/n5988 ), .IN1(\b/n5985 ), .SEL(msg[109]), .F(
        \b/n5989 ) );
  MUX \b/U6080  ( .IN0(\b/n5987 ), .IN1(\b/n5986 ), .SEL(msg[111]), .F(
        \b/n5988 ) );
  MUX \b/U6079  ( .IN0(\b/n5822 ), .IN1(n705), .SEL(msg[106]), .F(\b/n5987 )
         );
  MUX \b/U6078  ( .IN0(\b/n146 ), .IN1(\b/n165 ), .SEL(msg[106]), .F(\b/n5986 ) );
  MUX \b/U6077  ( .IN0(\b/n5981 ), .IN1(\b/n5982 ), .SEL(msg[111]), .F(
        \b/n5985 ) );
  NAND \b/U6076  ( .A(\b/n5983 ), .B(\b/n5984 ), .Z(\b/n5982 ) );
  MUX \b/U6075  ( .IN0(\b/n191 ), .IN1(\b/n5980 ), .SEL(msg[106]), .F(
        \b/n5981 ) );
  MUX \b/U6074  ( .IN0(\b/n166 ), .IN1(\b/n208 ), .SEL(msg[105]), .F(\b/n5980 ) );
  MUX \b/U6073  ( .IN0(\b/n5978 ), .IN1(\b/n5969 ), .SEL(msg[104]), .F(
        \b/n5979 ) );
  MUX \b/U6072  ( .IN0(\b/n5977 ), .IN1(\b/n5973 ), .SEL(msg[109]), .F(
        \b/n5978 ) );
  MUX \b/U6071  ( .IN0(\b/n5975 ), .IN1(\b/n5974 ), .SEL(msg[111]), .F(
        \b/n5977 ) );
  NAND \b/U6070  ( .A(\b/n156 ), .B(\b/n5976 ), .Z(\b/n5975 ) );
  MUX \b/U6069  ( .IN0(\b/n207 ), .IN1(\b/n169 ), .SEL(msg[106]), .F(\b/n5974 ) );
  MUX \b/U6068  ( .IN0(\b/n5972 ), .IN1(\b/n5970 ), .SEL(msg[111]), .F(
        \b/n5973 ) );
  MUX \b/U6067  ( .IN0(\b/n5813 ), .IN1(\b/n5971 ), .SEL(msg[106]), .F(
        \b/n5972 ) );
  AND \b/U6066  ( .A(msg[105]), .B(\b/n156 ), .Z(\b/n5971 ) );
  MUX \b/U6065  ( .IN0(\b/n161 ), .IN1(\b/n5832 ), .SEL(msg[106]), .F(
        \b/n5970 ) );
  MUX \b/U6064  ( .IN0(\b/n5968 ), .IN1(\b/n5962 ), .SEL(msg[109]), .F(
        \b/n5969 ) );
  MUX \b/U6063  ( .IN0(\b/n5967 ), .IN1(\b/n5965 ), .SEL(msg[111]), .F(
        \b/n5968 ) );
  MUX \b/U6062  ( .IN0(\b/n5966 ), .IN1(\b/n5802 ), .SEL(\b/n5850 ), .F(
        \b/n5967 ) );
  MUX \b/U6061  ( .IN0(msg[107]), .IN1(msg[108]), .SEL(msg[106]), .F(\b/n5966 ) );
  MUX \b/U6060  ( .IN0(\b/n5832 ), .IN1(\b/n5963 ), .SEL(msg[106]), .F(
        \b/n5965 ) );
  NAND \b/U6059  ( .A(\b/n5802 ), .B(\b/n5964 ), .Z(\b/n5963 ) );
  MUX \b/U6058  ( .IN0(\b/n5959 ), .IN1(\b/n5960 ), .SEL(msg[111]), .F(
        \b/n5962 ) );
  AND \b/U6057  ( .A(\b/n189 ), .B(\b/n5961 ), .Z(\b/n5960 ) );
  MUX \b/U6056  ( .IN0(\b/n170 ), .IN1(\b/n5803 ), .SEL(msg[106]), .F(
        \b/n5959 ) );
  MUX \b/U6055  ( .IN0(\b/n5958 ), .IN1(\b/n5942 ), .SEL(msg[110]), .F(
        shift_row_out[74]) );
  MUX \b/U6054  ( .IN0(\b/n5957 ), .IN1(\b/n5949 ), .SEL(msg[104]), .F(
        \b/n5958 ) );
  MUX \b/U6053  ( .IN0(\b/n5956 ), .IN1(\b/n5952 ), .SEL(msg[109]), .F(
        \b/n5957 ) );
  MUX \b/U6052  ( .IN0(\b/n5955 ), .IN1(\b/n5953 ), .SEL(msg[106]), .F(
        \b/n5956 ) );
  MUX \b/U6051  ( .IN0(\b/n178 ), .IN1(\b/n5954 ), .SEL(msg[111]), .F(
        \b/n5955 ) );
  MUX \b/U6050  ( .IN0(\b/n5810 ), .IN1(\b/n156 ), .SEL(msg[105]), .F(
        \b/n5954 ) );
  MUX \b/U6049  ( .IN0(\b/n5849 ), .IN1(\b/n196 ), .SEL(msg[111]), .F(
        \b/n5953 ) );
  MUX \b/U6048  ( .IN0(\b/n5951 ), .IN1(\b/n5950 ), .SEL(msg[106]), .F(
        \b/n5952 ) );
  MUX \b/U6047  ( .IN0(\b/n5803 ), .IN1(\b/n163 ), .SEL(msg[111]), .F(
        \b/n5951 ) );
  MUX \b/U6046  ( .IN0(\b/n199 ), .IN1(\b/n5836 ), .SEL(msg[111]), .F(
        \b/n5950 ) );
  MUX \b/U6045  ( .IN0(\b/n5948 ), .IN1(\b/n5944 ), .SEL(msg[109]), .F(
        \b/n5949 ) );
  MUX \b/U6044  ( .IN0(\b/n5945 ), .IN1(\b/n145 ), .SEL(msg[106]), .F(
        \b/n5948 ) );
  NAND \b/U6043  ( .A(\b/n5946 ), .B(\b/n5947 ), .Z(\b/n5945 ) );
  MUX \b/U6042  ( .IN0(n707), .IN1(\b/n5943 ), .SEL(\b/n5848 ), .F(\b/n5944 )
         );
  MUX \b/U6041  ( .IN0(\b/n177 ), .IN1(\b/n5815 ), .SEL(msg[106]), .F(
        \b/n5943 ) );
  MUX \b/U6040  ( .IN0(\b/n5941 ), .IN1(\b/n5933 ), .SEL(msg[104]), .F(
        \b/n5942 ) );
  MUX \b/U6039  ( .IN0(\b/n5940 ), .IN1(\b/n5937 ), .SEL(msg[109]), .F(
        \b/n5941 ) );
  MUX \b/U6038  ( .IN0(\b/n5939 ), .IN1(\b/n5938 ), .SEL(msg[106]), .F(
        \b/n5940 ) );
  MUX \b/U6037  ( .IN0(\b/n205 ), .IN1(msg[105]), .SEL(msg[111]), .F(\b/n5939 ) );
  MUX \b/U6036  ( .IN0(n710), .IN1(\b/n5816 ), .SEL(msg[111]), .F(\b/n5938 )
         );
  MUX \b/U6035  ( .IN0(\b/n5936 ), .IN1(\b/n5935 ), .SEL(msg[106]), .F(
        \b/n5937 ) );
  MUX \b/U6034  ( .IN0(\b/n210 ), .IN1(\b/n204 ), .SEL(msg[111]), .F(\b/n5936 ) );
  MUX \b/U6033  ( .IN0(n710), .IN1(\b/n5934 ), .SEL(msg[111]), .F(\b/n5935 )
         );
  MUX \b/U6032  ( .IN0(\b/n156 ), .IN1(\b/n193 ), .SEL(msg[105]), .F(\b/n5934 ) );
  MUX \b/U6031  ( .IN0(\b/n5932 ), .IN1(\b/n5926 ), .SEL(msg[109]), .F(
        \b/n5933 ) );
  MUX \b/U6030  ( .IN0(\b/n5929 ), .IN1(\b/n5928 ), .SEL(msg[106]), .F(
        \b/n5932 ) );
  NAND \b/U6029  ( .A(\b/n5930 ), .B(\b/n5931 ), .Z(\b/n5929 ) );
  MUX \b/U6028  ( .IN0(\b/n5802 ), .IN1(\b/n5927 ), .SEL(n708), .F(\b/n5928 )
         );
  MUX \b/U6027  ( .IN0(msg[107]), .IN1(\b/n166 ), .SEL(msg[111]), .F(\b/n5927 ) );
  MUX \b/U6026  ( .IN0(\b/n5925 ), .IN1(\b/n5924 ), .SEL(msg[106]), .F(
        \b/n5926 ) );
  MUX \b/U6025  ( .IN0(\b/n5847 ), .IN1(\b/n164 ), .SEL(msg[111]), .F(
        \b/n5925 ) );
  MUX \b/U6024  ( .IN0(\b/n5843 ), .IN1(\b/n5923 ), .SEL(msg[111]), .F(
        \b/n5924 ) );
  MUX \b/U6023  ( .IN0(\b/n5805 ), .IN1(\b/n5810 ), .SEL(msg[105]), .F(
        \b/n5923 ) );
  MUX \b/U6022  ( .IN0(\b/n5922 ), .IN1(\b/n5904 ), .SEL(msg[110]), .F(
        shift_row_out[73]) );
  MUX \b/U6021  ( .IN0(\b/n5921 ), .IN1(\b/n5912 ), .SEL(msg[104]), .F(
        \b/n5922 ) );
  MUX \b/U6020  ( .IN0(\b/n5920 ), .IN1(\b/n5916 ), .SEL(msg[109]), .F(
        \b/n5921 ) );
  MUX \b/U6019  ( .IN0(\b/n5919 ), .IN1(\b/n5918 ), .SEL(msg[106]), .F(
        \b/n5920 ) );
  MUX \b/U6018  ( .IN0(\b/n201 ), .IN1(n712), .SEL(msg[111]), .F(\b/n5919 ) );
  MUX \b/U6017  ( .IN0(\b/n5917 ), .IN1(n706), .SEL(msg[111]), .F(\b/n5918 )
         );
  NAND \b/U6016  ( .A(\b/n213 ), .B(\b/n172 ), .Z(\b/n5917 ) );
  MUX \b/U6015  ( .IN0(\b/n5915 ), .IN1(\b/n5914 ), .SEL(msg[106]), .F(
        \b/n5916 ) );
  MUX \b/U6014  ( .IN0(\b/n149 ), .IN1(\b/n5817 ), .SEL(msg[111]), .F(
        \b/n5915 ) );
  MUX \b/U6013  ( .IN0(\b/n5807 ), .IN1(\b/n5913 ), .SEL(msg[111]), .F(
        \b/n5914 ) );
  AND \b/U6012  ( .A(msg[105]), .B(msg[108]), .Z(\b/n5913 ) );
  MUX \b/U6011  ( .IN0(\b/n5911 ), .IN1(\b/n5908 ), .SEL(msg[109]), .F(
        \b/n5912 ) );
  MUX \b/U6010  ( .IN0(\b/n5910 ), .IN1(\b/n5909 ), .SEL(msg[106]), .F(
        \b/n5911 ) );
  MUX \b/U6009  ( .IN0(\b/n5846 ), .IN1(\b/n210 ), .SEL(msg[111]), .F(
        \b/n5910 ) );
  MUX \b/U6008  ( .IN0(\b/n185 ), .IN1(\b/n5815 ), .SEL(msg[111]), .F(
        \b/n5909 ) );
  MUX \b/U6007  ( .IN0(\b/n5905 ), .IN1(\b/n5906 ), .SEL(msg[106]), .F(
        \b/n5908 ) );
  AND \b/U6006  ( .A(\b/n5907 ), .B(\b/n5862 ), .Z(\b/n5906 ) );
  MUX \b/U6005  ( .IN0(\b/n5821 ), .IN1(\b/n5810 ), .SEL(msg[111]), .F(
        \b/n5905 ) );
  MUX \b/U6004  ( .IN0(\b/n5903 ), .IN1(\b/n5895 ), .SEL(msg[104]), .F(
        \b/n5904 ) );
  MUX \b/U6003  ( .IN0(\b/n5902 ), .IN1(\b/n5898 ), .SEL(msg[109]), .F(
        \b/n5903 ) );
  MUX \b/U6002  ( .IN0(\b/n5901 ), .IN1(\b/n5900 ), .SEL(msg[106]), .F(
        \b/n5902 ) );
  MUX \b/U6001  ( .IN0(\b/n5809 ), .IN1(\b/n174 ), .SEL(msg[111]), .F(
        \b/n5901 ) );
  MUX \b/U6000  ( .IN0(\b/n5899 ), .IN1(\b/n158 ), .SEL(msg[111]), .F(
        \b/n5900 ) );
  MUX \b/U5999  ( .IN0(\b/n5807 ), .IN1(\b/n166 ), .SEL(msg[105]), .F(
        \b/n5899 ) );
  MUX \b/U5998  ( .IN0(\b/n5897 ), .IN1(\b/n5896 ), .SEL(msg[106]), .F(
        \b/n5898 ) );
  MUX \b/U5997  ( .IN0(\b/n205 ), .IN1(\b/n183 ), .SEL(msg[111]), .F(\b/n5897 ) );
  MUX \b/U5996  ( .IN0(\b/n201 ), .IN1(\b/n161 ), .SEL(msg[111]), .F(\b/n5896 ) );
  MUX \b/U5995  ( .IN0(\b/n5894 ), .IN1(\b/n5889 ), .SEL(msg[109]), .F(
        \b/n5895 ) );
  MUX \b/U5994  ( .IN0(\b/n5893 ), .IN1(\b/n5890 ), .SEL(msg[106]), .F(
        \b/n5894 ) );
  MUX \b/U5993  ( .IN0(\b/n5891 ), .IN1(\b/n5892 ), .SEL(msg[111]), .F(
        \b/n5893 ) );
  NAND \b/U5992  ( .A(\b/n5810 ), .B(\b/n5882 ), .Z(\b/n5892 ) );
  MUX \b/U5991  ( .IN0(\b/n5810 ), .IN1(\b/n166 ), .SEL(msg[105]), .F(
        \b/n5891 ) );
  MUX \b/U5990  ( .IN0(\b/n5827 ), .IN1(\b/n5825 ), .SEL(msg[111]), .F(
        \b/n5890 ) );
  MUX \b/U5989  ( .IN0(\b/n5845 ), .IN1(\b/n5888 ), .SEL(msg[106]), .F(
        \b/n5889 ) );
  MUX \b/U5988  ( .IN0(\b/n172 ), .IN1(\b/n204 ), .SEL(msg[111]), .F(\b/n5888 ) );
  MUX \b/U5987  ( .IN0(\b/n5887 ), .IN1(\b/n5870 ), .SEL(msg[110]), .F(
        shift_row_out[72]) );
  MUX \b/U5986  ( .IN0(\b/n5886 ), .IN1(\b/n5878 ), .SEL(msg[104]), .F(
        \b/n5887 ) );
  MUX \b/U5985  ( .IN0(\b/n5885 ), .IN1(\b/n5883 ), .SEL(msg[106]), .F(
        \b/n5886 ) );
  MUX \b/U5984  ( .IN0(\b/n146 ), .IN1(\b/n5884 ), .SEL(msg[111]), .F(
        \b/n5885 ) );
  MUX \b/U5983  ( .IN0(\b/n199 ), .IN1(\b/n202 ), .SEL(msg[109]), .F(\b/n5884 ) );
  MUX \b/U5982  ( .IN0(\b/n5880 ), .IN1(\b/n5879 ), .SEL(msg[111]), .F(
        \b/n5883 ) );
  NAND \b/U5981  ( .A(\b/n5881 ), .B(\b/n5882 ), .Z(\b/n5880 ) );
  MUX \b/U5980  ( .IN0(\b/n198 ), .IN1(\b/n213 ), .SEL(msg[109]), .F(\b/n5879 ) );
  MUX \b/U5979  ( .IN0(\b/n5877 ), .IN1(\b/n5873 ), .SEL(msg[106]), .F(
        \b/n5878 ) );
  MUX \b/U5978  ( .IN0(\b/n5876 ), .IN1(\b/n5874 ), .SEL(msg[111]), .F(
        \b/n5877 ) );
  MUX \b/U5977  ( .IN0(\b/n5875 ), .IN1(\b/n151 ), .SEL(msg[109]), .F(
        \b/n5876 ) );
  NAND \b/U5976  ( .A(\b/n213 ), .B(\b/n5802 ), .Z(\b/n5875 ) );
  MUX \b/U5974  ( .IN0(\b/n5872 ), .IN1(\b/n5871 ), .SEL(msg[111]), .F(
        \b/n5873 ) );
  MUX \b/U5973  ( .IN0(n707), .IN1(\b/n148 ), .SEL(msg[109]), .F(\b/n5872 ) );
  MUX \b/U5972  ( .IN0(\b/n200 ), .IN1(\b/n156 ), .SEL(msg[109]), .F(\b/n5871 ) );
  MUX \b/U5971  ( .IN0(\b/n5869 ), .IN1(\b/n5859 ), .SEL(msg[104]), .F(
        \b/n5870 ) );
  MUX \b/U5970  ( .IN0(\b/n5868 ), .IN1(\b/n5864 ), .SEL(msg[106]), .F(
        \b/n5869 ) );
  MUX \b/U5969  ( .IN0(\b/n5867 ), .IN1(\b/n5866 ), .SEL(msg[111]), .F(
        \b/n5868 ) );
  MUX \b/U5968  ( .IN0(n705), .IN1(\b/n152 ), .SEL(msg[109]), .F(\b/n5867 ) );
  MUX \b/U5967  ( .IN0(\b/n5865 ), .IN1(\b/n189 ), .SEL(msg[109]), .F(
        \b/n5866 ) );
  NAND \b/U5966  ( .A(\b/n5801 ), .B(\b/n5803 ), .Z(\b/n5865 ) );
  MUX \b/U5965  ( .IN0(\b/n5863 ), .IN1(\b/n5860 ), .SEL(msg[111]), .F(
        \b/n5864 ) );
  MUX \b/U5964  ( .IN0(\b/n159 ), .IN1(\b/n5861 ), .SEL(msg[109]), .F(
        \b/n5863 ) );
  NAND \b/U5963  ( .A(\b/n5805 ), .B(\b/n5862 ), .Z(\b/n5861 ) );
  MUX \b/U5962  ( .IN0(\b/n5820 ), .IN1(\b/n5811 ), .SEL(msg[109]), .F(
        \b/n5860 ) );
  MUX \b/U5961  ( .IN0(\b/n5858 ), .IN1(\b/n5854 ), .SEL(msg[106]), .F(
        \b/n5859 ) );
  MUX \b/U5960  ( .IN0(\b/n5856 ), .IN1(\b/n5855 ), .SEL(msg[111]), .F(
        \b/n5858 ) );
  NAND \b/U5959  ( .A(\b/n5857 ), .B(\b/n5844 ), .Z(\b/n5856 ) );
  MUX \b/U5958  ( .IN0(msg[107]), .IN1(\b/n5836 ), .SEL(msg[109]), .F(
        \b/n5855 ) );
  MUX \b/U5957  ( .IN0(\b/n5853 ), .IN1(\b/n5852 ), .SEL(msg[111]), .F(
        \b/n5854 ) );
  MUX \b/U5956  ( .IN0(\b/n164 ), .IN1(\b/n180 ), .SEL(msg[109]), .F(\b/n5853 ) );
  MUX \b/U5955  ( .IN0(\b/n197 ), .IN1(\b/n185 ), .SEL(msg[109]), .F(\b/n5852 ) );
  XOR \b/U5954  ( .A(\b/n5802 ), .B(msg[105]), .Z(\b/n5851 ) );
  XOR \b/U5953  ( .A(msg[105]), .B(msg[106]), .Z(\b/n5850 ) );
  XOR \b/U5952  ( .A(msg[105]), .B(msg[107]), .Z(\b/n5849 ) );
  XOR \b/U5951  ( .A(msg[106]), .B(msg[111]), .Z(\b/n5848 ) );
  XOR \b/U5950  ( .A(\b/n213 ), .B(\b/n156 ), .Z(\b/n5847 ) );
  XOR \b/U5949  ( .A(msg[105]), .B(\b/n202 ), .Z(\b/n5846 ) );
  XOR \b/U5947  ( .A(msg[105]), .B(msg[109]), .Z(\b/n5844 ) );
  NAND \b/U5946  ( .A(msg[105]), .B(msg[107]), .Z(\b/n5843 ) );
  MUX \b/U5945  ( .IN0(\b/n5802 ), .IN1(\b/n156 ), .SEL(msg[105]), .F(
        \b/n5842 ) );
  MUX \b/U5943  ( .IN0(msg[107]), .IN1(\b/n193 ), .SEL(msg[105]), .F(\b/n5840 ) );
  MUX \b/U5942  ( .IN0(\b/n172 ), .IN1(\b/n193 ), .SEL(msg[105]), .F(\b/n5839 ) );
  MUX \b/U5941  ( .IN0(\b/n5805 ), .IN1(\b/n5807 ), .SEL(msg[105]), .F(
        \b/n5838 ) );
  MUX \b/U5940  ( .IN0(msg[108]), .IN1(\b/n172 ), .SEL(msg[105]), .F(\b/n5837 ) );
  OR \b/U5939  ( .A(msg[105]), .B(msg[108]), .Z(\b/n5836 ) );
  NAND \b/U5937  ( .A(\b/n193 ), .B(\b/n213 ), .Z(\b/n5834 ) );
  MUX \b/U5936  ( .IN0(\b/n193 ), .IN1(msg[108]), .SEL(msg[105]), .F(\b/n5833 ) );
  MUX \b/U5935  ( .IN0(\b/n5801 ), .IN1(\b/n5810 ), .SEL(msg[105]), .F(
        \b/n5832 ) );
  MUX \b/U5934  ( .IN0(\b/n208 ), .IN1(msg[108]), .SEL(msg[105]), .F(\b/n5831 ) );
  MUX \b/U5933  ( .IN0(\b/n166 ), .IN1(\b/n193 ), .SEL(msg[105]), .F(\b/n5830 ) );
  MUX \b/U5932  ( .IN0(\b/n5801 ), .IN1(msg[108]), .SEL(msg[105]), .F(
        \b/n5829 ) );
  MUX \b/U5931  ( .IN0(\b/n183 ), .IN1(\b/n172 ), .SEL(msg[105]), .F(\b/n5828 ) );
  XOR \b/U5930  ( .A(\b/n166 ), .B(msg[105]), .Z(\b/n5827 ) );
  MUX \b/U5929  ( .IN0(\b/n5807 ), .IN1(\b/n183 ), .SEL(msg[105]), .F(
        \b/n5826 ) );
  NANDN \b/U5928  ( .B(msg[105]), .A(msg[107]), .Z(\b/n5825 ) );
  MUX \b/U5927  ( .IN0(\b/n156 ), .IN1(msg[107]), .SEL(msg[105]), .F(\b/n5824 ) );
  NAND \b/U5925  ( .A(\b/n5805 ), .B(\b/n213 ), .Z(\b/n5822 ) );
  MUX \b/U5924  ( .IN0(msg[108]), .IN1(\b/n5802 ), .SEL(msg[105]), .F(
        \b/n5821 ) );
  MUX \b/U5923  ( .IN0(\b/n183 ), .IN1(msg[107]), .SEL(msg[105]), .F(\b/n5820 ) );
  MUX \b/U5921  ( .IN0(msg[108]), .IN1(\b/n202 ), .SEL(msg[105]), .F(\b/n5818 ) );
  MUX \b/U5920  ( .IN0(\b/n156 ), .IN1(\b/n208 ), .SEL(msg[105]), .F(\b/n5817 ) );
  NAND \b/U5919  ( .A(\b/n5803 ), .B(\b/n156 ), .Z(\b/n5816 ) );
  MUX \b/U5918  ( .IN0(\b/n5802 ), .IN1(\b/n5810 ), .SEL(msg[105]), .F(
        \b/n5815 ) );
  NAND \b/U5917  ( .A(\b/n5814 ), .B(\b/n5801 ), .Z(\b/n5813 ) );
  MUX \b/U5916  ( .IN0(\b/n5805 ), .IN1(\b/n208 ), .SEL(msg[105]), .F(
        \b/n5812 ) );
  MUX \b/U5915  ( .IN0(\b/n208 ), .IN1(\b/n172 ), .SEL(msg[105]), .F(\b/n5811 ) );
  NANDN \b/U5914  ( .B(msg[107]), .A(msg[108]), .Z(\b/n5810 ) );
  MUX \b/U5913  ( .IN0(\b/n5805 ), .IN1(msg[107]), .SEL(msg[105]), .F(
        \b/n5809 ) );
  OR \b/U5912  ( .A(msg[107]), .B(msg[108]), .Z(\b/n5805 ) );
  MUX \b/U5911  ( .IN0(\b/n156 ), .IN1(\b/n172 ), .SEL(msg[105]), .F(\b/n5808 ) );
  XOR \b/U5910  ( .A(\b/n166 ), .B(msg[107]), .Z(\b/n5807 ) );
  NANDN \b/U5909  ( .B(msg[107]), .A(msg[105]), .Z(\b/n5806 ) );
  NAND \b/U5908  ( .A(\b/n5805 ), .B(\b/n5803 ), .Z(\b/n5804 ) );
  NAND \b/U5907  ( .A(msg[105]), .B(\b/n5802 ), .Z(\b/n5803 ) );
  NANDN \b/U5906  ( .B(msg[108]), .A(msg[107]), .Z(\b/n5802 ) );
  NAND \b/U5905  ( .A(msg[107]), .B(msg[108]), .Z(\b/n5801 ) );
  MUX \b/U5904  ( .IN0(msg[100]), .IN1(\b/n5443 ), .SEL(msg[97]), .F(\b/n5800 ) );
  MUX \b/U5903  ( .IN0(msg[100]), .IN1(\b/n5444 ), .SEL(msg[97]), .F(\b/n5799 ) );
  MUX \b/U5902  ( .IN0(\b/n5446 ), .IN1(\b/n5449 ), .SEL(msg[97]), .F(
        \b/n5798 ) );
  MUX \b/U5901  ( .IN0(\b/n5468 ), .IN1(\b/n240 ), .SEL(msg[97]), .F(\b/n5797 ) );
  MUX \b/U5899  ( .IN0(\b/n5444 ), .IN1(\b/n5443 ), .SEL(msg[98]), .F(
        \b/n5614 ) );
  MUX \b/U5898  ( .IN0(\b/n5445 ), .IN1(\b/n283 ), .SEL(msg[98]), .F(\b/n5615 ) );
  MUX \b/U5897  ( .IN0(\b/n275 ), .IN1(\b/n220 ), .SEL(msg[97]), .F(\b/n5580 )
         );
  MUX \b/U5896  ( .IN0(\b/n5475 ), .IN1(\b/n5783 ), .SEL(msg[103]), .F(
        \b/n5795 ) );
  MUX \b/U5895  ( .IN0(\b/n5449 ), .IN1(\b/n5443 ), .SEL(msg[97]), .F(
        \b/n5786 ) );
  MUX \b/U5894  ( .IN0(\b/n278 ), .IN1(\b/n5468 ), .SEL(msg[97]), .F(\b/n5794 ) );
  MUX \b/U5893  ( .IN0(msg[99]), .IN1(\b/n240 ), .SEL(msg[97]), .F(\b/n5793 )
         );
  MUX \b/U5892  ( .IN0(\b/n5444 ), .IN1(\b/n278 ), .SEL(msg[97]), .F(\b/n5792 ) );
  MUX \b/U5891  ( .IN0(msg[100]), .IN1(\b/n5468 ), .SEL(msg[97]), .F(\b/n5791 ) );
  MUX \b/U5890  ( .IN0(\b/n250 ), .IN1(\b/n227 ), .SEL(msg[101]), .F(\b/n5498 ) );
  MUX \b/U5889  ( .IN0(\b/n5446 ), .IN1(\b/n220 ), .SEL(msg[97]), .F(\b/n5790 ) );
  NANDN \b/U5886  ( .B(\b/n5451 ), .A(msg[103]), .Z(\b/n5757 ) );
  NAND \b/U5885  ( .A(msg[103]), .B(\b/n224 ), .Z(\b/n5723 ) );
  NAND \b/U5884  ( .A(msg[103]), .B(\b/n260 ), .Z(\b/n5675 ) );
  NAND \b/U5883  ( .A(msg[103]), .B(\b/n5779 ), .Z(\b/n5701 ) );
  NAND \b/U5882  ( .A(msg[103]), .B(\b/n5703 ), .Z(\b/n5663 ) );
  NAND \b/U5880  ( .A(\b/n283 ), .B(\b/n240 ), .Z(\b/n5785 ) );
  NAND \b/U5879  ( .A(msg[103]), .B(\b/n5782 ), .Z(\b/n5777 ) );
  NAND \b/U5878  ( .A(n704), .B(msg[103]), .Z(\b/n5763 ) );
  NAND \b/U5876  ( .A(msg[98]), .B(\b/n5444 ), .Z(\b/n5628 ) );
  NAND \b/U5875  ( .A(msg[97]), .B(\b/n240 ), .Z(\b/n5572 ) );
  NAND \b/U5874  ( .A(msg[103]), .B(\b/n5786 ), .Z(\b/n5571 ) );
  NAND \b/U5873  ( .A(\b/n5785 ), .B(msg[103]), .Z(\b/n5579 ) );
  NAND \b/U5871  ( .A(\b/n5444 ), .B(\b/n5605 ), .Z(\b/n5783 ) );
  NANDN \b/U5870  ( .B(\b/n275 ), .A(\b/n283 ), .Z(\b/n5782 ) );
  NAND \b/U5867  ( .A(msg[97]), .B(\b/n5449 ), .Z(\b/n5605 ) );
  NAND \b/U5866  ( .A(\b/n5444 ), .B(msg[97]), .Z(\b/n5512 ) );
  NAND \b/U5865  ( .A(\b/n275 ), .B(\b/n283 ), .Z(\b/n5779 ) );
  ANDN \b/U5862  ( .A(msg[98]), .B(msg[97]), .Z(\b/n5633 ) );
  AND \b/U5861  ( .A(\b/n5777 ), .B(\b/n5446 ), .Z(\b/n5539 ) );
  MUX \b/U5860  ( .IN0(\b/n5776 ), .IN1(\b/n5760 ), .SEL(msg[96]), .F(
        shift_row_out[103]) );
  MUX \b/U5859  ( .IN0(\b/n5775 ), .IN1(\b/n5768 ), .SEL(msg[102]), .F(
        \b/n5776 ) );
  MUX \b/U5858  ( .IN0(\b/n5774 ), .IN1(\b/n5771 ), .SEL(msg[98]), .F(
        \b/n5775 ) );
  MUX \b/U5857  ( .IN0(\b/n5773 ), .IN1(\b/n5772 ), .SEL(msg[101]), .F(
        \b/n5774 ) );
  MUX \b/U5856  ( .IN0(msg[100]), .IN1(\b/n228 ), .SEL(msg[103]), .F(\b/n5773 ) );
  MUX \b/U5855  ( .IN0(\b/n5511 ), .IN1(\b/n224 ), .SEL(msg[103]), .F(
        \b/n5772 ) );
  MUX \b/U5854  ( .IN0(\b/n5770 ), .IN1(\b/n5769 ), .SEL(msg[101]), .F(
        \b/n5771 ) );
  MUX \b/U5853  ( .IN0(\b/n5445 ), .IN1(\b/n232 ), .SEL(msg[103]), .F(
        \b/n5770 ) );
  MUX \b/U5852  ( .IN0(\b/n5457 ), .IN1(\b/n5466 ), .SEL(msg[103]), .F(
        \b/n5769 ) );
  MUX \b/U5851  ( .IN0(\b/n5767 ), .IN1(\b/n5764 ), .SEL(msg[98]), .F(
        \b/n5768 ) );
  MUX \b/U5850  ( .IN0(\b/n5766 ), .IN1(\b/n5765 ), .SEL(msg[101]), .F(
        \b/n5767 ) );
  MUX \b/U5849  ( .IN0(\b/n279 ), .IN1(\b/n241 ), .SEL(msg[103]), .F(\b/n5766 ) );
  MUX \b/U5848  ( .IN0(\b/n5468 ), .IN1(\b/n5443 ), .SEL(msg[103]), .F(
        \b/n5765 ) );
  MUX \b/U5847  ( .IN0(\b/n5762 ), .IN1(\b/n5761 ), .SEL(msg[101]), .F(
        \b/n5764 ) );
  NAND \b/U5846  ( .A(\b/n5572 ), .B(\b/n5763 ), .Z(\b/n5762 ) );
  MUX \b/U5845  ( .IN0(\b/n242 ), .IN1(\b/n5481 ), .SEL(msg[103]), .F(
        \b/n5761 ) );
  MUX \b/U5844  ( .IN0(\b/n5759 ), .IN1(\b/n5751 ), .SEL(msg[102]), .F(
        \b/n5760 ) );
  MUX \b/U5843  ( .IN0(\b/n5758 ), .IN1(\b/n5754 ), .SEL(msg[98]), .F(
        \b/n5759 ) );
  MUX \b/U5842  ( .IN0(\b/n5755 ), .IN1(\b/n5756 ), .SEL(msg[101]), .F(
        \b/n5758 ) );
  AND \b/U5841  ( .A(\b/n226 ), .B(\b/n5757 ), .Z(\b/n5756 ) );
  MUX \b/U5840  ( .IN0(\b/n5480 ), .IN1(\b/n5454 ), .SEL(msg[103]), .F(
        \b/n5755 ) );
  MUX \b/U5839  ( .IN0(\b/n5753 ), .IN1(\b/n5752 ), .SEL(msg[101]), .F(
        \b/n5754 ) );
  MUX \b/U5838  ( .IN0(\b/n260 ), .IN1(\b/n5476 ), .SEL(msg[103]), .F(
        \b/n5753 ) );
  MUX \b/U5837  ( .IN0(\b/n5461 ), .IN1(n703), .SEL(msg[103]), .F(\b/n5752 )
         );
  MUX \b/U5836  ( .IN0(\b/n5750 ), .IN1(\b/n5747 ), .SEL(msg[98]), .F(
        \b/n5751 ) );
  MUX \b/U5835  ( .IN0(\b/n5749 ), .IN1(\b/n5748 ), .SEL(msg[101]), .F(
        \b/n5750 ) );
  MUX \b/U5834  ( .IN0(\b/n5485 ), .IN1(\b/n5470 ), .SEL(msg[103]), .F(
        \b/n5749 ) );
  MUX \b/U5833  ( .IN0(\b/n5447 ), .IN1(\b/n5492 ), .SEL(msg[103]), .F(
        \b/n5748 ) );
  MUX \b/U5832  ( .IN0(\b/n5746 ), .IN1(\b/n5745 ), .SEL(msg[101]), .F(
        \b/n5747 ) );
  MUX \b/U5831  ( .IN0(\b/n239 ), .IN1(\b/n5444 ), .SEL(msg[103]), .F(
        \b/n5746 ) );
  MUX \b/U5830  ( .IN0(\b/n5478 ), .IN1(\b/n5744 ), .SEL(msg[103]), .F(
        \b/n5745 ) );
  MUX \b/U5829  ( .IN0(\b/n278 ), .IN1(\b/n220 ), .SEL(msg[97]), .F(\b/n5744 )
         );
  MUX \b/U5828  ( .IN0(\b/n5743 ), .IN1(\b/n5726 ), .SEL(msg[96]), .F(
        shift_row_out[102]) );
  MUX \b/U5827  ( .IN0(\b/n5742 ), .IN1(\b/n5733 ), .SEL(msg[102]), .F(
        \b/n5743 ) );
  MUX \b/U5826  ( .IN0(\b/n5741 ), .IN1(\b/n5737 ), .SEL(msg[98]), .F(
        \b/n5742 ) );
  MUX \b/U5825  ( .IN0(\b/n5740 ), .IN1(\b/n5738 ), .SEL(msg[101]), .F(
        \b/n5741 ) );
  MUX \b/U5824  ( .IN0(\b/n5739 ), .IN1(\b/n5458 ), .SEL(msg[103]), .F(
        \b/n5740 ) );
  MUX \b/U5823  ( .IN0(\b/n278 ), .IN1(\b/n5443 ), .SEL(msg[97]), .F(\b/n5739 ) );
  MUX \b/U5822  ( .IN0(n702), .IN1(\b/n5523 ), .SEL(msg[103]), .F(\b/n5738 )
         );
  MUX \b/U5821  ( .IN0(\b/n5736 ), .IN1(\b/n5734 ), .SEL(msg[101]), .F(
        \b/n5737 ) );
  MUX \b/U5820  ( .IN0(\b/n5735 ), .IN1(\b/n243 ), .SEL(msg[103]), .F(
        \b/n5736 ) );
  MUX \b/U5819  ( .IN0(\b/n5443 ), .IN1(\b/n5446 ), .SEL(msg[97]), .F(
        \b/n5735 ) );
  MUX \b/U5818  ( .IN0(\b/n5482 ), .IN1(\b/n5489 ), .SEL(msg[103]), .F(
        \b/n5734 ) );
  MUX \b/U5817  ( .IN0(\b/n5732 ), .IN1(\b/n5729 ), .SEL(msg[98]), .F(
        \b/n5733 ) );
  MUX \b/U5816  ( .IN0(\b/n5731 ), .IN1(\b/n5730 ), .SEL(msg[101]), .F(
        \b/n5732 ) );
  MUX \b/U5815  ( .IN0(\b/n258 ), .IN1(\b/n5452 ), .SEL(msg[103]), .F(
        \b/n5731 ) );
  MUX \b/U5814  ( .IN0(\b/n5472 ), .IN1(\b/n274 ), .SEL(msg[103]), .F(
        \b/n5730 ) );
  MUX \b/U5813  ( .IN0(\b/n5728 ), .IN1(\b/n5727 ), .SEL(msg[101]), .F(
        \b/n5729 ) );
  MUX \b/U5812  ( .IN0(\b/n5457 ), .IN1(n703), .SEL(msg[103]), .F(\b/n5728 )
         );
  MUX \b/U5811  ( .IN0(\b/n228 ), .IN1(\b/n241 ), .SEL(msg[103]), .F(\b/n5727 ) );
  MUX \b/U5810  ( .IN0(\b/n5725 ), .IN1(\b/n5717 ), .SEL(msg[102]), .F(
        \b/n5726 ) );
  MUX \b/U5809  ( .IN0(\b/n5724 ), .IN1(\b/n5720 ), .SEL(msg[98]), .F(
        \b/n5725 ) );
  MUX \b/U5808  ( .IN0(\b/n5722 ), .IN1(\b/n5721 ), .SEL(msg[101]), .F(
        \b/n5724 ) );
  AND \b/U5807  ( .A(\b/n272 ), .B(\b/n5723 ), .Z(\b/n5722 ) );
  MUX \b/U5806  ( .IN0(\b/n249 ), .IN1(\b/n5449 ), .SEL(msg[103]), .F(
        \b/n5721 ) );
  MUX \b/U5805  ( .IN0(\b/n5719 ), .IN1(\b/n5718 ), .SEL(msg[101]), .F(
        \b/n5720 ) );
  MUX \b/U5804  ( .IN0(\b/n5556 ), .IN1(msg[99]), .SEL(msg[103]), .F(\b/n5719 ) );
  MUX \b/U5802  ( .IN0(\b/n5716 ), .IN1(\b/n5712 ), .SEL(msg[98]), .F(
        \b/n5717 ) );
  MUX \b/U5801  ( .IN0(\b/n5715 ), .IN1(\b/n5714 ), .SEL(msg[101]), .F(
        \b/n5716 ) );
  MUX \b/U5800  ( .IN0(\b/n5462 ), .IN1(\b/n241 ), .SEL(msg[103]), .F(
        \b/n5715 ) );
  MUX \b/U5799  ( .IN0(\b/n220 ), .IN1(\b/n5713 ), .SEL(msg[103]), .F(
        \b/n5714 ) );
  MUX \b/U5798  ( .IN0(\b/n250 ), .IN1(\b/n262 ), .SEL(msg[97]), .F(\b/n5713 )
         );
  MUX \b/U5797  ( .IN0(\b/n5711 ), .IN1(\b/n5709 ), .SEL(msg[101]), .F(
        \b/n5712 ) );
  MUX \b/U5796  ( .IN0(\b/n5710 ), .IN1(\b/n5483 ), .SEL(msg[103]), .F(
        \b/n5711 ) );
  NANDN \b/U5795  ( .B(msg[100]), .A(msg[97]), .Z(\b/n5710 ) );
  MUX \b/U5794  ( .IN0(\b/n218 ), .IN1(\b/n5458 ), .SEL(msg[103]), .F(
        \b/n5709 ) );
  NANDN \b/U5793  ( .B(\b/n275 ), .A(msg[97]), .Z(\b/n5458 ) );
  MUX \b/U5792  ( .IN0(\b/n5708 ), .IN1(\b/n5688 ), .SEL(msg[96]), .F(
        shift_row_out[101]) );
  MUX \b/U5791  ( .IN0(\b/n5707 ), .IN1(\b/n5697 ), .SEL(msg[102]), .F(
        \b/n5708 ) );
  MUX \b/U5790  ( .IN0(\b/n5706 ), .IN1(\b/n5702 ), .SEL(msg[98]), .F(
        \b/n5707 ) );
  MUX \b/U5789  ( .IN0(\b/n5705 ), .IN1(\b/n5704 ), .SEL(msg[101]), .F(
        \b/n5706 ) );
  MUX \b/U5788  ( .IN0(\b/n5444 ), .IN1(\b/n242 ), .SEL(msg[103]), .F(
        \b/n5705 ) );
  MUX \b/U5787  ( .IN0(\b/n277 ), .IN1(\b/n5703 ), .SEL(msg[103]), .F(
        \b/n5704 ) );
  NAND \b/U5786  ( .A(\b/n262 ), .B(\b/n283 ), .Z(\b/n5703 ) );
  MUX \b/U5785  ( .IN0(\b/n5700 ), .IN1(\b/n5699 ), .SEL(msg[101]), .F(
        \b/n5702 ) );
  AND \b/U5784  ( .A(\b/n5474 ), .B(\b/n5701 ), .Z(\b/n5700 ) );
  MUX \b/U5783  ( .IN0(\b/n5444 ), .IN1(\b/n5698 ), .SEL(msg[103]), .F(
        \b/n5699 ) );
  NAND \b/U5782  ( .A(\b/n5443 ), .B(\b/n5512 ), .Z(\b/n5698 ) );
  MUX \b/U5781  ( .IN0(\b/n5696 ), .IN1(\b/n5692 ), .SEL(msg[98]), .F(
        \b/n5697 ) );
  MUX \b/U5780  ( .IN0(\b/n5695 ), .IN1(\b/n5693 ), .SEL(msg[101]), .F(
        \b/n5696 ) );
  MUX \b/U5779  ( .IN0(\b/n5457 ), .IN1(\b/n5694 ), .SEL(msg[103]), .F(
        \b/n5695 ) );
  NAND \b/U5778  ( .A(msg[97]), .B(\b/n227 ), .Z(\b/n5694 ) );
  MUX \b/U5777  ( .IN0(\b/n5483 ), .IN1(\b/n229 ), .SEL(msg[103]), .F(
        \b/n5693 ) );
  MUX \b/U5776  ( .IN0(\b/n5691 ), .IN1(\b/n5690 ), .SEL(msg[101]), .F(
        \b/n5692 ) );
  MUX \b/U5775  ( .IN0(\b/n275 ), .IN1(\b/n280 ), .SEL(msg[103]), .F(\b/n5691 ) );
  MUX \b/U5774  ( .IN0(\b/n5689 ), .IN1(\b/n5446 ), .SEL(n701), .F(\b/n5690 )
         );
  AND \b/U5773  ( .A(msg[103]), .B(msg[99]), .Z(\b/n5689 ) );
  MUX \b/U5772  ( .IN0(\b/n5687 ), .IN1(\b/n5677 ), .SEL(msg[102]), .F(
        \b/n5688 ) );
  MUX \b/U5771  ( .IN0(\b/n5686 ), .IN1(\b/n5683 ), .SEL(msg[98]), .F(
        \b/n5687 ) );
  MUX \b/U5770  ( .IN0(\b/n5685 ), .IN1(\b/n5684 ), .SEL(msg[101]), .F(
        \b/n5686 ) );
  MUX \b/U5769  ( .IN0(\b/n5464 ), .IN1(\b/n269 ), .SEL(msg[103]), .F(
        \b/n5685 ) );
  MUX \b/U5768  ( .IN0(\b/n237 ), .IN1(n700), .SEL(msg[103]), .F(\b/n5684 ) );
  MUX \b/U5767  ( .IN0(\b/n5682 ), .IN1(\b/n5680 ), .SEL(msg[101]), .F(
        \b/n5683 ) );
  MUX \b/U5766  ( .IN0(\b/n5489 ), .IN1(\b/n5681 ), .SEL(msg[103]), .F(
        \b/n5682 ) );
  MUX \b/U5765  ( .IN0(\b/n240 ), .IN1(\b/n262 ), .SEL(msg[97]), .F(\b/n5681 )
         );
  MUX \b/U5764  ( .IN0(\b/n5679 ), .IN1(\b/n5678 ), .SEL(msg[103]), .F(
        \b/n5680 ) );
  AND \b/U5763  ( .A(\b/n5468 ), .B(\b/n5523 ), .Z(\b/n5679 ) );
  MUX \b/U5762  ( .IN0(\b/n227 ), .IN1(\b/n275 ), .SEL(msg[97]), .F(\b/n5678 )
         );
  MUX \b/U5761  ( .IN0(\b/n5676 ), .IN1(\b/n5672 ), .SEL(msg[98]), .F(
        \b/n5677 ) );
  MUX \b/U5760  ( .IN0(\b/n5673 ), .IN1(\b/n5674 ), .SEL(msg[101]), .F(
        \b/n5676 ) );
  AND \b/U5759  ( .A(\b/n5675 ), .B(\b/n5572 ), .Z(\b/n5674 ) );
  MUX \b/U5758  ( .IN0(\b/n5604 ), .IN1(\b/n5446 ), .SEL(msg[103]), .F(
        \b/n5673 ) );
  MUX \b/U5757  ( .IN0(\b/n5671 ), .IN1(\b/n5670 ), .SEL(msg[101]), .F(
        \b/n5672 ) );
  MUX \b/U5756  ( .IN0(n699), .IN1(\b/n270 ), .SEL(msg[103]), .F(\b/n5671 ) );
  MUX \b/U5755  ( .IN0(\b/n276 ), .IN1(\b/n240 ), .SEL(msg[103]), .F(\b/n5670 ) );
  MUX \b/U5754  ( .IN0(\b/n5669 ), .IN1(\b/n5654 ), .SEL(msg[96]), .F(
        shift_row_out[100]) );
  MUX \b/U5753  ( .IN0(\b/n5668 ), .IN1(\b/n5660 ), .SEL(msg[102]), .F(
        \b/n5669 ) );
  MUX \b/U5752  ( .IN0(\b/n5667 ), .IN1(\b/n5664 ), .SEL(msg[98]), .F(
        \b/n5668 ) );
  MUX \b/U5751  ( .IN0(\b/n5666 ), .IN1(\b/n5665 ), .SEL(msg[101]), .F(
        \b/n5667 ) );
  MUX \b/U5750  ( .IN0(\b/n251 ), .IN1(\b/n244 ), .SEL(msg[103]), .F(\b/n5666 ) );
  MUX \b/U5749  ( .IN0(\b/n5473 ), .IN1(\b/n266 ), .SEL(msg[103]), .F(
        \b/n5665 ) );
  MUX \b/U5748  ( .IN0(\b/n5661 ), .IN1(\b/n5662 ), .SEL(msg[101]), .F(
        \b/n5664 ) );
  AND \b/U5747  ( .A(\b/n5474 ), .B(\b/n5663 ), .Z(\b/n5662 ) );
  MUX \b/U5746  ( .IN0(\b/n5523 ), .IN1(\b/n5489 ), .SEL(msg[103]), .F(
        \b/n5661 ) );
  NAND \b/U5745  ( .A(msg[97]), .B(\b/n5443 ), .Z(\b/n5523 ) );
  MUX \b/U5744  ( .IN0(\b/n5659 ), .IN1(\b/n5656 ), .SEL(msg[98]), .F(
        \b/n5660 ) );
  MUX \b/U5743  ( .IN0(\b/n5658 ), .IN1(\b/n5657 ), .SEL(msg[101]), .F(
        \b/n5659 ) );
  MUX \b/U5742  ( .IN0(\b/n5466 ), .IN1(\b/n249 ), .SEL(msg[103]), .F(
        \b/n5658 ) );
  MUX \b/U5741  ( .IN0(n698), .IN1(\b/n251 ), .SEL(msg[103]), .F(\b/n5657 ) );
  MUX \b/U5740  ( .IN0(\b/n5448 ), .IN1(\b/n5655 ), .SEL(msg[101]), .F(
        \b/n5656 ) );
  MUX \b/U5739  ( .IN0(\b/n5479 ), .IN1(\b/n5480 ), .SEL(msg[103]), .F(
        \b/n5655 ) );
  MUX \b/U5738  ( .IN0(\b/n5653 ), .IN1(\b/n5645 ), .SEL(msg[102]), .F(
        \b/n5654 ) );
  MUX \b/U5737  ( .IN0(\b/n5652 ), .IN1(\b/n5648 ), .SEL(msg[98]), .F(
        \b/n5653 ) );
  MUX \b/U5736  ( .IN0(\b/n5651 ), .IN1(\b/n5650 ), .SEL(msg[101]), .F(
        \b/n5652 ) );
  MUX \b/U5735  ( .IN0(\b/n272 ), .IN1(\b/n253 ), .SEL(msg[103]), .F(\b/n5651 ) );
  MUX \b/U5734  ( .IN0(\b/n5467 ), .IN1(\b/n5649 ), .SEL(msg[103]), .F(
        \b/n5650 ) );
  AND \b/U5733  ( .A(\b/n5444 ), .B(\b/n283 ), .Z(\b/n5649 ) );
  MUX \b/U5732  ( .IN0(\b/n5647 ), .IN1(\b/n5646 ), .SEL(msg[101]), .F(
        \b/n5648 ) );
  MUX \b/U5731  ( .IN0(\b/n275 ), .IN1(\b/n5444 ), .SEL(msg[103]), .F(
        \b/n5647 ) );
  MUX \b/U5730  ( .IN0(\b/n226 ), .IN1(\b/n247 ), .SEL(msg[103]), .F(\b/n5646 ) );
  MUX \b/U5729  ( .IN0(\b/n5644 ), .IN1(\b/n5642 ), .SEL(msg[98]), .F(
        \b/n5645 ) );
  MUX \b/U5728  ( .IN0(\b/n5643 ), .IN1(\b/n215 ), .SEL(msg[101]), .F(
        \b/n5644 ) );
  MUX \b/U5727  ( .IN0(\b/n239 ), .IN1(\b/n5450 ), .SEL(msg[103]), .F(
        \b/n5643 ) );
  MUX \b/U5726  ( .IN0(\b/n5641 ), .IN1(\b/n5640 ), .SEL(msg[101]), .F(
        \b/n5642 ) );
  MUX \b/U5725  ( .IN0(\b/n240 ), .IN1(\b/n5470 ), .SEL(msg[103]), .F(
        \b/n5641 ) );
  MUX \b/U5724  ( .IN0(\b/n219 ), .IN1(\b/n5444 ), .SEL(msg[103]), .F(
        \b/n5640 ) );
  MUX \b/U5723  ( .IN0(\b/n5639 ), .IN1(\b/n5621 ), .SEL(msg[96]), .F(
        shift_row_out[99]) );
  MUX \b/U5722  ( .IN0(\b/n5638 ), .IN1(\b/n5630 ), .SEL(msg[102]), .F(
        \b/n5639 ) );
  MUX \b/U5721  ( .IN0(\b/n5637 ), .IN1(\b/n5634 ), .SEL(msg[101]), .F(
        \b/n5638 ) );
  MUX \b/U5720  ( .IN0(\b/n5636 ), .IN1(\b/n5635 ), .SEL(msg[103]), .F(
        \b/n5637 ) );
  MUX \b/U5719  ( .IN0(\b/n5462 ), .IN1(\b/n247 ), .SEL(msg[98]), .F(\b/n5636 ) );
  MUX \b/U5718  ( .IN0(n700), .IN1(\b/n271 ), .SEL(msg[98]), .F(\b/n5635 ) );
  MUX \b/U5717  ( .IN0(\b/n5632 ), .IN1(\b/n5631 ), .SEL(msg[103]), .F(
        \b/n5634 ) );
  AND \b/U5716  ( .A(\b/n5633 ), .B(msg[100]), .Z(\b/n5632 ) );
  MUX \b/U5715  ( .IN0(\b/n233 ), .IN1(\b/n5475 ), .SEL(msg[98]), .F(\b/n5631 ) );
  MUX \b/U5714  ( .IN0(\b/n5629 ), .IN1(\b/n5625 ), .SEL(msg[101]), .F(
        \b/n5630 ) );
  MUX \b/U5713  ( .IN0(\b/n5627 ), .IN1(\b/n5626 ), .SEL(msg[103]), .F(
        \b/n5629 ) );
  NAND \b/U5712  ( .A(\b/n275 ), .B(\b/n5628 ), .Z(\b/n5627 ) );
  MUX \b/U5711  ( .IN0(\b/n270 ), .IN1(\b/n224 ), .SEL(msg[98]), .F(\b/n5626 )
         );
  MUX \b/U5710  ( .IN0(\b/n5624 ), .IN1(\b/n5622 ), .SEL(msg[103]), .F(
        \b/n5625 ) );
  MUX \b/U5709  ( .IN0(\b/n5457 ), .IN1(\b/n5623 ), .SEL(msg[98]), .F(
        \b/n5624 ) );
  AND \b/U5708  ( .A(msg[97]), .B(\b/n275 ), .Z(\b/n5623 ) );
  MUX \b/U5707  ( .IN0(\b/n259 ), .IN1(\b/n5474 ), .SEL(msg[98]), .F(\b/n5622 ) );
  MUX \b/U5706  ( .IN0(\b/n5620 ), .IN1(\b/n5610 ), .SEL(msg[102]), .F(
        \b/n5621 ) );
  MUX \b/U5705  ( .IN0(\b/n5619 ), .IN1(\b/n5616 ), .SEL(msg[101]), .F(
        \b/n5620 ) );
  MUX \b/U5704  ( .IN0(\b/n5618 ), .IN1(\b/n5617 ), .SEL(msg[103]), .F(
        \b/n5619 ) );
  MUX \b/U5703  ( .IN0(\b/n5464 ), .IN1(n697), .SEL(msg[98]), .F(\b/n5618 ) );
  MUX \b/U5702  ( .IN0(\b/n221 ), .IN1(\b/n219 ), .SEL(msg[98]), .F(\b/n5617 )
         );
  MUX \b/U5701  ( .IN0(\b/n5612 ), .IN1(\b/n5613 ), .SEL(msg[103]), .F(
        \b/n5616 ) );
  NAND \b/U5700  ( .A(\b/n5614 ), .B(\b/n5615 ), .Z(\b/n5613 ) );
  MUX \b/U5699  ( .IN0(\b/n248 ), .IN1(\b/n5611 ), .SEL(msg[98]), .F(\b/n5612 ) );
  MUX \b/U5698  ( .IN0(\b/n220 ), .IN1(\b/n278 ), .SEL(msg[97]), .F(\b/n5611 )
         );
  MUX \b/U5697  ( .IN0(\b/n5609 ), .IN1(\b/n5603 ), .SEL(msg[101]), .F(
        \b/n5610 ) );
  MUX \b/U5696  ( .IN0(\b/n5608 ), .IN1(\b/n5606 ), .SEL(msg[103]), .F(
        \b/n5609 ) );
  MUX \b/U5695  ( .IN0(\b/n5607 ), .IN1(\b/n5446 ), .SEL(\b/n5491 ), .F(
        \b/n5608 ) );
  MUX \b/U5694  ( .IN0(msg[99]), .IN1(msg[100]), .SEL(msg[98]), .F(\b/n5607 )
         );
  MUX \b/U5693  ( .IN0(\b/n5474 ), .IN1(\b/n5604 ), .SEL(msg[98]), .F(
        \b/n5606 ) );
  NAND \b/U5692  ( .A(\b/n5446 ), .B(\b/n5605 ), .Z(\b/n5604 ) );
  MUX \b/U5691  ( .IN0(\b/n5600 ), .IN1(\b/n5601 ), .SEL(msg[103]), .F(
        \b/n5603 ) );
  AND \b/U5690  ( .A(\b/n236 ), .B(\b/n5602 ), .Z(\b/n5601 ) );
  MUX \b/U5689  ( .IN0(\b/n225 ), .IN1(\b/n5445 ), .SEL(msg[98]), .F(\b/n5600 ) );
  MUX \b/U5688  ( .IN0(\b/n5599 ), .IN1(\b/n5583 ), .SEL(msg[96]), .F(
        shift_row_out[98]) );
  MUX \b/U5687  ( .IN0(\b/n5598 ), .IN1(\b/n5590 ), .SEL(msg[102]), .F(
        \b/n5599 ) );
  MUX \b/U5686  ( .IN0(\b/n5597 ), .IN1(\b/n5593 ), .SEL(msg[98]), .F(
        \b/n5598 ) );
  MUX \b/U5685  ( .IN0(\b/n5596 ), .IN1(\b/n5594 ), .SEL(msg[101]), .F(
        \b/n5597 ) );
  MUX \b/U5684  ( .IN0(\b/n233 ), .IN1(\b/n5595 ), .SEL(msg[103]), .F(
        \b/n5596 ) );
  MUX \b/U5683  ( .IN0(\b/n5444 ), .IN1(\b/n275 ), .SEL(msg[97]), .F(\b/n5595 ) );
  MUX \b/U5682  ( .IN0(\b/n5445 ), .IN1(\b/n216 ), .SEL(msg[103]), .F(
        \b/n5594 ) );
  MUX \b/U5681  ( .IN0(\b/n5592 ), .IN1(\b/n5591 ), .SEL(msg[101]), .F(
        \b/n5593 ) );
  MUX \b/U5680  ( .IN0(\b/n5490 ), .IN1(\b/n243 ), .SEL(msg[103]), .F(
        \b/n5592 ) );
  MUX \b/U5679  ( .IN0(\b/n257 ), .IN1(\b/n5478 ), .SEL(msg[103]), .F(
        \b/n5591 ) );
  MUX \b/U5678  ( .IN0(\b/n5589 ), .IN1(\b/n5586 ), .SEL(msg[98]), .F(
        \b/n5590 ) );
  MUX \b/U5677  ( .IN0(\b/n5588 ), .IN1(\b/n5587 ), .SEL(msg[101]), .F(
        \b/n5589 ) );
  MUX \b/U5676  ( .IN0(\b/n244 ), .IN1(msg[97]), .SEL(msg[103]), .F(\b/n5588 )
         );
  MUX \b/U5675  ( .IN0(\b/n281 ), .IN1(\b/n242 ), .SEL(msg[103]), .F(\b/n5587 ) );
  MUX \b/U5674  ( .IN0(n702), .IN1(\b/n5585 ), .SEL(msg[103]), .F(\b/n5586 )
         );
  MUX \b/U5673  ( .IN0(\b/n5460 ), .IN1(\b/n5584 ), .SEL(msg[101]), .F(
        \b/n5585 ) );
  MUX \b/U5672  ( .IN0(\b/n275 ), .IN1(\b/n250 ), .SEL(msg[97]), .F(\b/n5584 )
         );
  MUX \b/U5671  ( .IN0(\b/n5582 ), .IN1(\b/n5574 ), .SEL(msg[102]), .F(
        \b/n5583 ) );
  MUX \b/U5670  ( .IN0(\b/n5581 ), .IN1(\b/n5576 ), .SEL(msg[98]), .F(
        \b/n5582 ) );
  MUX \b/U5669  ( .IN0(\b/n5578 ), .IN1(\b/n5577 ), .SEL(msg[101]), .F(
        \b/n5581 ) );
  NAND \b/U5668  ( .A(\b/n5579 ), .B(\b/n5580 ), .Z(\b/n5578 ) );
  MUX \b/U5667  ( .IN0(n699), .IN1(\b/n232 ), .SEL(msg[103]), .F(\b/n5577 ) );
  MUX \b/U5666  ( .IN0(\b/n215 ), .IN1(\b/n5575 ), .SEL(msg[101]), .F(
        \b/n5576 ) );
  MUX \b/U5665  ( .IN0(\b/n5459 ), .IN1(n699), .SEL(msg[103]), .F(\b/n5575 )
         );
  MUX \b/U5664  ( .IN0(\b/n5573 ), .IN1(\b/n5568 ), .SEL(msg[98]), .F(
        \b/n5574 ) );
  MUX \b/U5663  ( .IN0(\b/n5570 ), .IN1(\b/n5569 ), .SEL(msg[101]), .F(
        \b/n5573 ) );
  NAND \b/U5662  ( .A(\b/n5571 ), .B(\b/n5572 ), .Z(\b/n5570 ) );
  MUX \b/U5661  ( .IN0(\b/n5489 ), .IN1(\b/n217 ), .SEL(msg[103]), .F(
        \b/n5569 ) );
  MUX \b/U5660  ( .IN0(\b/n5567 ), .IN1(\b/n5565 ), .SEL(msg[101]), .F(
        \b/n5568 ) );
  MUX \b/U5659  ( .IN0(\b/n5446 ), .IN1(\b/n5566 ), .SEL(n701), .F(\b/n5567 )
         );
  MUX \b/U5658  ( .IN0(msg[99]), .IN1(\b/n220 ), .SEL(msg[103]), .F(\b/n5566 )
         );
  MUX \b/U5657  ( .IN0(\b/n5447 ), .IN1(\b/n5564 ), .SEL(msg[103]), .F(
        \b/n5565 ) );
  MUX \b/U5656  ( .IN0(\b/n5449 ), .IN1(\b/n5444 ), .SEL(msg[97]), .F(
        \b/n5564 ) );
  MUX \b/U5655  ( .IN0(\b/n5563 ), .IN1(\b/n5545 ), .SEL(msg[96]), .F(
        shift_row_out[97]) );
  MUX \b/U5654  ( .IN0(\b/n5562 ), .IN1(\b/n5553 ), .SEL(msg[102]), .F(
        \b/n5563 ) );
  MUX \b/U5653  ( .IN0(\b/n5561 ), .IN1(\b/n5558 ), .SEL(msg[98]), .F(
        \b/n5562 ) );
  MUX \b/U5652  ( .IN0(\b/n5560 ), .IN1(\b/n5559 ), .SEL(msg[101]), .F(
        \b/n5561 ) );
  MUX \b/U5651  ( .IN0(\b/n238 ), .IN1(n704), .SEL(msg[103]), .F(\b/n5560 ) );
  MUX \b/U5650  ( .IN0(\b/n272 ), .IN1(\b/n5461 ), .SEL(msg[103]), .F(
        \b/n5559 ) );
  MUX \b/U5649  ( .IN0(\b/n5557 ), .IN1(\b/n5555 ), .SEL(msg[101]), .F(
        \b/n5558 ) );
  MUX \b/U5648  ( .IN0(\b/n5556 ), .IN1(n698), .SEL(msg[103]), .F(\b/n5557 )
         );
  NAND \b/U5647  ( .A(\b/n283 ), .B(\b/n227 ), .Z(\b/n5556 ) );
  MUX \b/U5646  ( .IN0(\b/n5468 ), .IN1(\b/n5554 ), .SEL(msg[103]), .F(
        \b/n5555 ) );
  AND \b/U5645  ( .A(msg[97]), .B(msg[100]), .Z(\b/n5554 ) );
  MUX \b/U5644  ( .IN0(\b/n5552 ), .IN1(\b/n5549 ), .SEL(msg[98]), .F(
        \b/n5553 ) );
  MUX \b/U5643  ( .IN0(\b/n5551 ), .IN1(\b/n5550 ), .SEL(msg[101]), .F(
        \b/n5552 ) );
  MUX \b/U5642  ( .IN0(\b/n5452 ), .IN1(\b/n229 ), .SEL(msg[103]), .F(
        \b/n5551 ) );
  MUX \b/U5641  ( .IN0(\b/n244 ), .IN1(\b/n262 ), .SEL(msg[103]), .F(\b/n5550 ) );
  MUX \b/U5640  ( .IN0(\b/n5548 ), .IN1(\b/n5546 ), .SEL(msg[101]), .F(
        \b/n5549 ) );
  MUX \b/U5639  ( .IN0(\b/n5547 ), .IN1(\b/n276 ), .SEL(msg[103]), .F(
        \b/n5548 ) );
  MUX \b/U5638  ( .IN0(\b/n5468 ), .IN1(\b/n220 ), .SEL(msg[97]), .F(\b/n5547 ) );
  MUX \b/U5637  ( .IN0(\b/n238 ), .IN1(\b/n259 ), .SEL(msg[103]), .F(\b/n5546 ) );
  MUX \b/U5636  ( .IN0(\b/n5544 ), .IN1(\b/n5536 ), .SEL(msg[102]), .F(
        \b/n5545 ) );
  MUX \b/U5635  ( .IN0(\b/n5543 ), .IN1(\b/n5540 ), .SEL(msg[98]), .F(
        \b/n5544 ) );
  MUX \b/U5634  ( .IN0(\b/n5542 ), .IN1(\b/n5541 ), .SEL(msg[101]), .F(
        \b/n5543 ) );
  MUX \b/U5633  ( .IN0(\b/n5488 ), .IN1(\b/n281 ), .SEL(msg[103]), .F(
        \b/n5542 ) );
  MUX \b/U5632  ( .IN0(\b/n5463 ), .IN1(\b/n5444 ), .SEL(msg[103]), .F(
        \b/n5541 ) );
  MUX \b/U5631  ( .IN0(\b/n5537 ), .IN1(\b/n5538 ), .SEL(msg[101]), .F(
        \b/n5540 ) );
  AND \b/U5630  ( .A(\b/n5539 ), .B(\b/n5512 ), .Z(\b/n5538 ) );
  MUX \b/U5629  ( .IN0(\b/n264 ), .IN1(\b/n5459 ), .SEL(msg[103]), .F(
        \b/n5537 ) );
  MUX \b/U5628  ( .IN0(\b/n5535 ), .IN1(\b/n5531 ), .SEL(msg[98]), .F(
        \b/n5536 ) );
  MUX \b/U5627  ( .IN0(\b/n5534 ), .IN1(\b/n5487 ), .SEL(msg[101]), .F(
        \b/n5535 ) );
  MUX \b/U5626  ( .IN0(\b/n5532 ), .IN1(\b/n5533 ), .SEL(msg[103]), .F(
        \b/n5534 ) );
  NAND \b/U5625  ( .A(\b/n5444 ), .B(\b/n5523 ), .Z(\b/n5533 ) );
  MUX \b/U5624  ( .IN0(\b/n5444 ), .IN1(\b/n220 ), .SEL(msg[97]), .F(\b/n5532 ) );
  MUX \b/U5623  ( .IN0(\b/n5530 ), .IN1(\b/n5529 ), .SEL(msg[101]), .F(
        \b/n5531 ) );
  MUX \b/U5622  ( .IN0(\b/n5471 ), .IN1(\b/n5469 ), .SEL(msg[103]), .F(
        \b/n5530 ) );
  MUX \b/U5621  ( .IN0(\b/n227 ), .IN1(\b/n242 ), .SEL(msg[103]), .F(\b/n5529 ) );
  MUX \b/U5620  ( .IN0(\b/n5528 ), .IN1(\b/n5509 ), .SEL(msg[96]), .F(
        shift_row_out[96]) );
  MUX \b/U5619  ( .IN0(\b/n5527 ), .IN1(\b/n5519 ), .SEL(msg[102]), .F(
        \b/n5528 ) );
  MUX \b/U5618  ( .IN0(\b/n5526 ), .IN1(\b/n5524 ), .SEL(msg[98]), .F(
        \b/n5527 ) );
  MUX \b/U5617  ( .IN0(\b/n221 ), .IN1(\b/n5525 ), .SEL(msg[103]), .F(
        \b/n5526 ) );
  MUX \b/U5616  ( .IN0(\b/n257 ), .IN1(\b/n240 ), .SEL(msg[101]), .F(\b/n5525 ) );
  MUX \b/U5615  ( .IN0(\b/n5521 ), .IN1(\b/n5520 ), .SEL(msg[103]), .F(
        \b/n5524 ) );
  NAND \b/U5614  ( .A(\b/n5522 ), .B(\b/n5523 ), .Z(\b/n5521 ) );
  MUX \b/U5613  ( .IN0(\b/n256 ), .IN1(\b/n283 ), .SEL(msg[101]), .F(\b/n5520 ) );
  MUX \b/U5612  ( .IN0(\b/n5518 ), .IN1(\b/n5514 ), .SEL(msg[98]), .F(
        \b/n5519 ) );
  MUX \b/U5611  ( .IN0(\b/n5517 ), .IN1(\b/n5516 ), .SEL(msg[103]), .F(
        \b/n5518 ) );
  MUX \b/U5610  ( .IN0(n697), .IN1(\b/n273 ), .SEL(msg[101]), .F(\b/n5517 ) );
  MUX \b/U5609  ( .IN0(\b/n5515 ), .IN1(\b/n236 ), .SEL(msg[101]), .F(
        \b/n5516 ) );
  NAND \b/U5608  ( .A(\b/n5443 ), .B(\b/n5445 ), .Z(\b/n5515 ) );
  MUX \b/U5607  ( .IN0(\b/n5513 ), .IN1(\b/n5510 ), .SEL(msg[103]), .F(
        \b/n5514 ) );
  MUX \b/U5606  ( .IN0(\b/n277 ), .IN1(\b/n5511 ), .SEL(msg[101]), .F(
        \b/n5513 ) );
  NAND \b/U5605  ( .A(\b/n5449 ), .B(\b/n5512 ), .Z(\b/n5511 ) );
  MUX \b/U5604  ( .IN0(\b/n265 ), .IN1(\b/n5453 ), .SEL(msg[101]), .F(
        \b/n5510 ) );
  MUX \b/U5603  ( .IN0(\b/n5508 ), .IN1(\b/n5500 ), .SEL(msg[102]), .F(
        \b/n5509 ) );
  MUX \b/U5602  ( .IN0(\b/n5507 ), .IN1(\b/n5503 ), .SEL(msg[98]), .F(
        \b/n5508 ) );
  MUX \b/U5601  ( .IN0(\b/n5506 ), .IN1(\b/n5504 ), .SEL(msg[103]), .F(
        \b/n5507 ) );
  MUX \b/U5600  ( .IN0(\b/n5505 ), .IN1(\b/n235 ), .SEL(msg[101]), .F(
        \b/n5506 ) );
  NAND \b/U5599  ( .A(\b/n283 ), .B(\b/n5446 ), .Z(\b/n5505 ) );
  MUX \b/U5597  ( .IN0(\b/n5502 ), .IN1(\b/n5501 ), .SEL(msg[103]), .F(
        \b/n5503 ) );
  MUX \b/U5596  ( .IN0(n699), .IN1(\b/n271 ), .SEL(msg[101]), .F(\b/n5502 ) );
  MUX \b/U5595  ( .IN0(\b/n237 ), .IN1(\b/n275 ), .SEL(msg[101]), .F(\b/n5501 ) );
  MUX \b/U5594  ( .IN0(\b/n5499 ), .IN1(\b/n5495 ), .SEL(msg[98]), .F(
        \b/n5500 ) );
  MUX \b/U5593  ( .IN0(\b/n5497 ), .IN1(\b/n5496 ), .SEL(msg[103]), .F(
        \b/n5499 ) );
  NAND \b/U5592  ( .A(\b/n5498 ), .B(\b/n5486 ), .Z(\b/n5497 ) );
  MUX \b/U5591  ( .IN0(msg[99]), .IN1(\b/n5478 ), .SEL(msg[101]), .F(\b/n5496 ) );
  MUX \b/U5590  ( .IN0(\b/n5494 ), .IN1(\b/n5493 ), .SEL(msg[103]), .F(
        \b/n5495 ) );
  MUX \b/U5589  ( .IN0(\b/n217 ), .IN1(\b/n5456 ), .SEL(msg[101]), .F(
        \b/n5494 ) );
  MUX \b/U5588  ( .IN0(\b/n255 ), .IN1(\b/n264 ), .SEL(msg[101]), .F(\b/n5493 ) );
  XOR \b/U5587  ( .A(\b/n5446 ), .B(msg[97]), .Z(\b/n5492 ) );
  XOR \b/U5586  ( .A(msg[97]), .B(msg[98]), .Z(\b/n5491 ) );
  XOR \b/U5585  ( .A(msg[97]), .B(msg[99]), .Z(\b/n5490 ) );
  XOR \b/U5584  ( .A(\b/n283 ), .B(\b/n275 ), .Z(\b/n5489 ) );
  XOR \b/U5583  ( .A(msg[97]), .B(\b/n240 ), .Z(\b/n5488 ) );
  XOR \b/U5581  ( .A(\b/n278 ), .B(msg[100]), .Z(\b/n5468 ) );
  XOR \b/U5580  ( .A(msg[101]), .B(msg[97]), .Z(\b/n5486 ) );
  MUX \b/U5579  ( .IN0(\b/n5446 ), .IN1(\b/n275 ), .SEL(msg[97]), .F(\b/n5485 ) );
  MUX \b/U5577  ( .IN0(\b/n227 ), .IN1(\b/n250 ), .SEL(msg[97]), .F(\b/n5483 )
         );
  MUX \b/U5576  ( .IN0(msg[99]), .IN1(\b/n250 ), .SEL(msg[97]), .F(\b/n5482 )
         );
  MUX \b/U5575  ( .IN0(\b/n5449 ), .IN1(\b/n5468 ), .SEL(msg[97]), .F(
        \b/n5481 ) );
  MUX \b/U5574  ( .IN0(msg[100]), .IN1(\b/n227 ), .SEL(msg[97]), .F(\b/n5480 )
         );
  NAND \b/U5573  ( .A(\b/n250 ), .B(\b/n283 ), .Z(\b/n5479 ) );
  OR \b/U5572  ( .A(msg[100]), .B(msg[97]), .Z(\b/n5478 ) );
  MUX \b/U5570  ( .IN0(\b/n250 ), .IN1(msg[100]), .SEL(msg[97]), .F(\b/n5476 )
         );
  MUX \b/U5569  ( .IN0(\b/n278 ), .IN1(msg[100]), .SEL(msg[97]), .F(\b/n5475 )
         );
  MUX \b/U5568  ( .IN0(\b/n5443 ), .IN1(\b/n5444 ), .SEL(msg[97]), .F(
        \b/n5474 ) );
  MUX \b/U5567  ( .IN0(\b/n220 ), .IN1(\b/n250 ), .SEL(msg[97]), .F(\b/n5473 )
         );
  MUX \b/U5566  ( .IN0(\b/n5443 ), .IN1(msg[100]), .SEL(msg[97]), .F(\b/n5472 ) );
  XOR \b/U5565  ( .A(\b/n283 ), .B(msg[100]), .Z(\b/n5471 ) );
  MUX \b/U5564  ( .IN0(\b/n262 ), .IN1(\b/n227 ), .SEL(msg[97]), .F(\b/n5470 )
         );
  NANDN \b/U5563  ( .B(msg[97]), .A(msg[99]), .Z(\b/n5469 ) );
  MUX \b/U5562  ( .IN0(\b/n5468 ), .IN1(\b/n262 ), .SEL(msg[97]), .F(\b/n5467 ) );
  MUX \b/U5561  ( .IN0(\b/n275 ), .IN1(msg[99]), .SEL(msg[97]), .F(\b/n5466 )
         );
  NAND \b/U5559  ( .A(\b/n5449 ), .B(\b/n283 ), .Z(\b/n5464 ) );
  MUX \b/U5558  ( .IN0(msg[100]), .IN1(\b/n5446 ), .SEL(msg[97]), .F(\b/n5463 ) );
  MUX \b/U5557  ( .IN0(msg[100]), .IN1(\b/n240 ), .SEL(msg[97]), .F(\b/n5462 )
         );
  MUX \b/U5556  ( .IN0(\b/n275 ), .IN1(\b/n278 ), .SEL(msg[97]), .F(\b/n5461 )
         );
  NAND \b/U5555  ( .A(\b/n5445 ), .B(\b/n275 ), .Z(\b/n5460 ) );
  MUX \b/U5554  ( .IN0(\b/n5446 ), .IN1(\b/n5444 ), .SEL(msg[97]), .F(
        \b/n5459 ) );
  NAND \b/U5553  ( .A(\b/n5458 ), .B(\b/n5443 ), .Z(\b/n5457 ) );
  MUX \b/U5552  ( .IN0(\b/n5446 ), .IN1(\b/n278 ), .SEL(msg[97]), .F(\b/n5456 ) );
  NANDN \b/U5550  ( .B(msg[100]), .A(msg[99]), .Z(\b/n5446 ) );
  MUX \b/U5549  ( .IN0(\b/n5449 ), .IN1(\b/n278 ), .SEL(msg[97]), .F(\b/n5454 ) );
  MUX \b/U5548  ( .IN0(\b/n278 ), .IN1(\b/n227 ), .SEL(msg[97]), .F(\b/n5453 )
         );
  MUX \b/U5547  ( .IN0(\b/n5449 ), .IN1(msg[99]), .SEL(msg[97]), .F(\b/n5452 )
         );
  OR \b/U5546  ( .A(msg[100]), .B(msg[99]), .Z(\b/n5449 ) );
  MUX \b/U5545  ( .IN0(\b/n275 ), .IN1(\b/n227 ), .SEL(msg[97]), .F(\b/n5451 )
         );
  NANDN \b/U5544  ( .B(msg[99]), .A(msg[97]), .Z(\b/n5450 ) );
  NAND \b/U5543  ( .A(\b/n5449 ), .B(\b/n5445 ), .Z(\b/n5448 ) );
  NAND \b/U5542  ( .A(msg[97]), .B(msg[99]), .Z(\b/n5447 ) );
  NAND \b/U5541  ( .A(msg[97]), .B(\b/n5446 ), .Z(\b/n5445 ) );
  NANDN \b/U5540  ( .B(msg[99]), .A(msg[100]), .Z(\b/n5444 ) );
  NAND \b/U5539  ( .A(msg[100]), .B(msg[99]), .Z(\b/n5443 ) );
  MUX \b/U5538  ( .IN0(msg[92]), .IN1(\b/n5084 ), .SEL(msg[89]), .F(\b/n5442 )
         );
  MUX \b/U5537  ( .IN0(msg[92]), .IN1(\b/n5093 ), .SEL(msg[89]), .F(\b/n5441 )
         );
  MUX \b/U5536  ( .IN0(\b/n5085 ), .IN1(\b/n5088 ), .SEL(msg[89]), .F(
        \b/n5440 ) );
  MUX \b/U5535  ( .IN0(\b/n5090 ), .IN1(\b/n343 ), .SEL(msg[89]), .F(\b/n5439 ) );
  MUX \b/U5533  ( .IN0(\b/n5093 ), .IN1(\b/n5084 ), .SEL(msg[90]), .F(
        \b/n5266 ) );
  MUX \b/U5532  ( .IN0(\b/n5086 ), .IN1(\b/n354 ), .SEL(msg[90]), .F(\b/n5267 ) );
  MUX \b/U5531  ( .IN0(\b/n297 ), .IN1(\b/n307 ), .SEL(msg[89]), .F(\b/n5230 )
         );
  MUX \b/U5530  ( .IN0(\b/n5114 ), .IN1(\b/n5425 ), .SEL(msg[95]), .F(
        \b/n5437 ) );
  MUX \b/U5529  ( .IN0(\b/n5088 ), .IN1(\b/n5084 ), .SEL(msg[89]), .F(
        \b/n5428 ) );
  MUX \b/U5528  ( .IN0(\b/n349 ), .IN1(\b/n5090 ), .SEL(msg[89]), .F(\b/n5436 ) );
  MUX \b/U5527  ( .IN0(msg[91]), .IN1(\b/n343 ), .SEL(msg[89]), .F(\b/n5435 )
         );
  MUX \b/U5526  ( .IN0(\b/n5093 ), .IN1(\b/n349 ), .SEL(msg[89]), .F(\b/n5434 ) );
  MUX \b/U5525  ( .IN0(msg[92]), .IN1(\b/n5090 ), .SEL(msg[89]), .F(\b/n5433 )
         );
  MUX \b/U5524  ( .IN0(\b/n334 ), .IN1(\b/n313 ), .SEL(msg[93]), .F(\b/n5140 )
         );
  MUX \b/U5523  ( .IN0(\b/n5085 ), .IN1(\b/n307 ), .SEL(msg[89]), .F(\b/n5432 ) );
  NANDN \b/U5520  ( .B(\b/n5091 ), .A(msg[95]), .Z(\b/n5405 ) );
  NAND \b/U5519  ( .A(msg[95]), .B(\b/n310 ), .Z(\b/n5373 ) );
  NAND \b/U5518  ( .A(msg[95]), .B(\b/n322 ), .Z(\b/n5314 ) );
  NAND \b/U5517  ( .A(msg[95]), .B(\b/n5422 ), .Z(\b/n5347 ) );
  NAND \b/U5516  ( .A(msg[95]), .B(\b/n5342 ), .Z(\b/n5305 ) );
  NAND \b/U5514  ( .A(\b/n354 ), .B(\b/n343 ), .Z(\b/n5426 ) );
  NAND \b/U5513  ( .A(msg[95]), .B(\b/n5424 ), .Z(\b/n5419 ) );
  NAND \b/U5512  ( .A(n696), .B(msg[95]), .Z(\b/n5399 ) );
  NAND \b/U5510  ( .A(msg[90]), .B(\b/n5093 ), .Z(\b/n5259 ) );
  NAND \b/U5509  ( .A(\b/n343 ), .B(msg[89]), .Z(\b/n5214 ) );
  NAND \b/U5508  ( .A(msg[95]), .B(\b/n5428 ), .Z(\b/n5213 ) );
  NAND \b/U5506  ( .A(\b/n5426 ), .B(msg[95]), .Z(\b/n5229 ) );
  NAND \b/U5505  ( .A(\b/n5247 ), .B(\b/n5093 ), .Z(\b/n5425 ) );
  NANDN \b/U5504  ( .B(\b/n297 ), .A(\b/n354 ), .Z(\b/n5424 ) );
  NAND \b/U5502  ( .A(msg[89]), .B(\b/n5093 ), .Z(\b/n5145 ) );
  NAND \b/U5501  ( .A(\b/n297 ), .B(\b/n354 ), .Z(\b/n5422 ) );
  NAND \b/U5498  ( .A(msg[89]), .B(\b/n5088 ), .Z(\b/n5247 ) );
  ANDN \b/U5496  ( .A(msg[90]), .B(msg[89]), .Z(\b/n5275 ) );
  AND \b/U5495  ( .A(\b/n5085 ), .B(\b/n5419 ), .Z(\b/n5190 ) );
  MUX \b/U5494  ( .IN0(\b/n5418 ), .IN1(\b/n5402 ), .SEL(msg[94]), .F(
        shift_row_out[127]) );
  MUX \b/U5493  ( .IN0(\b/n5417 ), .IN1(\b/n5410 ), .SEL(msg[88]), .F(
        \b/n5418 ) );
  MUX \b/U5492  ( .IN0(\b/n5416 ), .IN1(\b/n5413 ), .SEL(msg[93]), .F(
        \b/n5417 ) );
  MUX \b/U5491  ( .IN0(\b/n5415 ), .IN1(\b/n5414 ), .SEL(msg[90]), .F(
        \b/n5416 ) );
  MUX \b/U5490  ( .IN0(msg[92]), .IN1(\b/n314 ), .SEL(msg[95]), .F(\b/n5415 )
         );
  MUX \b/U5489  ( .IN0(\b/n5086 ), .IN1(\b/n318 ), .SEL(msg[95]), .F(\b/n5414 ) );
  MUX \b/U5488  ( .IN0(\b/n5412 ), .IN1(\b/n5411 ), .SEL(msg[90]), .F(
        \b/n5413 ) );
  MUX \b/U5487  ( .IN0(\b/n5144 ), .IN1(\b/n310 ), .SEL(msg[95]), .F(\b/n5412 ) );
  MUX \b/U5486  ( .IN0(\b/n5096 ), .IN1(\b/n5107 ), .SEL(msg[95]), .F(
        \b/n5411 ) );
  MUX \b/U5485  ( .IN0(\b/n5409 ), .IN1(\b/n5406 ), .SEL(msg[93]), .F(
        \b/n5410 ) );
  MUX \b/U5484  ( .IN0(\b/n5408 ), .IN1(\b/n5407 ), .SEL(msg[90]), .F(
        \b/n5409 ) );
  MUX \b/U5483  ( .IN0(\b/n5120 ), .IN1(\b/n5095 ), .SEL(msg[95]), .F(
        \b/n5408 ) );
  MUX \b/U5482  ( .IN0(\b/n322 ), .IN1(\b/n5116 ), .SEL(msg[95]), .F(\b/n5407 ) );
  MUX \b/U5481  ( .IN0(\b/n5404 ), .IN1(\b/n5403 ), .SEL(msg[90]), .F(
        \b/n5406 ) );
  AND \b/U5480  ( .A(\b/n312 ), .B(\b/n5405 ), .Z(\b/n5404 ) );
  MUX \b/U5479  ( .IN0(\b/n5100 ), .IN1(n695), .SEL(msg[95]), .F(\b/n5403 ) );
  MUX \b/U5478  ( .IN0(\b/n5401 ), .IN1(\b/n5393 ), .SEL(msg[88]), .F(
        \b/n5402 ) );
  MUX \b/U5477  ( .IN0(\b/n5400 ), .IN1(\b/n5396 ), .SEL(msg[93]), .F(
        \b/n5401 ) );
  MUX \b/U5476  ( .IN0(\b/n5397 ), .IN1(\b/n5398 ), .SEL(msg[90]), .F(
        \b/n5400 ) );
  NAND \b/U5475  ( .A(\b/n5214 ), .B(\b/n5399 ), .Z(\b/n5398 ) );
  MUX \b/U5474  ( .IN0(\b/n352 ), .IN1(\b/n344 ), .SEL(msg[95]), .F(\b/n5397 )
         );
  MUX \b/U5473  ( .IN0(\b/n5395 ), .IN1(\b/n5394 ), .SEL(msg[90]), .F(
        \b/n5396 ) );
  MUX \b/U5472  ( .IN0(\b/n5090 ), .IN1(\b/n5084 ), .SEL(msg[95]), .F(
        \b/n5395 ) );
  MUX \b/U5471  ( .IN0(\b/n345 ), .IN1(\b/n5121 ), .SEL(msg[95]), .F(\b/n5394 ) );
  MUX \b/U5470  ( .IN0(\b/n5392 ), .IN1(\b/n5389 ), .SEL(msg[93]), .F(
        \b/n5393 ) );
  MUX \b/U5469  ( .IN0(\b/n5391 ), .IN1(\b/n5390 ), .SEL(msg[90]), .F(
        \b/n5392 ) );
  MUX \b/U5468  ( .IN0(\b/n5125 ), .IN1(\b/n5111 ), .SEL(msg[95]), .F(
        \b/n5391 ) );
  MUX \b/U5467  ( .IN0(\b/n298 ), .IN1(\b/n5093 ), .SEL(msg[95]), .F(\b/n5390 ) );
  MUX \b/U5466  ( .IN0(\b/n5388 ), .IN1(\b/n5387 ), .SEL(msg[90]), .F(
        \b/n5389 ) );
  MUX \b/U5465  ( .IN0(\b/n5126 ), .IN1(\b/n5134 ), .SEL(msg[95]), .F(
        \b/n5388 ) );
  MUX \b/U5464  ( .IN0(\b/n5119 ), .IN1(\b/n5386 ), .SEL(msg[95]), .F(
        \b/n5387 ) );
  MUX \b/U5463  ( .IN0(\b/n349 ), .IN1(\b/n307 ), .SEL(msg[89]), .F(\b/n5386 )
         );
  MUX \b/U5462  ( .IN0(\b/n5385 ), .IN1(\b/n5367 ), .SEL(msg[94]), .F(
        shift_row_out[126]) );
  MUX \b/U5461  ( .IN0(\b/n5384 ), .IN1(\b/n5375 ), .SEL(msg[88]), .F(
        \b/n5385 ) );
  MUX \b/U5460  ( .IN0(\b/n5383 ), .IN1(\b/n5378 ), .SEL(msg[93]), .F(
        \b/n5384 ) );
  MUX \b/U5459  ( .IN0(\b/n5382 ), .IN1(\b/n5380 ), .SEL(msg[90]), .F(
        \b/n5383 ) );
  MUX \b/U5458  ( .IN0(\b/n5381 ), .IN1(\b/n5097 ), .SEL(msg[95]), .F(
        \b/n5382 ) );
  MUX \b/U5457  ( .IN0(\b/n349 ), .IN1(\b/n5084 ), .SEL(msg[89]), .F(\b/n5381 ) );
  MUX \b/U5456  ( .IN0(\b/n5379 ), .IN1(\b/n337 ), .SEL(msg[95]), .F(\b/n5380 ) );
  MUX \b/U5455  ( .IN0(\b/n5084 ), .IN1(\b/n5085 ), .SEL(msg[89]), .F(
        \b/n5379 ) );
  MUX \b/U5454  ( .IN0(\b/n5377 ), .IN1(\b/n5376 ), .SEL(msg[90]), .F(
        \b/n5378 ) );
  MUX \b/U5453  ( .IN0(n694), .IN1(\b/n5165 ), .SEL(msg[95]), .F(\b/n5377 ) );
  MUX \b/U5452  ( .IN0(\b/n5123 ), .IN1(\b/n5130 ), .SEL(msg[95]), .F(
        \b/n5376 ) );
  MUX \b/U5451  ( .IN0(\b/n5374 ), .IN1(\b/n5370 ), .SEL(msg[93]), .F(
        \b/n5375 ) );
  MUX \b/U5450  ( .IN0(\b/n5372 ), .IN1(\b/n5371 ), .SEL(msg[90]), .F(
        \b/n5374 ) );
  AND \b/U5449  ( .A(\b/n290 ), .B(\b/n5373 ), .Z(\b/n5372 ) );
  MUX \b/U5448  ( .IN0(\b/n5200 ), .IN1(msg[91]), .SEL(msg[95]), .F(\b/n5371 )
         );
  MUX \b/U5447  ( .IN0(\b/n5369 ), .IN1(\b/n5368 ), .SEL(msg[90]), .F(
        \b/n5370 ) );
  MUX \b/U5446  ( .IN0(\b/n333 ), .IN1(\b/n5088 ), .SEL(msg[95]), .F(\b/n5369 ) );
  MUX \b/U5444  ( .IN0(\b/n5366 ), .IN1(\b/n5359 ), .SEL(msg[88]), .F(
        \b/n5367 ) );
  MUX \b/U5443  ( .IN0(\b/n5365 ), .IN1(\b/n5362 ), .SEL(msg[93]), .F(
        \b/n5366 ) );
  MUX \b/U5442  ( .IN0(\b/n5364 ), .IN1(\b/n5363 ), .SEL(msg[90]), .F(
        \b/n5365 ) );
  MUX \b/U5441  ( .IN0(\b/n329 ), .IN1(\b/n5092 ), .SEL(msg[95]), .F(\b/n5364 ) );
  MUX \b/U5440  ( .IN0(\b/n5096 ), .IN1(n695), .SEL(msg[95]), .F(\b/n5363 ) );
  MUX \b/U5439  ( .IN0(\b/n5361 ), .IN1(\b/n5360 ), .SEL(msg[90]), .F(
        \b/n5362 ) );
  MUX \b/U5438  ( .IN0(\b/n5112 ), .IN1(\b/n294 ), .SEL(msg[95]), .F(\b/n5361 ) );
  MUX \b/U5437  ( .IN0(\b/n314 ), .IN1(\b/n344 ), .SEL(msg[95]), .F(\b/n5360 )
         );
  MUX \b/U5436  ( .IN0(\b/n5358 ), .IN1(\b/n5354 ), .SEL(msg[93]), .F(
        \b/n5359 ) );
  MUX \b/U5435  ( .IN0(\b/n5357 ), .IN1(\b/n5356 ), .SEL(msg[90]), .F(
        \b/n5358 ) );
  MUX \b/U5434  ( .IN0(\b/n5101 ), .IN1(\b/n344 ), .SEL(msg[95]), .F(\b/n5357 ) );
  MUX \b/U5433  ( .IN0(\b/n5355 ), .IN1(\b/n5122 ), .SEL(msg[95]), .F(
        \b/n5356 ) );
  NANDN \b/U5432  ( .B(msg[92]), .A(msg[89]), .Z(\b/n5355 ) );
  MUX \b/U5431  ( .IN0(\b/n5353 ), .IN1(\b/n5351 ), .SEL(msg[90]), .F(
        \b/n5354 ) );
  MUX \b/U5430  ( .IN0(\b/n307 ), .IN1(\b/n5352 ), .SEL(msg[95]), .F(\b/n5353 ) );
  MUX \b/U5429  ( .IN0(\b/n334 ), .IN1(\b/n324 ), .SEL(msg[89]), .F(\b/n5352 )
         );
  MUX \b/U5428  ( .IN0(\b/n296 ), .IN1(\b/n5097 ), .SEL(msg[95]), .F(\b/n5351 ) );
  NANDN \b/U5427  ( .B(\b/n297 ), .A(msg[89]), .Z(\b/n5097 ) );
  MUX \b/U5426  ( .IN0(\b/n5350 ), .IN1(\b/n5329 ), .SEL(msg[94]), .F(
        shift_row_out[125]) );
  MUX \b/U5425  ( .IN0(\b/n5349 ), .IN1(\b/n5339 ), .SEL(msg[88]), .F(
        \b/n5350 ) );
  MUX \b/U5424  ( .IN0(\b/n5348 ), .IN1(\b/n5344 ), .SEL(msg[93]), .F(
        \b/n5349 ) );
  MUX \b/U5423  ( .IN0(\b/n5345 ), .IN1(\b/n5346 ), .SEL(msg[90]), .F(
        \b/n5348 ) );
  AND \b/U5422  ( .A(\b/n5115 ), .B(\b/n5347 ), .Z(\b/n5346 ) );
  MUX \b/U5421  ( .IN0(\b/n5093 ), .IN1(\b/n345 ), .SEL(msg[95]), .F(\b/n5345 ) );
  MUX \b/U5420  ( .IN0(\b/n5343 ), .IN1(\b/n5341 ), .SEL(msg[90]), .F(
        \b/n5344 ) );
  MUX \b/U5419  ( .IN0(\b/n300 ), .IN1(\b/n5342 ), .SEL(msg[95]), .F(\b/n5343 ) );
  NAND \b/U5418  ( .A(\b/n324 ), .B(\b/n354 ), .Z(\b/n5342 ) );
  MUX \b/U5417  ( .IN0(\b/n5093 ), .IN1(\b/n5340 ), .SEL(msg[95]), .F(
        \b/n5341 ) );
  NAND \b/U5416  ( .A(\b/n5084 ), .B(\b/n5145 ), .Z(\b/n5340 ) );
  MUX \b/U5415  ( .IN0(\b/n5338 ), .IN1(\b/n5334 ), .SEL(msg[93]), .F(
        \b/n5339 ) );
  MUX \b/U5414  ( .IN0(\b/n5337 ), .IN1(\b/n5336 ), .SEL(msg[90]), .F(
        \b/n5338 ) );
  MUX \b/U5413  ( .IN0(\b/n5105 ), .IN1(\b/n347 ), .SEL(msg[95]), .F(\b/n5337 ) );
  MUX \b/U5412  ( .IN0(\b/n5130 ), .IN1(\b/n5335 ), .SEL(msg[95]), .F(
        \b/n5336 ) );
  MUX \b/U5411  ( .IN0(\b/n343 ), .IN1(\b/n324 ), .SEL(msg[89]), .F(\b/n5335 )
         );
  MUX \b/U5410  ( .IN0(\b/n5333 ), .IN1(\b/n5332 ), .SEL(msg[90]), .F(
        \b/n5334 ) );
  MUX \b/U5409  ( .IN0(\b/n341 ), .IN1(n693), .SEL(msg[95]), .F(\b/n5333 ) );
  MUX \b/U5408  ( .IN0(\b/n5331 ), .IN1(\b/n5330 ), .SEL(msg[95]), .F(
        \b/n5332 ) );
  AND \b/U5407  ( .A(\b/n5090 ), .B(\b/n5165 ), .Z(\b/n5331 ) );
  MUX \b/U5406  ( .IN0(\b/n313 ), .IN1(\b/n297 ), .SEL(msg[89]), .F(\b/n5330 )
         );
  MUX \b/U5405  ( .IN0(\b/n5328 ), .IN1(\b/n5319 ), .SEL(msg[88]), .F(
        \b/n5329 ) );
  MUX \b/U5404  ( .IN0(\b/n5327 ), .IN1(\b/n5323 ), .SEL(msg[93]), .F(
        \b/n5328 ) );
  MUX \b/U5403  ( .IN0(\b/n5326 ), .IN1(\b/n5324 ), .SEL(msg[90]), .F(
        \b/n5327 ) );
  MUX \b/U5402  ( .IN0(\b/n5096 ), .IN1(\b/n5325 ), .SEL(msg[95]), .F(
        \b/n5326 ) );
  NAND \b/U5401  ( .A(msg[89]), .B(\b/n313 ), .Z(\b/n5325 ) );
  MUX \b/U5400  ( .IN0(\b/n297 ), .IN1(\b/n350 ), .SEL(msg[95]), .F(\b/n5324 )
         );
  MUX \b/U5399  ( .IN0(\b/n5322 ), .IN1(\b/n5321 ), .SEL(msg[90]), .F(
        \b/n5323 ) );
  MUX \b/U5398  ( .IN0(\b/n5122 ), .IN1(\b/n315 ), .SEL(msg[95]), .F(\b/n5322 ) );
  MUX \b/U5397  ( .IN0(\b/n5320 ), .IN1(\b/n5085 ), .SEL(n692), .F(\b/n5321 )
         );
  AND \b/U5396  ( .A(msg[95]), .B(msg[91]), .Z(\b/n5320 ) );
  MUX \b/U5395  ( .IN0(\b/n5318 ), .IN1(\b/n5315 ), .SEL(msg[93]), .F(
        \b/n5319 ) );
  MUX \b/U5394  ( .IN0(\b/n5317 ), .IN1(\b/n5316 ), .SEL(msg[90]), .F(
        \b/n5318 ) );
  MUX \b/U5393  ( .IN0(\b/n5246 ), .IN1(\b/n5085 ), .SEL(msg[95]), .F(
        \b/n5317 ) );
  MUX \b/U5392  ( .IN0(n691), .IN1(\b/n348 ), .SEL(msg[95]), .F(\b/n5316 ) );
  MUX \b/U5391  ( .IN0(\b/n5313 ), .IN1(\b/n5312 ), .SEL(msg[90]), .F(
        \b/n5315 ) );
  AND \b/U5390  ( .A(\b/n5314 ), .B(\b/n5214 ), .Z(\b/n5313 ) );
  MUX \b/U5389  ( .IN0(\b/n299 ), .IN1(\b/n343 ), .SEL(msg[95]), .F(\b/n5312 )
         );
  MUX \b/U5388  ( .IN0(\b/n5311 ), .IN1(\b/n5294 ), .SEL(msg[94]), .F(
        shift_row_out[124]) );
  MUX \b/U5387  ( .IN0(\b/n5310 ), .IN1(\b/n5302 ), .SEL(msg[88]), .F(
        \b/n5311 ) );
  MUX \b/U5386  ( .IN0(\b/n5309 ), .IN1(\b/n5306 ), .SEL(msg[93]), .F(
        \b/n5310 ) );
  MUX \b/U5385  ( .IN0(\b/n5308 ), .IN1(\b/n5307 ), .SEL(msg[90]), .F(
        \b/n5309 ) );
  MUX \b/U5384  ( .IN0(\b/n325 ), .IN1(\b/n346 ), .SEL(msg[95]), .F(\b/n5308 )
         );
  MUX \b/U5383  ( .IN0(\b/n5165 ), .IN1(\b/n5130 ), .SEL(msg[95]), .F(
        \b/n5307 ) );
  NAND \b/U5382  ( .A(msg[89]), .B(\b/n5084 ), .Z(\b/n5165 ) );
  MUX \b/U5381  ( .IN0(\b/n5303 ), .IN1(\b/n5304 ), .SEL(msg[90]), .F(
        \b/n5306 ) );
  AND \b/U5380  ( .A(\b/n5115 ), .B(\b/n5305 ), .Z(\b/n5304 ) );
  MUX \b/U5379  ( .IN0(\b/n5113 ), .IN1(\b/n328 ), .SEL(msg[95]), .F(\b/n5303 ) );
  MUX \b/U5378  ( .IN0(\b/n5301 ), .IN1(\b/n5298 ), .SEL(msg[93]), .F(
        \b/n5302 ) );
  MUX \b/U5377  ( .IN0(\b/n5300 ), .IN1(\b/n5299 ), .SEL(msg[90]), .F(
        \b/n5301 ) );
  MUX \b/U5376  ( .IN0(\b/n290 ), .IN1(\b/n336 ), .SEL(msg[95]), .F(\b/n5300 )
         );
  MUX \b/U5375  ( .IN0(\b/n297 ), .IN1(\b/n5093 ), .SEL(msg[95]), .F(\b/n5299 ) );
  MUX \b/U5374  ( .IN0(\b/n5297 ), .IN1(\b/n5295 ), .SEL(msg[90]), .F(
        \b/n5298 ) );
  MUX \b/U5373  ( .IN0(\b/n5109 ), .IN1(\b/n5296 ), .SEL(msg[95]), .F(
        \b/n5297 ) );
  AND \b/U5372  ( .A(\b/n5093 ), .B(\b/n354 ), .Z(\b/n5296 ) );
  MUX \b/U5371  ( .IN0(\b/n312 ), .IN1(\b/n331 ), .SEL(msg[95]), .F(\b/n5295 )
         );
  MUX \b/U5370  ( .IN0(\b/n5293 ), .IN1(\b/n5287 ), .SEL(msg[88]), .F(
        \b/n5294 ) );
  MUX \b/U5369  ( .IN0(\b/n5292 ), .IN1(\b/n5290 ), .SEL(msg[93]), .F(
        \b/n5293 ) );
  MUX \b/U5368  ( .IN0(\b/n5291 ), .IN1(\b/n5087 ), .SEL(msg[90]), .F(
        \b/n5292 ) );
  MUX \b/U5367  ( .IN0(\b/n5107 ), .IN1(\b/n333 ), .SEL(msg[95]), .F(\b/n5291 ) );
  MUX \b/U5366  ( .IN0(\b/n5289 ), .IN1(\b/n5288 ), .SEL(msg[90]), .F(
        \b/n5290 ) );
  MUX \b/U5365  ( .IN0(n690), .IN1(\b/n325 ), .SEL(msg[95]), .F(\b/n5289 ) );
  MUX \b/U5364  ( .IN0(\b/n5117 ), .IN1(\b/n5120 ), .SEL(msg[95]), .F(
        \b/n5288 ) );
  MUX \b/U5363  ( .IN0(\b/n5286 ), .IN1(\b/n5283 ), .SEL(msg[93]), .F(
        \b/n5287 ) );
  MUX \b/U5362  ( .IN0(\b/n5285 ), .IN1(\b/n5284 ), .SEL(msg[90]), .F(
        \b/n5286 ) );
  MUX \b/U5361  ( .IN0(\b/n298 ), .IN1(\b/n5089 ), .SEL(msg[95]), .F(\b/n5285 ) );
  MUX \b/U5360  ( .IN0(\b/n343 ), .IN1(\b/n5111 ), .SEL(msg[95]), .F(\b/n5284 ) );
  MUX \b/U5359  ( .IN0(\b/n286 ), .IN1(\b/n5282 ), .SEL(msg[90]), .F(\b/n5283 ) );
  MUX \b/U5358  ( .IN0(\b/n306 ), .IN1(\b/n5093 ), .SEL(msg[95]), .F(\b/n5282 ) );
  MUX \b/U5357  ( .IN0(\b/n5281 ), .IN1(\b/n5262 ), .SEL(msg[94]), .F(
        shift_row_out[123]) );
  MUX \b/U5356  ( .IN0(\b/n5280 ), .IN1(\b/n5272 ), .SEL(msg[88]), .F(
        \b/n5281 ) );
  MUX \b/U5355  ( .IN0(\b/n5279 ), .IN1(\b/n5276 ), .SEL(msg[93]), .F(
        \b/n5280 ) );
  MUX \b/U5354  ( .IN0(\b/n5278 ), .IN1(\b/n5277 ), .SEL(msg[95]), .F(
        \b/n5279 ) );
  MUX \b/U5353  ( .IN0(\b/n5101 ), .IN1(\b/n331 ), .SEL(msg[90]), .F(\b/n5278 ) );
  MUX \b/U5352  ( .IN0(n693), .IN1(\b/n289 ), .SEL(msg[90]), .F(\b/n5277 ) );
  MUX \b/U5351  ( .IN0(\b/n5274 ), .IN1(\b/n5273 ), .SEL(msg[95]), .F(
        \b/n5276 ) );
  AND \b/U5350  ( .A(\b/n5275 ), .B(msg[92]), .Z(\b/n5274 ) );
  MUX \b/U5349  ( .IN0(\b/n319 ), .IN1(\b/n5114 ), .SEL(msg[90]), .F(\b/n5273 ) );
  MUX \b/U5348  ( .IN0(\b/n5271 ), .IN1(\b/n5268 ), .SEL(msg[93]), .F(
        \b/n5272 ) );
  MUX \b/U5347  ( .IN0(\b/n5270 ), .IN1(\b/n5269 ), .SEL(msg[95]), .F(
        \b/n5271 ) );
  MUX \b/U5346  ( .IN0(\b/n5105 ), .IN1(n689), .SEL(msg[90]), .F(\b/n5270 ) );
  MUX \b/U5345  ( .IN0(\b/n287 ), .IN1(\b/n306 ), .SEL(msg[90]), .F(\b/n5269 )
         );
  MUX \b/U5344  ( .IN0(\b/n5264 ), .IN1(\b/n5265 ), .SEL(msg[95]), .F(
        \b/n5268 ) );
  NAND \b/U5343  ( .A(\b/n5266 ), .B(\b/n5267 ), .Z(\b/n5265 ) );
  MUX \b/U5342  ( .IN0(\b/n332 ), .IN1(\b/n5263 ), .SEL(msg[90]), .F(\b/n5264 ) );
  MUX \b/U5341  ( .IN0(\b/n307 ), .IN1(\b/n349 ), .SEL(msg[89]), .F(\b/n5263 )
         );
  MUX \b/U5340  ( .IN0(\b/n5261 ), .IN1(\b/n5252 ), .SEL(msg[88]), .F(
        \b/n5262 ) );
  MUX \b/U5339  ( .IN0(\b/n5260 ), .IN1(\b/n5256 ), .SEL(msg[93]), .F(
        \b/n5261 ) );
  MUX \b/U5338  ( .IN0(\b/n5258 ), .IN1(\b/n5257 ), .SEL(msg[95]), .F(
        \b/n5260 ) );
  NAND \b/U5337  ( .A(\b/n297 ), .B(\b/n5259 ), .Z(\b/n5258 ) );
  MUX \b/U5336  ( .IN0(\b/n348 ), .IN1(\b/n310 ), .SEL(msg[90]), .F(\b/n5257 )
         );
  MUX \b/U5335  ( .IN0(\b/n5255 ), .IN1(\b/n5253 ), .SEL(msg[95]), .F(
        \b/n5256 ) );
  MUX \b/U5334  ( .IN0(\b/n5096 ), .IN1(\b/n5254 ), .SEL(msg[90]), .F(
        \b/n5255 ) );
  AND \b/U5333  ( .A(msg[89]), .B(\b/n297 ), .Z(\b/n5254 ) );
  MUX \b/U5332  ( .IN0(\b/n302 ), .IN1(\b/n5115 ), .SEL(msg[90]), .F(\b/n5253 ) );
  MUX \b/U5331  ( .IN0(\b/n5251 ), .IN1(\b/n5245 ), .SEL(msg[93]), .F(
        \b/n5252 ) );
  MUX \b/U5330  ( .IN0(\b/n5250 ), .IN1(\b/n5248 ), .SEL(msg[95]), .F(
        \b/n5251 ) );
  MUX \b/U5329  ( .IN0(\b/n5249 ), .IN1(\b/n5085 ), .SEL(\b/n5133 ), .F(
        \b/n5250 ) );
  MUX \b/U5328  ( .IN0(msg[91]), .IN1(msg[92]), .SEL(msg[90]), .F(\b/n5249 )
         );
  MUX \b/U5327  ( .IN0(\b/n5115 ), .IN1(\b/n5246 ), .SEL(msg[90]), .F(
        \b/n5248 ) );
  NAND \b/U5326  ( .A(\b/n5085 ), .B(\b/n5247 ), .Z(\b/n5246 ) );
  MUX \b/U5325  ( .IN0(\b/n5242 ), .IN1(\b/n5243 ), .SEL(msg[95]), .F(
        \b/n5245 ) );
  AND \b/U5324  ( .A(\b/n330 ), .B(\b/n5244 ), .Z(\b/n5243 ) );
  MUX \b/U5323  ( .IN0(\b/n311 ), .IN1(\b/n5086 ), .SEL(msg[90]), .F(\b/n5242 ) );
  MUX \b/U5322  ( .IN0(\b/n5241 ), .IN1(\b/n5225 ), .SEL(msg[94]), .F(
        shift_row_out[122]) );
  MUX \b/U5321  ( .IN0(\b/n5240 ), .IN1(\b/n5232 ), .SEL(msg[88]), .F(
        \b/n5241 ) );
  MUX \b/U5320  ( .IN0(\b/n5239 ), .IN1(\b/n5235 ), .SEL(msg[93]), .F(
        \b/n5240 ) );
  MUX \b/U5319  ( .IN0(\b/n5238 ), .IN1(\b/n5236 ), .SEL(msg[90]), .F(
        \b/n5239 ) );
  MUX \b/U5318  ( .IN0(\b/n319 ), .IN1(\b/n5237 ), .SEL(msg[95]), .F(\b/n5238 ) );
  MUX \b/U5317  ( .IN0(\b/n5093 ), .IN1(\b/n297 ), .SEL(msg[89]), .F(\b/n5237 ) );
  MUX \b/U5316  ( .IN0(\b/n5132 ), .IN1(\b/n337 ), .SEL(msg[95]), .F(\b/n5236 ) );
  MUX \b/U5315  ( .IN0(\b/n5234 ), .IN1(\b/n5233 ), .SEL(msg[90]), .F(
        \b/n5235 ) );
  MUX \b/U5314  ( .IN0(\b/n5086 ), .IN1(\b/n304 ), .SEL(msg[95]), .F(\b/n5234 ) );
  MUX \b/U5313  ( .IN0(\b/n340 ), .IN1(\b/n5119 ), .SEL(msg[95]), .F(\b/n5233 ) );
  MUX \b/U5312  ( .IN0(\b/n5231 ), .IN1(\b/n5227 ), .SEL(msg[93]), .F(
        \b/n5232 ) );
  MUX \b/U5311  ( .IN0(\b/n5228 ), .IN1(\b/n286 ), .SEL(msg[90]), .F(\b/n5231 ) );
  NAND \b/U5310  ( .A(\b/n5229 ), .B(\b/n5230 ), .Z(\b/n5228 ) );
  MUX \b/U5309  ( .IN0(n691), .IN1(\b/n5226 ), .SEL(\b/n5131 ), .F(\b/n5227 )
         );
  MUX \b/U5308  ( .IN0(\b/n318 ), .IN1(\b/n5098 ), .SEL(msg[90]), .F(\b/n5226 ) );
  MUX \b/U5307  ( .IN0(\b/n5224 ), .IN1(\b/n5216 ), .SEL(msg[88]), .F(
        \b/n5225 ) );
  MUX \b/U5306  ( .IN0(\b/n5223 ), .IN1(\b/n5220 ), .SEL(msg[93]), .F(
        \b/n5224 ) );
  MUX \b/U5305  ( .IN0(\b/n5222 ), .IN1(\b/n5221 ), .SEL(msg[90]), .F(
        \b/n5223 ) );
  MUX \b/U5304  ( .IN0(\b/n346 ), .IN1(msg[89]), .SEL(msg[95]), .F(\b/n5222 )
         );
  MUX \b/U5303  ( .IN0(n694), .IN1(\b/n5099 ), .SEL(msg[95]), .F(\b/n5221 ) );
  MUX \b/U5302  ( .IN0(\b/n5219 ), .IN1(\b/n5218 ), .SEL(msg[90]), .F(
        \b/n5220 ) );
  MUX \b/U5301  ( .IN0(\b/n351 ), .IN1(\b/n345 ), .SEL(msg[95]), .F(\b/n5219 )
         );
  MUX \b/U5300  ( .IN0(n694), .IN1(\b/n5217 ), .SEL(msg[95]), .F(\b/n5218 ) );
  MUX \b/U5299  ( .IN0(\b/n297 ), .IN1(\b/n334 ), .SEL(msg[89]), .F(\b/n5217 )
         );
  MUX \b/U5298  ( .IN0(\b/n5215 ), .IN1(\b/n5209 ), .SEL(msg[93]), .F(
        \b/n5216 ) );
  MUX \b/U5297  ( .IN0(\b/n5212 ), .IN1(\b/n5211 ), .SEL(msg[90]), .F(
        \b/n5215 ) );
  NAND \b/U5296  ( .A(\b/n5213 ), .B(\b/n5214 ), .Z(\b/n5212 ) );
  MUX \b/U5295  ( .IN0(\b/n5085 ), .IN1(\b/n5210 ), .SEL(n692), .F(\b/n5211 )
         );
  MUX \b/U5294  ( .IN0(msg[91]), .IN1(\b/n307 ), .SEL(msg[95]), .F(\b/n5210 )
         );
  MUX \b/U5293  ( .IN0(\b/n5208 ), .IN1(\b/n5207 ), .SEL(msg[90]), .F(
        \b/n5209 ) );
  MUX \b/U5292  ( .IN0(\b/n5130 ), .IN1(\b/n305 ), .SEL(msg[95]), .F(\b/n5208 ) );
  MUX \b/U5291  ( .IN0(\b/n5126 ), .IN1(\b/n5206 ), .SEL(msg[95]), .F(
        \b/n5207 ) );
  MUX \b/U5290  ( .IN0(\b/n5088 ), .IN1(\b/n5093 ), .SEL(msg[89]), .F(
        \b/n5206 ) );
  MUX \b/U5289  ( .IN0(\b/n5205 ), .IN1(\b/n5187 ), .SEL(msg[94]), .F(
        shift_row_out[121]) );
  MUX \b/U5288  ( .IN0(\b/n5204 ), .IN1(\b/n5195 ), .SEL(msg[88]), .F(
        \b/n5205 ) );
  MUX \b/U5287  ( .IN0(\b/n5203 ), .IN1(\b/n5199 ), .SEL(msg[93]), .F(
        \b/n5204 ) );
  MUX \b/U5286  ( .IN0(\b/n5202 ), .IN1(\b/n5201 ), .SEL(msg[90]), .F(
        \b/n5203 ) );
  MUX \b/U5285  ( .IN0(\b/n342 ), .IN1(n696), .SEL(msg[95]), .F(\b/n5202 ) );
  MUX \b/U5284  ( .IN0(\b/n5200 ), .IN1(n690), .SEL(msg[95]), .F(\b/n5201 ) );
  NAND \b/U5283  ( .A(\b/n354 ), .B(\b/n313 ), .Z(\b/n5200 ) );
  MUX \b/U5282  ( .IN0(\b/n5198 ), .IN1(\b/n5197 ), .SEL(msg[90]), .F(
        \b/n5199 ) );
  MUX \b/U5281  ( .IN0(\b/n290 ), .IN1(\b/n5100 ), .SEL(msg[95]), .F(\b/n5198 ) );
  MUX \b/U5280  ( .IN0(\b/n5090 ), .IN1(\b/n5196 ), .SEL(msg[95]), .F(
        \b/n5197 ) );
  AND \b/U5279  ( .A(msg[89]), .B(msg[92]), .Z(\b/n5196 ) );
  MUX \b/U5278  ( .IN0(\b/n5194 ), .IN1(\b/n5191 ), .SEL(msg[93]), .F(
        \b/n5195 ) );
  MUX \b/U5277  ( .IN0(\b/n5193 ), .IN1(\b/n5192 ), .SEL(msg[90]), .F(
        \b/n5194 ) );
  MUX \b/U5276  ( .IN0(\b/n5129 ), .IN1(\b/n351 ), .SEL(msg[95]), .F(\b/n5193 ) );
  MUX \b/U5275  ( .IN0(\b/n326 ), .IN1(\b/n5098 ), .SEL(msg[95]), .F(\b/n5192 ) );
  MUX \b/U5274  ( .IN0(\b/n5188 ), .IN1(\b/n5189 ), .SEL(msg[90]), .F(
        \b/n5191 ) );
  AND \b/U5273  ( .A(\b/n5190 ), .B(\b/n5145 ), .Z(\b/n5189 ) );
  MUX \b/U5272  ( .IN0(\b/n5104 ), .IN1(\b/n5093 ), .SEL(msg[95]), .F(
        \b/n5188 ) );
  MUX \b/U5271  ( .IN0(\b/n5186 ), .IN1(\b/n5178 ), .SEL(msg[88]), .F(
        \b/n5187 ) );
  MUX \b/U5270  ( .IN0(\b/n5185 ), .IN1(\b/n5181 ), .SEL(msg[93]), .F(
        \b/n5186 ) );
  MUX \b/U5269  ( .IN0(\b/n5184 ), .IN1(\b/n5183 ), .SEL(msg[90]), .F(
        \b/n5185 ) );
  MUX \b/U5268  ( .IN0(\b/n5092 ), .IN1(\b/n315 ), .SEL(msg[95]), .F(\b/n5184 ) );
  MUX \b/U5267  ( .IN0(\b/n5182 ), .IN1(\b/n299 ), .SEL(msg[95]), .F(\b/n5183 ) );
  MUX \b/U5266  ( .IN0(\b/n5090 ), .IN1(\b/n307 ), .SEL(msg[89]), .F(\b/n5182 ) );
  MUX \b/U5265  ( .IN0(\b/n5180 ), .IN1(\b/n5179 ), .SEL(msg[90]), .F(
        \b/n5181 ) );
  MUX \b/U5264  ( .IN0(\b/n346 ), .IN1(\b/n324 ), .SEL(msg[95]), .F(\b/n5180 )
         );
  MUX \b/U5263  ( .IN0(\b/n342 ), .IN1(\b/n302 ), .SEL(msg[95]), .F(\b/n5179 )
         );
  MUX \b/U5262  ( .IN0(\b/n5177 ), .IN1(\b/n5172 ), .SEL(msg[93]), .F(
        \b/n5178 ) );
  MUX \b/U5261  ( .IN0(\b/n5176 ), .IN1(\b/n5173 ), .SEL(msg[90]), .F(
        \b/n5177 ) );
  MUX \b/U5260  ( .IN0(\b/n5174 ), .IN1(\b/n5175 ), .SEL(msg[95]), .F(
        \b/n5176 ) );
  NAND \b/U5259  ( .A(\b/n5093 ), .B(\b/n5165 ), .Z(\b/n5175 ) );
  MUX \b/U5258  ( .IN0(\b/n5093 ), .IN1(\b/n307 ), .SEL(msg[89]), .F(\b/n5174 ) );
  MUX \b/U5257  ( .IN0(\b/n5110 ), .IN1(\b/n5108 ), .SEL(msg[95]), .F(
        \b/n5173 ) );
  MUX \b/U5256  ( .IN0(\b/n5128 ), .IN1(\b/n5171 ), .SEL(msg[90]), .F(
        \b/n5172 ) );
  MUX \b/U5255  ( .IN0(\b/n313 ), .IN1(\b/n345 ), .SEL(msg[95]), .F(\b/n5171 )
         );
  MUX \b/U5254  ( .IN0(\b/n5170 ), .IN1(\b/n5153 ), .SEL(msg[94]), .F(
        shift_row_out[120]) );
  MUX \b/U5253  ( .IN0(\b/n5169 ), .IN1(\b/n5161 ), .SEL(msg[88]), .F(
        \b/n5170 ) );
  MUX \b/U5252  ( .IN0(\b/n5168 ), .IN1(\b/n5166 ), .SEL(msg[90]), .F(
        \b/n5169 ) );
  MUX \b/U5251  ( .IN0(\b/n287 ), .IN1(\b/n5167 ), .SEL(msg[95]), .F(\b/n5168 ) );
  MUX \b/U5250  ( .IN0(\b/n340 ), .IN1(\b/n343 ), .SEL(msg[93]), .F(\b/n5167 )
         );
  MUX \b/U5249  ( .IN0(\b/n5163 ), .IN1(\b/n5162 ), .SEL(msg[95]), .F(
        \b/n5166 ) );
  NAND \b/U5248  ( .A(\b/n5164 ), .B(\b/n5165 ), .Z(\b/n5163 ) );
  MUX \b/U5247  ( .IN0(\b/n339 ), .IN1(\b/n354 ), .SEL(msg[93]), .F(\b/n5162 )
         );
  MUX \b/U5246  ( .IN0(\b/n5160 ), .IN1(\b/n5156 ), .SEL(msg[90]), .F(
        \b/n5161 ) );
  MUX \b/U5245  ( .IN0(\b/n5159 ), .IN1(\b/n5157 ), .SEL(msg[95]), .F(
        \b/n5160 ) );
  MUX \b/U5244  ( .IN0(\b/n5158 ), .IN1(\b/n292 ), .SEL(msg[93]), .F(\b/n5159 ) );
  NAND \b/U5243  ( .A(\b/n354 ), .B(\b/n5085 ), .Z(\b/n5158 ) );
  MUX \b/U5241  ( .IN0(\b/n5155 ), .IN1(\b/n5154 ), .SEL(msg[95]), .F(
        \b/n5156 ) );
  MUX \b/U5240  ( .IN0(n691), .IN1(\b/n289 ), .SEL(msg[93]), .F(\b/n5155 ) );
  MUX \b/U5239  ( .IN0(\b/n341 ), .IN1(\b/n297 ), .SEL(msg[93]), .F(\b/n5154 )
         );
  MUX \b/U5238  ( .IN0(\b/n5152 ), .IN1(\b/n5142 ), .SEL(msg[88]), .F(
        \b/n5153 ) );
  MUX \b/U5237  ( .IN0(\b/n5151 ), .IN1(\b/n5147 ), .SEL(msg[90]), .F(
        \b/n5152 ) );
  MUX \b/U5236  ( .IN0(\b/n5150 ), .IN1(\b/n5149 ), .SEL(msg[95]), .F(
        \b/n5151 ) );
  MUX \b/U5235  ( .IN0(n689), .IN1(\b/n293 ), .SEL(msg[93]), .F(\b/n5150 ) );
  MUX \b/U5234  ( .IN0(\b/n5148 ), .IN1(\b/n330 ), .SEL(msg[93]), .F(\b/n5149 ) );
  NAND \b/U5233  ( .A(\b/n5084 ), .B(\b/n5086 ), .Z(\b/n5148 ) );
  MUX \b/U5232  ( .IN0(\b/n5146 ), .IN1(\b/n5143 ), .SEL(msg[95]), .F(
        \b/n5147 ) );
  MUX \b/U5231  ( .IN0(\b/n300 ), .IN1(\b/n5144 ), .SEL(msg[93]), .F(\b/n5146 ) );
  NAND \b/U5230  ( .A(\b/n5088 ), .B(\b/n5145 ), .Z(\b/n5144 ) );
  MUX \b/U5229  ( .IN0(\b/n5103 ), .IN1(\b/n5094 ), .SEL(msg[93]), .F(
        \b/n5143 ) );
  MUX \b/U5228  ( .IN0(\b/n5141 ), .IN1(\b/n5137 ), .SEL(msg[90]), .F(
        \b/n5142 ) );
  MUX \b/U5227  ( .IN0(\b/n5139 ), .IN1(\b/n5138 ), .SEL(msg[95]), .F(
        \b/n5141 ) );
  NAND \b/U5226  ( .A(\b/n5140 ), .B(\b/n5127 ), .Z(\b/n5139 ) );
  MUX \b/U5225  ( .IN0(msg[91]), .IN1(\b/n5119 ), .SEL(msg[93]), .F(\b/n5138 )
         );
  MUX \b/U5224  ( .IN0(\b/n5136 ), .IN1(\b/n5135 ), .SEL(msg[95]), .F(
        \b/n5137 ) );
  MUX \b/U5223  ( .IN0(\b/n305 ), .IN1(\b/n321 ), .SEL(msg[93]), .F(\b/n5136 )
         );
  MUX \b/U5222  ( .IN0(\b/n338 ), .IN1(\b/n326 ), .SEL(msg[93]), .F(\b/n5135 )
         );
  XOR \b/U5221  ( .A(\b/n5085 ), .B(msg[89]), .Z(\b/n5134 ) );
  XOR \b/U5220  ( .A(msg[89]), .B(msg[90]), .Z(\b/n5133 ) );
  XOR \b/U5219  ( .A(msg[89]), .B(msg[91]), .Z(\b/n5132 ) );
  XOR \b/U5218  ( .A(msg[90]), .B(msg[95]), .Z(\b/n5131 ) );
  XOR \b/U5217  ( .A(\b/n354 ), .B(\b/n297 ), .Z(\b/n5130 ) );
  XOR \b/U5216  ( .A(msg[89]), .B(\b/n343 ), .Z(\b/n5129 ) );
  XOR \b/U5214  ( .A(msg[89]), .B(msg[93]), .Z(\b/n5127 ) );
  NAND \b/U5213  ( .A(msg[89]), .B(msg[91]), .Z(\b/n5126 ) );
  MUX \b/U5212  ( .IN0(\b/n5085 ), .IN1(\b/n297 ), .SEL(msg[89]), .F(\b/n5125 ) );
  MUX \b/U5210  ( .IN0(msg[91]), .IN1(\b/n334 ), .SEL(msg[89]), .F(\b/n5123 )
         );
  MUX \b/U5209  ( .IN0(\b/n313 ), .IN1(\b/n334 ), .SEL(msg[89]), .F(\b/n5122 )
         );
  MUX \b/U5208  ( .IN0(\b/n5088 ), .IN1(\b/n5090 ), .SEL(msg[89]), .F(
        \b/n5121 ) );
  MUX \b/U5207  ( .IN0(msg[92]), .IN1(\b/n313 ), .SEL(msg[89]), .F(\b/n5120 )
         );
  OR \b/U5206  ( .A(msg[89]), .B(msg[92]), .Z(\b/n5119 ) );
  NAND \b/U5204  ( .A(\b/n334 ), .B(\b/n354 ), .Z(\b/n5117 ) );
  MUX \b/U5203  ( .IN0(\b/n334 ), .IN1(msg[92]), .SEL(msg[89]), .F(\b/n5116 )
         );
  MUX \b/U5202  ( .IN0(\b/n5084 ), .IN1(\b/n5093 ), .SEL(msg[89]), .F(
        \b/n5115 ) );
  MUX \b/U5201  ( .IN0(\b/n349 ), .IN1(msg[92]), .SEL(msg[89]), .F(\b/n5114 )
         );
  MUX \b/U5200  ( .IN0(\b/n307 ), .IN1(\b/n334 ), .SEL(msg[89]), .F(\b/n5113 )
         );
  MUX \b/U5199  ( .IN0(\b/n5084 ), .IN1(msg[92]), .SEL(msg[89]), .F(\b/n5112 )
         );
  MUX \b/U5198  ( .IN0(\b/n324 ), .IN1(\b/n313 ), .SEL(msg[89]), .F(\b/n5111 )
         );
  XOR \b/U5197  ( .A(\b/n307 ), .B(msg[89]), .Z(\b/n5110 ) );
  MUX \b/U5196  ( .IN0(\b/n5090 ), .IN1(\b/n324 ), .SEL(msg[89]), .F(\b/n5109 ) );
  NANDN \b/U5195  ( .B(msg[89]), .A(msg[91]), .Z(\b/n5108 ) );
  MUX \b/U5194  ( .IN0(\b/n297 ), .IN1(msg[91]), .SEL(msg[89]), .F(\b/n5107 )
         );
  NAND \b/U5192  ( .A(\b/n5088 ), .B(\b/n354 ), .Z(\b/n5105 ) );
  MUX \b/U5191  ( .IN0(msg[92]), .IN1(\b/n5085 ), .SEL(msg[89]), .F(\b/n5104 )
         );
  MUX \b/U5190  ( .IN0(\b/n324 ), .IN1(msg[91]), .SEL(msg[89]), .F(\b/n5103 )
         );
  MUX \b/U5188  ( .IN0(msg[92]), .IN1(\b/n343 ), .SEL(msg[89]), .F(\b/n5101 )
         );
  MUX \b/U5187  ( .IN0(\b/n297 ), .IN1(\b/n349 ), .SEL(msg[89]), .F(\b/n5100 )
         );
  NAND \b/U5186  ( .A(\b/n5086 ), .B(\b/n297 ), .Z(\b/n5099 ) );
  MUX \b/U5185  ( .IN0(\b/n5085 ), .IN1(\b/n5093 ), .SEL(msg[89]), .F(
        \b/n5098 ) );
  NAND \b/U5184  ( .A(\b/n5097 ), .B(\b/n5084 ), .Z(\b/n5096 ) );
  MUX \b/U5183  ( .IN0(\b/n5088 ), .IN1(\b/n349 ), .SEL(msg[89]), .F(\b/n5095 ) );
  MUX \b/U5182  ( .IN0(\b/n349 ), .IN1(\b/n313 ), .SEL(msg[89]), .F(\b/n5094 )
         );
  NANDN \b/U5181  ( .B(msg[91]), .A(msg[92]), .Z(\b/n5093 ) );
  MUX \b/U5180  ( .IN0(\b/n5088 ), .IN1(msg[91]), .SEL(msg[89]), .F(\b/n5092 )
         );
  OR \b/U5179  ( .A(msg[91]), .B(msg[92]), .Z(\b/n5088 ) );
  MUX \b/U5178  ( .IN0(\b/n297 ), .IN1(\b/n313 ), .SEL(msg[89]), .F(\b/n5091 )
         );
  XOR \b/U5177  ( .A(\b/n307 ), .B(msg[91]), .Z(\b/n5090 ) );
  NANDN \b/U5176  ( .B(msg[91]), .A(msg[89]), .Z(\b/n5089 ) );
  NAND \b/U5175  ( .A(\b/n5088 ), .B(\b/n5086 ), .Z(\b/n5087 ) );
  NAND \b/U5174  ( .A(msg[89]), .B(\b/n5085 ), .Z(\b/n5086 ) );
  NANDN \b/U5173  ( .B(msg[92]), .A(msg[91]), .Z(\b/n5085 ) );
  NAND \b/U5172  ( .A(msg[91]), .B(msg[92]), .Z(\b/n5084 ) );
  MUX \b/U5171  ( .IN0(msg[84]), .IN1(\b/n4725 ), .SEL(msg[81]), .F(\b/n5083 )
         );
  MUX \b/U5170  ( .IN0(msg[84]), .IN1(\b/n4734 ), .SEL(msg[81]), .F(\b/n5082 )
         );
  MUX \b/U5169  ( .IN0(\b/n4726 ), .IN1(\b/n4729 ), .SEL(msg[81]), .F(
        \b/n5081 ) );
  MUX \b/U5168  ( .IN0(\b/n4731 ), .IN1(\b/n414 ), .SEL(msg[81]), .F(\b/n5080 ) );
  MUX \b/U5166  ( .IN0(\b/n4734 ), .IN1(\b/n4725 ), .SEL(msg[82]), .F(
        \b/n4907 ) );
  MUX \b/U5165  ( .IN0(\b/n4727 ), .IN1(\b/n425 ), .SEL(msg[82]), .F(\b/n4908 ) );
  MUX \b/U5164  ( .IN0(\b/n368 ), .IN1(\b/n378 ), .SEL(msg[81]), .F(\b/n4871 )
         );
  MUX \b/U5163  ( .IN0(\b/n4755 ), .IN1(\b/n5066 ), .SEL(msg[87]), .F(
        \b/n5078 ) );
  MUX \b/U5162  ( .IN0(\b/n4729 ), .IN1(\b/n4725 ), .SEL(msg[81]), .F(
        \b/n5069 ) );
  MUX \b/U5161  ( .IN0(\b/n420 ), .IN1(\b/n4731 ), .SEL(msg[81]), .F(\b/n5077 ) );
  MUX \b/U5160  ( .IN0(msg[83]), .IN1(\b/n414 ), .SEL(msg[81]), .F(\b/n5076 )
         );
  MUX \b/U5159  ( .IN0(\b/n4734 ), .IN1(\b/n420 ), .SEL(msg[81]), .F(\b/n5075 ) );
  MUX \b/U5158  ( .IN0(msg[84]), .IN1(\b/n4731 ), .SEL(msg[81]), .F(\b/n5074 )
         );
  MUX \b/U5157  ( .IN0(\b/n405 ), .IN1(\b/n384 ), .SEL(msg[85]), .F(\b/n4781 )
         );
  MUX \b/U5156  ( .IN0(\b/n4726 ), .IN1(\b/n378 ), .SEL(msg[81]), .F(\b/n5073 ) );
  NANDN \b/U5153  ( .B(\b/n4732 ), .A(msg[87]), .Z(\b/n5046 ) );
  NAND \b/U5152  ( .A(msg[87]), .B(\b/n381 ), .Z(\b/n5014 ) );
  NAND \b/U5151  ( .A(msg[87]), .B(\b/n393 ), .Z(\b/n4955 ) );
  NAND \b/U5150  ( .A(msg[87]), .B(\b/n5063 ), .Z(\b/n4988 ) );
  NAND \b/U5149  ( .A(msg[87]), .B(\b/n4983 ), .Z(\b/n4946 ) );
  NAND \b/U5147  ( .A(\b/n425 ), .B(\b/n414 ), .Z(\b/n5067 ) );
  NAND \b/U5146  ( .A(msg[87]), .B(\b/n5065 ), .Z(\b/n5060 ) );
  NAND \b/U5145  ( .A(n688), .B(msg[87]), .Z(\b/n5040 ) );
  NAND \b/U5143  ( .A(msg[82]), .B(\b/n4734 ), .Z(\b/n4900 ) );
  NAND \b/U5142  ( .A(\b/n414 ), .B(msg[81]), .Z(\b/n4855 ) );
  NAND \b/U5141  ( .A(msg[87]), .B(\b/n5069 ), .Z(\b/n4854 ) );
  NAND \b/U5139  ( .A(\b/n5067 ), .B(msg[87]), .Z(\b/n4870 ) );
  NAND \b/U5138  ( .A(\b/n4888 ), .B(\b/n4734 ), .Z(\b/n5066 ) );
  NANDN \b/U5137  ( .B(\b/n368 ), .A(\b/n425 ), .Z(\b/n5065 ) );
  NAND \b/U5135  ( .A(msg[81]), .B(\b/n4734 ), .Z(\b/n4786 ) );
  NAND \b/U5134  ( .A(\b/n368 ), .B(\b/n425 ), .Z(\b/n5063 ) );
  NAND \b/U5131  ( .A(msg[81]), .B(\b/n4729 ), .Z(\b/n4888 ) );
  ANDN \b/U5129  ( .A(msg[82]), .B(msg[81]), .Z(\b/n4916 ) );
  AND \b/U5128  ( .A(\b/n4726 ), .B(\b/n5060 ), .Z(\b/n4831 ) );
  MUX \b/U5127  ( .IN0(\b/n5059 ), .IN1(\b/n5043 ), .SEL(msg[86]), .F(
        shift_row_out[23]) );
  MUX \b/U5126  ( .IN0(\b/n5058 ), .IN1(\b/n5051 ), .SEL(msg[80]), .F(
        \b/n5059 ) );
  MUX \b/U5125  ( .IN0(\b/n5057 ), .IN1(\b/n5054 ), .SEL(msg[85]), .F(
        \b/n5058 ) );
  MUX \b/U5124  ( .IN0(\b/n5056 ), .IN1(\b/n5055 ), .SEL(msg[82]), .F(
        \b/n5057 ) );
  MUX \b/U5123  ( .IN0(msg[84]), .IN1(\b/n385 ), .SEL(msg[87]), .F(\b/n5056 )
         );
  MUX \b/U5122  ( .IN0(\b/n4727 ), .IN1(\b/n389 ), .SEL(msg[87]), .F(\b/n5055 ) );
  MUX \b/U5121  ( .IN0(\b/n5053 ), .IN1(\b/n5052 ), .SEL(msg[82]), .F(
        \b/n5054 ) );
  MUX \b/U5120  ( .IN0(\b/n4785 ), .IN1(\b/n381 ), .SEL(msg[87]), .F(\b/n5053 ) );
  MUX \b/U5119  ( .IN0(\b/n4737 ), .IN1(\b/n4748 ), .SEL(msg[87]), .F(
        \b/n5052 ) );
  MUX \b/U5118  ( .IN0(\b/n5050 ), .IN1(\b/n5047 ), .SEL(msg[85]), .F(
        \b/n5051 ) );
  MUX \b/U5117  ( .IN0(\b/n5049 ), .IN1(\b/n5048 ), .SEL(msg[82]), .F(
        \b/n5050 ) );
  MUX \b/U5116  ( .IN0(\b/n4761 ), .IN1(\b/n4736 ), .SEL(msg[87]), .F(
        \b/n5049 ) );
  MUX \b/U5115  ( .IN0(\b/n393 ), .IN1(\b/n4757 ), .SEL(msg[87]), .F(\b/n5048 ) );
  MUX \b/U5114  ( .IN0(\b/n5045 ), .IN1(\b/n5044 ), .SEL(msg[82]), .F(
        \b/n5047 ) );
  AND \b/U5113  ( .A(\b/n383 ), .B(\b/n5046 ), .Z(\b/n5045 ) );
  MUX \b/U5112  ( .IN0(\b/n4741 ), .IN1(n687), .SEL(msg[87]), .F(\b/n5044 ) );
  MUX \b/U5111  ( .IN0(\b/n5042 ), .IN1(\b/n5034 ), .SEL(msg[80]), .F(
        \b/n5043 ) );
  MUX \b/U5110  ( .IN0(\b/n5041 ), .IN1(\b/n5037 ), .SEL(msg[85]), .F(
        \b/n5042 ) );
  MUX \b/U5109  ( .IN0(\b/n5038 ), .IN1(\b/n5039 ), .SEL(msg[82]), .F(
        \b/n5041 ) );
  NAND \b/U5108  ( .A(\b/n4855 ), .B(\b/n5040 ), .Z(\b/n5039 ) );
  MUX \b/U5107  ( .IN0(\b/n423 ), .IN1(\b/n415 ), .SEL(msg[87]), .F(\b/n5038 )
         );
  MUX \b/U5106  ( .IN0(\b/n5036 ), .IN1(\b/n5035 ), .SEL(msg[82]), .F(
        \b/n5037 ) );
  MUX \b/U5105  ( .IN0(\b/n4731 ), .IN1(\b/n4725 ), .SEL(msg[87]), .F(
        \b/n5036 ) );
  MUX \b/U5104  ( .IN0(\b/n416 ), .IN1(\b/n4762 ), .SEL(msg[87]), .F(\b/n5035 ) );
  MUX \b/U5103  ( .IN0(\b/n5033 ), .IN1(\b/n5030 ), .SEL(msg[85]), .F(
        \b/n5034 ) );
  MUX \b/U5102  ( .IN0(\b/n5032 ), .IN1(\b/n5031 ), .SEL(msg[82]), .F(
        \b/n5033 ) );
  MUX \b/U5101  ( .IN0(\b/n4766 ), .IN1(\b/n4752 ), .SEL(msg[87]), .F(
        \b/n5032 ) );
  MUX \b/U5100  ( .IN0(\b/n369 ), .IN1(\b/n4734 ), .SEL(msg[87]), .F(\b/n5031 ) );
  MUX \b/U5099  ( .IN0(\b/n5029 ), .IN1(\b/n5028 ), .SEL(msg[82]), .F(
        \b/n5030 ) );
  MUX \b/U5098  ( .IN0(\b/n4767 ), .IN1(\b/n4775 ), .SEL(msg[87]), .F(
        \b/n5029 ) );
  MUX \b/U5097  ( .IN0(\b/n4760 ), .IN1(\b/n5027 ), .SEL(msg[87]), .F(
        \b/n5028 ) );
  MUX \b/U5096  ( .IN0(\b/n420 ), .IN1(\b/n378 ), .SEL(msg[81]), .F(\b/n5027 )
         );
  MUX \b/U5095  ( .IN0(\b/n5026 ), .IN1(\b/n5008 ), .SEL(msg[86]), .F(
        shift_row_out[22]) );
  MUX \b/U5094  ( .IN0(\b/n5025 ), .IN1(\b/n5016 ), .SEL(msg[80]), .F(
        \b/n5026 ) );
  MUX \b/U5093  ( .IN0(\b/n5024 ), .IN1(\b/n5019 ), .SEL(msg[85]), .F(
        \b/n5025 ) );
  MUX \b/U5092  ( .IN0(\b/n5023 ), .IN1(\b/n5021 ), .SEL(msg[82]), .F(
        \b/n5024 ) );
  MUX \b/U5091  ( .IN0(\b/n5022 ), .IN1(\b/n4738 ), .SEL(msg[87]), .F(
        \b/n5023 ) );
  MUX \b/U5090  ( .IN0(\b/n420 ), .IN1(\b/n4725 ), .SEL(msg[81]), .F(\b/n5022 ) );
  MUX \b/U5089  ( .IN0(\b/n5020 ), .IN1(\b/n408 ), .SEL(msg[87]), .F(\b/n5021 ) );
  MUX \b/U5088  ( .IN0(\b/n4725 ), .IN1(\b/n4726 ), .SEL(msg[81]), .F(
        \b/n5020 ) );
  MUX \b/U5087  ( .IN0(\b/n5018 ), .IN1(\b/n5017 ), .SEL(msg[82]), .F(
        \b/n5019 ) );
  MUX \b/U5086  ( .IN0(n686), .IN1(\b/n4806 ), .SEL(msg[87]), .F(\b/n5018 ) );
  MUX \b/U5085  ( .IN0(\b/n4764 ), .IN1(\b/n4771 ), .SEL(msg[87]), .F(
        \b/n5017 ) );
  MUX \b/U5084  ( .IN0(\b/n5015 ), .IN1(\b/n5011 ), .SEL(msg[85]), .F(
        \b/n5016 ) );
  MUX \b/U5083  ( .IN0(\b/n5013 ), .IN1(\b/n5012 ), .SEL(msg[82]), .F(
        \b/n5015 ) );
  AND \b/U5082  ( .A(\b/n361 ), .B(\b/n5014 ), .Z(\b/n5013 ) );
  MUX \b/U5081  ( .IN0(\b/n4841 ), .IN1(msg[83]), .SEL(msg[87]), .F(\b/n5012 )
         );
  MUX \b/U5080  ( .IN0(\b/n5010 ), .IN1(\b/n5009 ), .SEL(msg[82]), .F(
        \b/n5011 ) );
  MUX \b/U5079  ( .IN0(\b/n404 ), .IN1(\b/n4729 ), .SEL(msg[87]), .F(\b/n5010 ) );
  MUX \b/U5077  ( .IN0(\b/n5007 ), .IN1(\b/n5000 ), .SEL(msg[80]), .F(
        \b/n5008 ) );
  MUX \b/U5076  ( .IN0(\b/n5006 ), .IN1(\b/n5003 ), .SEL(msg[85]), .F(
        \b/n5007 ) );
  MUX \b/U5075  ( .IN0(\b/n5005 ), .IN1(\b/n5004 ), .SEL(msg[82]), .F(
        \b/n5006 ) );
  MUX \b/U5074  ( .IN0(\b/n400 ), .IN1(\b/n4733 ), .SEL(msg[87]), .F(\b/n5005 ) );
  MUX \b/U5073  ( .IN0(\b/n4737 ), .IN1(n687), .SEL(msg[87]), .F(\b/n5004 ) );
  MUX \b/U5072  ( .IN0(\b/n5002 ), .IN1(\b/n5001 ), .SEL(msg[82]), .F(
        \b/n5003 ) );
  MUX \b/U5071  ( .IN0(\b/n4753 ), .IN1(\b/n365 ), .SEL(msg[87]), .F(\b/n5002 ) );
  MUX \b/U5070  ( .IN0(\b/n385 ), .IN1(\b/n415 ), .SEL(msg[87]), .F(\b/n5001 )
         );
  MUX \b/U5069  ( .IN0(\b/n4999 ), .IN1(\b/n4995 ), .SEL(msg[85]), .F(
        \b/n5000 ) );
  MUX \b/U5068  ( .IN0(\b/n4998 ), .IN1(\b/n4997 ), .SEL(msg[82]), .F(
        \b/n4999 ) );
  MUX \b/U5067  ( .IN0(\b/n4742 ), .IN1(\b/n415 ), .SEL(msg[87]), .F(\b/n4998 ) );
  MUX \b/U5066  ( .IN0(\b/n4996 ), .IN1(\b/n4763 ), .SEL(msg[87]), .F(
        \b/n4997 ) );
  NANDN \b/U5065  ( .B(msg[84]), .A(msg[81]), .Z(\b/n4996 ) );
  MUX \b/U5064  ( .IN0(\b/n4994 ), .IN1(\b/n4992 ), .SEL(msg[82]), .F(
        \b/n4995 ) );
  MUX \b/U5063  ( .IN0(\b/n378 ), .IN1(\b/n4993 ), .SEL(msg[87]), .F(\b/n4994 ) );
  MUX \b/U5062  ( .IN0(\b/n405 ), .IN1(\b/n395 ), .SEL(msg[81]), .F(\b/n4993 )
         );
  MUX \b/U5061  ( .IN0(\b/n367 ), .IN1(\b/n4738 ), .SEL(msg[87]), .F(\b/n4992 ) );
  NANDN \b/U5060  ( .B(\b/n368 ), .A(msg[81]), .Z(\b/n4738 ) );
  MUX \b/U5059  ( .IN0(\b/n4991 ), .IN1(\b/n4970 ), .SEL(msg[86]), .F(
        shift_row_out[21]) );
  MUX \b/U5058  ( .IN0(\b/n4990 ), .IN1(\b/n4980 ), .SEL(msg[80]), .F(
        \b/n4991 ) );
  MUX \b/U5057  ( .IN0(\b/n4989 ), .IN1(\b/n4985 ), .SEL(msg[85]), .F(
        \b/n4990 ) );
  MUX \b/U5056  ( .IN0(\b/n4986 ), .IN1(\b/n4987 ), .SEL(msg[82]), .F(
        \b/n4989 ) );
  AND \b/U5055  ( .A(\b/n4756 ), .B(\b/n4988 ), .Z(\b/n4987 ) );
  MUX \b/U5054  ( .IN0(\b/n4734 ), .IN1(\b/n416 ), .SEL(msg[87]), .F(\b/n4986 ) );
  MUX \b/U5053  ( .IN0(\b/n4984 ), .IN1(\b/n4982 ), .SEL(msg[82]), .F(
        \b/n4985 ) );
  MUX \b/U5052  ( .IN0(\b/n371 ), .IN1(\b/n4983 ), .SEL(msg[87]), .F(\b/n4984 ) );
  NAND \b/U5051  ( .A(\b/n395 ), .B(\b/n425 ), .Z(\b/n4983 ) );
  MUX \b/U5050  ( .IN0(\b/n4734 ), .IN1(\b/n4981 ), .SEL(msg[87]), .F(
        \b/n4982 ) );
  NAND \b/U5049  ( .A(\b/n4725 ), .B(\b/n4786 ), .Z(\b/n4981 ) );
  MUX \b/U5048  ( .IN0(\b/n4979 ), .IN1(\b/n4975 ), .SEL(msg[85]), .F(
        \b/n4980 ) );
  MUX \b/U5047  ( .IN0(\b/n4978 ), .IN1(\b/n4977 ), .SEL(msg[82]), .F(
        \b/n4979 ) );
  MUX \b/U5046  ( .IN0(\b/n4746 ), .IN1(\b/n418 ), .SEL(msg[87]), .F(\b/n4978 ) );
  MUX \b/U5045  ( .IN0(\b/n4771 ), .IN1(\b/n4976 ), .SEL(msg[87]), .F(
        \b/n4977 ) );
  MUX \b/U5044  ( .IN0(\b/n414 ), .IN1(\b/n395 ), .SEL(msg[81]), .F(\b/n4976 )
         );
  MUX \b/U5043  ( .IN0(\b/n4974 ), .IN1(\b/n4973 ), .SEL(msg[82]), .F(
        \b/n4975 ) );
  MUX \b/U5042  ( .IN0(\b/n412 ), .IN1(n685), .SEL(msg[87]), .F(\b/n4974 ) );
  MUX \b/U5041  ( .IN0(\b/n4972 ), .IN1(\b/n4971 ), .SEL(msg[87]), .F(
        \b/n4973 ) );
  AND \b/U5040  ( .A(\b/n4731 ), .B(\b/n4806 ), .Z(\b/n4972 ) );
  MUX \b/U5039  ( .IN0(\b/n384 ), .IN1(\b/n368 ), .SEL(msg[81]), .F(\b/n4971 )
         );
  MUX \b/U5038  ( .IN0(\b/n4969 ), .IN1(\b/n4960 ), .SEL(msg[80]), .F(
        \b/n4970 ) );
  MUX \b/U5037  ( .IN0(\b/n4968 ), .IN1(\b/n4964 ), .SEL(msg[85]), .F(
        \b/n4969 ) );
  MUX \b/U5036  ( .IN0(\b/n4967 ), .IN1(\b/n4965 ), .SEL(msg[82]), .F(
        \b/n4968 ) );
  MUX \b/U5035  ( .IN0(\b/n4737 ), .IN1(\b/n4966 ), .SEL(msg[87]), .F(
        \b/n4967 ) );
  NAND \b/U5034  ( .A(msg[81]), .B(\b/n384 ), .Z(\b/n4966 ) );
  MUX \b/U5033  ( .IN0(\b/n368 ), .IN1(\b/n421 ), .SEL(msg[87]), .F(\b/n4965 )
         );
  MUX \b/U5032  ( .IN0(\b/n4963 ), .IN1(\b/n4962 ), .SEL(msg[82]), .F(
        \b/n4964 ) );
  MUX \b/U5031  ( .IN0(\b/n4763 ), .IN1(\b/n386 ), .SEL(msg[87]), .F(\b/n4963 ) );
  MUX \b/U5030  ( .IN0(\b/n4961 ), .IN1(\b/n4726 ), .SEL(n684), .F(\b/n4962 )
         );
  AND \b/U5029  ( .A(msg[87]), .B(msg[83]), .Z(\b/n4961 ) );
  MUX \b/U5028  ( .IN0(\b/n4959 ), .IN1(\b/n4956 ), .SEL(msg[85]), .F(
        \b/n4960 ) );
  MUX \b/U5027  ( .IN0(\b/n4958 ), .IN1(\b/n4957 ), .SEL(msg[82]), .F(
        \b/n4959 ) );
  MUX \b/U5026  ( .IN0(\b/n4887 ), .IN1(\b/n4726 ), .SEL(msg[87]), .F(
        \b/n4958 ) );
  MUX \b/U5025  ( .IN0(n683), .IN1(\b/n419 ), .SEL(msg[87]), .F(\b/n4957 ) );
  MUX \b/U5024  ( .IN0(\b/n4954 ), .IN1(\b/n4953 ), .SEL(msg[82]), .F(
        \b/n4956 ) );
  AND \b/U5023  ( .A(\b/n4955 ), .B(\b/n4855 ), .Z(\b/n4954 ) );
  MUX \b/U5022  ( .IN0(\b/n370 ), .IN1(\b/n414 ), .SEL(msg[87]), .F(\b/n4953 )
         );
  MUX \b/U5021  ( .IN0(\b/n4952 ), .IN1(\b/n4935 ), .SEL(msg[86]), .F(
        shift_row_out[20]) );
  MUX \b/U5020  ( .IN0(\b/n4951 ), .IN1(\b/n4943 ), .SEL(msg[80]), .F(
        \b/n4952 ) );
  MUX \b/U5019  ( .IN0(\b/n4950 ), .IN1(\b/n4947 ), .SEL(msg[85]), .F(
        \b/n4951 ) );
  MUX \b/U5018  ( .IN0(\b/n4949 ), .IN1(\b/n4948 ), .SEL(msg[82]), .F(
        \b/n4950 ) );
  MUX \b/U5017  ( .IN0(\b/n396 ), .IN1(\b/n417 ), .SEL(msg[87]), .F(\b/n4949 )
         );
  MUX \b/U5016  ( .IN0(\b/n4806 ), .IN1(\b/n4771 ), .SEL(msg[87]), .F(
        \b/n4948 ) );
  NAND \b/U5015  ( .A(msg[81]), .B(\b/n4725 ), .Z(\b/n4806 ) );
  MUX \b/U5014  ( .IN0(\b/n4944 ), .IN1(\b/n4945 ), .SEL(msg[82]), .F(
        \b/n4947 ) );
  AND \b/U5013  ( .A(\b/n4756 ), .B(\b/n4946 ), .Z(\b/n4945 ) );
  MUX \b/U5012  ( .IN0(\b/n4754 ), .IN1(\b/n399 ), .SEL(msg[87]), .F(\b/n4944 ) );
  MUX \b/U5011  ( .IN0(\b/n4942 ), .IN1(\b/n4939 ), .SEL(msg[85]), .F(
        \b/n4943 ) );
  MUX \b/U5010  ( .IN0(\b/n4941 ), .IN1(\b/n4940 ), .SEL(msg[82]), .F(
        \b/n4942 ) );
  MUX \b/U5009  ( .IN0(\b/n361 ), .IN1(\b/n407 ), .SEL(msg[87]), .F(\b/n4941 )
         );
  MUX \b/U5008  ( .IN0(\b/n368 ), .IN1(\b/n4734 ), .SEL(msg[87]), .F(\b/n4940 ) );
  MUX \b/U5007  ( .IN0(\b/n4938 ), .IN1(\b/n4936 ), .SEL(msg[82]), .F(
        \b/n4939 ) );
  MUX \b/U5006  ( .IN0(\b/n4750 ), .IN1(\b/n4937 ), .SEL(msg[87]), .F(
        \b/n4938 ) );
  AND \b/U5005  ( .A(\b/n4734 ), .B(\b/n425 ), .Z(\b/n4937 ) );
  MUX \b/U5004  ( .IN0(\b/n383 ), .IN1(\b/n402 ), .SEL(msg[87]), .F(\b/n4936 )
         );
  MUX \b/U5003  ( .IN0(\b/n4934 ), .IN1(\b/n4928 ), .SEL(msg[80]), .F(
        \b/n4935 ) );
  MUX \b/U5002  ( .IN0(\b/n4933 ), .IN1(\b/n4931 ), .SEL(msg[85]), .F(
        \b/n4934 ) );
  MUX \b/U5001  ( .IN0(\b/n4932 ), .IN1(\b/n4728 ), .SEL(msg[82]), .F(
        \b/n4933 ) );
  MUX \b/U5000  ( .IN0(\b/n4748 ), .IN1(\b/n404 ), .SEL(msg[87]), .F(\b/n4932 ) );
  MUX \b/U4999  ( .IN0(\b/n4930 ), .IN1(\b/n4929 ), .SEL(msg[82]), .F(
        \b/n4931 ) );
  MUX \b/U4998  ( .IN0(n682), .IN1(\b/n396 ), .SEL(msg[87]), .F(\b/n4930 ) );
  MUX \b/U4997  ( .IN0(\b/n4758 ), .IN1(\b/n4761 ), .SEL(msg[87]), .F(
        \b/n4929 ) );
  MUX \b/U4996  ( .IN0(\b/n4927 ), .IN1(\b/n4924 ), .SEL(msg[85]), .F(
        \b/n4928 ) );
  MUX \b/U4995  ( .IN0(\b/n4926 ), .IN1(\b/n4925 ), .SEL(msg[82]), .F(
        \b/n4927 ) );
  MUX \b/U4994  ( .IN0(\b/n369 ), .IN1(\b/n4730 ), .SEL(msg[87]), .F(\b/n4926 ) );
  MUX \b/U4993  ( .IN0(\b/n414 ), .IN1(\b/n4752 ), .SEL(msg[87]), .F(\b/n4925 ) );
  MUX \b/U4992  ( .IN0(\b/n357 ), .IN1(\b/n4923 ), .SEL(msg[82]), .F(\b/n4924 ) );
  MUX \b/U4991  ( .IN0(\b/n377 ), .IN1(\b/n4734 ), .SEL(msg[87]), .F(\b/n4923 ) );
  MUX \b/U4990  ( .IN0(\b/n4922 ), .IN1(\b/n4903 ), .SEL(msg[86]), .F(
        shift_row_out[19]) );
  MUX \b/U4989  ( .IN0(\b/n4921 ), .IN1(\b/n4913 ), .SEL(msg[80]), .F(
        \b/n4922 ) );
  MUX \b/U4988  ( .IN0(\b/n4920 ), .IN1(\b/n4917 ), .SEL(msg[85]), .F(
        \b/n4921 ) );
  MUX \b/U4987  ( .IN0(\b/n4919 ), .IN1(\b/n4918 ), .SEL(msg[87]), .F(
        \b/n4920 ) );
  MUX \b/U4986  ( .IN0(\b/n4742 ), .IN1(\b/n402 ), .SEL(msg[82]), .F(\b/n4919 ) );
  MUX \b/U4985  ( .IN0(n685), .IN1(\b/n360 ), .SEL(msg[82]), .F(\b/n4918 ) );
  MUX \b/U4984  ( .IN0(\b/n4915 ), .IN1(\b/n4914 ), .SEL(msg[87]), .F(
        \b/n4917 ) );
  AND \b/U4983  ( .A(\b/n4916 ), .B(msg[84]), .Z(\b/n4915 ) );
  MUX \b/U4982  ( .IN0(\b/n390 ), .IN1(\b/n4755 ), .SEL(msg[82]), .F(\b/n4914 ) );
  MUX \b/U4981  ( .IN0(\b/n4912 ), .IN1(\b/n4909 ), .SEL(msg[85]), .F(
        \b/n4913 ) );
  MUX \b/U4980  ( .IN0(\b/n4911 ), .IN1(\b/n4910 ), .SEL(msg[87]), .F(
        \b/n4912 ) );
  MUX \b/U4979  ( .IN0(\b/n4746 ), .IN1(n681), .SEL(msg[82]), .F(\b/n4911 ) );
  MUX \b/U4978  ( .IN0(\b/n358 ), .IN1(\b/n377 ), .SEL(msg[82]), .F(\b/n4910 )
         );
  MUX \b/U4977  ( .IN0(\b/n4905 ), .IN1(\b/n4906 ), .SEL(msg[87]), .F(
        \b/n4909 ) );
  NAND \b/U4976  ( .A(\b/n4907 ), .B(\b/n4908 ), .Z(\b/n4906 ) );
  MUX \b/U4975  ( .IN0(\b/n403 ), .IN1(\b/n4904 ), .SEL(msg[82]), .F(\b/n4905 ) );
  MUX \b/U4974  ( .IN0(\b/n378 ), .IN1(\b/n420 ), .SEL(msg[81]), .F(\b/n4904 )
         );
  MUX \b/U4973  ( .IN0(\b/n4902 ), .IN1(\b/n4893 ), .SEL(msg[80]), .F(
        \b/n4903 ) );
  MUX \b/U4972  ( .IN0(\b/n4901 ), .IN1(\b/n4897 ), .SEL(msg[85]), .F(
        \b/n4902 ) );
  MUX \b/U4971  ( .IN0(\b/n4899 ), .IN1(\b/n4898 ), .SEL(msg[87]), .F(
        \b/n4901 ) );
  NAND \b/U4970  ( .A(\b/n368 ), .B(\b/n4900 ), .Z(\b/n4899 ) );
  MUX \b/U4969  ( .IN0(\b/n419 ), .IN1(\b/n381 ), .SEL(msg[82]), .F(\b/n4898 )
         );
  MUX \b/U4968  ( .IN0(\b/n4896 ), .IN1(\b/n4894 ), .SEL(msg[87]), .F(
        \b/n4897 ) );
  MUX \b/U4967  ( .IN0(\b/n4737 ), .IN1(\b/n4895 ), .SEL(msg[82]), .F(
        \b/n4896 ) );
  AND \b/U4966  ( .A(msg[81]), .B(\b/n368 ), .Z(\b/n4895 ) );
  MUX \b/U4965  ( .IN0(\b/n373 ), .IN1(\b/n4756 ), .SEL(msg[82]), .F(\b/n4894 ) );
  MUX \b/U4964  ( .IN0(\b/n4892 ), .IN1(\b/n4886 ), .SEL(msg[85]), .F(
        \b/n4893 ) );
  MUX \b/U4963  ( .IN0(\b/n4891 ), .IN1(\b/n4889 ), .SEL(msg[87]), .F(
        \b/n4892 ) );
  MUX \b/U4962  ( .IN0(\b/n4890 ), .IN1(\b/n4726 ), .SEL(\b/n4774 ), .F(
        \b/n4891 ) );
  MUX \b/U4961  ( .IN0(msg[83]), .IN1(msg[84]), .SEL(msg[82]), .F(\b/n4890 )
         );
  MUX \b/U4960  ( .IN0(\b/n4756 ), .IN1(\b/n4887 ), .SEL(msg[82]), .F(
        \b/n4889 ) );
  NAND \b/U4959  ( .A(\b/n4726 ), .B(\b/n4888 ), .Z(\b/n4887 ) );
  MUX \b/U4958  ( .IN0(\b/n4883 ), .IN1(\b/n4884 ), .SEL(msg[87]), .F(
        \b/n4886 ) );
  AND \b/U4957  ( .A(\b/n401 ), .B(\b/n4885 ), .Z(\b/n4884 ) );
  MUX \b/U4956  ( .IN0(\b/n382 ), .IN1(\b/n4727 ), .SEL(msg[82]), .F(\b/n4883 ) );
  MUX \b/U4955  ( .IN0(\b/n4882 ), .IN1(\b/n4866 ), .SEL(msg[86]), .F(
        shift_row_out[18]) );
  MUX \b/U4954  ( .IN0(\b/n4881 ), .IN1(\b/n4873 ), .SEL(msg[80]), .F(
        \b/n4882 ) );
  MUX \b/U4953  ( .IN0(\b/n4880 ), .IN1(\b/n4876 ), .SEL(msg[85]), .F(
        \b/n4881 ) );
  MUX \b/U4952  ( .IN0(\b/n4879 ), .IN1(\b/n4877 ), .SEL(msg[82]), .F(
        \b/n4880 ) );
  MUX \b/U4951  ( .IN0(\b/n390 ), .IN1(\b/n4878 ), .SEL(msg[87]), .F(\b/n4879 ) );
  MUX \b/U4950  ( .IN0(\b/n4734 ), .IN1(\b/n368 ), .SEL(msg[81]), .F(\b/n4878 ) );
  MUX \b/U4949  ( .IN0(\b/n4773 ), .IN1(\b/n408 ), .SEL(msg[87]), .F(\b/n4877 ) );
  MUX \b/U4948  ( .IN0(\b/n4875 ), .IN1(\b/n4874 ), .SEL(msg[82]), .F(
        \b/n4876 ) );
  MUX \b/U4947  ( .IN0(\b/n4727 ), .IN1(\b/n375 ), .SEL(msg[87]), .F(\b/n4875 ) );
  MUX \b/U4946  ( .IN0(\b/n411 ), .IN1(\b/n4760 ), .SEL(msg[87]), .F(\b/n4874 ) );
  MUX \b/U4945  ( .IN0(\b/n4872 ), .IN1(\b/n4868 ), .SEL(msg[85]), .F(
        \b/n4873 ) );
  MUX \b/U4944  ( .IN0(\b/n4869 ), .IN1(\b/n357 ), .SEL(msg[82]), .F(\b/n4872 ) );
  NAND \b/U4943  ( .A(\b/n4870 ), .B(\b/n4871 ), .Z(\b/n4869 ) );
  MUX \b/U4942  ( .IN0(n683), .IN1(\b/n4867 ), .SEL(\b/n4772 ), .F(\b/n4868 )
         );
  MUX \b/U4941  ( .IN0(\b/n389 ), .IN1(\b/n4739 ), .SEL(msg[82]), .F(\b/n4867 ) );
  MUX \b/U4940  ( .IN0(\b/n4865 ), .IN1(\b/n4857 ), .SEL(msg[80]), .F(
        \b/n4866 ) );
  MUX \b/U4939  ( .IN0(\b/n4864 ), .IN1(\b/n4861 ), .SEL(msg[85]), .F(
        \b/n4865 ) );
  MUX \b/U4938  ( .IN0(\b/n4863 ), .IN1(\b/n4862 ), .SEL(msg[82]), .F(
        \b/n4864 ) );
  MUX \b/U4937  ( .IN0(\b/n417 ), .IN1(msg[81]), .SEL(msg[87]), .F(\b/n4863 )
         );
  MUX \b/U4936  ( .IN0(n686), .IN1(\b/n4740 ), .SEL(msg[87]), .F(\b/n4862 ) );
  MUX \b/U4935  ( .IN0(\b/n4860 ), .IN1(\b/n4859 ), .SEL(msg[82]), .F(
        \b/n4861 ) );
  MUX \b/U4934  ( .IN0(\b/n422 ), .IN1(\b/n416 ), .SEL(msg[87]), .F(\b/n4860 )
         );
  MUX \b/U4933  ( .IN0(n686), .IN1(\b/n4858 ), .SEL(msg[87]), .F(\b/n4859 ) );
  MUX \b/U4932  ( .IN0(\b/n368 ), .IN1(\b/n405 ), .SEL(msg[81]), .F(\b/n4858 )
         );
  MUX \b/U4931  ( .IN0(\b/n4856 ), .IN1(\b/n4850 ), .SEL(msg[85]), .F(
        \b/n4857 ) );
  MUX \b/U4930  ( .IN0(\b/n4853 ), .IN1(\b/n4852 ), .SEL(msg[82]), .F(
        \b/n4856 ) );
  NAND \b/U4929  ( .A(\b/n4854 ), .B(\b/n4855 ), .Z(\b/n4853 ) );
  MUX \b/U4928  ( .IN0(\b/n4726 ), .IN1(\b/n4851 ), .SEL(n684), .F(\b/n4852 )
         );
  MUX \b/U4927  ( .IN0(msg[83]), .IN1(\b/n378 ), .SEL(msg[87]), .F(\b/n4851 )
         );
  MUX \b/U4926  ( .IN0(\b/n4849 ), .IN1(\b/n4848 ), .SEL(msg[82]), .F(
        \b/n4850 ) );
  MUX \b/U4925  ( .IN0(\b/n4771 ), .IN1(\b/n376 ), .SEL(msg[87]), .F(\b/n4849 ) );
  MUX \b/U4924  ( .IN0(\b/n4767 ), .IN1(\b/n4847 ), .SEL(msg[87]), .F(
        \b/n4848 ) );
  MUX \b/U4923  ( .IN0(\b/n4729 ), .IN1(\b/n4734 ), .SEL(msg[81]), .F(
        \b/n4847 ) );
  MUX \b/U4922  ( .IN0(\b/n4846 ), .IN1(\b/n4828 ), .SEL(msg[86]), .F(
        shift_row_out[17]) );
  MUX \b/U4921  ( .IN0(\b/n4845 ), .IN1(\b/n4836 ), .SEL(msg[80]), .F(
        \b/n4846 ) );
  MUX \b/U4920  ( .IN0(\b/n4844 ), .IN1(\b/n4840 ), .SEL(msg[85]), .F(
        \b/n4845 ) );
  MUX \b/U4919  ( .IN0(\b/n4843 ), .IN1(\b/n4842 ), .SEL(msg[82]), .F(
        \b/n4844 ) );
  MUX \b/U4918  ( .IN0(\b/n413 ), .IN1(n688), .SEL(msg[87]), .F(\b/n4843 ) );
  MUX \b/U4917  ( .IN0(\b/n4841 ), .IN1(n682), .SEL(msg[87]), .F(\b/n4842 ) );
  NAND \b/U4916  ( .A(\b/n425 ), .B(\b/n384 ), .Z(\b/n4841 ) );
  MUX \b/U4915  ( .IN0(\b/n4839 ), .IN1(\b/n4838 ), .SEL(msg[82]), .F(
        \b/n4840 ) );
  MUX \b/U4914  ( .IN0(\b/n361 ), .IN1(\b/n4741 ), .SEL(msg[87]), .F(\b/n4839 ) );
  MUX \b/U4913  ( .IN0(\b/n4731 ), .IN1(\b/n4837 ), .SEL(msg[87]), .F(
        \b/n4838 ) );
  AND \b/U4912  ( .A(msg[81]), .B(msg[84]), .Z(\b/n4837 ) );
  MUX \b/U4911  ( .IN0(\b/n4835 ), .IN1(\b/n4832 ), .SEL(msg[85]), .F(
        \b/n4836 ) );
  MUX \b/U4910  ( .IN0(\b/n4834 ), .IN1(\b/n4833 ), .SEL(msg[82]), .F(
        \b/n4835 ) );
  MUX \b/U4909  ( .IN0(\b/n4770 ), .IN1(\b/n422 ), .SEL(msg[87]), .F(\b/n4834 ) );
  MUX \b/U4908  ( .IN0(\b/n397 ), .IN1(\b/n4739 ), .SEL(msg[87]), .F(\b/n4833 ) );
  MUX \b/U4907  ( .IN0(\b/n4829 ), .IN1(\b/n4830 ), .SEL(msg[82]), .F(
        \b/n4832 ) );
  AND \b/U4906  ( .A(\b/n4831 ), .B(\b/n4786 ), .Z(\b/n4830 ) );
  MUX \b/U4905  ( .IN0(\b/n4745 ), .IN1(\b/n4734 ), .SEL(msg[87]), .F(
        \b/n4829 ) );
  MUX \b/U4904  ( .IN0(\b/n4827 ), .IN1(\b/n4819 ), .SEL(msg[80]), .F(
        \b/n4828 ) );
  MUX \b/U4903  ( .IN0(\b/n4826 ), .IN1(\b/n4822 ), .SEL(msg[85]), .F(
        \b/n4827 ) );
  MUX \b/U4902  ( .IN0(\b/n4825 ), .IN1(\b/n4824 ), .SEL(msg[82]), .F(
        \b/n4826 ) );
  MUX \b/U4901  ( .IN0(\b/n4733 ), .IN1(\b/n386 ), .SEL(msg[87]), .F(\b/n4825 ) );
  MUX \b/U4900  ( .IN0(\b/n4823 ), .IN1(\b/n370 ), .SEL(msg[87]), .F(\b/n4824 ) );
  MUX \b/U4899  ( .IN0(\b/n4731 ), .IN1(\b/n378 ), .SEL(msg[81]), .F(\b/n4823 ) );
  MUX \b/U4898  ( .IN0(\b/n4821 ), .IN1(\b/n4820 ), .SEL(msg[82]), .F(
        \b/n4822 ) );
  MUX \b/U4897  ( .IN0(\b/n417 ), .IN1(\b/n395 ), .SEL(msg[87]), .F(\b/n4821 )
         );
  MUX \b/U4896  ( .IN0(\b/n413 ), .IN1(\b/n373 ), .SEL(msg[87]), .F(\b/n4820 )
         );
  MUX \b/U4895  ( .IN0(\b/n4818 ), .IN1(\b/n4813 ), .SEL(msg[85]), .F(
        \b/n4819 ) );
  MUX \b/U4894  ( .IN0(\b/n4817 ), .IN1(\b/n4814 ), .SEL(msg[82]), .F(
        \b/n4818 ) );
  MUX \b/U4893  ( .IN0(\b/n4815 ), .IN1(\b/n4816 ), .SEL(msg[87]), .F(
        \b/n4817 ) );
  NAND \b/U4892  ( .A(\b/n4734 ), .B(\b/n4806 ), .Z(\b/n4816 ) );
  MUX \b/U4891  ( .IN0(\b/n4734 ), .IN1(\b/n378 ), .SEL(msg[81]), .F(\b/n4815 ) );
  MUX \b/U4890  ( .IN0(\b/n4751 ), .IN1(\b/n4749 ), .SEL(msg[87]), .F(
        \b/n4814 ) );
  MUX \b/U4889  ( .IN0(\b/n4769 ), .IN1(\b/n4812 ), .SEL(msg[82]), .F(
        \b/n4813 ) );
  MUX \b/U4888  ( .IN0(\b/n384 ), .IN1(\b/n416 ), .SEL(msg[87]), .F(\b/n4812 )
         );
  MUX \b/U4887  ( .IN0(\b/n4811 ), .IN1(\b/n4794 ), .SEL(msg[86]), .F(
        shift_row_out[16]) );
  MUX \b/U4886  ( .IN0(\b/n4810 ), .IN1(\b/n4802 ), .SEL(msg[80]), .F(
        \b/n4811 ) );
  MUX \b/U4885  ( .IN0(\b/n4809 ), .IN1(\b/n4807 ), .SEL(msg[82]), .F(
        \b/n4810 ) );
  MUX \b/U4884  ( .IN0(\b/n358 ), .IN1(\b/n4808 ), .SEL(msg[87]), .F(\b/n4809 ) );
  MUX \b/U4883  ( .IN0(\b/n411 ), .IN1(\b/n414 ), .SEL(msg[85]), .F(\b/n4808 )
         );
  MUX \b/U4882  ( .IN0(\b/n4804 ), .IN1(\b/n4803 ), .SEL(msg[87]), .F(
        \b/n4807 ) );
  NAND \b/U4881  ( .A(\b/n4805 ), .B(\b/n4806 ), .Z(\b/n4804 ) );
  MUX \b/U4880  ( .IN0(\b/n410 ), .IN1(\b/n425 ), .SEL(msg[85]), .F(\b/n4803 )
         );
  MUX \b/U4879  ( .IN0(\b/n4801 ), .IN1(\b/n4797 ), .SEL(msg[82]), .F(
        \b/n4802 ) );
  MUX \b/U4878  ( .IN0(\b/n4800 ), .IN1(\b/n4798 ), .SEL(msg[87]), .F(
        \b/n4801 ) );
  MUX \b/U4877  ( .IN0(\b/n4799 ), .IN1(\b/n363 ), .SEL(msg[85]), .F(\b/n4800 ) );
  NAND \b/U4876  ( .A(\b/n425 ), .B(\b/n4726 ), .Z(\b/n4799 ) );
  MUX \b/U4874  ( .IN0(\b/n4796 ), .IN1(\b/n4795 ), .SEL(msg[87]), .F(
        \b/n4797 ) );
  MUX \b/U4873  ( .IN0(n683), .IN1(\b/n360 ), .SEL(msg[85]), .F(\b/n4796 ) );
  MUX \b/U4872  ( .IN0(\b/n412 ), .IN1(\b/n368 ), .SEL(msg[85]), .F(\b/n4795 )
         );
  MUX \b/U4871  ( .IN0(\b/n4793 ), .IN1(\b/n4783 ), .SEL(msg[80]), .F(
        \b/n4794 ) );
  MUX \b/U4870  ( .IN0(\b/n4792 ), .IN1(\b/n4788 ), .SEL(msg[82]), .F(
        \b/n4793 ) );
  MUX \b/U4869  ( .IN0(\b/n4791 ), .IN1(\b/n4790 ), .SEL(msg[87]), .F(
        \b/n4792 ) );
  MUX \b/U4868  ( .IN0(n681), .IN1(\b/n364 ), .SEL(msg[85]), .F(\b/n4791 ) );
  MUX \b/U4867  ( .IN0(\b/n4789 ), .IN1(\b/n401 ), .SEL(msg[85]), .F(\b/n4790 ) );
  NAND \b/U4866  ( .A(\b/n4725 ), .B(\b/n4727 ), .Z(\b/n4789 ) );
  MUX \b/U4865  ( .IN0(\b/n4787 ), .IN1(\b/n4784 ), .SEL(msg[87]), .F(
        \b/n4788 ) );
  MUX \b/U4864  ( .IN0(\b/n371 ), .IN1(\b/n4785 ), .SEL(msg[85]), .F(\b/n4787 ) );
  NAND \b/U4863  ( .A(\b/n4729 ), .B(\b/n4786 ), .Z(\b/n4785 ) );
  MUX \b/U4862  ( .IN0(\b/n4744 ), .IN1(\b/n4735 ), .SEL(msg[85]), .F(
        \b/n4784 ) );
  MUX \b/U4861  ( .IN0(\b/n4782 ), .IN1(\b/n4778 ), .SEL(msg[82]), .F(
        \b/n4783 ) );
  MUX \b/U4860  ( .IN0(\b/n4780 ), .IN1(\b/n4779 ), .SEL(msg[87]), .F(
        \b/n4782 ) );
  NAND \b/U4859  ( .A(\b/n4781 ), .B(\b/n4768 ), .Z(\b/n4780 ) );
  MUX \b/U4858  ( .IN0(msg[83]), .IN1(\b/n4760 ), .SEL(msg[85]), .F(\b/n4779 )
         );
  MUX \b/U4857  ( .IN0(\b/n4777 ), .IN1(\b/n4776 ), .SEL(msg[87]), .F(
        \b/n4778 ) );
  MUX \b/U4856  ( .IN0(\b/n376 ), .IN1(\b/n392 ), .SEL(msg[85]), .F(\b/n4777 )
         );
  MUX \b/U4855  ( .IN0(\b/n409 ), .IN1(\b/n397 ), .SEL(msg[85]), .F(\b/n4776 )
         );
  XOR \b/U4854  ( .A(\b/n4726 ), .B(msg[81]), .Z(\b/n4775 ) );
  XOR \b/U4853  ( .A(msg[81]), .B(msg[82]), .Z(\b/n4774 ) );
  XOR \b/U4852  ( .A(msg[81]), .B(msg[83]), .Z(\b/n4773 ) );
  XOR \b/U4851  ( .A(msg[82]), .B(msg[87]), .Z(\b/n4772 ) );
  XOR \b/U4850  ( .A(\b/n425 ), .B(\b/n368 ), .Z(\b/n4771 ) );
  XOR \b/U4849  ( .A(msg[81]), .B(\b/n414 ), .Z(\b/n4770 ) );
  XOR \b/U4847  ( .A(msg[81]), .B(msg[85]), .Z(\b/n4768 ) );
  NAND \b/U4846  ( .A(msg[81]), .B(msg[83]), .Z(\b/n4767 ) );
  MUX \b/U4845  ( .IN0(\b/n4726 ), .IN1(\b/n368 ), .SEL(msg[81]), .F(\b/n4766 ) );
  MUX \b/U4843  ( .IN0(msg[83]), .IN1(\b/n405 ), .SEL(msg[81]), .F(\b/n4764 )
         );
  MUX \b/U4842  ( .IN0(\b/n384 ), .IN1(\b/n405 ), .SEL(msg[81]), .F(\b/n4763 )
         );
  MUX \b/U4841  ( .IN0(\b/n4729 ), .IN1(\b/n4731 ), .SEL(msg[81]), .F(
        \b/n4762 ) );
  MUX \b/U4840  ( .IN0(msg[84]), .IN1(\b/n384 ), .SEL(msg[81]), .F(\b/n4761 )
         );
  OR \b/U4839  ( .A(msg[81]), .B(msg[84]), .Z(\b/n4760 ) );
  NAND \b/U4837  ( .A(\b/n405 ), .B(\b/n425 ), .Z(\b/n4758 ) );
  MUX \b/U4836  ( .IN0(\b/n405 ), .IN1(msg[84]), .SEL(msg[81]), .F(\b/n4757 )
         );
  MUX \b/U4835  ( .IN0(\b/n4725 ), .IN1(\b/n4734 ), .SEL(msg[81]), .F(
        \b/n4756 ) );
  MUX \b/U4834  ( .IN0(\b/n420 ), .IN1(msg[84]), .SEL(msg[81]), .F(\b/n4755 )
         );
  MUX \b/U4833  ( .IN0(\b/n378 ), .IN1(\b/n405 ), .SEL(msg[81]), .F(\b/n4754 )
         );
  MUX \b/U4832  ( .IN0(\b/n4725 ), .IN1(msg[84]), .SEL(msg[81]), .F(\b/n4753 )
         );
  MUX \b/U4831  ( .IN0(\b/n395 ), .IN1(\b/n384 ), .SEL(msg[81]), .F(\b/n4752 )
         );
  XOR \b/U4830  ( .A(\b/n378 ), .B(msg[81]), .Z(\b/n4751 ) );
  MUX \b/U4829  ( .IN0(\b/n4731 ), .IN1(\b/n395 ), .SEL(msg[81]), .F(\b/n4750 ) );
  NANDN \b/U4828  ( .B(msg[81]), .A(msg[83]), .Z(\b/n4749 ) );
  MUX \b/U4827  ( .IN0(\b/n368 ), .IN1(msg[83]), .SEL(msg[81]), .F(\b/n4748 )
         );
  NAND \b/U4825  ( .A(\b/n4729 ), .B(\b/n425 ), .Z(\b/n4746 ) );
  MUX \b/U4824  ( .IN0(msg[84]), .IN1(\b/n4726 ), .SEL(msg[81]), .F(\b/n4745 )
         );
  MUX \b/U4823  ( .IN0(\b/n395 ), .IN1(msg[83]), .SEL(msg[81]), .F(\b/n4744 )
         );
  MUX \b/U4821  ( .IN0(msg[84]), .IN1(\b/n414 ), .SEL(msg[81]), .F(\b/n4742 )
         );
  MUX \b/U4820  ( .IN0(\b/n368 ), .IN1(\b/n420 ), .SEL(msg[81]), .F(\b/n4741 )
         );
  NAND \b/U4819  ( .A(\b/n4727 ), .B(\b/n368 ), .Z(\b/n4740 ) );
  MUX \b/U4818  ( .IN0(\b/n4726 ), .IN1(\b/n4734 ), .SEL(msg[81]), .F(
        \b/n4739 ) );
  NAND \b/U4817  ( .A(\b/n4738 ), .B(\b/n4725 ), .Z(\b/n4737 ) );
  MUX \b/U4816  ( .IN0(\b/n4729 ), .IN1(\b/n420 ), .SEL(msg[81]), .F(\b/n4736 ) );
  MUX \b/U4815  ( .IN0(\b/n420 ), .IN1(\b/n384 ), .SEL(msg[81]), .F(\b/n4735 )
         );
  NANDN \b/U4814  ( .B(msg[83]), .A(msg[84]), .Z(\b/n4734 ) );
  MUX \b/U4813  ( .IN0(\b/n4729 ), .IN1(msg[83]), .SEL(msg[81]), .F(\b/n4733 )
         );
  OR \b/U4812  ( .A(msg[83]), .B(msg[84]), .Z(\b/n4729 ) );
  MUX \b/U4811  ( .IN0(\b/n368 ), .IN1(\b/n384 ), .SEL(msg[81]), .F(\b/n4732 )
         );
  XOR \b/U4810  ( .A(\b/n378 ), .B(msg[83]), .Z(\b/n4731 ) );
  NANDN \b/U4809  ( .B(msg[83]), .A(msg[81]), .Z(\b/n4730 ) );
  NAND \b/U4808  ( .A(\b/n4729 ), .B(\b/n4727 ), .Z(\b/n4728 ) );
  NAND \b/U4807  ( .A(msg[81]), .B(\b/n4726 ), .Z(\b/n4727 ) );
  NANDN \b/U4806  ( .B(msg[84]), .A(msg[83]), .Z(\b/n4726 ) );
  NAND \b/U4805  ( .A(msg[83]), .B(msg[84]), .Z(\b/n4725 ) );
  MUX \b/U4804  ( .IN0(msg[76]), .IN1(\b/n4366 ), .SEL(msg[73]), .F(\b/n4724 )
         );
  MUX \b/U4803  ( .IN0(msg[76]), .IN1(\b/n4375 ), .SEL(msg[73]), .F(\b/n4723 )
         );
  MUX \b/U4802  ( .IN0(\b/n4367 ), .IN1(\b/n4370 ), .SEL(msg[73]), .F(
        \b/n4722 ) );
  MUX \b/U4801  ( .IN0(\b/n4372 ), .IN1(\b/n485 ), .SEL(msg[73]), .F(\b/n4721 ) );
  MUX \b/U4799  ( .IN0(\b/n4375 ), .IN1(\b/n4366 ), .SEL(msg[74]), .F(
        \b/n4548 ) );
  MUX \b/U4798  ( .IN0(\b/n4368 ), .IN1(\b/n496 ), .SEL(msg[74]), .F(\b/n4549 ) );
  MUX \b/U4797  ( .IN0(\b/n439 ), .IN1(\b/n449 ), .SEL(msg[73]), .F(\b/n4512 )
         );
  MUX \b/U4796  ( .IN0(\b/n4396 ), .IN1(\b/n4707 ), .SEL(msg[79]), .F(
        \b/n4719 ) );
  MUX \b/U4795  ( .IN0(\b/n4370 ), .IN1(\b/n4366 ), .SEL(msg[73]), .F(
        \b/n4710 ) );
  MUX \b/U4794  ( .IN0(\b/n491 ), .IN1(\b/n4372 ), .SEL(msg[73]), .F(\b/n4718 ) );
  MUX \b/U4793  ( .IN0(msg[75]), .IN1(\b/n485 ), .SEL(msg[73]), .F(\b/n4717 )
         );
  MUX \b/U4792  ( .IN0(\b/n4375 ), .IN1(\b/n491 ), .SEL(msg[73]), .F(\b/n4716 ) );
  MUX \b/U4791  ( .IN0(msg[76]), .IN1(\b/n4372 ), .SEL(msg[73]), .F(\b/n4715 )
         );
  MUX \b/U4790  ( .IN0(\b/n476 ), .IN1(\b/n455 ), .SEL(msg[77]), .F(\b/n4422 )
         );
  MUX \b/U4789  ( .IN0(\b/n4367 ), .IN1(\b/n449 ), .SEL(msg[73]), .F(\b/n4714 ) );
  NANDN \b/U4786  ( .B(\b/n4373 ), .A(msg[79]), .Z(\b/n4687 ) );
  NAND \b/U4785  ( .A(msg[79]), .B(\b/n452 ), .Z(\b/n4655 ) );
  NAND \b/U4784  ( .A(msg[79]), .B(\b/n464 ), .Z(\b/n4596 ) );
  NAND \b/U4783  ( .A(msg[79]), .B(\b/n4704 ), .Z(\b/n4629 ) );
  NAND \b/U4782  ( .A(msg[79]), .B(\b/n4624 ), .Z(\b/n4587 ) );
  NAND \b/U4780  ( .A(\b/n496 ), .B(\b/n485 ), .Z(\b/n4708 ) );
  NAND \b/U4779  ( .A(msg[79]), .B(\b/n4706 ), .Z(\b/n4701 ) );
  NAND \b/U4778  ( .A(n680), .B(msg[79]), .Z(\b/n4681 ) );
  NAND \b/U4776  ( .A(msg[74]), .B(\b/n4375 ), .Z(\b/n4541 ) );
  NAND \b/U4775  ( .A(\b/n485 ), .B(msg[73]), .Z(\b/n4496 ) );
  NAND \b/U4774  ( .A(msg[79]), .B(\b/n4710 ), .Z(\b/n4495 ) );
  NAND \b/U4772  ( .A(\b/n4708 ), .B(msg[79]), .Z(\b/n4511 ) );
  NAND \b/U4771  ( .A(\b/n4529 ), .B(\b/n4375 ), .Z(\b/n4707 ) );
  NANDN \b/U4770  ( .B(\b/n439 ), .A(\b/n496 ), .Z(\b/n4706 ) );
  NAND \b/U4768  ( .A(msg[73]), .B(\b/n4375 ), .Z(\b/n4427 ) );
  NAND \b/U4767  ( .A(\b/n439 ), .B(\b/n496 ), .Z(\b/n4704 ) );
  NAND \b/U4764  ( .A(msg[73]), .B(\b/n4370 ), .Z(\b/n4529 ) );
  ANDN \b/U4762  ( .A(msg[74]), .B(msg[73]), .Z(\b/n4557 ) );
  AND \b/U4761  ( .A(\b/n4367 ), .B(\b/n4701 ), .Z(\b/n4472 ) );
  MUX \b/U4760  ( .IN0(\b/n4700 ), .IN1(\b/n4684 ), .SEL(msg[78]), .F(
        shift_row_out[47]) );
  MUX \b/U4759  ( .IN0(\b/n4699 ), .IN1(\b/n4692 ), .SEL(msg[72]), .F(
        \b/n4700 ) );
  MUX \b/U4758  ( .IN0(\b/n4698 ), .IN1(\b/n4695 ), .SEL(msg[77]), .F(
        \b/n4699 ) );
  MUX \b/U4757  ( .IN0(\b/n4697 ), .IN1(\b/n4696 ), .SEL(msg[74]), .F(
        \b/n4698 ) );
  MUX \b/U4756  ( .IN0(msg[76]), .IN1(\b/n456 ), .SEL(msg[79]), .F(\b/n4697 )
         );
  MUX \b/U4755  ( .IN0(\b/n4368 ), .IN1(\b/n460 ), .SEL(msg[79]), .F(\b/n4696 ) );
  MUX \b/U4754  ( .IN0(\b/n4694 ), .IN1(\b/n4693 ), .SEL(msg[74]), .F(
        \b/n4695 ) );
  MUX \b/U4753  ( .IN0(\b/n4426 ), .IN1(\b/n452 ), .SEL(msg[79]), .F(\b/n4694 ) );
  MUX \b/U4752  ( .IN0(\b/n4378 ), .IN1(\b/n4389 ), .SEL(msg[79]), .F(
        \b/n4693 ) );
  MUX \b/U4751  ( .IN0(\b/n4691 ), .IN1(\b/n4688 ), .SEL(msg[77]), .F(
        \b/n4692 ) );
  MUX \b/U4750  ( .IN0(\b/n4690 ), .IN1(\b/n4689 ), .SEL(msg[74]), .F(
        \b/n4691 ) );
  MUX \b/U4749  ( .IN0(\b/n4402 ), .IN1(\b/n4377 ), .SEL(msg[79]), .F(
        \b/n4690 ) );
  MUX \b/U4748  ( .IN0(\b/n464 ), .IN1(\b/n4398 ), .SEL(msg[79]), .F(\b/n4689 ) );
  MUX \b/U4747  ( .IN0(\b/n4686 ), .IN1(\b/n4685 ), .SEL(msg[74]), .F(
        \b/n4688 ) );
  AND \b/U4746  ( .A(\b/n454 ), .B(\b/n4687 ), .Z(\b/n4686 ) );
  MUX \b/U4745  ( .IN0(\b/n4382 ), .IN1(n679), .SEL(msg[79]), .F(\b/n4685 ) );
  MUX \b/U4744  ( .IN0(\b/n4683 ), .IN1(\b/n4675 ), .SEL(msg[72]), .F(
        \b/n4684 ) );
  MUX \b/U4743  ( .IN0(\b/n4682 ), .IN1(\b/n4678 ), .SEL(msg[77]), .F(
        \b/n4683 ) );
  MUX \b/U4742  ( .IN0(\b/n4679 ), .IN1(\b/n4680 ), .SEL(msg[74]), .F(
        \b/n4682 ) );
  NAND \b/U4741  ( .A(\b/n4496 ), .B(\b/n4681 ), .Z(\b/n4680 ) );
  MUX \b/U4740  ( .IN0(\b/n494 ), .IN1(\b/n486 ), .SEL(msg[79]), .F(\b/n4679 )
         );
  MUX \b/U4739  ( .IN0(\b/n4677 ), .IN1(\b/n4676 ), .SEL(msg[74]), .F(
        \b/n4678 ) );
  MUX \b/U4738  ( .IN0(\b/n4372 ), .IN1(\b/n4366 ), .SEL(msg[79]), .F(
        \b/n4677 ) );
  MUX \b/U4737  ( .IN0(\b/n487 ), .IN1(\b/n4403 ), .SEL(msg[79]), .F(\b/n4676 ) );
  MUX \b/U4736  ( .IN0(\b/n4674 ), .IN1(\b/n4671 ), .SEL(msg[77]), .F(
        \b/n4675 ) );
  MUX \b/U4735  ( .IN0(\b/n4673 ), .IN1(\b/n4672 ), .SEL(msg[74]), .F(
        \b/n4674 ) );
  MUX \b/U4734  ( .IN0(\b/n4407 ), .IN1(\b/n4393 ), .SEL(msg[79]), .F(
        \b/n4673 ) );
  MUX \b/U4733  ( .IN0(\b/n440 ), .IN1(\b/n4375 ), .SEL(msg[79]), .F(\b/n4672 ) );
  MUX \b/U4732  ( .IN0(\b/n4670 ), .IN1(\b/n4669 ), .SEL(msg[74]), .F(
        \b/n4671 ) );
  MUX \b/U4731  ( .IN0(\b/n4408 ), .IN1(\b/n4416 ), .SEL(msg[79]), .F(
        \b/n4670 ) );
  MUX \b/U4730  ( .IN0(\b/n4401 ), .IN1(\b/n4668 ), .SEL(msg[79]), .F(
        \b/n4669 ) );
  MUX \b/U4729  ( .IN0(\b/n491 ), .IN1(\b/n449 ), .SEL(msg[73]), .F(\b/n4668 )
         );
  MUX \b/U4728  ( .IN0(\b/n4667 ), .IN1(\b/n4649 ), .SEL(msg[78]), .F(
        shift_row_out[46]) );
  MUX \b/U4727  ( .IN0(\b/n4666 ), .IN1(\b/n4657 ), .SEL(msg[72]), .F(
        \b/n4667 ) );
  MUX \b/U4726  ( .IN0(\b/n4665 ), .IN1(\b/n4660 ), .SEL(msg[77]), .F(
        \b/n4666 ) );
  MUX \b/U4725  ( .IN0(\b/n4664 ), .IN1(\b/n4662 ), .SEL(msg[74]), .F(
        \b/n4665 ) );
  MUX \b/U4724  ( .IN0(\b/n4663 ), .IN1(\b/n4379 ), .SEL(msg[79]), .F(
        \b/n4664 ) );
  MUX \b/U4723  ( .IN0(\b/n491 ), .IN1(\b/n4366 ), .SEL(msg[73]), .F(\b/n4663 ) );
  MUX \b/U4722  ( .IN0(\b/n4661 ), .IN1(\b/n479 ), .SEL(msg[79]), .F(\b/n4662 ) );
  MUX \b/U4721  ( .IN0(\b/n4366 ), .IN1(\b/n4367 ), .SEL(msg[73]), .F(
        \b/n4661 ) );
  MUX \b/U4720  ( .IN0(\b/n4659 ), .IN1(\b/n4658 ), .SEL(msg[74]), .F(
        \b/n4660 ) );
  MUX \b/U4719  ( .IN0(n678), .IN1(\b/n4447 ), .SEL(msg[79]), .F(\b/n4659 ) );
  MUX \b/U4718  ( .IN0(\b/n4405 ), .IN1(\b/n4412 ), .SEL(msg[79]), .F(
        \b/n4658 ) );
  MUX \b/U4717  ( .IN0(\b/n4656 ), .IN1(\b/n4652 ), .SEL(msg[77]), .F(
        \b/n4657 ) );
  MUX \b/U4716  ( .IN0(\b/n4654 ), .IN1(\b/n4653 ), .SEL(msg[74]), .F(
        \b/n4656 ) );
  AND \b/U4715  ( .A(\b/n432 ), .B(\b/n4655 ), .Z(\b/n4654 ) );
  MUX \b/U4714  ( .IN0(\b/n4482 ), .IN1(msg[75]), .SEL(msg[79]), .F(\b/n4653 )
         );
  MUX \b/U4713  ( .IN0(\b/n4651 ), .IN1(\b/n4650 ), .SEL(msg[74]), .F(
        \b/n4652 ) );
  MUX \b/U4712  ( .IN0(\b/n475 ), .IN1(\b/n4370 ), .SEL(msg[79]), .F(\b/n4651 ) );
  MUX \b/U4710  ( .IN0(\b/n4648 ), .IN1(\b/n4641 ), .SEL(msg[72]), .F(
        \b/n4649 ) );
  MUX \b/U4709  ( .IN0(\b/n4647 ), .IN1(\b/n4644 ), .SEL(msg[77]), .F(
        \b/n4648 ) );
  MUX \b/U4708  ( .IN0(\b/n4646 ), .IN1(\b/n4645 ), .SEL(msg[74]), .F(
        \b/n4647 ) );
  MUX \b/U4707  ( .IN0(\b/n471 ), .IN1(\b/n4374 ), .SEL(msg[79]), .F(\b/n4646 ) );
  MUX \b/U4706  ( .IN0(\b/n4378 ), .IN1(n679), .SEL(msg[79]), .F(\b/n4645 ) );
  MUX \b/U4705  ( .IN0(\b/n4643 ), .IN1(\b/n4642 ), .SEL(msg[74]), .F(
        \b/n4644 ) );
  MUX \b/U4704  ( .IN0(\b/n4394 ), .IN1(\b/n436 ), .SEL(msg[79]), .F(\b/n4643 ) );
  MUX \b/U4703  ( .IN0(\b/n456 ), .IN1(\b/n486 ), .SEL(msg[79]), .F(\b/n4642 )
         );
  MUX \b/U4702  ( .IN0(\b/n4640 ), .IN1(\b/n4636 ), .SEL(msg[77]), .F(
        \b/n4641 ) );
  MUX \b/U4701  ( .IN0(\b/n4639 ), .IN1(\b/n4638 ), .SEL(msg[74]), .F(
        \b/n4640 ) );
  MUX \b/U4700  ( .IN0(\b/n4383 ), .IN1(\b/n486 ), .SEL(msg[79]), .F(\b/n4639 ) );
  MUX \b/U4699  ( .IN0(\b/n4637 ), .IN1(\b/n4404 ), .SEL(msg[79]), .F(
        \b/n4638 ) );
  NANDN \b/U4698  ( .B(msg[76]), .A(msg[73]), .Z(\b/n4637 ) );
  MUX \b/U4697  ( .IN0(\b/n4635 ), .IN1(\b/n4633 ), .SEL(msg[74]), .F(
        \b/n4636 ) );
  MUX \b/U4696  ( .IN0(\b/n449 ), .IN1(\b/n4634 ), .SEL(msg[79]), .F(\b/n4635 ) );
  MUX \b/U4695  ( .IN0(\b/n476 ), .IN1(\b/n466 ), .SEL(msg[73]), .F(\b/n4634 )
         );
  MUX \b/U4694  ( .IN0(\b/n438 ), .IN1(\b/n4379 ), .SEL(msg[79]), .F(\b/n4633 ) );
  NANDN \b/U4693  ( .B(\b/n439 ), .A(msg[73]), .Z(\b/n4379 ) );
  MUX \b/U4692  ( .IN0(\b/n4632 ), .IN1(\b/n4611 ), .SEL(msg[78]), .F(
        shift_row_out[45]) );
  MUX \b/U4691  ( .IN0(\b/n4631 ), .IN1(\b/n4621 ), .SEL(msg[72]), .F(
        \b/n4632 ) );
  MUX \b/U4690  ( .IN0(\b/n4630 ), .IN1(\b/n4626 ), .SEL(msg[77]), .F(
        \b/n4631 ) );
  MUX \b/U4689  ( .IN0(\b/n4627 ), .IN1(\b/n4628 ), .SEL(msg[74]), .F(
        \b/n4630 ) );
  AND \b/U4688  ( .A(\b/n4397 ), .B(\b/n4629 ), .Z(\b/n4628 ) );
  MUX \b/U4687  ( .IN0(\b/n4375 ), .IN1(\b/n487 ), .SEL(msg[79]), .F(\b/n4627 ) );
  MUX \b/U4686  ( .IN0(\b/n4625 ), .IN1(\b/n4623 ), .SEL(msg[74]), .F(
        \b/n4626 ) );
  MUX \b/U4685  ( .IN0(\b/n442 ), .IN1(\b/n4624 ), .SEL(msg[79]), .F(\b/n4625 ) );
  NAND \b/U4684  ( .A(\b/n466 ), .B(\b/n496 ), .Z(\b/n4624 ) );
  MUX \b/U4683  ( .IN0(\b/n4375 ), .IN1(\b/n4622 ), .SEL(msg[79]), .F(
        \b/n4623 ) );
  NAND \b/U4682  ( .A(\b/n4366 ), .B(\b/n4427 ), .Z(\b/n4622 ) );
  MUX \b/U4681  ( .IN0(\b/n4620 ), .IN1(\b/n4616 ), .SEL(msg[77]), .F(
        \b/n4621 ) );
  MUX \b/U4680  ( .IN0(\b/n4619 ), .IN1(\b/n4618 ), .SEL(msg[74]), .F(
        \b/n4620 ) );
  MUX \b/U4679  ( .IN0(\b/n4387 ), .IN1(\b/n489 ), .SEL(msg[79]), .F(\b/n4619 ) );
  MUX \b/U4678  ( .IN0(\b/n4412 ), .IN1(\b/n4617 ), .SEL(msg[79]), .F(
        \b/n4618 ) );
  MUX \b/U4677  ( .IN0(\b/n485 ), .IN1(\b/n466 ), .SEL(msg[73]), .F(\b/n4617 )
         );
  MUX \b/U4676  ( .IN0(\b/n4615 ), .IN1(\b/n4614 ), .SEL(msg[74]), .F(
        \b/n4616 ) );
  MUX \b/U4675  ( .IN0(\b/n483 ), .IN1(n677), .SEL(msg[79]), .F(\b/n4615 ) );
  MUX \b/U4674  ( .IN0(\b/n4613 ), .IN1(\b/n4612 ), .SEL(msg[79]), .F(
        \b/n4614 ) );
  AND \b/U4673  ( .A(\b/n4372 ), .B(\b/n4447 ), .Z(\b/n4613 ) );
  MUX \b/U4672  ( .IN0(\b/n455 ), .IN1(\b/n439 ), .SEL(msg[73]), .F(\b/n4612 )
         );
  MUX \b/U4671  ( .IN0(\b/n4610 ), .IN1(\b/n4601 ), .SEL(msg[72]), .F(
        \b/n4611 ) );
  MUX \b/U4670  ( .IN0(\b/n4609 ), .IN1(\b/n4605 ), .SEL(msg[77]), .F(
        \b/n4610 ) );
  MUX \b/U4669  ( .IN0(\b/n4608 ), .IN1(\b/n4606 ), .SEL(msg[74]), .F(
        \b/n4609 ) );
  MUX \b/U4668  ( .IN0(\b/n4378 ), .IN1(\b/n4607 ), .SEL(msg[79]), .F(
        \b/n4608 ) );
  NAND \b/U4667  ( .A(msg[73]), .B(\b/n455 ), .Z(\b/n4607 ) );
  MUX \b/U4666  ( .IN0(\b/n439 ), .IN1(\b/n492 ), .SEL(msg[79]), .F(\b/n4606 )
         );
  MUX \b/U4665  ( .IN0(\b/n4604 ), .IN1(\b/n4603 ), .SEL(msg[74]), .F(
        \b/n4605 ) );
  MUX \b/U4664  ( .IN0(\b/n4404 ), .IN1(\b/n457 ), .SEL(msg[79]), .F(\b/n4604 ) );
  MUX \b/U4663  ( .IN0(\b/n4602 ), .IN1(\b/n4367 ), .SEL(n676), .F(\b/n4603 )
         );
  AND \b/U4662  ( .A(msg[79]), .B(msg[75]), .Z(\b/n4602 ) );
  MUX \b/U4661  ( .IN0(\b/n4600 ), .IN1(\b/n4597 ), .SEL(msg[77]), .F(
        \b/n4601 ) );
  MUX \b/U4660  ( .IN0(\b/n4599 ), .IN1(\b/n4598 ), .SEL(msg[74]), .F(
        \b/n4600 ) );
  MUX \b/U4659  ( .IN0(\b/n4528 ), .IN1(\b/n4367 ), .SEL(msg[79]), .F(
        \b/n4599 ) );
  MUX \b/U4658  ( .IN0(n675), .IN1(\b/n490 ), .SEL(msg[79]), .F(\b/n4598 ) );
  MUX \b/U4657  ( .IN0(\b/n4595 ), .IN1(\b/n4594 ), .SEL(msg[74]), .F(
        \b/n4597 ) );
  AND \b/U4656  ( .A(\b/n4596 ), .B(\b/n4496 ), .Z(\b/n4595 ) );
  MUX \b/U4655  ( .IN0(\b/n441 ), .IN1(\b/n485 ), .SEL(msg[79]), .F(\b/n4594 )
         );
  MUX \b/U4654  ( .IN0(\b/n4593 ), .IN1(\b/n4576 ), .SEL(msg[78]), .F(
        shift_row_out[44]) );
  MUX \b/U4653  ( .IN0(\b/n4592 ), .IN1(\b/n4584 ), .SEL(msg[72]), .F(
        \b/n4593 ) );
  MUX \b/U4652  ( .IN0(\b/n4591 ), .IN1(\b/n4588 ), .SEL(msg[77]), .F(
        \b/n4592 ) );
  MUX \b/U4651  ( .IN0(\b/n4590 ), .IN1(\b/n4589 ), .SEL(msg[74]), .F(
        \b/n4591 ) );
  MUX \b/U4650  ( .IN0(\b/n467 ), .IN1(\b/n488 ), .SEL(msg[79]), .F(\b/n4590 )
         );
  MUX \b/U4649  ( .IN0(\b/n4447 ), .IN1(\b/n4412 ), .SEL(msg[79]), .F(
        \b/n4589 ) );
  NAND \b/U4648  ( .A(msg[73]), .B(\b/n4366 ), .Z(\b/n4447 ) );
  MUX \b/U4647  ( .IN0(\b/n4585 ), .IN1(\b/n4586 ), .SEL(msg[74]), .F(
        \b/n4588 ) );
  AND \b/U4646  ( .A(\b/n4397 ), .B(\b/n4587 ), .Z(\b/n4586 ) );
  MUX \b/U4645  ( .IN0(\b/n4395 ), .IN1(\b/n470 ), .SEL(msg[79]), .F(\b/n4585 ) );
  MUX \b/U4644  ( .IN0(\b/n4583 ), .IN1(\b/n4580 ), .SEL(msg[77]), .F(
        \b/n4584 ) );
  MUX \b/U4643  ( .IN0(\b/n4582 ), .IN1(\b/n4581 ), .SEL(msg[74]), .F(
        \b/n4583 ) );
  MUX \b/U4642  ( .IN0(\b/n432 ), .IN1(\b/n478 ), .SEL(msg[79]), .F(\b/n4582 )
         );
  MUX \b/U4641  ( .IN0(\b/n439 ), .IN1(\b/n4375 ), .SEL(msg[79]), .F(\b/n4581 ) );
  MUX \b/U4640  ( .IN0(\b/n4579 ), .IN1(\b/n4577 ), .SEL(msg[74]), .F(
        \b/n4580 ) );
  MUX \b/U4639  ( .IN0(\b/n4391 ), .IN1(\b/n4578 ), .SEL(msg[79]), .F(
        \b/n4579 ) );
  AND \b/U4638  ( .A(\b/n4375 ), .B(\b/n496 ), .Z(\b/n4578 ) );
  MUX \b/U4637  ( .IN0(\b/n454 ), .IN1(\b/n473 ), .SEL(msg[79]), .F(\b/n4577 )
         );
  MUX \b/U4636  ( .IN0(\b/n4575 ), .IN1(\b/n4569 ), .SEL(msg[72]), .F(
        \b/n4576 ) );
  MUX \b/U4635  ( .IN0(\b/n4574 ), .IN1(\b/n4572 ), .SEL(msg[77]), .F(
        \b/n4575 ) );
  MUX \b/U4634  ( .IN0(\b/n4573 ), .IN1(\b/n4369 ), .SEL(msg[74]), .F(
        \b/n4574 ) );
  MUX \b/U4633  ( .IN0(\b/n4389 ), .IN1(\b/n475 ), .SEL(msg[79]), .F(\b/n4573 ) );
  MUX \b/U4632  ( .IN0(\b/n4571 ), .IN1(\b/n4570 ), .SEL(msg[74]), .F(
        \b/n4572 ) );
  MUX \b/U4631  ( .IN0(n674), .IN1(\b/n467 ), .SEL(msg[79]), .F(\b/n4571 ) );
  MUX \b/U4630  ( .IN0(\b/n4399 ), .IN1(\b/n4402 ), .SEL(msg[79]), .F(
        \b/n4570 ) );
  MUX \b/U4629  ( .IN0(\b/n4568 ), .IN1(\b/n4565 ), .SEL(msg[77]), .F(
        \b/n4569 ) );
  MUX \b/U4628  ( .IN0(\b/n4567 ), .IN1(\b/n4566 ), .SEL(msg[74]), .F(
        \b/n4568 ) );
  MUX \b/U4627  ( .IN0(\b/n440 ), .IN1(\b/n4371 ), .SEL(msg[79]), .F(\b/n4567 ) );
  MUX \b/U4626  ( .IN0(\b/n485 ), .IN1(\b/n4393 ), .SEL(msg[79]), .F(\b/n4566 ) );
  MUX \b/U4625  ( .IN0(\b/n428 ), .IN1(\b/n4564 ), .SEL(msg[74]), .F(\b/n4565 ) );
  MUX \b/U4624  ( .IN0(\b/n448 ), .IN1(\b/n4375 ), .SEL(msg[79]), .F(\b/n4564 ) );
  MUX \b/U4623  ( .IN0(\b/n4563 ), .IN1(\b/n4544 ), .SEL(msg[78]), .F(
        shift_row_out[43]) );
  MUX \b/U4622  ( .IN0(\b/n4562 ), .IN1(\b/n4554 ), .SEL(msg[72]), .F(
        \b/n4563 ) );
  MUX \b/U4621  ( .IN0(\b/n4561 ), .IN1(\b/n4558 ), .SEL(msg[77]), .F(
        \b/n4562 ) );
  MUX \b/U4620  ( .IN0(\b/n4560 ), .IN1(\b/n4559 ), .SEL(msg[79]), .F(
        \b/n4561 ) );
  MUX \b/U4619  ( .IN0(\b/n4383 ), .IN1(\b/n473 ), .SEL(msg[74]), .F(\b/n4560 ) );
  MUX \b/U4618  ( .IN0(n677), .IN1(\b/n431 ), .SEL(msg[74]), .F(\b/n4559 ) );
  MUX \b/U4617  ( .IN0(\b/n4556 ), .IN1(\b/n4555 ), .SEL(msg[79]), .F(
        \b/n4558 ) );
  AND \b/U4616  ( .A(\b/n4557 ), .B(msg[76]), .Z(\b/n4556 ) );
  MUX \b/U4615  ( .IN0(\b/n461 ), .IN1(\b/n4396 ), .SEL(msg[74]), .F(\b/n4555 ) );
  MUX \b/U4614  ( .IN0(\b/n4553 ), .IN1(\b/n4550 ), .SEL(msg[77]), .F(
        \b/n4554 ) );
  MUX \b/U4613  ( .IN0(\b/n4552 ), .IN1(\b/n4551 ), .SEL(msg[79]), .F(
        \b/n4553 ) );
  MUX \b/U4612  ( .IN0(\b/n4387 ), .IN1(n673), .SEL(msg[74]), .F(\b/n4552 ) );
  MUX \b/U4611  ( .IN0(\b/n429 ), .IN1(\b/n448 ), .SEL(msg[74]), .F(\b/n4551 )
         );
  MUX \b/U4610  ( .IN0(\b/n4546 ), .IN1(\b/n4547 ), .SEL(msg[79]), .F(
        \b/n4550 ) );
  NAND \b/U4609  ( .A(\b/n4548 ), .B(\b/n4549 ), .Z(\b/n4547 ) );
  MUX \b/U4608  ( .IN0(\b/n474 ), .IN1(\b/n4545 ), .SEL(msg[74]), .F(\b/n4546 ) );
  MUX \b/U4607  ( .IN0(\b/n449 ), .IN1(\b/n491 ), .SEL(msg[73]), .F(\b/n4545 )
         );
  MUX \b/U4606  ( .IN0(\b/n4543 ), .IN1(\b/n4534 ), .SEL(msg[72]), .F(
        \b/n4544 ) );
  MUX \b/U4605  ( .IN0(\b/n4542 ), .IN1(\b/n4538 ), .SEL(msg[77]), .F(
        \b/n4543 ) );
  MUX \b/U4604  ( .IN0(\b/n4540 ), .IN1(\b/n4539 ), .SEL(msg[79]), .F(
        \b/n4542 ) );
  NAND \b/U4603  ( .A(\b/n439 ), .B(\b/n4541 ), .Z(\b/n4540 ) );
  MUX \b/U4602  ( .IN0(\b/n490 ), .IN1(\b/n452 ), .SEL(msg[74]), .F(\b/n4539 )
         );
  MUX \b/U4601  ( .IN0(\b/n4537 ), .IN1(\b/n4535 ), .SEL(msg[79]), .F(
        \b/n4538 ) );
  MUX \b/U4600  ( .IN0(\b/n4378 ), .IN1(\b/n4536 ), .SEL(msg[74]), .F(
        \b/n4537 ) );
  AND \b/U4599  ( .A(msg[73]), .B(\b/n439 ), .Z(\b/n4536 ) );
  MUX \b/U4598  ( .IN0(\b/n444 ), .IN1(\b/n4397 ), .SEL(msg[74]), .F(\b/n4535 ) );
  MUX \b/U4597  ( .IN0(\b/n4533 ), .IN1(\b/n4527 ), .SEL(msg[77]), .F(
        \b/n4534 ) );
  MUX \b/U4596  ( .IN0(\b/n4532 ), .IN1(\b/n4530 ), .SEL(msg[79]), .F(
        \b/n4533 ) );
  MUX \b/U4595  ( .IN0(\b/n4531 ), .IN1(\b/n4367 ), .SEL(\b/n4415 ), .F(
        \b/n4532 ) );
  MUX \b/U4594  ( .IN0(msg[75]), .IN1(msg[76]), .SEL(msg[74]), .F(\b/n4531 )
         );
  MUX \b/U4593  ( .IN0(\b/n4397 ), .IN1(\b/n4528 ), .SEL(msg[74]), .F(
        \b/n4530 ) );
  NAND \b/U4592  ( .A(\b/n4367 ), .B(\b/n4529 ), .Z(\b/n4528 ) );
  MUX \b/U4591  ( .IN0(\b/n4524 ), .IN1(\b/n4525 ), .SEL(msg[79]), .F(
        \b/n4527 ) );
  AND \b/U4590  ( .A(\b/n472 ), .B(\b/n4526 ), .Z(\b/n4525 ) );
  MUX \b/U4589  ( .IN0(\b/n453 ), .IN1(\b/n4368 ), .SEL(msg[74]), .F(\b/n4524 ) );
  MUX \b/U4588  ( .IN0(\b/n4523 ), .IN1(\b/n4507 ), .SEL(msg[78]), .F(
        shift_row_out[42]) );
  MUX \b/U4587  ( .IN0(\b/n4522 ), .IN1(\b/n4514 ), .SEL(msg[72]), .F(
        \b/n4523 ) );
  MUX \b/U4586  ( .IN0(\b/n4521 ), .IN1(\b/n4517 ), .SEL(msg[77]), .F(
        \b/n4522 ) );
  MUX \b/U4585  ( .IN0(\b/n4520 ), .IN1(\b/n4518 ), .SEL(msg[74]), .F(
        \b/n4521 ) );
  MUX \b/U4584  ( .IN0(\b/n461 ), .IN1(\b/n4519 ), .SEL(msg[79]), .F(\b/n4520 ) );
  MUX \b/U4583  ( .IN0(\b/n4375 ), .IN1(\b/n439 ), .SEL(msg[73]), .F(\b/n4519 ) );
  MUX \b/U4582  ( .IN0(\b/n4414 ), .IN1(\b/n479 ), .SEL(msg[79]), .F(\b/n4518 ) );
  MUX \b/U4581  ( .IN0(\b/n4516 ), .IN1(\b/n4515 ), .SEL(msg[74]), .F(
        \b/n4517 ) );
  MUX \b/U4580  ( .IN0(\b/n4368 ), .IN1(\b/n446 ), .SEL(msg[79]), .F(\b/n4516 ) );
  MUX \b/U4579  ( .IN0(\b/n482 ), .IN1(\b/n4401 ), .SEL(msg[79]), .F(\b/n4515 ) );
  MUX \b/U4578  ( .IN0(\b/n4513 ), .IN1(\b/n4509 ), .SEL(msg[77]), .F(
        \b/n4514 ) );
  MUX \b/U4577  ( .IN0(\b/n4510 ), .IN1(\b/n428 ), .SEL(msg[74]), .F(\b/n4513 ) );
  NAND \b/U4576  ( .A(\b/n4511 ), .B(\b/n4512 ), .Z(\b/n4510 ) );
  MUX \b/U4575  ( .IN0(n675), .IN1(\b/n4508 ), .SEL(\b/n4413 ), .F(\b/n4509 )
         );
  MUX \b/U4574  ( .IN0(\b/n460 ), .IN1(\b/n4380 ), .SEL(msg[74]), .F(\b/n4508 ) );
  MUX \b/U4573  ( .IN0(\b/n4506 ), .IN1(\b/n4498 ), .SEL(msg[72]), .F(
        \b/n4507 ) );
  MUX \b/U4572  ( .IN0(\b/n4505 ), .IN1(\b/n4502 ), .SEL(msg[77]), .F(
        \b/n4506 ) );
  MUX \b/U4571  ( .IN0(\b/n4504 ), .IN1(\b/n4503 ), .SEL(msg[74]), .F(
        \b/n4505 ) );
  MUX \b/U4570  ( .IN0(\b/n488 ), .IN1(msg[73]), .SEL(msg[79]), .F(\b/n4504 )
         );
  MUX \b/U4569  ( .IN0(n678), .IN1(\b/n4381 ), .SEL(msg[79]), .F(\b/n4503 ) );
  MUX \b/U4568  ( .IN0(\b/n4501 ), .IN1(\b/n4500 ), .SEL(msg[74]), .F(
        \b/n4502 ) );
  MUX \b/U4567  ( .IN0(\b/n493 ), .IN1(\b/n487 ), .SEL(msg[79]), .F(\b/n4501 )
         );
  MUX \b/U4566  ( .IN0(n678), .IN1(\b/n4499 ), .SEL(msg[79]), .F(\b/n4500 ) );
  MUX \b/U4565  ( .IN0(\b/n439 ), .IN1(\b/n476 ), .SEL(msg[73]), .F(\b/n4499 )
         );
  MUX \b/U4564  ( .IN0(\b/n4497 ), .IN1(\b/n4491 ), .SEL(msg[77]), .F(
        \b/n4498 ) );
  MUX \b/U4563  ( .IN0(\b/n4494 ), .IN1(\b/n4493 ), .SEL(msg[74]), .F(
        \b/n4497 ) );
  NAND \b/U4562  ( .A(\b/n4495 ), .B(\b/n4496 ), .Z(\b/n4494 ) );
  MUX \b/U4561  ( .IN0(\b/n4367 ), .IN1(\b/n4492 ), .SEL(n676), .F(\b/n4493 )
         );
  MUX \b/U4560  ( .IN0(msg[75]), .IN1(\b/n449 ), .SEL(msg[79]), .F(\b/n4492 )
         );
  MUX \b/U4559  ( .IN0(\b/n4490 ), .IN1(\b/n4489 ), .SEL(msg[74]), .F(
        \b/n4491 ) );
  MUX \b/U4558  ( .IN0(\b/n4412 ), .IN1(\b/n447 ), .SEL(msg[79]), .F(\b/n4490 ) );
  MUX \b/U4557  ( .IN0(\b/n4408 ), .IN1(\b/n4488 ), .SEL(msg[79]), .F(
        \b/n4489 ) );
  MUX \b/U4556  ( .IN0(\b/n4370 ), .IN1(\b/n4375 ), .SEL(msg[73]), .F(
        \b/n4488 ) );
  MUX \b/U4555  ( .IN0(\b/n4487 ), .IN1(\b/n4469 ), .SEL(msg[78]), .F(
        shift_row_out[41]) );
  MUX \b/U4554  ( .IN0(\b/n4486 ), .IN1(\b/n4477 ), .SEL(msg[72]), .F(
        \b/n4487 ) );
  MUX \b/U4553  ( .IN0(\b/n4485 ), .IN1(\b/n4481 ), .SEL(msg[77]), .F(
        \b/n4486 ) );
  MUX \b/U4552  ( .IN0(\b/n4484 ), .IN1(\b/n4483 ), .SEL(msg[74]), .F(
        \b/n4485 ) );
  MUX \b/U4551  ( .IN0(\b/n484 ), .IN1(n680), .SEL(msg[79]), .F(\b/n4484 ) );
  MUX \b/U4550  ( .IN0(\b/n4482 ), .IN1(n674), .SEL(msg[79]), .F(\b/n4483 ) );
  NAND \b/U4549  ( .A(\b/n496 ), .B(\b/n455 ), .Z(\b/n4482 ) );
  MUX \b/U4548  ( .IN0(\b/n4480 ), .IN1(\b/n4479 ), .SEL(msg[74]), .F(
        \b/n4481 ) );
  MUX \b/U4547  ( .IN0(\b/n432 ), .IN1(\b/n4382 ), .SEL(msg[79]), .F(\b/n4480 ) );
  MUX \b/U4546  ( .IN0(\b/n4372 ), .IN1(\b/n4478 ), .SEL(msg[79]), .F(
        \b/n4479 ) );
  AND \b/U4545  ( .A(msg[73]), .B(msg[76]), .Z(\b/n4478 ) );
  MUX \b/U4544  ( .IN0(\b/n4476 ), .IN1(\b/n4473 ), .SEL(msg[77]), .F(
        \b/n4477 ) );
  MUX \b/U4543  ( .IN0(\b/n4475 ), .IN1(\b/n4474 ), .SEL(msg[74]), .F(
        \b/n4476 ) );
  MUX \b/U4542  ( .IN0(\b/n4411 ), .IN1(\b/n493 ), .SEL(msg[79]), .F(\b/n4475 ) );
  MUX \b/U4541  ( .IN0(\b/n468 ), .IN1(\b/n4380 ), .SEL(msg[79]), .F(\b/n4474 ) );
  MUX \b/U4540  ( .IN0(\b/n4470 ), .IN1(\b/n4471 ), .SEL(msg[74]), .F(
        \b/n4473 ) );
  AND \b/U4539  ( .A(\b/n4472 ), .B(\b/n4427 ), .Z(\b/n4471 ) );
  MUX \b/U4538  ( .IN0(\b/n4386 ), .IN1(\b/n4375 ), .SEL(msg[79]), .F(
        \b/n4470 ) );
  MUX \b/U4537  ( .IN0(\b/n4468 ), .IN1(\b/n4460 ), .SEL(msg[72]), .F(
        \b/n4469 ) );
  MUX \b/U4536  ( .IN0(\b/n4467 ), .IN1(\b/n4463 ), .SEL(msg[77]), .F(
        \b/n4468 ) );
  MUX \b/U4535  ( .IN0(\b/n4466 ), .IN1(\b/n4465 ), .SEL(msg[74]), .F(
        \b/n4467 ) );
  MUX \b/U4534  ( .IN0(\b/n4374 ), .IN1(\b/n457 ), .SEL(msg[79]), .F(\b/n4466 ) );
  MUX \b/U4533  ( .IN0(\b/n4464 ), .IN1(\b/n441 ), .SEL(msg[79]), .F(\b/n4465 ) );
  MUX \b/U4532  ( .IN0(\b/n4372 ), .IN1(\b/n449 ), .SEL(msg[73]), .F(\b/n4464 ) );
  MUX \b/U4531  ( .IN0(\b/n4462 ), .IN1(\b/n4461 ), .SEL(msg[74]), .F(
        \b/n4463 ) );
  MUX \b/U4530  ( .IN0(\b/n488 ), .IN1(\b/n466 ), .SEL(msg[79]), .F(\b/n4462 )
         );
  MUX \b/U4529  ( .IN0(\b/n484 ), .IN1(\b/n444 ), .SEL(msg[79]), .F(\b/n4461 )
         );
  MUX \b/U4528  ( .IN0(\b/n4459 ), .IN1(\b/n4454 ), .SEL(msg[77]), .F(
        \b/n4460 ) );
  MUX \b/U4527  ( .IN0(\b/n4458 ), .IN1(\b/n4455 ), .SEL(msg[74]), .F(
        \b/n4459 ) );
  MUX \b/U4526  ( .IN0(\b/n4456 ), .IN1(\b/n4457 ), .SEL(msg[79]), .F(
        \b/n4458 ) );
  NAND \b/U4525  ( .A(\b/n4375 ), .B(\b/n4447 ), .Z(\b/n4457 ) );
  MUX \b/U4524  ( .IN0(\b/n4375 ), .IN1(\b/n449 ), .SEL(msg[73]), .F(\b/n4456 ) );
  MUX \b/U4523  ( .IN0(\b/n4392 ), .IN1(\b/n4390 ), .SEL(msg[79]), .F(
        \b/n4455 ) );
  MUX \b/U4522  ( .IN0(\b/n4410 ), .IN1(\b/n4453 ), .SEL(msg[74]), .F(
        \b/n4454 ) );
  MUX \b/U4521  ( .IN0(\b/n455 ), .IN1(\b/n487 ), .SEL(msg[79]), .F(\b/n4453 )
         );
  MUX \b/U4520  ( .IN0(\b/n4452 ), .IN1(\b/n4435 ), .SEL(msg[78]), .F(
        shift_row_out[40]) );
  MUX \b/U4519  ( .IN0(\b/n4451 ), .IN1(\b/n4443 ), .SEL(msg[72]), .F(
        \b/n4452 ) );
  MUX \b/U4518  ( .IN0(\b/n4450 ), .IN1(\b/n4448 ), .SEL(msg[74]), .F(
        \b/n4451 ) );
  MUX \b/U4517  ( .IN0(\b/n429 ), .IN1(\b/n4449 ), .SEL(msg[79]), .F(\b/n4450 ) );
  MUX \b/U4516  ( .IN0(\b/n482 ), .IN1(\b/n485 ), .SEL(msg[77]), .F(\b/n4449 )
         );
  MUX \b/U4515  ( .IN0(\b/n4445 ), .IN1(\b/n4444 ), .SEL(msg[79]), .F(
        \b/n4448 ) );
  NAND \b/U4514  ( .A(\b/n4446 ), .B(\b/n4447 ), .Z(\b/n4445 ) );
  MUX \b/U4513  ( .IN0(\b/n481 ), .IN1(\b/n496 ), .SEL(msg[77]), .F(\b/n4444 )
         );
  MUX \b/U4512  ( .IN0(\b/n4442 ), .IN1(\b/n4438 ), .SEL(msg[74]), .F(
        \b/n4443 ) );
  MUX \b/U4511  ( .IN0(\b/n4441 ), .IN1(\b/n4439 ), .SEL(msg[79]), .F(
        \b/n4442 ) );
  MUX \b/U4510  ( .IN0(\b/n4440 ), .IN1(\b/n434 ), .SEL(msg[77]), .F(\b/n4441 ) );
  NAND \b/U4509  ( .A(\b/n496 ), .B(\b/n4367 ), .Z(\b/n4440 ) );
  MUX \b/U4507  ( .IN0(\b/n4437 ), .IN1(\b/n4436 ), .SEL(msg[79]), .F(
        \b/n4438 ) );
  MUX \b/U4506  ( .IN0(n675), .IN1(\b/n431 ), .SEL(msg[77]), .F(\b/n4437 ) );
  MUX \b/U4505  ( .IN0(\b/n483 ), .IN1(\b/n439 ), .SEL(msg[77]), .F(\b/n4436 )
         );
  MUX \b/U4504  ( .IN0(\b/n4434 ), .IN1(\b/n4424 ), .SEL(msg[72]), .F(
        \b/n4435 ) );
  MUX \b/U4503  ( .IN0(\b/n4433 ), .IN1(\b/n4429 ), .SEL(msg[74]), .F(
        \b/n4434 ) );
  MUX \b/U4502  ( .IN0(\b/n4432 ), .IN1(\b/n4431 ), .SEL(msg[79]), .F(
        \b/n4433 ) );
  MUX \b/U4501  ( .IN0(n673), .IN1(\b/n435 ), .SEL(msg[77]), .F(\b/n4432 ) );
  MUX \b/U4500  ( .IN0(\b/n4430 ), .IN1(\b/n472 ), .SEL(msg[77]), .F(\b/n4431 ) );
  NAND \b/U4499  ( .A(\b/n4366 ), .B(\b/n4368 ), .Z(\b/n4430 ) );
  MUX \b/U4498  ( .IN0(\b/n4428 ), .IN1(\b/n4425 ), .SEL(msg[79]), .F(
        \b/n4429 ) );
  MUX \b/U4497  ( .IN0(\b/n442 ), .IN1(\b/n4426 ), .SEL(msg[77]), .F(\b/n4428 ) );
  NAND \b/U4496  ( .A(\b/n4370 ), .B(\b/n4427 ), .Z(\b/n4426 ) );
  MUX \b/U4495  ( .IN0(\b/n4385 ), .IN1(\b/n4376 ), .SEL(msg[77]), .F(
        \b/n4425 ) );
  MUX \b/U4494  ( .IN0(\b/n4423 ), .IN1(\b/n4419 ), .SEL(msg[74]), .F(
        \b/n4424 ) );
  MUX \b/U4493  ( .IN0(\b/n4421 ), .IN1(\b/n4420 ), .SEL(msg[79]), .F(
        \b/n4423 ) );
  NAND \b/U4492  ( .A(\b/n4422 ), .B(\b/n4409 ), .Z(\b/n4421 ) );
  MUX \b/U4491  ( .IN0(msg[75]), .IN1(\b/n4401 ), .SEL(msg[77]), .F(\b/n4420 )
         );
  MUX \b/U4490  ( .IN0(\b/n4418 ), .IN1(\b/n4417 ), .SEL(msg[79]), .F(
        \b/n4419 ) );
  MUX \b/U4489  ( .IN0(\b/n447 ), .IN1(\b/n463 ), .SEL(msg[77]), .F(\b/n4418 )
         );
  MUX \b/U4488  ( .IN0(\b/n480 ), .IN1(\b/n468 ), .SEL(msg[77]), .F(\b/n4417 )
         );
  XOR \b/U4487  ( .A(\b/n4367 ), .B(msg[73]), .Z(\b/n4416 ) );
  XOR \b/U4486  ( .A(msg[73]), .B(msg[74]), .Z(\b/n4415 ) );
  XOR \b/U4485  ( .A(msg[73]), .B(msg[75]), .Z(\b/n4414 ) );
  XOR \b/U4484  ( .A(msg[74]), .B(msg[79]), .Z(\b/n4413 ) );
  XOR \b/U4483  ( .A(\b/n496 ), .B(\b/n439 ), .Z(\b/n4412 ) );
  XOR \b/U4482  ( .A(msg[73]), .B(\b/n485 ), .Z(\b/n4411 ) );
  XOR \b/U4480  ( .A(msg[73]), .B(msg[77]), .Z(\b/n4409 ) );
  NAND \b/U4479  ( .A(msg[73]), .B(msg[75]), .Z(\b/n4408 ) );
  MUX \b/U4478  ( .IN0(\b/n4367 ), .IN1(\b/n439 ), .SEL(msg[73]), .F(\b/n4407 ) );
  MUX \b/U4476  ( .IN0(msg[75]), .IN1(\b/n476 ), .SEL(msg[73]), .F(\b/n4405 )
         );
  MUX \b/U4475  ( .IN0(\b/n455 ), .IN1(\b/n476 ), .SEL(msg[73]), .F(\b/n4404 )
         );
  MUX \b/U4474  ( .IN0(\b/n4370 ), .IN1(\b/n4372 ), .SEL(msg[73]), .F(
        \b/n4403 ) );
  MUX \b/U4473  ( .IN0(msg[76]), .IN1(\b/n455 ), .SEL(msg[73]), .F(\b/n4402 )
         );
  OR \b/U4472  ( .A(msg[73]), .B(msg[76]), .Z(\b/n4401 ) );
  NAND \b/U4470  ( .A(\b/n476 ), .B(\b/n496 ), .Z(\b/n4399 ) );
  MUX \b/U4469  ( .IN0(\b/n476 ), .IN1(msg[76]), .SEL(msg[73]), .F(\b/n4398 )
         );
  MUX \b/U4468  ( .IN0(\b/n4366 ), .IN1(\b/n4375 ), .SEL(msg[73]), .F(
        \b/n4397 ) );
  MUX \b/U4467  ( .IN0(\b/n491 ), .IN1(msg[76]), .SEL(msg[73]), .F(\b/n4396 )
         );
  MUX \b/U4466  ( .IN0(\b/n449 ), .IN1(\b/n476 ), .SEL(msg[73]), .F(\b/n4395 )
         );
  MUX \b/U4465  ( .IN0(\b/n4366 ), .IN1(msg[76]), .SEL(msg[73]), .F(\b/n4394 )
         );
  MUX \b/U4464  ( .IN0(\b/n466 ), .IN1(\b/n455 ), .SEL(msg[73]), .F(\b/n4393 )
         );
  XOR \b/U4463  ( .A(\b/n449 ), .B(msg[73]), .Z(\b/n4392 ) );
  MUX \b/U4462  ( .IN0(\b/n4372 ), .IN1(\b/n466 ), .SEL(msg[73]), .F(\b/n4391 ) );
  NANDN \b/U4461  ( .B(msg[73]), .A(msg[75]), .Z(\b/n4390 ) );
  MUX \b/U4460  ( .IN0(\b/n439 ), .IN1(msg[75]), .SEL(msg[73]), .F(\b/n4389 )
         );
  NAND \b/U4458  ( .A(\b/n4370 ), .B(\b/n496 ), .Z(\b/n4387 ) );
  MUX \b/U4457  ( .IN0(msg[76]), .IN1(\b/n4367 ), .SEL(msg[73]), .F(\b/n4386 )
         );
  MUX \b/U4456  ( .IN0(\b/n466 ), .IN1(msg[75]), .SEL(msg[73]), .F(\b/n4385 )
         );
  MUX \b/U4454  ( .IN0(msg[76]), .IN1(\b/n485 ), .SEL(msg[73]), .F(\b/n4383 )
         );
  MUX \b/U4453  ( .IN0(\b/n439 ), .IN1(\b/n491 ), .SEL(msg[73]), .F(\b/n4382 )
         );
  NAND \b/U4452  ( .A(\b/n4368 ), .B(\b/n439 ), .Z(\b/n4381 ) );
  MUX \b/U4451  ( .IN0(\b/n4367 ), .IN1(\b/n4375 ), .SEL(msg[73]), .F(
        \b/n4380 ) );
  NAND \b/U4450  ( .A(\b/n4379 ), .B(\b/n4366 ), .Z(\b/n4378 ) );
  MUX \b/U4449  ( .IN0(\b/n4370 ), .IN1(\b/n491 ), .SEL(msg[73]), .F(\b/n4377 ) );
  MUX \b/U4448  ( .IN0(\b/n491 ), .IN1(\b/n455 ), .SEL(msg[73]), .F(\b/n4376 )
         );
  NANDN \b/U4447  ( .B(msg[75]), .A(msg[76]), .Z(\b/n4375 ) );
  MUX \b/U4446  ( .IN0(\b/n4370 ), .IN1(msg[75]), .SEL(msg[73]), .F(\b/n4374 )
         );
  OR \b/U4445  ( .A(msg[75]), .B(msg[76]), .Z(\b/n4370 ) );
  MUX \b/U4444  ( .IN0(\b/n439 ), .IN1(\b/n455 ), .SEL(msg[73]), .F(\b/n4373 )
         );
  XOR \b/U4443  ( .A(\b/n449 ), .B(msg[75]), .Z(\b/n4372 ) );
  NANDN \b/U4442  ( .B(msg[75]), .A(msg[73]), .Z(\b/n4371 ) );
  NAND \b/U4441  ( .A(\b/n4370 ), .B(\b/n4368 ), .Z(\b/n4369 ) );
  NAND \b/U4440  ( .A(msg[73]), .B(\b/n4367 ), .Z(\b/n4368 ) );
  NANDN \b/U4439  ( .B(msg[76]), .A(msg[75]), .Z(\b/n4367 ) );
  NAND \b/U4438  ( .A(msg[75]), .B(msg[76]), .Z(\b/n4366 ) );
  MUX \b/U4437  ( .IN0(msg[68]), .IN1(\b/n4007 ), .SEL(msg[65]), .F(\b/n4365 )
         );
  MUX \b/U4436  ( .IN0(msg[68]), .IN1(\b/n4016 ), .SEL(msg[65]), .F(\b/n4364 )
         );
  MUX \b/U4435  ( .IN0(\b/n4008 ), .IN1(\b/n4011 ), .SEL(msg[65]), .F(
        \b/n4363 ) );
  MUX \b/U4434  ( .IN0(\b/n4013 ), .IN1(\b/n556 ), .SEL(msg[65]), .F(\b/n4362 ) );
  MUX \b/U4432  ( .IN0(\b/n4016 ), .IN1(\b/n4007 ), .SEL(msg[66]), .F(
        \b/n4189 ) );
  MUX \b/U4431  ( .IN0(\b/n4009 ), .IN1(\b/n567 ), .SEL(msg[66]), .F(\b/n4190 ) );
  MUX \b/U4430  ( .IN0(\b/n510 ), .IN1(\b/n520 ), .SEL(msg[65]), .F(\b/n4153 )
         );
  MUX \b/U4429  ( .IN0(\b/n4037 ), .IN1(\b/n4348 ), .SEL(msg[71]), .F(
        \b/n4360 ) );
  MUX \b/U4428  ( .IN0(\b/n4011 ), .IN1(\b/n4007 ), .SEL(msg[65]), .F(
        \b/n4351 ) );
  MUX \b/U4427  ( .IN0(\b/n562 ), .IN1(\b/n4013 ), .SEL(msg[65]), .F(\b/n4359 ) );
  MUX \b/U4426  ( .IN0(msg[67]), .IN1(\b/n556 ), .SEL(msg[65]), .F(\b/n4358 )
         );
  MUX \b/U4425  ( .IN0(\b/n4016 ), .IN1(\b/n562 ), .SEL(msg[65]), .F(\b/n4357 ) );
  MUX \b/U4424  ( .IN0(msg[68]), .IN1(\b/n4013 ), .SEL(msg[65]), .F(\b/n4356 )
         );
  MUX \b/U4423  ( .IN0(\b/n547 ), .IN1(\b/n526 ), .SEL(msg[69]), .F(\b/n4063 )
         );
  MUX \b/U4422  ( .IN0(\b/n4008 ), .IN1(\b/n520 ), .SEL(msg[65]), .F(\b/n4355 ) );
  NANDN \b/U4419  ( .B(\b/n4014 ), .A(msg[71]), .Z(\b/n4328 ) );
  NAND \b/U4418  ( .A(msg[71]), .B(\b/n523 ), .Z(\b/n4296 ) );
  NAND \b/U4417  ( .A(msg[71]), .B(\b/n535 ), .Z(\b/n4237 ) );
  NAND \b/U4416  ( .A(msg[71]), .B(\b/n4345 ), .Z(\b/n4270 ) );
  NAND \b/U4415  ( .A(msg[71]), .B(\b/n4265 ), .Z(\b/n4228 ) );
  NAND \b/U4413  ( .A(\b/n567 ), .B(\b/n556 ), .Z(\b/n4349 ) );
  NAND \b/U4412  ( .A(msg[71]), .B(\b/n4347 ), .Z(\b/n4342 ) );
  NAND \b/U4411  ( .A(n672), .B(msg[71]), .Z(\b/n4322 ) );
  NAND \b/U4409  ( .A(msg[66]), .B(\b/n4016 ), .Z(\b/n4182 ) );
  NAND \b/U4408  ( .A(\b/n556 ), .B(msg[65]), .Z(\b/n4137 ) );
  NAND \b/U4407  ( .A(msg[71]), .B(\b/n4351 ), .Z(\b/n4136 ) );
  NAND \b/U4405  ( .A(\b/n4349 ), .B(msg[71]), .Z(\b/n4152 ) );
  NAND \b/U4404  ( .A(\b/n4170 ), .B(\b/n4016 ), .Z(\b/n4348 ) );
  NANDN \b/U4403  ( .B(\b/n510 ), .A(\b/n567 ), .Z(\b/n4347 ) );
  NAND \b/U4401  ( .A(msg[65]), .B(\b/n4016 ), .Z(\b/n4068 ) );
  NAND \b/U4400  ( .A(\b/n510 ), .B(\b/n567 ), .Z(\b/n4345 ) );
  NAND \b/U4397  ( .A(msg[65]), .B(\b/n4011 ), .Z(\b/n4170 ) );
  ANDN \b/U4395  ( .A(msg[66]), .B(msg[65]), .Z(\b/n4198 ) );
  AND \b/U4394  ( .A(\b/n4008 ), .B(\b/n4342 ), .Z(\b/n4113 ) );
  MUX \b/U4393  ( .IN0(\b/n4341 ), .IN1(\b/n4325 ), .SEL(msg[70]), .F(
        shift_row_out[71]) );
  MUX \b/U4392  ( .IN0(\b/n4340 ), .IN1(\b/n4333 ), .SEL(msg[64]), .F(
        \b/n4341 ) );
  MUX \b/U4391  ( .IN0(\b/n4339 ), .IN1(\b/n4336 ), .SEL(msg[69]), .F(
        \b/n4340 ) );
  MUX \b/U4390  ( .IN0(\b/n4338 ), .IN1(\b/n4337 ), .SEL(msg[66]), .F(
        \b/n4339 ) );
  MUX \b/U4389  ( .IN0(msg[68]), .IN1(\b/n527 ), .SEL(msg[71]), .F(\b/n4338 )
         );
  MUX \b/U4388  ( .IN0(\b/n4009 ), .IN1(\b/n531 ), .SEL(msg[71]), .F(\b/n4337 ) );
  MUX \b/U4387  ( .IN0(\b/n4335 ), .IN1(\b/n4334 ), .SEL(msg[66]), .F(
        \b/n4336 ) );
  MUX \b/U4386  ( .IN0(\b/n4067 ), .IN1(\b/n523 ), .SEL(msg[71]), .F(\b/n4335 ) );
  MUX \b/U4385  ( .IN0(\b/n4019 ), .IN1(\b/n4030 ), .SEL(msg[71]), .F(
        \b/n4334 ) );
  MUX \b/U4384  ( .IN0(\b/n4332 ), .IN1(\b/n4329 ), .SEL(msg[69]), .F(
        \b/n4333 ) );
  MUX \b/U4383  ( .IN0(\b/n4331 ), .IN1(\b/n4330 ), .SEL(msg[66]), .F(
        \b/n4332 ) );
  MUX \b/U4382  ( .IN0(\b/n4043 ), .IN1(\b/n4018 ), .SEL(msg[71]), .F(
        \b/n4331 ) );
  MUX \b/U4381  ( .IN0(\b/n535 ), .IN1(\b/n4039 ), .SEL(msg[71]), .F(\b/n4330 ) );
  MUX \b/U4380  ( .IN0(\b/n4327 ), .IN1(\b/n4326 ), .SEL(msg[66]), .F(
        \b/n4329 ) );
  AND \b/U4379  ( .A(\b/n525 ), .B(\b/n4328 ), .Z(\b/n4327 ) );
  MUX \b/U4378  ( .IN0(\b/n4023 ), .IN1(n671), .SEL(msg[71]), .F(\b/n4326 ) );
  MUX \b/U4377  ( .IN0(\b/n4324 ), .IN1(\b/n4316 ), .SEL(msg[64]), .F(
        \b/n4325 ) );
  MUX \b/U4376  ( .IN0(\b/n4323 ), .IN1(\b/n4319 ), .SEL(msg[69]), .F(
        \b/n4324 ) );
  MUX \b/U4375  ( .IN0(\b/n4320 ), .IN1(\b/n4321 ), .SEL(msg[66]), .F(
        \b/n4323 ) );
  NAND \b/U4374  ( .A(\b/n4137 ), .B(\b/n4322 ), .Z(\b/n4321 ) );
  MUX \b/U4373  ( .IN0(\b/n565 ), .IN1(\b/n557 ), .SEL(msg[71]), .F(\b/n4320 )
         );
  MUX \b/U4372  ( .IN0(\b/n4318 ), .IN1(\b/n4317 ), .SEL(msg[66]), .F(
        \b/n4319 ) );
  MUX \b/U4371  ( .IN0(\b/n4013 ), .IN1(\b/n4007 ), .SEL(msg[71]), .F(
        \b/n4318 ) );
  MUX \b/U4370  ( .IN0(\b/n558 ), .IN1(\b/n4044 ), .SEL(msg[71]), .F(\b/n4317 ) );
  MUX \b/U4369  ( .IN0(\b/n4315 ), .IN1(\b/n4312 ), .SEL(msg[69]), .F(
        \b/n4316 ) );
  MUX \b/U4368  ( .IN0(\b/n4314 ), .IN1(\b/n4313 ), .SEL(msg[66]), .F(
        \b/n4315 ) );
  MUX \b/U4367  ( .IN0(\b/n4048 ), .IN1(\b/n4034 ), .SEL(msg[71]), .F(
        \b/n4314 ) );
  MUX \b/U4366  ( .IN0(\b/n511 ), .IN1(\b/n4016 ), .SEL(msg[71]), .F(\b/n4313 ) );
  MUX \b/U4365  ( .IN0(\b/n4311 ), .IN1(\b/n4310 ), .SEL(msg[66]), .F(
        \b/n4312 ) );
  MUX \b/U4364  ( .IN0(\b/n4049 ), .IN1(\b/n4057 ), .SEL(msg[71]), .F(
        \b/n4311 ) );
  MUX \b/U4363  ( .IN0(\b/n4042 ), .IN1(\b/n4309 ), .SEL(msg[71]), .F(
        \b/n4310 ) );
  MUX \b/U4362  ( .IN0(\b/n562 ), .IN1(\b/n520 ), .SEL(msg[65]), .F(\b/n4309 )
         );
  MUX \b/U4361  ( .IN0(\b/n4308 ), .IN1(\b/n4290 ), .SEL(msg[70]), .F(
        shift_row_out[70]) );
  MUX \b/U4360  ( .IN0(\b/n4307 ), .IN1(\b/n4298 ), .SEL(msg[64]), .F(
        \b/n4308 ) );
  MUX \b/U4359  ( .IN0(\b/n4306 ), .IN1(\b/n4301 ), .SEL(msg[69]), .F(
        \b/n4307 ) );
  MUX \b/U4358  ( .IN0(\b/n4305 ), .IN1(\b/n4303 ), .SEL(msg[66]), .F(
        \b/n4306 ) );
  MUX \b/U4357  ( .IN0(\b/n4304 ), .IN1(\b/n4020 ), .SEL(msg[71]), .F(
        \b/n4305 ) );
  MUX \b/U4356  ( .IN0(\b/n562 ), .IN1(\b/n4007 ), .SEL(msg[65]), .F(\b/n4304 ) );
  MUX \b/U4355  ( .IN0(\b/n4302 ), .IN1(\b/n550 ), .SEL(msg[71]), .F(\b/n4303 ) );
  MUX \b/U4354  ( .IN0(\b/n4007 ), .IN1(\b/n4008 ), .SEL(msg[65]), .F(
        \b/n4302 ) );
  MUX \b/U4353  ( .IN0(\b/n4300 ), .IN1(\b/n4299 ), .SEL(msg[66]), .F(
        \b/n4301 ) );
  MUX \b/U4352  ( .IN0(n670), .IN1(\b/n4088 ), .SEL(msg[71]), .F(\b/n4300 ) );
  MUX \b/U4351  ( .IN0(\b/n4046 ), .IN1(\b/n4053 ), .SEL(msg[71]), .F(
        \b/n4299 ) );
  MUX \b/U4350  ( .IN0(\b/n4297 ), .IN1(\b/n4293 ), .SEL(msg[69]), .F(
        \b/n4298 ) );
  MUX \b/U4349  ( .IN0(\b/n4295 ), .IN1(\b/n4294 ), .SEL(msg[66]), .F(
        \b/n4297 ) );
  AND \b/U4348  ( .A(\b/n503 ), .B(\b/n4296 ), .Z(\b/n4295 ) );
  MUX \b/U4347  ( .IN0(\b/n4123 ), .IN1(msg[67]), .SEL(msg[71]), .F(\b/n4294 )
         );
  MUX \b/U4346  ( .IN0(\b/n4292 ), .IN1(\b/n4291 ), .SEL(msg[66]), .F(
        \b/n4293 ) );
  MUX \b/U4345  ( .IN0(\b/n546 ), .IN1(\b/n4011 ), .SEL(msg[71]), .F(\b/n4292 ) );
  MUX \b/U4343  ( .IN0(\b/n4289 ), .IN1(\b/n4282 ), .SEL(msg[64]), .F(
        \b/n4290 ) );
  MUX \b/U4342  ( .IN0(\b/n4288 ), .IN1(\b/n4285 ), .SEL(msg[69]), .F(
        \b/n4289 ) );
  MUX \b/U4341  ( .IN0(\b/n4287 ), .IN1(\b/n4286 ), .SEL(msg[66]), .F(
        \b/n4288 ) );
  MUX \b/U4340  ( .IN0(\b/n542 ), .IN1(\b/n4015 ), .SEL(msg[71]), .F(\b/n4287 ) );
  MUX \b/U4339  ( .IN0(\b/n4019 ), .IN1(n671), .SEL(msg[71]), .F(\b/n4286 ) );
  MUX \b/U4338  ( .IN0(\b/n4284 ), .IN1(\b/n4283 ), .SEL(msg[66]), .F(
        \b/n4285 ) );
  MUX \b/U4337  ( .IN0(\b/n4035 ), .IN1(\b/n507 ), .SEL(msg[71]), .F(\b/n4284 ) );
  MUX \b/U4336  ( .IN0(\b/n527 ), .IN1(\b/n557 ), .SEL(msg[71]), .F(\b/n4283 )
         );
  MUX \b/U4335  ( .IN0(\b/n4281 ), .IN1(\b/n4277 ), .SEL(msg[69]), .F(
        \b/n4282 ) );
  MUX \b/U4334  ( .IN0(\b/n4280 ), .IN1(\b/n4279 ), .SEL(msg[66]), .F(
        \b/n4281 ) );
  MUX \b/U4333  ( .IN0(\b/n4024 ), .IN1(\b/n557 ), .SEL(msg[71]), .F(\b/n4280 ) );
  MUX \b/U4332  ( .IN0(\b/n4278 ), .IN1(\b/n4045 ), .SEL(msg[71]), .F(
        \b/n4279 ) );
  NANDN \b/U4331  ( .B(msg[68]), .A(msg[65]), .Z(\b/n4278 ) );
  MUX \b/U4330  ( .IN0(\b/n4276 ), .IN1(\b/n4274 ), .SEL(msg[66]), .F(
        \b/n4277 ) );
  MUX \b/U4329  ( .IN0(\b/n520 ), .IN1(\b/n4275 ), .SEL(msg[71]), .F(\b/n4276 ) );
  MUX \b/U4328  ( .IN0(\b/n547 ), .IN1(\b/n537 ), .SEL(msg[65]), .F(\b/n4275 )
         );
  MUX \b/U4327  ( .IN0(\b/n509 ), .IN1(\b/n4020 ), .SEL(msg[71]), .F(\b/n4274 ) );
  NANDN \b/U4326  ( .B(\b/n510 ), .A(msg[65]), .Z(\b/n4020 ) );
  MUX \b/U4325  ( .IN0(\b/n4273 ), .IN1(\b/n4252 ), .SEL(msg[70]), .F(
        shift_row_out[69]) );
  MUX \b/U4324  ( .IN0(\b/n4272 ), .IN1(\b/n4262 ), .SEL(msg[64]), .F(
        \b/n4273 ) );
  MUX \b/U4323  ( .IN0(\b/n4271 ), .IN1(\b/n4267 ), .SEL(msg[69]), .F(
        \b/n4272 ) );
  MUX \b/U4322  ( .IN0(\b/n4268 ), .IN1(\b/n4269 ), .SEL(msg[66]), .F(
        \b/n4271 ) );
  AND \b/U4321  ( .A(\b/n4038 ), .B(\b/n4270 ), .Z(\b/n4269 ) );
  MUX \b/U4320  ( .IN0(\b/n4016 ), .IN1(\b/n558 ), .SEL(msg[71]), .F(\b/n4268 ) );
  MUX \b/U4319  ( .IN0(\b/n4266 ), .IN1(\b/n4264 ), .SEL(msg[66]), .F(
        \b/n4267 ) );
  MUX \b/U4318  ( .IN0(\b/n513 ), .IN1(\b/n4265 ), .SEL(msg[71]), .F(\b/n4266 ) );
  NAND \b/U4317  ( .A(\b/n537 ), .B(\b/n567 ), .Z(\b/n4265 ) );
  MUX \b/U4316  ( .IN0(\b/n4016 ), .IN1(\b/n4263 ), .SEL(msg[71]), .F(
        \b/n4264 ) );
  NAND \b/U4315  ( .A(\b/n4007 ), .B(\b/n4068 ), .Z(\b/n4263 ) );
  MUX \b/U4314  ( .IN0(\b/n4261 ), .IN1(\b/n4257 ), .SEL(msg[69]), .F(
        \b/n4262 ) );
  MUX \b/U4313  ( .IN0(\b/n4260 ), .IN1(\b/n4259 ), .SEL(msg[66]), .F(
        \b/n4261 ) );
  MUX \b/U4312  ( .IN0(\b/n4028 ), .IN1(\b/n560 ), .SEL(msg[71]), .F(\b/n4260 ) );
  MUX \b/U4311  ( .IN0(\b/n4053 ), .IN1(\b/n4258 ), .SEL(msg[71]), .F(
        \b/n4259 ) );
  MUX \b/U4310  ( .IN0(\b/n556 ), .IN1(\b/n537 ), .SEL(msg[65]), .F(\b/n4258 )
         );
  MUX \b/U4309  ( .IN0(\b/n4256 ), .IN1(\b/n4255 ), .SEL(msg[66]), .F(
        \b/n4257 ) );
  MUX \b/U4308  ( .IN0(\b/n554 ), .IN1(n669), .SEL(msg[71]), .F(\b/n4256 ) );
  MUX \b/U4307  ( .IN0(\b/n4254 ), .IN1(\b/n4253 ), .SEL(msg[71]), .F(
        \b/n4255 ) );
  AND \b/U4306  ( .A(\b/n4013 ), .B(\b/n4088 ), .Z(\b/n4254 ) );
  MUX \b/U4305  ( .IN0(\b/n526 ), .IN1(\b/n510 ), .SEL(msg[65]), .F(\b/n4253 )
         );
  MUX \b/U4304  ( .IN0(\b/n4251 ), .IN1(\b/n4242 ), .SEL(msg[64]), .F(
        \b/n4252 ) );
  MUX \b/U4303  ( .IN0(\b/n4250 ), .IN1(\b/n4246 ), .SEL(msg[69]), .F(
        \b/n4251 ) );
  MUX \b/U4302  ( .IN0(\b/n4249 ), .IN1(\b/n4247 ), .SEL(msg[66]), .F(
        \b/n4250 ) );
  MUX \b/U4301  ( .IN0(\b/n4019 ), .IN1(\b/n4248 ), .SEL(msg[71]), .F(
        \b/n4249 ) );
  NAND \b/U4300  ( .A(msg[65]), .B(\b/n526 ), .Z(\b/n4248 ) );
  MUX \b/U4299  ( .IN0(\b/n510 ), .IN1(\b/n563 ), .SEL(msg[71]), .F(\b/n4247 )
         );
  MUX \b/U4298  ( .IN0(\b/n4245 ), .IN1(\b/n4244 ), .SEL(msg[66]), .F(
        \b/n4246 ) );
  MUX \b/U4297  ( .IN0(\b/n4045 ), .IN1(\b/n528 ), .SEL(msg[71]), .F(\b/n4245 ) );
  MUX \b/U4296  ( .IN0(\b/n4243 ), .IN1(\b/n4008 ), .SEL(n668), .F(\b/n4244 )
         );
  AND \b/U4295  ( .A(msg[71]), .B(msg[67]), .Z(\b/n4243 ) );
  MUX \b/U4294  ( .IN0(\b/n4241 ), .IN1(\b/n4238 ), .SEL(msg[69]), .F(
        \b/n4242 ) );
  MUX \b/U4293  ( .IN0(\b/n4240 ), .IN1(\b/n4239 ), .SEL(msg[66]), .F(
        \b/n4241 ) );
  MUX \b/U4292  ( .IN0(\b/n4169 ), .IN1(\b/n4008 ), .SEL(msg[71]), .F(
        \b/n4240 ) );
  MUX \b/U4291  ( .IN0(n667), .IN1(\b/n561 ), .SEL(msg[71]), .F(\b/n4239 ) );
  MUX \b/U4290  ( .IN0(\b/n4236 ), .IN1(\b/n4235 ), .SEL(msg[66]), .F(
        \b/n4238 ) );
  AND \b/U4289  ( .A(\b/n4237 ), .B(\b/n4137 ), .Z(\b/n4236 ) );
  MUX \b/U4288  ( .IN0(\b/n512 ), .IN1(\b/n556 ), .SEL(msg[71]), .F(\b/n4235 )
         );
  MUX \b/U4287  ( .IN0(\b/n4234 ), .IN1(\b/n4217 ), .SEL(msg[70]), .F(
        shift_row_out[68]) );
  MUX \b/U4286  ( .IN0(\b/n4233 ), .IN1(\b/n4225 ), .SEL(msg[64]), .F(
        \b/n4234 ) );
  MUX \b/U4285  ( .IN0(\b/n4232 ), .IN1(\b/n4229 ), .SEL(msg[69]), .F(
        \b/n4233 ) );
  MUX \b/U4284  ( .IN0(\b/n4231 ), .IN1(\b/n4230 ), .SEL(msg[66]), .F(
        \b/n4232 ) );
  MUX \b/U4283  ( .IN0(\b/n538 ), .IN1(\b/n559 ), .SEL(msg[71]), .F(\b/n4231 )
         );
  MUX \b/U4282  ( .IN0(\b/n4088 ), .IN1(\b/n4053 ), .SEL(msg[71]), .F(
        \b/n4230 ) );
  NAND \b/U4281  ( .A(msg[65]), .B(\b/n4007 ), .Z(\b/n4088 ) );
  MUX \b/U4280  ( .IN0(\b/n4226 ), .IN1(\b/n4227 ), .SEL(msg[66]), .F(
        \b/n4229 ) );
  AND \b/U4279  ( .A(\b/n4038 ), .B(\b/n4228 ), .Z(\b/n4227 ) );
  MUX \b/U4278  ( .IN0(\b/n4036 ), .IN1(\b/n541 ), .SEL(msg[71]), .F(\b/n4226 ) );
  MUX \b/U4277  ( .IN0(\b/n4224 ), .IN1(\b/n4221 ), .SEL(msg[69]), .F(
        \b/n4225 ) );
  MUX \b/U4276  ( .IN0(\b/n4223 ), .IN1(\b/n4222 ), .SEL(msg[66]), .F(
        \b/n4224 ) );
  MUX \b/U4275  ( .IN0(\b/n503 ), .IN1(\b/n549 ), .SEL(msg[71]), .F(\b/n4223 )
         );
  MUX \b/U4274  ( .IN0(\b/n510 ), .IN1(\b/n4016 ), .SEL(msg[71]), .F(\b/n4222 ) );
  MUX \b/U4273  ( .IN0(\b/n4220 ), .IN1(\b/n4218 ), .SEL(msg[66]), .F(
        \b/n4221 ) );
  MUX \b/U4272  ( .IN0(\b/n4032 ), .IN1(\b/n4219 ), .SEL(msg[71]), .F(
        \b/n4220 ) );
  AND \b/U4271  ( .A(\b/n4016 ), .B(\b/n567 ), .Z(\b/n4219 ) );
  MUX \b/U4270  ( .IN0(\b/n525 ), .IN1(\b/n544 ), .SEL(msg[71]), .F(\b/n4218 )
         );
  MUX \b/U4269  ( .IN0(\b/n4216 ), .IN1(\b/n4210 ), .SEL(msg[64]), .F(
        \b/n4217 ) );
  MUX \b/U4268  ( .IN0(\b/n4215 ), .IN1(\b/n4213 ), .SEL(msg[69]), .F(
        \b/n4216 ) );
  MUX \b/U4267  ( .IN0(\b/n4214 ), .IN1(\b/n4010 ), .SEL(msg[66]), .F(
        \b/n4215 ) );
  MUX \b/U4266  ( .IN0(\b/n4030 ), .IN1(\b/n546 ), .SEL(msg[71]), .F(\b/n4214 ) );
  MUX \b/U4265  ( .IN0(\b/n4212 ), .IN1(\b/n4211 ), .SEL(msg[66]), .F(
        \b/n4213 ) );
  MUX \b/U4264  ( .IN0(n666), .IN1(\b/n538 ), .SEL(msg[71]), .F(\b/n4212 ) );
  MUX \b/U4263  ( .IN0(\b/n4040 ), .IN1(\b/n4043 ), .SEL(msg[71]), .F(
        \b/n4211 ) );
  MUX \b/U4262  ( .IN0(\b/n4209 ), .IN1(\b/n4206 ), .SEL(msg[69]), .F(
        \b/n4210 ) );
  MUX \b/U4261  ( .IN0(\b/n4208 ), .IN1(\b/n4207 ), .SEL(msg[66]), .F(
        \b/n4209 ) );
  MUX \b/U4260  ( .IN0(\b/n511 ), .IN1(\b/n4012 ), .SEL(msg[71]), .F(\b/n4208 ) );
  MUX \b/U4259  ( .IN0(\b/n556 ), .IN1(\b/n4034 ), .SEL(msg[71]), .F(\b/n4207 ) );
  MUX \b/U4258  ( .IN0(\b/n499 ), .IN1(\b/n4205 ), .SEL(msg[66]), .F(\b/n4206 ) );
  MUX \b/U4257  ( .IN0(\b/n519 ), .IN1(\b/n4016 ), .SEL(msg[71]), .F(\b/n4205 ) );
  MUX \b/U4256  ( .IN0(\b/n4204 ), .IN1(\b/n4185 ), .SEL(msg[70]), .F(
        shift_row_out[67]) );
  MUX \b/U4255  ( .IN0(\b/n4203 ), .IN1(\b/n4195 ), .SEL(msg[64]), .F(
        \b/n4204 ) );
  MUX \b/U4254  ( .IN0(\b/n4202 ), .IN1(\b/n4199 ), .SEL(msg[69]), .F(
        \b/n4203 ) );
  MUX \b/U4253  ( .IN0(\b/n4201 ), .IN1(\b/n4200 ), .SEL(msg[71]), .F(
        \b/n4202 ) );
  MUX \b/U4252  ( .IN0(\b/n4024 ), .IN1(\b/n544 ), .SEL(msg[66]), .F(\b/n4201 ) );
  MUX \b/U4251  ( .IN0(n669), .IN1(\b/n502 ), .SEL(msg[66]), .F(\b/n4200 ) );
  MUX \b/U4250  ( .IN0(\b/n4197 ), .IN1(\b/n4196 ), .SEL(msg[71]), .F(
        \b/n4199 ) );
  AND \b/U4249  ( .A(\b/n4198 ), .B(msg[68]), .Z(\b/n4197 ) );
  MUX \b/U4248  ( .IN0(\b/n532 ), .IN1(\b/n4037 ), .SEL(msg[66]), .F(\b/n4196 ) );
  MUX \b/U4247  ( .IN0(\b/n4194 ), .IN1(\b/n4191 ), .SEL(msg[69]), .F(
        \b/n4195 ) );
  MUX \b/U4246  ( .IN0(\b/n4193 ), .IN1(\b/n4192 ), .SEL(msg[71]), .F(
        \b/n4194 ) );
  MUX \b/U4245  ( .IN0(\b/n4028 ), .IN1(n665), .SEL(msg[66]), .F(\b/n4193 ) );
  MUX \b/U4244  ( .IN0(\b/n500 ), .IN1(\b/n519 ), .SEL(msg[66]), .F(\b/n4192 )
         );
  MUX \b/U4243  ( .IN0(\b/n4187 ), .IN1(\b/n4188 ), .SEL(msg[71]), .F(
        \b/n4191 ) );
  NAND \b/U4242  ( .A(\b/n4189 ), .B(\b/n4190 ), .Z(\b/n4188 ) );
  MUX \b/U4241  ( .IN0(\b/n545 ), .IN1(\b/n4186 ), .SEL(msg[66]), .F(\b/n4187 ) );
  MUX \b/U4240  ( .IN0(\b/n520 ), .IN1(\b/n562 ), .SEL(msg[65]), .F(\b/n4186 )
         );
  MUX \b/U4239  ( .IN0(\b/n4184 ), .IN1(\b/n4175 ), .SEL(msg[64]), .F(
        \b/n4185 ) );
  MUX \b/U4238  ( .IN0(\b/n4183 ), .IN1(\b/n4179 ), .SEL(msg[69]), .F(
        \b/n4184 ) );
  MUX \b/U4237  ( .IN0(\b/n4181 ), .IN1(\b/n4180 ), .SEL(msg[71]), .F(
        \b/n4183 ) );
  NAND \b/U4236  ( .A(\b/n510 ), .B(\b/n4182 ), .Z(\b/n4181 ) );
  MUX \b/U4235  ( .IN0(\b/n561 ), .IN1(\b/n523 ), .SEL(msg[66]), .F(\b/n4180 )
         );
  MUX \b/U4234  ( .IN0(\b/n4178 ), .IN1(\b/n4176 ), .SEL(msg[71]), .F(
        \b/n4179 ) );
  MUX \b/U4233  ( .IN0(\b/n4019 ), .IN1(\b/n4177 ), .SEL(msg[66]), .F(
        \b/n4178 ) );
  AND \b/U4232  ( .A(msg[65]), .B(\b/n510 ), .Z(\b/n4177 ) );
  MUX \b/U4231  ( .IN0(\b/n515 ), .IN1(\b/n4038 ), .SEL(msg[66]), .F(\b/n4176 ) );
  MUX \b/U4230  ( .IN0(\b/n4174 ), .IN1(\b/n4168 ), .SEL(msg[69]), .F(
        \b/n4175 ) );
  MUX \b/U4229  ( .IN0(\b/n4173 ), .IN1(\b/n4171 ), .SEL(msg[71]), .F(
        \b/n4174 ) );
  MUX \b/U4228  ( .IN0(\b/n4172 ), .IN1(\b/n4008 ), .SEL(\b/n4056 ), .F(
        \b/n4173 ) );
  MUX \b/U4227  ( .IN0(msg[67]), .IN1(msg[68]), .SEL(msg[66]), .F(\b/n4172 )
         );
  MUX \b/U4226  ( .IN0(\b/n4038 ), .IN1(\b/n4169 ), .SEL(msg[66]), .F(
        \b/n4171 ) );
  NAND \b/U4225  ( .A(\b/n4008 ), .B(\b/n4170 ), .Z(\b/n4169 ) );
  MUX \b/U4224  ( .IN0(\b/n4165 ), .IN1(\b/n4166 ), .SEL(msg[71]), .F(
        \b/n4168 ) );
  AND \b/U4223  ( .A(\b/n543 ), .B(\b/n4167 ), .Z(\b/n4166 ) );
  MUX \b/U4222  ( .IN0(\b/n524 ), .IN1(\b/n4009 ), .SEL(msg[66]), .F(\b/n4165 ) );
  MUX \b/U4221  ( .IN0(\b/n4164 ), .IN1(\b/n4148 ), .SEL(msg[70]), .F(
        shift_row_out[66]) );
  MUX \b/U4220  ( .IN0(\b/n4163 ), .IN1(\b/n4155 ), .SEL(msg[64]), .F(
        \b/n4164 ) );
  MUX \b/U4219  ( .IN0(\b/n4162 ), .IN1(\b/n4158 ), .SEL(msg[69]), .F(
        \b/n4163 ) );
  MUX \b/U4218  ( .IN0(\b/n4161 ), .IN1(\b/n4159 ), .SEL(msg[66]), .F(
        \b/n4162 ) );
  MUX \b/U4217  ( .IN0(\b/n532 ), .IN1(\b/n4160 ), .SEL(msg[71]), .F(\b/n4161 ) );
  MUX \b/U4216  ( .IN0(\b/n4016 ), .IN1(\b/n510 ), .SEL(msg[65]), .F(\b/n4160 ) );
  MUX \b/U4215  ( .IN0(\b/n4055 ), .IN1(\b/n550 ), .SEL(msg[71]), .F(\b/n4159 ) );
  MUX \b/U4214  ( .IN0(\b/n4157 ), .IN1(\b/n4156 ), .SEL(msg[66]), .F(
        \b/n4158 ) );
  MUX \b/U4213  ( .IN0(\b/n4009 ), .IN1(\b/n517 ), .SEL(msg[71]), .F(\b/n4157 ) );
  MUX \b/U4212  ( .IN0(\b/n553 ), .IN1(\b/n4042 ), .SEL(msg[71]), .F(\b/n4156 ) );
  MUX \b/U4211  ( .IN0(\b/n4154 ), .IN1(\b/n4150 ), .SEL(msg[69]), .F(
        \b/n4155 ) );
  MUX \b/U4210  ( .IN0(\b/n4151 ), .IN1(\b/n499 ), .SEL(msg[66]), .F(\b/n4154 ) );
  NAND \b/U4209  ( .A(\b/n4152 ), .B(\b/n4153 ), .Z(\b/n4151 ) );
  MUX \b/U4208  ( .IN0(n667), .IN1(\b/n4149 ), .SEL(\b/n4054 ), .F(\b/n4150 )
         );
  MUX \b/U4207  ( .IN0(\b/n531 ), .IN1(\b/n4021 ), .SEL(msg[66]), .F(\b/n4149 ) );
  MUX \b/U4206  ( .IN0(\b/n4147 ), .IN1(\b/n4139 ), .SEL(msg[64]), .F(
        \b/n4148 ) );
  MUX \b/U4205  ( .IN0(\b/n4146 ), .IN1(\b/n4143 ), .SEL(msg[69]), .F(
        \b/n4147 ) );
  MUX \b/U4204  ( .IN0(\b/n4145 ), .IN1(\b/n4144 ), .SEL(msg[66]), .F(
        \b/n4146 ) );
  MUX \b/U4203  ( .IN0(\b/n559 ), .IN1(msg[65]), .SEL(msg[71]), .F(\b/n4145 )
         );
  MUX \b/U4202  ( .IN0(n670), .IN1(\b/n4022 ), .SEL(msg[71]), .F(\b/n4144 ) );
  MUX \b/U4201  ( .IN0(\b/n4142 ), .IN1(\b/n4141 ), .SEL(msg[66]), .F(
        \b/n4143 ) );
  MUX \b/U4200  ( .IN0(\b/n564 ), .IN1(\b/n558 ), .SEL(msg[71]), .F(\b/n4142 )
         );
  MUX \b/U4199  ( .IN0(n670), .IN1(\b/n4140 ), .SEL(msg[71]), .F(\b/n4141 ) );
  MUX \b/U4198  ( .IN0(\b/n510 ), .IN1(\b/n547 ), .SEL(msg[65]), .F(\b/n4140 )
         );
  MUX \b/U4197  ( .IN0(\b/n4138 ), .IN1(\b/n4132 ), .SEL(msg[69]), .F(
        \b/n4139 ) );
  MUX \b/U4196  ( .IN0(\b/n4135 ), .IN1(\b/n4134 ), .SEL(msg[66]), .F(
        \b/n4138 ) );
  NAND \b/U4195  ( .A(\b/n4136 ), .B(\b/n4137 ), .Z(\b/n4135 ) );
  MUX \b/U4194  ( .IN0(\b/n4008 ), .IN1(\b/n4133 ), .SEL(n668), .F(\b/n4134 )
         );
  MUX \b/U4193  ( .IN0(msg[67]), .IN1(\b/n520 ), .SEL(msg[71]), .F(\b/n4133 )
         );
  MUX \b/U4192  ( .IN0(\b/n4131 ), .IN1(\b/n4130 ), .SEL(msg[66]), .F(
        \b/n4132 ) );
  MUX \b/U4191  ( .IN0(\b/n4053 ), .IN1(\b/n518 ), .SEL(msg[71]), .F(\b/n4131 ) );
  MUX \b/U4190  ( .IN0(\b/n4049 ), .IN1(\b/n4129 ), .SEL(msg[71]), .F(
        \b/n4130 ) );
  MUX \b/U4189  ( .IN0(\b/n4011 ), .IN1(\b/n4016 ), .SEL(msg[65]), .F(
        \b/n4129 ) );
  MUX \b/U4188  ( .IN0(\b/n4128 ), .IN1(\b/n4110 ), .SEL(msg[70]), .F(
        shift_row_out[65]) );
  MUX \b/U4187  ( .IN0(\b/n4127 ), .IN1(\b/n4118 ), .SEL(msg[64]), .F(
        \b/n4128 ) );
  MUX \b/U4186  ( .IN0(\b/n4126 ), .IN1(\b/n4122 ), .SEL(msg[69]), .F(
        \b/n4127 ) );
  MUX \b/U4185  ( .IN0(\b/n4125 ), .IN1(\b/n4124 ), .SEL(msg[66]), .F(
        \b/n4126 ) );
  MUX \b/U4184  ( .IN0(\b/n555 ), .IN1(n672), .SEL(msg[71]), .F(\b/n4125 ) );
  MUX \b/U4183  ( .IN0(\b/n4123 ), .IN1(n666), .SEL(msg[71]), .F(\b/n4124 ) );
  NAND \b/U4182  ( .A(\b/n567 ), .B(\b/n526 ), .Z(\b/n4123 ) );
  MUX \b/U4181  ( .IN0(\b/n4121 ), .IN1(\b/n4120 ), .SEL(msg[66]), .F(
        \b/n4122 ) );
  MUX \b/U4180  ( .IN0(\b/n503 ), .IN1(\b/n4023 ), .SEL(msg[71]), .F(\b/n4121 ) );
  MUX \b/U4179  ( .IN0(\b/n4013 ), .IN1(\b/n4119 ), .SEL(msg[71]), .F(
        \b/n4120 ) );
  AND \b/U4178  ( .A(msg[65]), .B(msg[68]), .Z(\b/n4119 ) );
  MUX \b/U4177  ( .IN0(\b/n4117 ), .IN1(\b/n4114 ), .SEL(msg[69]), .F(
        \b/n4118 ) );
  MUX \b/U4176  ( .IN0(\b/n4116 ), .IN1(\b/n4115 ), .SEL(msg[66]), .F(
        \b/n4117 ) );
  MUX \b/U4175  ( .IN0(\b/n4052 ), .IN1(\b/n564 ), .SEL(msg[71]), .F(\b/n4116 ) );
  MUX \b/U4174  ( .IN0(\b/n539 ), .IN1(\b/n4021 ), .SEL(msg[71]), .F(\b/n4115 ) );
  MUX \b/U4173  ( .IN0(\b/n4111 ), .IN1(\b/n4112 ), .SEL(msg[66]), .F(
        \b/n4114 ) );
  AND \b/U4172  ( .A(\b/n4113 ), .B(\b/n4068 ), .Z(\b/n4112 ) );
  MUX \b/U4171  ( .IN0(\b/n4027 ), .IN1(\b/n4016 ), .SEL(msg[71]), .F(
        \b/n4111 ) );
  MUX \b/U4170  ( .IN0(\b/n4109 ), .IN1(\b/n4101 ), .SEL(msg[64]), .F(
        \b/n4110 ) );
  MUX \b/U4169  ( .IN0(\b/n4108 ), .IN1(\b/n4104 ), .SEL(msg[69]), .F(
        \b/n4109 ) );
  MUX \b/U4168  ( .IN0(\b/n4107 ), .IN1(\b/n4106 ), .SEL(msg[66]), .F(
        \b/n4108 ) );
  MUX \b/U4167  ( .IN0(\b/n4015 ), .IN1(\b/n528 ), .SEL(msg[71]), .F(\b/n4107 ) );
  MUX \b/U4166  ( .IN0(\b/n4105 ), .IN1(\b/n512 ), .SEL(msg[71]), .F(\b/n4106 ) );
  MUX \b/U4165  ( .IN0(\b/n4013 ), .IN1(\b/n520 ), .SEL(msg[65]), .F(\b/n4105 ) );
  MUX \b/U4164  ( .IN0(\b/n4103 ), .IN1(\b/n4102 ), .SEL(msg[66]), .F(
        \b/n4104 ) );
  MUX \b/U4163  ( .IN0(\b/n559 ), .IN1(\b/n537 ), .SEL(msg[71]), .F(\b/n4103 )
         );
  MUX \b/U4162  ( .IN0(\b/n555 ), .IN1(\b/n515 ), .SEL(msg[71]), .F(\b/n4102 )
         );
  MUX \b/U4161  ( .IN0(\b/n4100 ), .IN1(\b/n4095 ), .SEL(msg[69]), .F(
        \b/n4101 ) );
  MUX \b/U4160  ( .IN0(\b/n4099 ), .IN1(\b/n4096 ), .SEL(msg[66]), .F(
        \b/n4100 ) );
  MUX \b/U4159  ( .IN0(\b/n4097 ), .IN1(\b/n4098 ), .SEL(msg[71]), .F(
        \b/n4099 ) );
  NAND \b/U4158  ( .A(\b/n4016 ), .B(\b/n4088 ), .Z(\b/n4098 ) );
  MUX \b/U4157  ( .IN0(\b/n4016 ), .IN1(\b/n520 ), .SEL(msg[65]), .F(\b/n4097 ) );
  MUX \b/U4156  ( .IN0(\b/n4033 ), .IN1(\b/n4031 ), .SEL(msg[71]), .F(
        \b/n4096 ) );
  MUX \b/U4155  ( .IN0(\b/n4051 ), .IN1(\b/n4094 ), .SEL(msg[66]), .F(
        \b/n4095 ) );
  MUX \b/U4154  ( .IN0(\b/n526 ), .IN1(\b/n558 ), .SEL(msg[71]), .F(\b/n4094 )
         );
  MUX \b/U4153  ( .IN0(\b/n4093 ), .IN1(\b/n4076 ), .SEL(msg[70]), .F(
        shift_row_out[64]) );
  MUX \b/U4152  ( .IN0(\b/n4092 ), .IN1(\b/n4084 ), .SEL(msg[64]), .F(
        \b/n4093 ) );
  MUX \b/U4151  ( .IN0(\b/n4091 ), .IN1(\b/n4089 ), .SEL(msg[66]), .F(
        \b/n4092 ) );
  MUX \b/U4150  ( .IN0(\b/n500 ), .IN1(\b/n4090 ), .SEL(msg[71]), .F(\b/n4091 ) );
  MUX \b/U4149  ( .IN0(\b/n553 ), .IN1(\b/n556 ), .SEL(msg[69]), .F(\b/n4090 )
         );
  MUX \b/U4148  ( .IN0(\b/n4086 ), .IN1(\b/n4085 ), .SEL(msg[71]), .F(
        \b/n4089 ) );
  NAND \b/U4147  ( .A(\b/n4087 ), .B(\b/n4088 ), .Z(\b/n4086 ) );
  MUX \b/U4146  ( .IN0(\b/n552 ), .IN1(\b/n567 ), .SEL(msg[69]), .F(\b/n4085 )
         );
  MUX \b/U4145  ( .IN0(\b/n4083 ), .IN1(\b/n4079 ), .SEL(msg[66]), .F(
        \b/n4084 ) );
  MUX \b/U4144  ( .IN0(\b/n4082 ), .IN1(\b/n4080 ), .SEL(msg[71]), .F(
        \b/n4083 ) );
  MUX \b/U4143  ( .IN0(\b/n4081 ), .IN1(\b/n505 ), .SEL(msg[69]), .F(\b/n4082 ) );
  NAND \b/U4142  ( .A(\b/n567 ), .B(\b/n4008 ), .Z(\b/n4081 ) );
  MUX \b/U4140  ( .IN0(\b/n4078 ), .IN1(\b/n4077 ), .SEL(msg[71]), .F(
        \b/n4079 ) );
  MUX \b/U4139  ( .IN0(n667), .IN1(\b/n502 ), .SEL(msg[69]), .F(\b/n4078 ) );
  MUX \b/U4138  ( .IN0(\b/n554 ), .IN1(\b/n510 ), .SEL(msg[69]), .F(\b/n4077 )
         );
  MUX \b/U4137  ( .IN0(\b/n4075 ), .IN1(\b/n4065 ), .SEL(msg[64]), .F(
        \b/n4076 ) );
  MUX \b/U4136  ( .IN0(\b/n4074 ), .IN1(\b/n4070 ), .SEL(msg[66]), .F(
        \b/n4075 ) );
  MUX \b/U4135  ( .IN0(\b/n4073 ), .IN1(\b/n4072 ), .SEL(msg[71]), .F(
        \b/n4074 ) );
  MUX \b/U4134  ( .IN0(n665), .IN1(\b/n506 ), .SEL(msg[69]), .F(\b/n4073 ) );
  MUX \b/U4133  ( .IN0(\b/n4071 ), .IN1(\b/n543 ), .SEL(msg[69]), .F(\b/n4072 ) );
  NAND \b/U4132  ( .A(\b/n4007 ), .B(\b/n4009 ), .Z(\b/n4071 ) );
  MUX \b/U4131  ( .IN0(\b/n4069 ), .IN1(\b/n4066 ), .SEL(msg[71]), .F(
        \b/n4070 ) );
  MUX \b/U4130  ( .IN0(\b/n513 ), .IN1(\b/n4067 ), .SEL(msg[69]), .F(\b/n4069 ) );
  NAND \b/U4129  ( .A(\b/n4011 ), .B(\b/n4068 ), .Z(\b/n4067 ) );
  MUX \b/U4128  ( .IN0(\b/n4026 ), .IN1(\b/n4017 ), .SEL(msg[69]), .F(
        \b/n4066 ) );
  MUX \b/U4127  ( .IN0(\b/n4064 ), .IN1(\b/n4060 ), .SEL(msg[66]), .F(
        \b/n4065 ) );
  MUX \b/U4126  ( .IN0(\b/n4062 ), .IN1(\b/n4061 ), .SEL(msg[71]), .F(
        \b/n4064 ) );
  NAND \b/U4125  ( .A(\b/n4063 ), .B(\b/n4050 ), .Z(\b/n4062 ) );
  MUX \b/U4124  ( .IN0(msg[67]), .IN1(\b/n4042 ), .SEL(msg[69]), .F(\b/n4061 )
         );
  MUX \b/U4123  ( .IN0(\b/n4059 ), .IN1(\b/n4058 ), .SEL(msg[71]), .F(
        \b/n4060 ) );
  MUX \b/U4122  ( .IN0(\b/n518 ), .IN1(\b/n534 ), .SEL(msg[69]), .F(\b/n4059 )
         );
  MUX \b/U4121  ( .IN0(\b/n551 ), .IN1(\b/n539 ), .SEL(msg[69]), .F(\b/n4058 )
         );
  XOR \b/U4120  ( .A(\b/n4008 ), .B(msg[65]), .Z(\b/n4057 ) );
  XOR \b/U4119  ( .A(msg[65]), .B(msg[66]), .Z(\b/n4056 ) );
  XOR \b/U4118  ( .A(msg[65]), .B(msg[67]), .Z(\b/n4055 ) );
  XOR \b/U4117  ( .A(msg[66]), .B(msg[71]), .Z(\b/n4054 ) );
  XOR \b/U4116  ( .A(\b/n567 ), .B(\b/n510 ), .Z(\b/n4053 ) );
  XOR \b/U4115  ( .A(msg[65]), .B(\b/n556 ), .Z(\b/n4052 ) );
  XOR \b/U4113  ( .A(msg[65]), .B(msg[69]), .Z(\b/n4050 ) );
  NAND \b/U4112  ( .A(msg[65]), .B(msg[67]), .Z(\b/n4049 ) );
  MUX \b/U4111  ( .IN0(\b/n4008 ), .IN1(\b/n510 ), .SEL(msg[65]), .F(\b/n4048 ) );
  MUX \b/U4109  ( .IN0(msg[67]), .IN1(\b/n547 ), .SEL(msg[65]), .F(\b/n4046 )
         );
  MUX \b/U4108  ( .IN0(\b/n526 ), .IN1(\b/n547 ), .SEL(msg[65]), .F(\b/n4045 )
         );
  MUX \b/U4107  ( .IN0(\b/n4011 ), .IN1(\b/n4013 ), .SEL(msg[65]), .F(
        \b/n4044 ) );
  MUX \b/U4106  ( .IN0(msg[68]), .IN1(\b/n526 ), .SEL(msg[65]), .F(\b/n4043 )
         );
  OR \b/U4105  ( .A(msg[65]), .B(msg[68]), .Z(\b/n4042 ) );
  NAND \b/U4103  ( .A(\b/n547 ), .B(\b/n567 ), .Z(\b/n4040 ) );
  MUX \b/U4102  ( .IN0(\b/n547 ), .IN1(msg[68]), .SEL(msg[65]), .F(\b/n4039 )
         );
  MUX \b/U4101  ( .IN0(\b/n4007 ), .IN1(\b/n4016 ), .SEL(msg[65]), .F(
        \b/n4038 ) );
  MUX \b/U4100  ( .IN0(\b/n562 ), .IN1(msg[68]), .SEL(msg[65]), .F(\b/n4037 )
         );
  MUX \b/U4099  ( .IN0(\b/n520 ), .IN1(\b/n547 ), .SEL(msg[65]), .F(\b/n4036 )
         );
  MUX \b/U4098  ( .IN0(\b/n4007 ), .IN1(msg[68]), .SEL(msg[65]), .F(\b/n4035 )
         );
  MUX \b/U4097  ( .IN0(\b/n537 ), .IN1(\b/n526 ), .SEL(msg[65]), .F(\b/n4034 )
         );
  XOR \b/U4096  ( .A(\b/n520 ), .B(msg[65]), .Z(\b/n4033 ) );
  MUX \b/U4095  ( .IN0(\b/n4013 ), .IN1(\b/n537 ), .SEL(msg[65]), .F(\b/n4032 ) );
  NANDN \b/U4094  ( .B(msg[65]), .A(msg[67]), .Z(\b/n4031 ) );
  MUX \b/U4093  ( .IN0(\b/n510 ), .IN1(msg[67]), .SEL(msg[65]), .F(\b/n4030 )
         );
  NAND \b/U4091  ( .A(\b/n4011 ), .B(\b/n567 ), .Z(\b/n4028 ) );
  MUX \b/U4090  ( .IN0(msg[68]), .IN1(\b/n4008 ), .SEL(msg[65]), .F(\b/n4027 )
         );
  MUX \b/U4089  ( .IN0(\b/n537 ), .IN1(msg[67]), .SEL(msg[65]), .F(\b/n4026 )
         );
  MUX \b/U4087  ( .IN0(msg[68]), .IN1(\b/n556 ), .SEL(msg[65]), .F(\b/n4024 )
         );
  MUX \b/U4086  ( .IN0(\b/n510 ), .IN1(\b/n562 ), .SEL(msg[65]), .F(\b/n4023 )
         );
  NAND \b/U4085  ( .A(\b/n4009 ), .B(\b/n510 ), .Z(\b/n4022 ) );
  MUX \b/U4084  ( .IN0(\b/n4008 ), .IN1(\b/n4016 ), .SEL(msg[65]), .F(
        \b/n4021 ) );
  NAND \b/U4083  ( .A(\b/n4020 ), .B(\b/n4007 ), .Z(\b/n4019 ) );
  MUX \b/U4082  ( .IN0(\b/n4011 ), .IN1(\b/n562 ), .SEL(msg[65]), .F(\b/n4018 ) );
  MUX \b/U4081  ( .IN0(\b/n562 ), .IN1(\b/n526 ), .SEL(msg[65]), .F(\b/n4017 )
         );
  NANDN \b/U4080  ( .B(msg[67]), .A(msg[68]), .Z(\b/n4016 ) );
  MUX \b/U4079  ( .IN0(\b/n4011 ), .IN1(msg[67]), .SEL(msg[65]), .F(\b/n4015 )
         );
  OR \b/U4078  ( .A(msg[67]), .B(msg[68]), .Z(\b/n4011 ) );
  MUX \b/U4077  ( .IN0(\b/n510 ), .IN1(\b/n526 ), .SEL(msg[65]), .F(\b/n4014 )
         );
  XOR \b/U4076  ( .A(\b/n520 ), .B(msg[67]), .Z(\b/n4013 ) );
  NANDN \b/U4075  ( .B(msg[67]), .A(msg[65]), .Z(\b/n4012 ) );
  NAND \b/U4074  ( .A(\b/n4011 ), .B(\b/n4009 ), .Z(\b/n4010 ) );
  NAND \b/U4073  ( .A(msg[65]), .B(\b/n4008 ), .Z(\b/n4009 ) );
  NANDN \b/U4072  ( .B(msg[68]), .A(msg[67]), .Z(\b/n4008 ) );
  NAND \b/U4071  ( .A(msg[67]), .B(msg[68]), .Z(\b/n4007 ) );
  MUX \b/U4070  ( .IN0(msg[60]), .IN1(\b/n3648 ), .SEL(msg[57]), .F(\b/n4006 )
         );
  MUX \b/U4069  ( .IN0(msg[60]), .IN1(\b/n3657 ), .SEL(msg[57]), .F(\b/n4005 )
         );
  MUX \b/U4068  ( .IN0(\b/n3649 ), .IN1(\b/n3652 ), .SEL(msg[57]), .F(
        \b/n4004 ) );
  MUX \b/U4067  ( .IN0(\b/n3654 ), .IN1(\b/n627 ), .SEL(msg[57]), .F(\b/n4003 ) );
  MUX \b/U4065  ( .IN0(\b/n3657 ), .IN1(\b/n3648 ), .SEL(msg[58]), .F(
        \b/n3830 ) );
  MUX \b/U4064  ( .IN0(\b/n3650 ), .IN1(\b/n638 ), .SEL(msg[58]), .F(\b/n3831 ) );
  MUX \b/U4063  ( .IN0(\b/n581 ), .IN1(\b/n591 ), .SEL(msg[57]), .F(\b/n3794 )
         );
  MUX \b/U4062  ( .IN0(\b/n3678 ), .IN1(\b/n3989 ), .SEL(msg[63]), .F(
        \b/n4001 ) );
  MUX \b/U4061  ( .IN0(\b/n3652 ), .IN1(\b/n3648 ), .SEL(msg[57]), .F(
        \b/n3992 ) );
  MUX \b/U4060  ( .IN0(\b/n633 ), .IN1(\b/n3654 ), .SEL(msg[57]), .F(\b/n4000 ) );
  MUX \b/U4059  ( .IN0(msg[59]), .IN1(\b/n627 ), .SEL(msg[57]), .F(\b/n3999 )
         );
  MUX \b/U4058  ( .IN0(\b/n3657 ), .IN1(\b/n633 ), .SEL(msg[57]), .F(\b/n3998 ) );
  MUX \b/U4057  ( .IN0(msg[60]), .IN1(\b/n3654 ), .SEL(msg[57]), .F(\b/n3997 )
         );
  MUX \b/U4056  ( .IN0(\b/n618 ), .IN1(\b/n597 ), .SEL(msg[61]), .F(\b/n3704 )
         );
  MUX \b/U4055  ( .IN0(\b/n3649 ), .IN1(\b/n591 ), .SEL(msg[57]), .F(\b/n3996 ) );
  NANDN \b/U4052  ( .B(\b/n3655 ), .A(msg[63]), .Z(\b/n3969 ) );
  NAND \b/U4051  ( .A(msg[63]), .B(\b/n594 ), .Z(\b/n3937 ) );
  NAND \b/U4050  ( .A(msg[63]), .B(\b/n606 ), .Z(\b/n3878 ) );
  NAND \b/U4049  ( .A(msg[63]), .B(\b/n3986 ), .Z(\b/n3911 ) );
  NAND \b/U4048  ( .A(msg[63]), .B(\b/n3906 ), .Z(\b/n3869 ) );
  NAND \b/U4046  ( .A(\b/n638 ), .B(\b/n627 ), .Z(\b/n3990 ) );
  NAND \b/U4045  ( .A(msg[63]), .B(\b/n3988 ), .Z(\b/n3983 ) );
  NAND \b/U4044  ( .A(n664), .B(msg[63]), .Z(\b/n3963 ) );
  NAND \b/U4042  ( .A(msg[58]), .B(\b/n3657 ), .Z(\b/n3823 ) );
  NAND \b/U4041  ( .A(\b/n627 ), .B(msg[57]), .Z(\b/n3778 ) );
  NAND \b/U4040  ( .A(msg[63]), .B(\b/n3992 ), .Z(\b/n3777 ) );
  NAND \b/U4038  ( .A(\b/n3990 ), .B(msg[63]), .Z(\b/n3793 ) );
  NAND \b/U4037  ( .A(\b/n3811 ), .B(\b/n3657 ), .Z(\b/n3989 ) );
  NANDN \b/U4036  ( .B(\b/n581 ), .A(\b/n638 ), .Z(\b/n3988 ) );
  NAND \b/U4034  ( .A(msg[57]), .B(\b/n3657 ), .Z(\b/n3709 ) );
  NAND \b/U4033  ( .A(\b/n581 ), .B(\b/n638 ), .Z(\b/n3986 ) );
  NAND \b/U4030  ( .A(msg[57]), .B(\b/n3652 ), .Z(\b/n3811 ) );
  ANDN \b/U4028  ( .A(msg[58]), .B(msg[57]), .Z(\b/n3839 ) );
  AND \b/U4027  ( .A(\b/n3649 ), .B(\b/n3983 ), .Z(\b/n3754 ) );
  MUX \b/U4026  ( .IN0(\b/n3982 ), .IN1(\b/n3966 ), .SEL(msg[62]), .F(
        shift_row_out[95]) );
  MUX \b/U4025  ( .IN0(\b/n3981 ), .IN1(\b/n3974 ), .SEL(msg[56]), .F(
        \b/n3982 ) );
  MUX \b/U4024  ( .IN0(\b/n3980 ), .IN1(\b/n3977 ), .SEL(msg[61]), .F(
        \b/n3981 ) );
  MUX \b/U4023  ( .IN0(\b/n3979 ), .IN1(\b/n3978 ), .SEL(msg[58]), .F(
        \b/n3980 ) );
  MUX \b/U4022  ( .IN0(msg[60]), .IN1(\b/n598 ), .SEL(msg[63]), .F(\b/n3979 )
         );
  MUX \b/U4021  ( .IN0(\b/n3650 ), .IN1(\b/n602 ), .SEL(msg[63]), .F(\b/n3978 ) );
  MUX \b/U4020  ( .IN0(\b/n3976 ), .IN1(\b/n3975 ), .SEL(msg[58]), .F(
        \b/n3977 ) );
  MUX \b/U4019  ( .IN0(\b/n3708 ), .IN1(\b/n594 ), .SEL(msg[63]), .F(\b/n3976 ) );
  MUX \b/U4018  ( .IN0(\b/n3660 ), .IN1(\b/n3671 ), .SEL(msg[63]), .F(
        \b/n3975 ) );
  MUX \b/U4017  ( .IN0(\b/n3973 ), .IN1(\b/n3970 ), .SEL(msg[61]), .F(
        \b/n3974 ) );
  MUX \b/U4016  ( .IN0(\b/n3972 ), .IN1(\b/n3971 ), .SEL(msg[58]), .F(
        \b/n3973 ) );
  MUX \b/U4015  ( .IN0(\b/n3684 ), .IN1(\b/n3659 ), .SEL(msg[63]), .F(
        \b/n3972 ) );
  MUX \b/U4014  ( .IN0(\b/n606 ), .IN1(\b/n3680 ), .SEL(msg[63]), .F(\b/n3971 ) );
  MUX \b/U4013  ( .IN0(\b/n3968 ), .IN1(\b/n3967 ), .SEL(msg[58]), .F(
        \b/n3970 ) );
  AND \b/U4012  ( .A(\b/n596 ), .B(\b/n3969 ), .Z(\b/n3968 ) );
  MUX \b/U4011  ( .IN0(\b/n3664 ), .IN1(n663), .SEL(msg[63]), .F(\b/n3967 ) );
  MUX \b/U4010  ( .IN0(\b/n3965 ), .IN1(\b/n3957 ), .SEL(msg[56]), .F(
        \b/n3966 ) );
  MUX \b/U4009  ( .IN0(\b/n3964 ), .IN1(\b/n3960 ), .SEL(msg[61]), .F(
        \b/n3965 ) );
  MUX \b/U4008  ( .IN0(\b/n3961 ), .IN1(\b/n3962 ), .SEL(msg[58]), .F(
        \b/n3964 ) );
  NAND \b/U4007  ( .A(\b/n3778 ), .B(\b/n3963 ), .Z(\b/n3962 ) );
  MUX \b/U4006  ( .IN0(\b/n636 ), .IN1(\b/n628 ), .SEL(msg[63]), .F(\b/n3961 )
         );
  MUX \b/U4005  ( .IN0(\b/n3959 ), .IN1(\b/n3958 ), .SEL(msg[58]), .F(
        \b/n3960 ) );
  MUX \b/U4004  ( .IN0(\b/n3654 ), .IN1(\b/n3648 ), .SEL(msg[63]), .F(
        \b/n3959 ) );
  MUX \b/U4003  ( .IN0(\b/n629 ), .IN1(\b/n3685 ), .SEL(msg[63]), .F(\b/n3958 ) );
  MUX \b/U4002  ( .IN0(\b/n3956 ), .IN1(\b/n3953 ), .SEL(msg[61]), .F(
        \b/n3957 ) );
  MUX \b/U4001  ( .IN0(\b/n3955 ), .IN1(\b/n3954 ), .SEL(msg[58]), .F(
        \b/n3956 ) );
  MUX \b/U4000  ( .IN0(\b/n3689 ), .IN1(\b/n3675 ), .SEL(msg[63]), .F(
        \b/n3955 ) );
  MUX \b/U3999  ( .IN0(\b/n582 ), .IN1(\b/n3657 ), .SEL(msg[63]), .F(\b/n3954 ) );
  MUX \b/U3998  ( .IN0(\b/n3952 ), .IN1(\b/n3951 ), .SEL(msg[58]), .F(
        \b/n3953 ) );
  MUX \b/U3997  ( .IN0(\b/n3690 ), .IN1(\b/n3698 ), .SEL(msg[63]), .F(
        \b/n3952 ) );
  MUX \b/U3996  ( .IN0(\b/n3683 ), .IN1(\b/n3950 ), .SEL(msg[63]), .F(
        \b/n3951 ) );
  MUX \b/U3995  ( .IN0(\b/n633 ), .IN1(\b/n591 ), .SEL(msg[57]), .F(\b/n3950 )
         );
  MUX \b/U3994  ( .IN0(\b/n3949 ), .IN1(\b/n3931 ), .SEL(msg[62]), .F(
        shift_row_out[94]) );
  MUX \b/U3993  ( .IN0(\b/n3948 ), .IN1(\b/n3939 ), .SEL(msg[56]), .F(
        \b/n3949 ) );
  MUX \b/U3992  ( .IN0(\b/n3947 ), .IN1(\b/n3942 ), .SEL(msg[61]), .F(
        \b/n3948 ) );
  MUX \b/U3991  ( .IN0(\b/n3946 ), .IN1(\b/n3944 ), .SEL(msg[58]), .F(
        \b/n3947 ) );
  MUX \b/U3990  ( .IN0(\b/n3945 ), .IN1(\b/n3661 ), .SEL(msg[63]), .F(
        \b/n3946 ) );
  MUX \b/U3989  ( .IN0(\b/n633 ), .IN1(\b/n3648 ), .SEL(msg[57]), .F(\b/n3945 ) );
  MUX \b/U3988  ( .IN0(\b/n3943 ), .IN1(\b/n621 ), .SEL(msg[63]), .F(\b/n3944 ) );
  MUX \b/U3987  ( .IN0(\b/n3648 ), .IN1(\b/n3649 ), .SEL(msg[57]), .F(
        \b/n3943 ) );
  MUX \b/U3986  ( .IN0(\b/n3941 ), .IN1(\b/n3940 ), .SEL(msg[58]), .F(
        \b/n3942 ) );
  MUX \b/U3985  ( .IN0(n662), .IN1(\b/n3729 ), .SEL(msg[63]), .F(\b/n3941 ) );
  MUX \b/U3984  ( .IN0(\b/n3687 ), .IN1(\b/n3694 ), .SEL(msg[63]), .F(
        \b/n3940 ) );
  MUX \b/U3983  ( .IN0(\b/n3938 ), .IN1(\b/n3934 ), .SEL(msg[61]), .F(
        \b/n3939 ) );
  MUX \b/U3982  ( .IN0(\b/n3936 ), .IN1(\b/n3935 ), .SEL(msg[58]), .F(
        \b/n3938 ) );
  AND \b/U3981  ( .A(\b/n574 ), .B(\b/n3937 ), .Z(\b/n3936 ) );
  MUX \b/U3980  ( .IN0(\b/n3764 ), .IN1(msg[59]), .SEL(msg[63]), .F(\b/n3935 )
         );
  MUX \b/U3979  ( .IN0(\b/n3933 ), .IN1(\b/n3932 ), .SEL(msg[58]), .F(
        \b/n3934 ) );
  MUX \b/U3978  ( .IN0(\b/n617 ), .IN1(\b/n3652 ), .SEL(msg[63]), .F(\b/n3933 ) );
  MUX \b/U3976  ( .IN0(\b/n3930 ), .IN1(\b/n3923 ), .SEL(msg[56]), .F(
        \b/n3931 ) );
  MUX \b/U3975  ( .IN0(\b/n3929 ), .IN1(\b/n3926 ), .SEL(msg[61]), .F(
        \b/n3930 ) );
  MUX \b/U3974  ( .IN0(\b/n3928 ), .IN1(\b/n3927 ), .SEL(msg[58]), .F(
        \b/n3929 ) );
  MUX \b/U3973  ( .IN0(\b/n613 ), .IN1(\b/n3656 ), .SEL(msg[63]), .F(\b/n3928 ) );
  MUX \b/U3972  ( .IN0(\b/n3660 ), .IN1(n663), .SEL(msg[63]), .F(\b/n3927 ) );
  MUX \b/U3971  ( .IN0(\b/n3925 ), .IN1(\b/n3924 ), .SEL(msg[58]), .F(
        \b/n3926 ) );
  MUX \b/U3970  ( .IN0(\b/n3676 ), .IN1(\b/n578 ), .SEL(msg[63]), .F(\b/n3925 ) );
  MUX \b/U3969  ( .IN0(\b/n598 ), .IN1(\b/n628 ), .SEL(msg[63]), .F(\b/n3924 )
         );
  MUX \b/U3968  ( .IN0(\b/n3922 ), .IN1(\b/n3918 ), .SEL(msg[61]), .F(
        \b/n3923 ) );
  MUX \b/U3967  ( .IN0(\b/n3921 ), .IN1(\b/n3920 ), .SEL(msg[58]), .F(
        \b/n3922 ) );
  MUX \b/U3966  ( .IN0(\b/n3665 ), .IN1(\b/n628 ), .SEL(msg[63]), .F(\b/n3921 ) );
  MUX \b/U3965  ( .IN0(\b/n3919 ), .IN1(\b/n3686 ), .SEL(msg[63]), .F(
        \b/n3920 ) );
  NANDN \b/U3964  ( .B(msg[60]), .A(msg[57]), .Z(\b/n3919 ) );
  MUX \b/U3963  ( .IN0(\b/n3917 ), .IN1(\b/n3915 ), .SEL(msg[58]), .F(
        \b/n3918 ) );
  MUX \b/U3962  ( .IN0(\b/n591 ), .IN1(\b/n3916 ), .SEL(msg[63]), .F(\b/n3917 ) );
  MUX \b/U3961  ( .IN0(\b/n618 ), .IN1(\b/n608 ), .SEL(msg[57]), .F(\b/n3916 )
         );
  MUX \b/U3960  ( .IN0(\b/n580 ), .IN1(\b/n3661 ), .SEL(msg[63]), .F(\b/n3915 ) );
  NANDN \b/U3959  ( .B(\b/n581 ), .A(msg[57]), .Z(\b/n3661 ) );
  MUX \b/U3958  ( .IN0(\b/n3914 ), .IN1(\b/n3893 ), .SEL(msg[62]), .F(
        shift_row_out[93]) );
  MUX \b/U3957  ( .IN0(\b/n3913 ), .IN1(\b/n3903 ), .SEL(msg[56]), .F(
        \b/n3914 ) );
  MUX \b/U3956  ( .IN0(\b/n3912 ), .IN1(\b/n3908 ), .SEL(msg[61]), .F(
        \b/n3913 ) );
  MUX \b/U3955  ( .IN0(\b/n3909 ), .IN1(\b/n3910 ), .SEL(msg[58]), .F(
        \b/n3912 ) );
  AND \b/U3954  ( .A(\b/n3679 ), .B(\b/n3911 ), .Z(\b/n3910 ) );
  MUX \b/U3953  ( .IN0(\b/n3657 ), .IN1(\b/n629 ), .SEL(msg[63]), .F(\b/n3909 ) );
  MUX \b/U3952  ( .IN0(\b/n3907 ), .IN1(\b/n3905 ), .SEL(msg[58]), .F(
        \b/n3908 ) );
  MUX \b/U3951  ( .IN0(\b/n584 ), .IN1(\b/n3906 ), .SEL(msg[63]), .F(\b/n3907 ) );
  NAND \b/U3950  ( .A(\b/n608 ), .B(\b/n638 ), .Z(\b/n3906 ) );
  MUX \b/U3949  ( .IN0(\b/n3657 ), .IN1(\b/n3904 ), .SEL(msg[63]), .F(
        \b/n3905 ) );
  NAND \b/U3948  ( .A(\b/n3648 ), .B(\b/n3709 ), .Z(\b/n3904 ) );
  MUX \b/U3947  ( .IN0(\b/n3902 ), .IN1(\b/n3898 ), .SEL(msg[61]), .F(
        \b/n3903 ) );
  MUX \b/U3946  ( .IN0(\b/n3901 ), .IN1(\b/n3900 ), .SEL(msg[58]), .F(
        \b/n3902 ) );
  MUX \b/U3945  ( .IN0(\b/n3669 ), .IN1(\b/n631 ), .SEL(msg[63]), .F(\b/n3901 ) );
  MUX \b/U3944  ( .IN0(\b/n3694 ), .IN1(\b/n3899 ), .SEL(msg[63]), .F(
        \b/n3900 ) );
  MUX \b/U3943  ( .IN0(\b/n627 ), .IN1(\b/n608 ), .SEL(msg[57]), .F(\b/n3899 )
         );
  MUX \b/U3942  ( .IN0(\b/n3897 ), .IN1(\b/n3896 ), .SEL(msg[58]), .F(
        \b/n3898 ) );
  MUX \b/U3941  ( .IN0(\b/n625 ), .IN1(n661), .SEL(msg[63]), .F(\b/n3897 ) );
  MUX \b/U3940  ( .IN0(\b/n3895 ), .IN1(\b/n3894 ), .SEL(msg[63]), .F(
        \b/n3896 ) );
  AND \b/U3939  ( .A(\b/n3654 ), .B(\b/n3729 ), .Z(\b/n3895 ) );
  MUX \b/U3938  ( .IN0(\b/n597 ), .IN1(\b/n581 ), .SEL(msg[57]), .F(\b/n3894 )
         );
  MUX \b/U3937  ( .IN0(\b/n3892 ), .IN1(\b/n3883 ), .SEL(msg[56]), .F(
        \b/n3893 ) );
  MUX \b/U3936  ( .IN0(\b/n3891 ), .IN1(\b/n3887 ), .SEL(msg[61]), .F(
        \b/n3892 ) );
  MUX \b/U3935  ( .IN0(\b/n3890 ), .IN1(\b/n3888 ), .SEL(msg[58]), .F(
        \b/n3891 ) );
  MUX \b/U3934  ( .IN0(\b/n3660 ), .IN1(\b/n3889 ), .SEL(msg[63]), .F(
        \b/n3890 ) );
  NAND \b/U3933  ( .A(msg[57]), .B(\b/n597 ), .Z(\b/n3889 ) );
  MUX \b/U3932  ( .IN0(\b/n581 ), .IN1(\b/n634 ), .SEL(msg[63]), .F(\b/n3888 )
         );
  MUX \b/U3931  ( .IN0(\b/n3886 ), .IN1(\b/n3885 ), .SEL(msg[58]), .F(
        \b/n3887 ) );
  MUX \b/U3930  ( .IN0(\b/n3686 ), .IN1(\b/n599 ), .SEL(msg[63]), .F(\b/n3886 ) );
  MUX \b/U3929  ( .IN0(\b/n3884 ), .IN1(\b/n3649 ), .SEL(n660), .F(\b/n3885 )
         );
  AND \b/U3928  ( .A(msg[63]), .B(msg[59]), .Z(\b/n3884 ) );
  MUX \b/U3927  ( .IN0(\b/n3882 ), .IN1(\b/n3879 ), .SEL(msg[61]), .F(
        \b/n3883 ) );
  MUX \b/U3926  ( .IN0(\b/n3881 ), .IN1(\b/n3880 ), .SEL(msg[58]), .F(
        \b/n3882 ) );
  MUX \b/U3925  ( .IN0(\b/n3810 ), .IN1(\b/n3649 ), .SEL(msg[63]), .F(
        \b/n3881 ) );
  MUX \b/U3924  ( .IN0(n659), .IN1(\b/n632 ), .SEL(msg[63]), .F(\b/n3880 ) );
  MUX \b/U3923  ( .IN0(\b/n3877 ), .IN1(\b/n3876 ), .SEL(msg[58]), .F(
        \b/n3879 ) );
  AND \b/U3922  ( .A(\b/n3878 ), .B(\b/n3778 ), .Z(\b/n3877 ) );
  MUX \b/U3921  ( .IN0(\b/n583 ), .IN1(\b/n627 ), .SEL(msg[63]), .F(\b/n3876 )
         );
  MUX \b/U3920  ( .IN0(\b/n3875 ), .IN1(\b/n3858 ), .SEL(msg[62]), .F(
        shift_row_out[92]) );
  MUX \b/U3919  ( .IN0(\b/n3874 ), .IN1(\b/n3866 ), .SEL(msg[56]), .F(
        \b/n3875 ) );
  MUX \b/U3918  ( .IN0(\b/n3873 ), .IN1(\b/n3870 ), .SEL(msg[61]), .F(
        \b/n3874 ) );
  MUX \b/U3917  ( .IN0(\b/n3872 ), .IN1(\b/n3871 ), .SEL(msg[58]), .F(
        \b/n3873 ) );
  MUX \b/U3916  ( .IN0(\b/n609 ), .IN1(\b/n630 ), .SEL(msg[63]), .F(\b/n3872 )
         );
  MUX \b/U3915  ( .IN0(\b/n3729 ), .IN1(\b/n3694 ), .SEL(msg[63]), .F(
        \b/n3871 ) );
  NAND \b/U3914  ( .A(msg[57]), .B(\b/n3648 ), .Z(\b/n3729 ) );
  MUX \b/U3913  ( .IN0(\b/n3867 ), .IN1(\b/n3868 ), .SEL(msg[58]), .F(
        \b/n3870 ) );
  AND \b/U3912  ( .A(\b/n3679 ), .B(\b/n3869 ), .Z(\b/n3868 ) );
  MUX \b/U3911  ( .IN0(\b/n3677 ), .IN1(\b/n612 ), .SEL(msg[63]), .F(\b/n3867 ) );
  MUX \b/U3910  ( .IN0(\b/n3865 ), .IN1(\b/n3862 ), .SEL(msg[61]), .F(
        \b/n3866 ) );
  MUX \b/U3909  ( .IN0(\b/n3864 ), .IN1(\b/n3863 ), .SEL(msg[58]), .F(
        \b/n3865 ) );
  MUX \b/U3908  ( .IN0(\b/n574 ), .IN1(\b/n620 ), .SEL(msg[63]), .F(\b/n3864 )
         );
  MUX \b/U3907  ( .IN0(\b/n581 ), .IN1(\b/n3657 ), .SEL(msg[63]), .F(\b/n3863 ) );
  MUX \b/U3906  ( .IN0(\b/n3861 ), .IN1(\b/n3859 ), .SEL(msg[58]), .F(
        \b/n3862 ) );
  MUX \b/U3905  ( .IN0(\b/n3673 ), .IN1(\b/n3860 ), .SEL(msg[63]), .F(
        \b/n3861 ) );
  AND \b/U3904  ( .A(\b/n3657 ), .B(\b/n638 ), .Z(\b/n3860 ) );
  MUX \b/U3903  ( .IN0(\b/n596 ), .IN1(\b/n615 ), .SEL(msg[63]), .F(\b/n3859 )
         );
  MUX \b/U3902  ( .IN0(\b/n3857 ), .IN1(\b/n3851 ), .SEL(msg[56]), .F(
        \b/n3858 ) );
  MUX \b/U3901  ( .IN0(\b/n3856 ), .IN1(\b/n3854 ), .SEL(msg[61]), .F(
        \b/n3857 ) );
  MUX \b/U3900  ( .IN0(\b/n3855 ), .IN1(\b/n3651 ), .SEL(msg[58]), .F(
        \b/n3856 ) );
  MUX \b/U3899  ( .IN0(\b/n3671 ), .IN1(\b/n617 ), .SEL(msg[63]), .F(\b/n3855 ) );
  MUX \b/U3898  ( .IN0(\b/n3853 ), .IN1(\b/n3852 ), .SEL(msg[58]), .F(
        \b/n3854 ) );
  MUX \b/U3897  ( .IN0(n658), .IN1(\b/n609 ), .SEL(msg[63]), .F(\b/n3853 ) );
  MUX \b/U3896  ( .IN0(\b/n3681 ), .IN1(\b/n3684 ), .SEL(msg[63]), .F(
        \b/n3852 ) );
  MUX \b/U3895  ( .IN0(\b/n3850 ), .IN1(\b/n3847 ), .SEL(msg[61]), .F(
        \b/n3851 ) );
  MUX \b/U3894  ( .IN0(\b/n3849 ), .IN1(\b/n3848 ), .SEL(msg[58]), .F(
        \b/n3850 ) );
  MUX \b/U3893  ( .IN0(\b/n582 ), .IN1(\b/n3653 ), .SEL(msg[63]), .F(\b/n3849 ) );
  MUX \b/U3892  ( .IN0(\b/n627 ), .IN1(\b/n3675 ), .SEL(msg[63]), .F(\b/n3848 ) );
  MUX \b/U3891  ( .IN0(\b/n570 ), .IN1(\b/n3846 ), .SEL(msg[58]), .F(\b/n3847 ) );
  MUX \b/U3890  ( .IN0(\b/n590 ), .IN1(\b/n3657 ), .SEL(msg[63]), .F(\b/n3846 ) );
  MUX \b/U3889  ( .IN0(\b/n3845 ), .IN1(\b/n3826 ), .SEL(msg[62]), .F(
        shift_row_out[91]) );
  MUX \b/U3888  ( .IN0(\b/n3844 ), .IN1(\b/n3836 ), .SEL(msg[56]), .F(
        \b/n3845 ) );
  MUX \b/U3887  ( .IN0(\b/n3843 ), .IN1(\b/n3840 ), .SEL(msg[61]), .F(
        \b/n3844 ) );
  MUX \b/U3886  ( .IN0(\b/n3842 ), .IN1(\b/n3841 ), .SEL(msg[63]), .F(
        \b/n3843 ) );
  MUX \b/U3885  ( .IN0(\b/n3665 ), .IN1(\b/n615 ), .SEL(msg[58]), .F(\b/n3842 ) );
  MUX \b/U3884  ( .IN0(n661), .IN1(\b/n573 ), .SEL(msg[58]), .F(\b/n3841 ) );
  MUX \b/U3883  ( .IN0(\b/n3838 ), .IN1(\b/n3837 ), .SEL(msg[63]), .F(
        \b/n3840 ) );
  AND \b/U3882  ( .A(\b/n3839 ), .B(msg[60]), .Z(\b/n3838 ) );
  MUX \b/U3881  ( .IN0(\b/n603 ), .IN1(\b/n3678 ), .SEL(msg[58]), .F(\b/n3837 ) );
  MUX \b/U3880  ( .IN0(\b/n3835 ), .IN1(\b/n3832 ), .SEL(msg[61]), .F(
        \b/n3836 ) );
  MUX \b/U3879  ( .IN0(\b/n3834 ), .IN1(\b/n3833 ), .SEL(msg[63]), .F(
        \b/n3835 ) );
  MUX \b/U3878  ( .IN0(\b/n3669 ), .IN1(n657), .SEL(msg[58]), .F(\b/n3834 ) );
  MUX \b/U3877  ( .IN0(\b/n571 ), .IN1(\b/n590 ), .SEL(msg[58]), .F(\b/n3833 )
         );
  MUX \b/U3876  ( .IN0(\b/n3828 ), .IN1(\b/n3829 ), .SEL(msg[63]), .F(
        \b/n3832 ) );
  NAND \b/U3875  ( .A(\b/n3830 ), .B(\b/n3831 ), .Z(\b/n3829 ) );
  MUX \b/U3874  ( .IN0(\b/n616 ), .IN1(\b/n3827 ), .SEL(msg[58]), .F(\b/n3828 ) );
  MUX \b/U3873  ( .IN0(\b/n591 ), .IN1(\b/n633 ), .SEL(msg[57]), .F(\b/n3827 )
         );
  MUX \b/U3872  ( .IN0(\b/n3825 ), .IN1(\b/n3816 ), .SEL(msg[56]), .F(
        \b/n3826 ) );
  MUX \b/U3871  ( .IN0(\b/n3824 ), .IN1(\b/n3820 ), .SEL(msg[61]), .F(
        \b/n3825 ) );
  MUX \b/U3870  ( .IN0(\b/n3822 ), .IN1(\b/n3821 ), .SEL(msg[63]), .F(
        \b/n3824 ) );
  NAND \b/U3869  ( .A(\b/n581 ), .B(\b/n3823 ), .Z(\b/n3822 ) );
  MUX \b/U3868  ( .IN0(\b/n632 ), .IN1(\b/n594 ), .SEL(msg[58]), .F(\b/n3821 )
         );
  MUX \b/U3867  ( .IN0(\b/n3819 ), .IN1(\b/n3817 ), .SEL(msg[63]), .F(
        \b/n3820 ) );
  MUX \b/U3866  ( .IN0(\b/n3660 ), .IN1(\b/n3818 ), .SEL(msg[58]), .F(
        \b/n3819 ) );
  AND \b/U3865  ( .A(msg[57]), .B(\b/n581 ), .Z(\b/n3818 ) );
  MUX \b/U3864  ( .IN0(\b/n586 ), .IN1(\b/n3679 ), .SEL(msg[58]), .F(\b/n3817 ) );
  MUX \b/U3863  ( .IN0(\b/n3815 ), .IN1(\b/n3809 ), .SEL(msg[61]), .F(
        \b/n3816 ) );
  MUX \b/U3862  ( .IN0(\b/n3814 ), .IN1(\b/n3812 ), .SEL(msg[63]), .F(
        \b/n3815 ) );
  MUX \b/U3861  ( .IN0(\b/n3813 ), .IN1(\b/n3649 ), .SEL(\b/n3697 ), .F(
        \b/n3814 ) );
  MUX \b/U3860  ( .IN0(msg[59]), .IN1(msg[60]), .SEL(msg[58]), .F(\b/n3813 )
         );
  MUX \b/U3859  ( .IN0(\b/n3679 ), .IN1(\b/n3810 ), .SEL(msg[58]), .F(
        \b/n3812 ) );
  NAND \b/U3858  ( .A(\b/n3649 ), .B(\b/n3811 ), .Z(\b/n3810 ) );
  MUX \b/U3857  ( .IN0(\b/n3806 ), .IN1(\b/n3807 ), .SEL(msg[63]), .F(
        \b/n3809 ) );
  AND \b/U3856  ( .A(\b/n614 ), .B(\b/n3808 ), .Z(\b/n3807 ) );
  MUX \b/U3855  ( .IN0(\b/n595 ), .IN1(\b/n3650 ), .SEL(msg[58]), .F(\b/n3806 ) );
  MUX \b/U3854  ( .IN0(\b/n3805 ), .IN1(\b/n3789 ), .SEL(msg[62]), .F(
        shift_row_out[90]) );
  MUX \b/U3853  ( .IN0(\b/n3804 ), .IN1(\b/n3796 ), .SEL(msg[56]), .F(
        \b/n3805 ) );
  MUX \b/U3852  ( .IN0(\b/n3803 ), .IN1(\b/n3799 ), .SEL(msg[61]), .F(
        \b/n3804 ) );
  MUX \b/U3851  ( .IN0(\b/n3802 ), .IN1(\b/n3800 ), .SEL(msg[58]), .F(
        \b/n3803 ) );
  MUX \b/U3850  ( .IN0(\b/n603 ), .IN1(\b/n3801 ), .SEL(msg[63]), .F(\b/n3802 ) );
  MUX \b/U3849  ( .IN0(\b/n3657 ), .IN1(\b/n581 ), .SEL(msg[57]), .F(\b/n3801 ) );
  MUX \b/U3848  ( .IN0(\b/n3696 ), .IN1(\b/n621 ), .SEL(msg[63]), .F(\b/n3800 ) );
  MUX \b/U3847  ( .IN0(\b/n3798 ), .IN1(\b/n3797 ), .SEL(msg[58]), .F(
        \b/n3799 ) );
  MUX \b/U3846  ( .IN0(\b/n3650 ), .IN1(\b/n588 ), .SEL(msg[63]), .F(\b/n3798 ) );
  MUX \b/U3845  ( .IN0(\b/n624 ), .IN1(\b/n3683 ), .SEL(msg[63]), .F(\b/n3797 ) );
  MUX \b/U3844  ( .IN0(\b/n3795 ), .IN1(\b/n3791 ), .SEL(msg[61]), .F(
        \b/n3796 ) );
  MUX \b/U3843  ( .IN0(\b/n3792 ), .IN1(\b/n570 ), .SEL(msg[58]), .F(\b/n3795 ) );
  NAND \b/U3842  ( .A(\b/n3793 ), .B(\b/n3794 ), .Z(\b/n3792 ) );
  MUX \b/U3841  ( .IN0(n659), .IN1(\b/n3790 ), .SEL(\b/n3695 ), .F(\b/n3791 )
         );
  MUX \b/U3840  ( .IN0(\b/n602 ), .IN1(\b/n3662 ), .SEL(msg[58]), .F(\b/n3790 ) );
  MUX \b/U3839  ( .IN0(\b/n3788 ), .IN1(\b/n3780 ), .SEL(msg[56]), .F(
        \b/n3789 ) );
  MUX \b/U3838  ( .IN0(\b/n3787 ), .IN1(\b/n3784 ), .SEL(msg[61]), .F(
        \b/n3788 ) );
  MUX \b/U3837  ( .IN0(\b/n3786 ), .IN1(\b/n3785 ), .SEL(msg[58]), .F(
        \b/n3787 ) );
  MUX \b/U3836  ( .IN0(\b/n630 ), .IN1(msg[57]), .SEL(msg[63]), .F(\b/n3786 )
         );
  MUX \b/U3835  ( .IN0(n662), .IN1(\b/n3663 ), .SEL(msg[63]), .F(\b/n3785 ) );
  MUX \b/U3834  ( .IN0(\b/n3783 ), .IN1(\b/n3782 ), .SEL(msg[58]), .F(
        \b/n3784 ) );
  MUX \b/U3833  ( .IN0(\b/n635 ), .IN1(\b/n629 ), .SEL(msg[63]), .F(\b/n3783 )
         );
  MUX \b/U3832  ( .IN0(n662), .IN1(\b/n3781 ), .SEL(msg[63]), .F(\b/n3782 ) );
  MUX \b/U3831  ( .IN0(\b/n581 ), .IN1(\b/n618 ), .SEL(msg[57]), .F(\b/n3781 )
         );
  MUX \b/U3830  ( .IN0(\b/n3779 ), .IN1(\b/n3773 ), .SEL(msg[61]), .F(
        \b/n3780 ) );
  MUX \b/U3829  ( .IN0(\b/n3776 ), .IN1(\b/n3775 ), .SEL(msg[58]), .F(
        \b/n3779 ) );
  NAND \b/U3828  ( .A(\b/n3777 ), .B(\b/n3778 ), .Z(\b/n3776 ) );
  MUX \b/U3827  ( .IN0(\b/n3649 ), .IN1(\b/n3774 ), .SEL(n660), .F(\b/n3775 )
         );
  MUX \b/U3826  ( .IN0(msg[59]), .IN1(\b/n591 ), .SEL(msg[63]), .F(\b/n3774 )
         );
  MUX \b/U3825  ( .IN0(\b/n3772 ), .IN1(\b/n3771 ), .SEL(msg[58]), .F(
        \b/n3773 ) );
  MUX \b/U3824  ( .IN0(\b/n3694 ), .IN1(\b/n589 ), .SEL(msg[63]), .F(\b/n3772 ) );
  MUX \b/U3823  ( .IN0(\b/n3690 ), .IN1(\b/n3770 ), .SEL(msg[63]), .F(
        \b/n3771 ) );
  MUX \b/U3822  ( .IN0(\b/n3652 ), .IN1(\b/n3657 ), .SEL(msg[57]), .F(
        \b/n3770 ) );
  MUX \b/U3821  ( .IN0(\b/n3769 ), .IN1(\b/n3751 ), .SEL(msg[62]), .F(
        shift_row_out[89]) );
  MUX \b/U3820  ( .IN0(\b/n3768 ), .IN1(\b/n3759 ), .SEL(msg[56]), .F(
        \b/n3769 ) );
  MUX \b/U3819  ( .IN0(\b/n3767 ), .IN1(\b/n3763 ), .SEL(msg[61]), .F(
        \b/n3768 ) );
  MUX \b/U3818  ( .IN0(\b/n3766 ), .IN1(\b/n3765 ), .SEL(msg[58]), .F(
        \b/n3767 ) );
  MUX \b/U3817  ( .IN0(\b/n626 ), .IN1(n664), .SEL(msg[63]), .F(\b/n3766 ) );
  MUX \b/U3816  ( .IN0(\b/n3764 ), .IN1(n658), .SEL(msg[63]), .F(\b/n3765 ) );
  NAND \b/U3815  ( .A(\b/n638 ), .B(\b/n597 ), .Z(\b/n3764 ) );
  MUX \b/U3814  ( .IN0(\b/n3762 ), .IN1(\b/n3761 ), .SEL(msg[58]), .F(
        \b/n3763 ) );
  MUX \b/U3813  ( .IN0(\b/n574 ), .IN1(\b/n3664 ), .SEL(msg[63]), .F(\b/n3762 ) );
  MUX \b/U3812  ( .IN0(\b/n3654 ), .IN1(\b/n3760 ), .SEL(msg[63]), .F(
        \b/n3761 ) );
  AND \b/U3811  ( .A(msg[57]), .B(msg[60]), .Z(\b/n3760 ) );
  MUX \b/U3810  ( .IN0(\b/n3758 ), .IN1(\b/n3755 ), .SEL(msg[61]), .F(
        \b/n3759 ) );
  MUX \b/U3809  ( .IN0(\b/n3757 ), .IN1(\b/n3756 ), .SEL(msg[58]), .F(
        \b/n3758 ) );
  MUX \b/U3808  ( .IN0(\b/n3693 ), .IN1(\b/n635 ), .SEL(msg[63]), .F(\b/n3757 ) );
  MUX \b/U3807  ( .IN0(\b/n610 ), .IN1(\b/n3662 ), .SEL(msg[63]), .F(\b/n3756 ) );
  MUX \b/U3806  ( .IN0(\b/n3752 ), .IN1(\b/n3753 ), .SEL(msg[58]), .F(
        \b/n3755 ) );
  AND \b/U3805  ( .A(\b/n3754 ), .B(\b/n3709 ), .Z(\b/n3753 ) );
  MUX \b/U3804  ( .IN0(\b/n3668 ), .IN1(\b/n3657 ), .SEL(msg[63]), .F(
        \b/n3752 ) );
  MUX \b/U3803  ( .IN0(\b/n3750 ), .IN1(\b/n3742 ), .SEL(msg[56]), .F(
        \b/n3751 ) );
  MUX \b/U3802  ( .IN0(\b/n3749 ), .IN1(\b/n3745 ), .SEL(msg[61]), .F(
        \b/n3750 ) );
  MUX \b/U3801  ( .IN0(\b/n3748 ), .IN1(\b/n3747 ), .SEL(msg[58]), .F(
        \b/n3749 ) );
  MUX \b/U3800  ( .IN0(\b/n3656 ), .IN1(\b/n599 ), .SEL(msg[63]), .F(\b/n3748 ) );
  MUX \b/U3799  ( .IN0(\b/n3746 ), .IN1(\b/n583 ), .SEL(msg[63]), .F(\b/n3747 ) );
  MUX \b/U3798  ( .IN0(\b/n3654 ), .IN1(\b/n591 ), .SEL(msg[57]), .F(\b/n3746 ) );
  MUX \b/U3797  ( .IN0(\b/n3744 ), .IN1(\b/n3743 ), .SEL(msg[58]), .F(
        \b/n3745 ) );
  MUX \b/U3796  ( .IN0(\b/n630 ), .IN1(\b/n608 ), .SEL(msg[63]), .F(\b/n3744 )
         );
  MUX \b/U3795  ( .IN0(\b/n626 ), .IN1(\b/n586 ), .SEL(msg[63]), .F(\b/n3743 )
         );
  MUX \b/U3794  ( .IN0(\b/n3741 ), .IN1(\b/n3736 ), .SEL(msg[61]), .F(
        \b/n3742 ) );
  MUX \b/U3793  ( .IN0(\b/n3740 ), .IN1(\b/n3737 ), .SEL(msg[58]), .F(
        \b/n3741 ) );
  MUX \b/U3792  ( .IN0(\b/n3738 ), .IN1(\b/n3739 ), .SEL(msg[63]), .F(
        \b/n3740 ) );
  NAND \b/U3791  ( .A(\b/n3657 ), .B(\b/n3729 ), .Z(\b/n3739 ) );
  MUX \b/U3790  ( .IN0(\b/n3657 ), .IN1(\b/n591 ), .SEL(msg[57]), .F(\b/n3738 ) );
  MUX \b/U3789  ( .IN0(\b/n3674 ), .IN1(\b/n3672 ), .SEL(msg[63]), .F(
        \b/n3737 ) );
  MUX \b/U3788  ( .IN0(\b/n3692 ), .IN1(\b/n3735 ), .SEL(msg[58]), .F(
        \b/n3736 ) );
  MUX \b/U3787  ( .IN0(\b/n597 ), .IN1(\b/n629 ), .SEL(msg[63]), .F(\b/n3735 )
         );
  MUX \b/U3786  ( .IN0(\b/n3734 ), .IN1(\b/n3717 ), .SEL(msg[62]), .F(
        shift_row_out[88]) );
  MUX \b/U3785  ( .IN0(\b/n3733 ), .IN1(\b/n3725 ), .SEL(msg[56]), .F(
        \b/n3734 ) );
  MUX \b/U3784  ( .IN0(\b/n3732 ), .IN1(\b/n3730 ), .SEL(msg[58]), .F(
        \b/n3733 ) );
  MUX \b/U3783  ( .IN0(\b/n571 ), .IN1(\b/n3731 ), .SEL(msg[63]), .F(\b/n3732 ) );
  MUX \b/U3782  ( .IN0(\b/n624 ), .IN1(\b/n627 ), .SEL(msg[61]), .F(\b/n3731 )
         );
  MUX \b/U3781  ( .IN0(\b/n3727 ), .IN1(\b/n3726 ), .SEL(msg[63]), .F(
        \b/n3730 ) );
  NAND \b/U3780  ( .A(\b/n3728 ), .B(\b/n3729 ), .Z(\b/n3727 ) );
  MUX \b/U3779  ( .IN0(\b/n623 ), .IN1(\b/n638 ), .SEL(msg[61]), .F(\b/n3726 )
         );
  MUX \b/U3778  ( .IN0(\b/n3724 ), .IN1(\b/n3720 ), .SEL(msg[58]), .F(
        \b/n3725 ) );
  MUX \b/U3777  ( .IN0(\b/n3723 ), .IN1(\b/n3721 ), .SEL(msg[63]), .F(
        \b/n3724 ) );
  MUX \b/U3776  ( .IN0(\b/n3722 ), .IN1(\b/n576 ), .SEL(msg[61]), .F(\b/n3723 ) );
  NAND \b/U3775  ( .A(\b/n638 ), .B(\b/n3649 ), .Z(\b/n3722 ) );
  MUX \b/U3773  ( .IN0(\b/n3719 ), .IN1(\b/n3718 ), .SEL(msg[63]), .F(
        \b/n3720 ) );
  MUX \b/U3772  ( .IN0(n659), .IN1(\b/n573 ), .SEL(msg[61]), .F(\b/n3719 ) );
  MUX \b/U3771  ( .IN0(\b/n625 ), .IN1(\b/n581 ), .SEL(msg[61]), .F(\b/n3718 )
         );
  MUX \b/U3770  ( .IN0(\b/n3716 ), .IN1(\b/n3706 ), .SEL(msg[56]), .F(
        \b/n3717 ) );
  MUX \b/U3769  ( .IN0(\b/n3715 ), .IN1(\b/n3711 ), .SEL(msg[58]), .F(
        \b/n3716 ) );
  MUX \b/U3768  ( .IN0(\b/n3714 ), .IN1(\b/n3713 ), .SEL(msg[63]), .F(
        \b/n3715 ) );
  MUX \b/U3767  ( .IN0(n657), .IN1(\b/n577 ), .SEL(msg[61]), .F(\b/n3714 ) );
  MUX \b/U3766  ( .IN0(\b/n3712 ), .IN1(\b/n614 ), .SEL(msg[61]), .F(\b/n3713 ) );
  NAND \b/U3765  ( .A(\b/n3648 ), .B(\b/n3650 ), .Z(\b/n3712 ) );
  MUX \b/U3764  ( .IN0(\b/n3710 ), .IN1(\b/n3707 ), .SEL(msg[63]), .F(
        \b/n3711 ) );
  MUX \b/U3763  ( .IN0(\b/n584 ), .IN1(\b/n3708 ), .SEL(msg[61]), .F(\b/n3710 ) );
  NAND \b/U3762  ( .A(\b/n3652 ), .B(\b/n3709 ), .Z(\b/n3708 ) );
  MUX \b/U3761  ( .IN0(\b/n3667 ), .IN1(\b/n3658 ), .SEL(msg[61]), .F(
        \b/n3707 ) );
  MUX \b/U3760  ( .IN0(\b/n3705 ), .IN1(\b/n3701 ), .SEL(msg[58]), .F(
        \b/n3706 ) );
  MUX \b/U3759  ( .IN0(\b/n3703 ), .IN1(\b/n3702 ), .SEL(msg[63]), .F(
        \b/n3705 ) );
  NAND \b/U3758  ( .A(\b/n3704 ), .B(\b/n3691 ), .Z(\b/n3703 ) );
  MUX \b/U3757  ( .IN0(msg[59]), .IN1(\b/n3683 ), .SEL(msg[61]), .F(\b/n3702 )
         );
  MUX \b/U3756  ( .IN0(\b/n3700 ), .IN1(\b/n3699 ), .SEL(msg[63]), .F(
        \b/n3701 ) );
  MUX \b/U3755  ( .IN0(\b/n589 ), .IN1(\b/n605 ), .SEL(msg[61]), .F(\b/n3700 )
         );
  MUX \b/U3754  ( .IN0(\b/n622 ), .IN1(\b/n610 ), .SEL(msg[61]), .F(\b/n3699 )
         );
  XOR \b/U3753  ( .A(\b/n3649 ), .B(msg[57]), .Z(\b/n3698 ) );
  XOR \b/U3752  ( .A(msg[57]), .B(msg[58]), .Z(\b/n3697 ) );
  XOR \b/U3751  ( .A(msg[57]), .B(msg[59]), .Z(\b/n3696 ) );
  XOR \b/U3750  ( .A(msg[58]), .B(msg[63]), .Z(\b/n3695 ) );
  XOR \b/U3749  ( .A(\b/n638 ), .B(\b/n581 ), .Z(\b/n3694 ) );
  XOR \b/U3748  ( .A(msg[57]), .B(\b/n627 ), .Z(\b/n3693 ) );
  XOR \b/U3746  ( .A(msg[57]), .B(msg[61]), .Z(\b/n3691 ) );
  NAND \b/U3745  ( .A(msg[57]), .B(msg[59]), .Z(\b/n3690 ) );
  MUX \b/U3744  ( .IN0(\b/n3649 ), .IN1(\b/n581 ), .SEL(msg[57]), .F(\b/n3689 ) );
  MUX \b/U3742  ( .IN0(msg[59]), .IN1(\b/n618 ), .SEL(msg[57]), .F(\b/n3687 )
         );
  MUX \b/U3741  ( .IN0(\b/n597 ), .IN1(\b/n618 ), .SEL(msg[57]), .F(\b/n3686 )
         );
  MUX \b/U3740  ( .IN0(\b/n3652 ), .IN1(\b/n3654 ), .SEL(msg[57]), .F(
        \b/n3685 ) );
  MUX \b/U3739  ( .IN0(msg[60]), .IN1(\b/n597 ), .SEL(msg[57]), .F(\b/n3684 )
         );
  OR \b/U3738  ( .A(msg[57]), .B(msg[60]), .Z(\b/n3683 ) );
  NAND \b/U3736  ( .A(\b/n618 ), .B(\b/n638 ), .Z(\b/n3681 ) );
  MUX \b/U3735  ( .IN0(\b/n618 ), .IN1(msg[60]), .SEL(msg[57]), .F(\b/n3680 )
         );
  MUX \b/U3734  ( .IN0(\b/n3648 ), .IN1(\b/n3657 ), .SEL(msg[57]), .F(
        \b/n3679 ) );
  MUX \b/U3733  ( .IN0(\b/n633 ), .IN1(msg[60]), .SEL(msg[57]), .F(\b/n3678 )
         );
  MUX \b/U3732  ( .IN0(\b/n591 ), .IN1(\b/n618 ), .SEL(msg[57]), .F(\b/n3677 )
         );
  MUX \b/U3731  ( .IN0(\b/n3648 ), .IN1(msg[60]), .SEL(msg[57]), .F(\b/n3676 )
         );
  MUX \b/U3730  ( .IN0(\b/n608 ), .IN1(\b/n597 ), .SEL(msg[57]), .F(\b/n3675 )
         );
  XOR \b/U3729  ( .A(\b/n591 ), .B(msg[57]), .Z(\b/n3674 ) );
  MUX \b/U3728  ( .IN0(\b/n3654 ), .IN1(\b/n608 ), .SEL(msg[57]), .F(\b/n3673 ) );
  NANDN \b/U3727  ( .B(msg[57]), .A(msg[59]), .Z(\b/n3672 ) );
  MUX \b/U3726  ( .IN0(\b/n581 ), .IN1(msg[59]), .SEL(msg[57]), .F(\b/n3671 )
         );
  NAND \b/U3724  ( .A(\b/n3652 ), .B(\b/n638 ), .Z(\b/n3669 ) );
  MUX \b/U3723  ( .IN0(msg[60]), .IN1(\b/n3649 ), .SEL(msg[57]), .F(\b/n3668 )
         );
  MUX \b/U3722  ( .IN0(\b/n608 ), .IN1(msg[59]), .SEL(msg[57]), .F(\b/n3667 )
         );
  MUX \b/U3720  ( .IN0(msg[60]), .IN1(\b/n627 ), .SEL(msg[57]), .F(\b/n3665 )
         );
  MUX \b/U3719  ( .IN0(\b/n581 ), .IN1(\b/n633 ), .SEL(msg[57]), .F(\b/n3664 )
         );
  NAND \b/U3718  ( .A(\b/n3650 ), .B(\b/n581 ), .Z(\b/n3663 ) );
  MUX \b/U3717  ( .IN0(\b/n3649 ), .IN1(\b/n3657 ), .SEL(msg[57]), .F(
        \b/n3662 ) );
  NAND \b/U3716  ( .A(\b/n3661 ), .B(\b/n3648 ), .Z(\b/n3660 ) );
  MUX \b/U3715  ( .IN0(\b/n3652 ), .IN1(\b/n633 ), .SEL(msg[57]), .F(\b/n3659 ) );
  MUX \b/U3714  ( .IN0(\b/n633 ), .IN1(\b/n597 ), .SEL(msg[57]), .F(\b/n3658 )
         );
  NANDN \b/U3713  ( .B(msg[59]), .A(msg[60]), .Z(\b/n3657 ) );
  MUX \b/U3712  ( .IN0(\b/n3652 ), .IN1(msg[59]), .SEL(msg[57]), .F(\b/n3656 )
         );
  OR \b/U3711  ( .A(msg[59]), .B(msg[60]), .Z(\b/n3652 ) );
  MUX \b/U3710  ( .IN0(\b/n581 ), .IN1(\b/n597 ), .SEL(msg[57]), .F(\b/n3655 )
         );
  XOR \b/U3709  ( .A(\b/n591 ), .B(msg[59]), .Z(\b/n3654 ) );
  NANDN \b/U3708  ( .B(msg[59]), .A(msg[57]), .Z(\b/n3653 ) );
  NAND \b/U3707  ( .A(\b/n3652 ), .B(\b/n3650 ), .Z(\b/n3651 ) );
  NAND \b/U3706  ( .A(msg[57]), .B(\b/n3649 ), .Z(\b/n3650 ) );
  NANDN \b/U3705  ( .B(msg[60]), .A(msg[59]), .Z(\b/n3649 ) );
  NAND \b/U3704  ( .A(msg[59]), .B(msg[60]), .Z(\b/n3648 ) );
  MUX \b/U3703  ( .IN0(msg[52]), .IN1(\b/n3289 ), .SEL(msg[49]), .F(\b/n3647 )
         );
  MUX \b/U3702  ( .IN0(msg[52]), .IN1(\b/n3298 ), .SEL(msg[49]), .F(\b/n3646 )
         );
  MUX \b/U3701  ( .IN0(\b/n3290 ), .IN1(\b/n3293 ), .SEL(msg[49]), .F(
        \b/n3645 ) );
  MUX \b/U3700  ( .IN0(\b/n3295 ), .IN1(\b/n698 ), .SEL(msg[49]), .F(\b/n3644 ) );
  MUX \b/U3698  ( .IN0(\b/n3298 ), .IN1(\b/n3289 ), .SEL(msg[50]), .F(
        \b/n3471 ) );
  MUX \b/U3697  ( .IN0(\b/n3291 ), .IN1(\b/n709 ), .SEL(msg[50]), .F(\b/n3472 ) );
  MUX \b/U3696  ( .IN0(\b/n652 ), .IN1(\b/n662 ), .SEL(msg[49]), .F(\b/n3435 )
         );
  MUX \b/U3695  ( .IN0(\b/n3319 ), .IN1(\b/n3630 ), .SEL(msg[55]), .F(
        \b/n3642 ) );
  MUX \b/U3694  ( .IN0(\b/n3293 ), .IN1(\b/n3289 ), .SEL(msg[49]), .F(
        \b/n3633 ) );
  MUX \b/U3693  ( .IN0(\b/n704 ), .IN1(\b/n3295 ), .SEL(msg[49]), .F(\b/n3641 ) );
  MUX \b/U3692  ( .IN0(msg[51]), .IN1(\b/n698 ), .SEL(msg[49]), .F(\b/n3640 )
         );
  MUX \b/U3691  ( .IN0(\b/n3298 ), .IN1(\b/n704 ), .SEL(msg[49]), .F(\b/n3639 ) );
  MUX \b/U3690  ( .IN0(msg[52]), .IN1(\b/n3295 ), .SEL(msg[49]), .F(\b/n3638 )
         );
  MUX \b/U3689  ( .IN0(\b/n689 ), .IN1(\b/n668 ), .SEL(msg[53]), .F(\b/n3345 )
         );
  MUX \b/U3688  ( .IN0(\b/n3290 ), .IN1(\b/n662 ), .SEL(msg[49]), .F(\b/n3637 ) );
  NANDN \b/U3685  ( .B(\b/n3296 ), .A(msg[55]), .Z(\b/n3610 ) );
  NAND \b/U3684  ( .A(msg[55]), .B(\b/n665 ), .Z(\b/n3578 ) );
  NAND \b/U3683  ( .A(msg[55]), .B(\b/n677 ), .Z(\b/n3519 ) );
  NAND \b/U3682  ( .A(msg[55]), .B(\b/n3627 ), .Z(\b/n3552 ) );
  NAND \b/U3681  ( .A(msg[55]), .B(\b/n3547 ), .Z(\b/n3510 ) );
  NAND \b/U3679  ( .A(\b/n709 ), .B(\b/n698 ), .Z(\b/n3631 ) );
  NAND \b/U3678  ( .A(msg[55]), .B(\b/n3629 ), .Z(\b/n3624 ) );
  NAND \b/U3677  ( .A(n656), .B(msg[55]), .Z(\b/n3604 ) );
  NAND \b/U3675  ( .A(msg[50]), .B(\b/n3298 ), .Z(\b/n3464 ) );
  NAND \b/U3674  ( .A(\b/n698 ), .B(msg[49]), .Z(\b/n3419 ) );
  NAND \b/U3673  ( .A(msg[55]), .B(\b/n3633 ), .Z(\b/n3418 ) );
  NAND \b/U3671  ( .A(\b/n3631 ), .B(msg[55]), .Z(\b/n3434 ) );
  NAND \b/U3670  ( .A(\b/n3452 ), .B(\b/n3298 ), .Z(\b/n3630 ) );
  NANDN \b/U3669  ( .B(\b/n652 ), .A(\b/n709 ), .Z(\b/n3629 ) );
  NAND \b/U3667  ( .A(msg[49]), .B(\b/n3298 ), .Z(\b/n3350 ) );
  NAND \b/U3666  ( .A(\b/n652 ), .B(\b/n709 ), .Z(\b/n3627 ) );
  NAND \b/U3663  ( .A(msg[49]), .B(\b/n3293 ), .Z(\b/n3452 ) );
  ANDN \b/U3661  ( .A(msg[50]), .B(msg[49]), .Z(\b/n3480 ) );
  AND \b/U3660  ( .A(\b/n3290 ), .B(\b/n3624 ), .Z(\b/n3395 ) );
  MUX \b/U3659  ( .IN0(\b/n3623 ), .IN1(\b/n3607 ), .SEL(msg[54]), .F(
        shift_row_out[119]) );
  MUX \b/U3658  ( .IN0(\b/n3622 ), .IN1(\b/n3615 ), .SEL(msg[48]), .F(
        \b/n3623 ) );
  MUX \b/U3657  ( .IN0(\b/n3621 ), .IN1(\b/n3618 ), .SEL(msg[53]), .F(
        \b/n3622 ) );
  MUX \b/U3656  ( .IN0(\b/n3620 ), .IN1(\b/n3619 ), .SEL(msg[50]), .F(
        \b/n3621 ) );
  MUX \b/U3655  ( .IN0(msg[52]), .IN1(\b/n669 ), .SEL(msg[55]), .F(\b/n3620 )
         );
  MUX \b/U3654  ( .IN0(\b/n3291 ), .IN1(\b/n673 ), .SEL(msg[55]), .F(\b/n3619 ) );
  MUX \b/U3653  ( .IN0(\b/n3617 ), .IN1(\b/n3616 ), .SEL(msg[50]), .F(
        \b/n3618 ) );
  MUX \b/U3652  ( .IN0(\b/n3349 ), .IN1(\b/n665 ), .SEL(msg[55]), .F(\b/n3617 ) );
  MUX \b/U3651  ( .IN0(\b/n3301 ), .IN1(\b/n3312 ), .SEL(msg[55]), .F(
        \b/n3616 ) );
  MUX \b/U3650  ( .IN0(\b/n3614 ), .IN1(\b/n3611 ), .SEL(msg[53]), .F(
        \b/n3615 ) );
  MUX \b/U3649  ( .IN0(\b/n3613 ), .IN1(\b/n3612 ), .SEL(msg[50]), .F(
        \b/n3614 ) );
  MUX \b/U3648  ( .IN0(\b/n3325 ), .IN1(\b/n3300 ), .SEL(msg[55]), .F(
        \b/n3613 ) );
  MUX \b/U3647  ( .IN0(\b/n677 ), .IN1(\b/n3321 ), .SEL(msg[55]), .F(\b/n3612 ) );
  MUX \b/U3646  ( .IN0(\b/n3609 ), .IN1(\b/n3608 ), .SEL(msg[50]), .F(
        \b/n3611 ) );
  AND \b/U3645  ( .A(\b/n667 ), .B(\b/n3610 ), .Z(\b/n3609 ) );
  MUX \b/U3644  ( .IN0(\b/n3305 ), .IN1(n655), .SEL(msg[55]), .F(\b/n3608 ) );
  MUX \b/U3643  ( .IN0(\b/n3606 ), .IN1(\b/n3598 ), .SEL(msg[48]), .F(
        \b/n3607 ) );
  MUX \b/U3642  ( .IN0(\b/n3605 ), .IN1(\b/n3601 ), .SEL(msg[53]), .F(
        \b/n3606 ) );
  MUX \b/U3641  ( .IN0(\b/n3602 ), .IN1(\b/n3603 ), .SEL(msg[50]), .F(
        \b/n3605 ) );
  NAND \b/U3640  ( .A(\b/n3419 ), .B(\b/n3604 ), .Z(\b/n3603 ) );
  MUX \b/U3639  ( .IN0(\b/n707 ), .IN1(\b/n699 ), .SEL(msg[55]), .F(\b/n3602 )
         );
  MUX \b/U3638  ( .IN0(\b/n3600 ), .IN1(\b/n3599 ), .SEL(msg[50]), .F(
        \b/n3601 ) );
  MUX \b/U3637  ( .IN0(\b/n3295 ), .IN1(\b/n3289 ), .SEL(msg[55]), .F(
        \b/n3600 ) );
  MUX \b/U3636  ( .IN0(\b/n700 ), .IN1(\b/n3326 ), .SEL(msg[55]), .F(\b/n3599 ) );
  MUX \b/U3635  ( .IN0(\b/n3597 ), .IN1(\b/n3594 ), .SEL(msg[53]), .F(
        \b/n3598 ) );
  MUX \b/U3634  ( .IN0(\b/n3596 ), .IN1(\b/n3595 ), .SEL(msg[50]), .F(
        \b/n3597 ) );
  MUX \b/U3633  ( .IN0(\b/n3330 ), .IN1(\b/n3316 ), .SEL(msg[55]), .F(
        \b/n3596 ) );
  MUX \b/U3632  ( .IN0(\b/n653 ), .IN1(\b/n3298 ), .SEL(msg[55]), .F(\b/n3595 ) );
  MUX \b/U3631  ( .IN0(\b/n3593 ), .IN1(\b/n3592 ), .SEL(msg[50]), .F(
        \b/n3594 ) );
  MUX \b/U3630  ( .IN0(\b/n3331 ), .IN1(\b/n3339 ), .SEL(msg[55]), .F(
        \b/n3593 ) );
  MUX \b/U3629  ( .IN0(\b/n3324 ), .IN1(\b/n3591 ), .SEL(msg[55]), .F(
        \b/n3592 ) );
  MUX \b/U3628  ( .IN0(\b/n704 ), .IN1(\b/n662 ), .SEL(msg[49]), .F(\b/n3591 )
         );
  MUX \b/U3627  ( .IN0(\b/n3590 ), .IN1(\b/n3572 ), .SEL(msg[54]), .F(
        shift_row_out[118]) );
  MUX \b/U3626  ( .IN0(\b/n3589 ), .IN1(\b/n3580 ), .SEL(msg[48]), .F(
        \b/n3590 ) );
  MUX \b/U3625  ( .IN0(\b/n3588 ), .IN1(\b/n3583 ), .SEL(msg[53]), .F(
        \b/n3589 ) );
  MUX \b/U3624  ( .IN0(\b/n3587 ), .IN1(\b/n3585 ), .SEL(msg[50]), .F(
        \b/n3588 ) );
  MUX \b/U3623  ( .IN0(\b/n3586 ), .IN1(\b/n3302 ), .SEL(msg[55]), .F(
        \b/n3587 ) );
  MUX \b/U3622  ( .IN0(\b/n704 ), .IN1(\b/n3289 ), .SEL(msg[49]), .F(\b/n3586 ) );
  MUX \b/U3621  ( .IN0(\b/n3584 ), .IN1(\b/n692 ), .SEL(msg[55]), .F(\b/n3585 ) );
  MUX \b/U3620  ( .IN0(\b/n3289 ), .IN1(\b/n3290 ), .SEL(msg[49]), .F(
        \b/n3584 ) );
  MUX \b/U3619  ( .IN0(\b/n3582 ), .IN1(\b/n3581 ), .SEL(msg[50]), .F(
        \b/n3583 ) );
  MUX \b/U3618  ( .IN0(n654), .IN1(\b/n3370 ), .SEL(msg[55]), .F(\b/n3582 ) );
  MUX \b/U3617  ( .IN0(\b/n3328 ), .IN1(\b/n3335 ), .SEL(msg[55]), .F(
        \b/n3581 ) );
  MUX \b/U3616  ( .IN0(\b/n3579 ), .IN1(\b/n3575 ), .SEL(msg[53]), .F(
        \b/n3580 ) );
  MUX \b/U3615  ( .IN0(\b/n3577 ), .IN1(\b/n3576 ), .SEL(msg[50]), .F(
        \b/n3579 ) );
  AND \b/U3614  ( .A(\b/n645 ), .B(\b/n3578 ), .Z(\b/n3577 ) );
  MUX \b/U3613  ( .IN0(\b/n3405 ), .IN1(msg[51]), .SEL(msg[55]), .F(\b/n3576 )
         );
  MUX \b/U3612  ( .IN0(\b/n3574 ), .IN1(\b/n3573 ), .SEL(msg[50]), .F(
        \b/n3575 ) );
  MUX \b/U3611  ( .IN0(\b/n688 ), .IN1(\b/n3293 ), .SEL(msg[55]), .F(\b/n3574 ) );
  MUX \b/U3609  ( .IN0(\b/n3571 ), .IN1(\b/n3564 ), .SEL(msg[48]), .F(
        \b/n3572 ) );
  MUX \b/U3608  ( .IN0(\b/n3570 ), .IN1(\b/n3567 ), .SEL(msg[53]), .F(
        \b/n3571 ) );
  MUX \b/U3607  ( .IN0(\b/n3569 ), .IN1(\b/n3568 ), .SEL(msg[50]), .F(
        \b/n3570 ) );
  MUX \b/U3606  ( .IN0(\b/n684 ), .IN1(\b/n3297 ), .SEL(msg[55]), .F(\b/n3569 ) );
  MUX \b/U3605  ( .IN0(\b/n3301 ), .IN1(n655), .SEL(msg[55]), .F(\b/n3568 ) );
  MUX \b/U3604  ( .IN0(\b/n3566 ), .IN1(\b/n3565 ), .SEL(msg[50]), .F(
        \b/n3567 ) );
  MUX \b/U3603  ( .IN0(\b/n3317 ), .IN1(\b/n649 ), .SEL(msg[55]), .F(\b/n3566 ) );
  MUX \b/U3602  ( .IN0(\b/n669 ), .IN1(\b/n699 ), .SEL(msg[55]), .F(\b/n3565 )
         );
  MUX \b/U3601  ( .IN0(\b/n3563 ), .IN1(\b/n3559 ), .SEL(msg[53]), .F(
        \b/n3564 ) );
  MUX \b/U3600  ( .IN0(\b/n3562 ), .IN1(\b/n3561 ), .SEL(msg[50]), .F(
        \b/n3563 ) );
  MUX \b/U3599  ( .IN0(\b/n3306 ), .IN1(\b/n699 ), .SEL(msg[55]), .F(\b/n3562 ) );
  MUX \b/U3598  ( .IN0(\b/n3560 ), .IN1(\b/n3327 ), .SEL(msg[55]), .F(
        \b/n3561 ) );
  NANDN \b/U3597  ( .B(msg[52]), .A(msg[49]), .Z(\b/n3560 ) );
  MUX \b/U3596  ( .IN0(\b/n3558 ), .IN1(\b/n3556 ), .SEL(msg[50]), .F(
        \b/n3559 ) );
  MUX \b/U3595  ( .IN0(\b/n662 ), .IN1(\b/n3557 ), .SEL(msg[55]), .F(\b/n3558 ) );
  MUX \b/U3594  ( .IN0(\b/n689 ), .IN1(\b/n679 ), .SEL(msg[49]), .F(\b/n3557 )
         );
  MUX \b/U3593  ( .IN0(\b/n651 ), .IN1(\b/n3302 ), .SEL(msg[55]), .F(\b/n3556 ) );
  NANDN \b/U3592  ( .B(\b/n652 ), .A(msg[49]), .Z(\b/n3302 ) );
  MUX \b/U3591  ( .IN0(\b/n3555 ), .IN1(\b/n3534 ), .SEL(msg[54]), .F(
        shift_row_out[117]) );
  MUX \b/U3590  ( .IN0(\b/n3554 ), .IN1(\b/n3544 ), .SEL(msg[48]), .F(
        \b/n3555 ) );
  MUX \b/U3589  ( .IN0(\b/n3553 ), .IN1(\b/n3549 ), .SEL(msg[53]), .F(
        \b/n3554 ) );
  MUX \b/U3588  ( .IN0(\b/n3550 ), .IN1(\b/n3551 ), .SEL(msg[50]), .F(
        \b/n3553 ) );
  AND \b/U3587  ( .A(\b/n3320 ), .B(\b/n3552 ), .Z(\b/n3551 ) );
  MUX \b/U3586  ( .IN0(\b/n3298 ), .IN1(\b/n700 ), .SEL(msg[55]), .F(\b/n3550 ) );
  MUX \b/U3585  ( .IN0(\b/n3548 ), .IN1(\b/n3546 ), .SEL(msg[50]), .F(
        \b/n3549 ) );
  MUX \b/U3584  ( .IN0(\b/n655 ), .IN1(\b/n3547 ), .SEL(msg[55]), .F(\b/n3548 ) );
  NAND \b/U3583  ( .A(\b/n679 ), .B(\b/n709 ), .Z(\b/n3547 ) );
  MUX \b/U3582  ( .IN0(\b/n3298 ), .IN1(\b/n3545 ), .SEL(msg[55]), .F(
        \b/n3546 ) );
  NAND \b/U3581  ( .A(\b/n3289 ), .B(\b/n3350 ), .Z(\b/n3545 ) );
  MUX \b/U3580  ( .IN0(\b/n3543 ), .IN1(\b/n3539 ), .SEL(msg[53]), .F(
        \b/n3544 ) );
  MUX \b/U3579  ( .IN0(\b/n3542 ), .IN1(\b/n3541 ), .SEL(msg[50]), .F(
        \b/n3543 ) );
  MUX \b/U3578  ( .IN0(\b/n3310 ), .IN1(\b/n702 ), .SEL(msg[55]), .F(\b/n3542 ) );
  MUX \b/U3577  ( .IN0(\b/n3335 ), .IN1(\b/n3540 ), .SEL(msg[55]), .F(
        \b/n3541 ) );
  MUX \b/U3576  ( .IN0(\b/n698 ), .IN1(\b/n679 ), .SEL(msg[49]), .F(\b/n3540 )
         );
  MUX \b/U3575  ( .IN0(\b/n3538 ), .IN1(\b/n3537 ), .SEL(msg[50]), .F(
        \b/n3539 ) );
  MUX \b/U3574  ( .IN0(\b/n696 ), .IN1(n653), .SEL(msg[55]), .F(\b/n3538 ) );
  MUX \b/U3573  ( .IN0(\b/n3536 ), .IN1(\b/n3535 ), .SEL(msg[55]), .F(
        \b/n3537 ) );
  AND \b/U3572  ( .A(\b/n3295 ), .B(\b/n3370 ), .Z(\b/n3536 ) );
  MUX \b/U3571  ( .IN0(\b/n668 ), .IN1(\b/n652 ), .SEL(msg[49]), .F(\b/n3535 )
         );
  MUX \b/U3570  ( .IN0(\b/n3533 ), .IN1(\b/n3524 ), .SEL(msg[48]), .F(
        \b/n3534 ) );
  MUX \b/U3569  ( .IN0(\b/n3532 ), .IN1(\b/n3528 ), .SEL(msg[53]), .F(
        \b/n3533 ) );
  MUX \b/U3568  ( .IN0(\b/n3531 ), .IN1(\b/n3529 ), .SEL(msg[50]), .F(
        \b/n3532 ) );
  MUX \b/U3567  ( .IN0(\b/n3301 ), .IN1(\b/n3530 ), .SEL(msg[55]), .F(
        \b/n3531 ) );
  NAND \b/U3566  ( .A(msg[49]), .B(\b/n668 ), .Z(\b/n3530 ) );
  MUX \b/U3565  ( .IN0(\b/n652 ), .IN1(\b/n705 ), .SEL(msg[55]), .F(\b/n3529 )
         );
  MUX \b/U3564  ( .IN0(\b/n3527 ), .IN1(\b/n3526 ), .SEL(msg[50]), .F(
        \b/n3528 ) );
  MUX \b/U3563  ( .IN0(\b/n3327 ), .IN1(\b/n670 ), .SEL(msg[55]), .F(\b/n3527 ) );
  MUX \b/U3562  ( .IN0(\b/n3525 ), .IN1(\b/n3290 ), .SEL(n652), .F(\b/n3526 )
         );
  AND \b/U3561  ( .A(msg[55]), .B(msg[51]), .Z(\b/n3525 ) );
  MUX \b/U3560  ( .IN0(\b/n3523 ), .IN1(\b/n3520 ), .SEL(msg[53]), .F(
        \b/n3524 ) );
  MUX \b/U3559  ( .IN0(\b/n3522 ), .IN1(\b/n3521 ), .SEL(msg[50]), .F(
        \b/n3523 ) );
  MUX \b/U3558  ( .IN0(\b/n3451 ), .IN1(\b/n3290 ), .SEL(msg[55]), .F(
        \b/n3522 ) );
  MUX \b/U3557  ( .IN0(n651), .IN1(\b/n703 ), .SEL(msg[55]), .F(\b/n3521 ) );
  MUX \b/U3556  ( .IN0(\b/n3518 ), .IN1(\b/n3517 ), .SEL(msg[50]), .F(
        \b/n3520 ) );
  AND \b/U3555  ( .A(\b/n3519 ), .B(\b/n3419 ), .Z(\b/n3518 ) );
  MUX \b/U3554  ( .IN0(\b/n654 ), .IN1(\b/n698 ), .SEL(msg[55]), .F(\b/n3517 )
         );
  MUX \b/U3553  ( .IN0(\b/n3516 ), .IN1(\b/n3499 ), .SEL(msg[54]), .F(
        shift_row_out[116]) );
  MUX \b/U3552  ( .IN0(\b/n3515 ), .IN1(\b/n3507 ), .SEL(msg[48]), .F(
        \b/n3516 ) );
  MUX \b/U3551  ( .IN0(\b/n3514 ), .IN1(\b/n3511 ), .SEL(msg[53]), .F(
        \b/n3515 ) );
  MUX \b/U3550  ( .IN0(\b/n3513 ), .IN1(\b/n3512 ), .SEL(msg[50]), .F(
        \b/n3514 ) );
  MUX \b/U3549  ( .IN0(\b/n680 ), .IN1(\b/n701 ), .SEL(msg[55]), .F(\b/n3513 )
         );
  MUX \b/U3548  ( .IN0(\b/n3370 ), .IN1(\b/n3335 ), .SEL(msg[55]), .F(
        \b/n3512 ) );
  NAND \b/U3547  ( .A(msg[49]), .B(\b/n3289 ), .Z(\b/n3370 ) );
  MUX \b/U3546  ( .IN0(\b/n3508 ), .IN1(\b/n3509 ), .SEL(msg[50]), .F(
        \b/n3511 ) );
  AND \b/U3545  ( .A(\b/n3320 ), .B(\b/n3510 ), .Z(\b/n3509 ) );
  MUX \b/U3544  ( .IN0(\b/n3318 ), .IN1(\b/n683 ), .SEL(msg[55]), .F(\b/n3508 ) );
  MUX \b/U3543  ( .IN0(\b/n3506 ), .IN1(\b/n3503 ), .SEL(msg[53]), .F(
        \b/n3507 ) );
  MUX \b/U3542  ( .IN0(\b/n3505 ), .IN1(\b/n3504 ), .SEL(msg[50]), .F(
        \b/n3506 ) );
  MUX \b/U3541  ( .IN0(\b/n645 ), .IN1(\b/n691 ), .SEL(msg[55]), .F(\b/n3505 )
         );
  MUX \b/U3540  ( .IN0(\b/n652 ), .IN1(\b/n3298 ), .SEL(msg[55]), .F(\b/n3504 ) );
  MUX \b/U3539  ( .IN0(\b/n3502 ), .IN1(\b/n3500 ), .SEL(msg[50]), .F(
        \b/n3503 ) );
  MUX \b/U3538  ( .IN0(\b/n3314 ), .IN1(\b/n3501 ), .SEL(msg[55]), .F(
        \b/n3502 ) );
  AND \b/U3537  ( .A(\b/n3298 ), .B(\b/n709 ), .Z(\b/n3501 ) );
  MUX \b/U3536  ( .IN0(\b/n667 ), .IN1(\b/n686 ), .SEL(msg[55]), .F(\b/n3500 )
         );
  MUX \b/U3535  ( .IN0(\b/n3498 ), .IN1(\b/n3492 ), .SEL(msg[48]), .F(
        \b/n3499 ) );
  MUX \b/U3534  ( .IN0(\b/n3497 ), .IN1(\b/n3495 ), .SEL(msg[53]), .F(
        \b/n3498 ) );
  MUX \b/U3533  ( .IN0(\b/n3496 ), .IN1(\b/n3292 ), .SEL(msg[50]), .F(
        \b/n3497 ) );
  MUX \b/U3532  ( .IN0(\b/n3312 ), .IN1(\b/n688 ), .SEL(msg[55]), .F(\b/n3496 ) );
  MUX \b/U3531  ( .IN0(\b/n3494 ), .IN1(\b/n3493 ), .SEL(msg[50]), .F(
        \b/n3495 ) );
  MUX \b/U3530  ( .IN0(n650), .IN1(\b/n680 ), .SEL(msg[55]), .F(\b/n3494 ) );
  MUX \b/U3529  ( .IN0(\b/n3322 ), .IN1(\b/n3325 ), .SEL(msg[55]), .F(
        \b/n3493 ) );
  MUX \b/U3528  ( .IN0(\b/n3491 ), .IN1(\b/n3488 ), .SEL(msg[53]), .F(
        \b/n3492 ) );
  MUX \b/U3527  ( .IN0(\b/n3490 ), .IN1(\b/n3489 ), .SEL(msg[50]), .F(
        \b/n3491 ) );
  MUX \b/U3526  ( .IN0(\b/n653 ), .IN1(\b/n3294 ), .SEL(msg[55]), .F(\b/n3490 ) );
  MUX \b/U3525  ( .IN0(\b/n698 ), .IN1(\b/n3316 ), .SEL(msg[55]), .F(\b/n3489 ) );
  MUX \b/U3524  ( .IN0(\b/n641 ), .IN1(\b/n3487 ), .SEL(msg[50]), .F(\b/n3488 ) );
  MUX \b/U3523  ( .IN0(\b/n661 ), .IN1(\b/n3298 ), .SEL(msg[55]), .F(\b/n3487 ) );
  MUX \b/U3522  ( .IN0(\b/n3486 ), .IN1(\b/n3467 ), .SEL(msg[54]), .F(
        shift_row_out[115]) );
  MUX \b/U3521  ( .IN0(\b/n3485 ), .IN1(\b/n3477 ), .SEL(msg[48]), .F(
        \b/n3486 ) );
  MUX \b/U3520  ( .IN0(\b/n3484 ), .IN1(\b/n3481 ), .SEL(msg[53]), .F(
        \b/n3485 ) );
  MUX \b/U3519  ( .IN0(\b/n3483 ), .IN1(\b/n3482 ), .SEL(msg[55]), .F(
        \b/n3484 ) );
  MUX \b/U3518  ( .IN0(\b/n3306 ), .IN1(\b/n686 ), .SEL(msg[50]), .F(\b/n3483 ) );
  MUX \b/U3517  ( .IN0(n653), .IN1(\b/n644 ), .SEL(msg[50]), .F(\b/n3482 ) );
  MUX \b/U3516  ( .IN0(\b/n3479 ), .IN1(\b/n3478 ), .SEL(msg[55]), .F(
        \b/n3481 ) );
  AND \b/U3515  ( .A(\b/n3480 ), .B(msg[52]), .Z(\b/n3479 ) );
  MUX \b/U3514  ( .IN0(\b/n674 ), .IN1(\b/n3319 ), .SEL(msg[50]), .F(\b/n3478 ) );
  MUX \b/U3513  ( .IN0(\b/n3476 ), .IN1(\b/n3473 ), .SEL(msg[53]), .F(
        \b/n3477 ) );
  MUX \b/U3512  ( .IN0(\b/n3475 ), .IN1(\b/n3474 ), .SEL(msg[55]), .F(
        \b/n3476 ) );
  MUX \b/U3511  ( .IN0(\b/n3310 ), .IN1(n649), .SEL(msg[50]), .F(\b/n3475 ) );
  MUX \b/U3510  ( .IN0(\b/n642 ), .IN1(\b/n661 ), .SEL(msg[50]), .F(\b/n3474 )
         );
  MUX \b/U3509  ( .IN0(\b/n3469 ), .IN1(\b/n3470 ), .SEL(msg[55]), .F(
        \b/n3473 ) );
  NAND \b/U3508  ( .A(\b/n3471 ), .B(\b/n3472 ), .Z(\b/n3470 ) );
  MUX \b/U3507  ( .IN0(\b/n687 ), .IN1(\b/n3468 ), .SEL(msg[50]), .F(\b/n3469 ) );
  MUX \b/U3506  ( .IN0(\b/n662 ), .IN1(\b/n704 ), .SEL(msg[49]), .F(\b/n3468 )
         );
  MUX \b/U3505  ( .IN0(\b/n3466 ), .IN1(\b/n3457 ), .SEL(msg[48]), .F(
        \b/n3467 ) );
  MUX \b/U3504  ( .IN0(\b/n3465 ), .IN1(\b/n3461 ), .SEL(msg[53]), .F(
        \b/n3466 ) );
  MUX \b/U3503  ( .IN0(\b/n3463 ), .IN1(\b/n3462 ), .SEL(msg[55]), .F(
        \b/n3465 ) );
  NAND \b/U3502  ( .A(\b/n652 ), .B(\b/n3464 ), .Z(\b/n3463 ) );
  MUX \b/U3501  ( .IN0(\b/n703 ), .IN1(\b/n665 ), .SEL(msg[50]), .F(\b/n3462 )
         );
  MUX \b/U3500  ( .IN0(\b/n3460 ), .IN1(\b/n3458 ), .SEL(msg[55]), .F(
        \b/n3461 ) );
  MUX \b/U3499  ( .IN0(\b/n3301 ), .IN1(\b/n3459 ), .SEL(msg[50]), .F(
        \b/n3460 ) );
  AND \b/U3498  ( .A(msg[49]), .B(\b/n652 ), .Z(\b/n3459 ) );
  MUX \b/U3497  ( .IN0(\b/n657 ), .IN1(\b/n3320 ), .SEL(msg[50]), .F(\b/n3458 ) );
  MUX \b/U3496  ( .IN0(\b/n3456 ), .IN1(\b/n3450 ), .SEL(msg[53]), .F(
        \b/n3457 ) );
  MUX \b/U3495  ( .IN0(\b/n3455 ), .IN1(\b/n3453 ), .SEL(msg[55]), .F(
        \b/n3456 ) );
  MUX \b/U3494  ( .IN0(\b/n3454 ), .IN1(\b/n3290 ), .SEL(\b/n3338 ), .F(
        \b/n3455 ) );
  MUX \b/U3493  ( .IN0(msg[51]), .IN1(msg[52]), .SEL(msg[50]), .F(\b/n3454 )
         );
  MUX \b/U3492  ( .IN0(\b/n3320 ), .IN1(\b/n3451 ), .SEL(msg[50]), .F(
        \b/n3453 ) );
  NAND \b/U3491  ( .A(\b/n3290 ), .B(\b/n3452 ), .Z(\b/n3451 ) );
  MUX \b/U3490  ( .IN0(\b/n3447 ), .IN1(\b/n3448 ), .SEL(msg[55]), .F(
        \b/n3450 ) );
  AND \b/U3489  ( .A(\b/n685 ), .B(\b/n3449 ), .Z(\b/n3448 ) );
  MUX \b/U3488  ( .IN0(\b/n666 ), .IN1(\b/n3291 ), .SEL(msg[50]), .F(\b/n3447 ) );
  MUX \b/U3487  ( .IN0(\b/n3446 ), .IN1(\b/n3430 ), .SEL(msg[54]), .F(
        shift_row_out[114]) );
  MUX \b/U3486  ( .IN0(\b/n3445 ), .IN1(\b/n3437 ), .SEL(msg[48]), .F(
        \b/n3446 ) );
  MUX \b/U3485  ( .IN0(\b/n3444 ), .IN1(\b/n3440 ), .SEL(msg[53]), .F(
        \b/n3445 ) );
  MUX \b/U3484  ( .IN0(\b/n3443 ), .IN1(\b/n3441 ), .SEL(msg[50]), .F(
        \b/n3444 ) );
  MUX \b/U3483  ( .IN0(\b/n674 ), .IN1(\b/n3442 ), .SEL(msg[55]), .F(\b/n3443 ) );
  MUX \b/U3482  ( .IN0(\b/n3298 ), .IN1(\b/n652 ), .SEL(msg[49]), .F(\b/n3442 ) );
  MUX \b/U3481  ( .IN0(\b/n3337 ), .IN1(\b/n692 ), .SEL(msg[55]), .F(\b/n3441 ) );
  MUX \b/U3480  ( .IN0(\b/n3439 ), .IN1(\b/n3438 ), .SEL(msg[50]), .F(
        \b/n3440 ) );
  MUX \b/U3479  ( .IN0(\b/n3291 ), .IN1(\b/n659 ), .SEL(msg[55]), .F(\b/n3439 ) );
  MUX \b/U3478  ( .IN0(\b/n695 ), .IN1(\b/n3324 ), .SEL(msg[55]), .F(\b/n3438 ) );
  MUX \b/U3477  ( .IN0(\b/n3436 ), .IN1(\b/n3432 ), .SEL(msg[53]), .F(
        \b/n3437 ) );
  MUX \b/U3476  ( .IN0(\b/n3433 ), .IN1(\b/n641 ), .SEL(msg[50]), .F(\b/n3436 ) );
  NAND \b/U3475  ( .A(\b/n3434 ), .B(\b/n3435 ), .Z(\b/n3433 ) );
  MUX \b/U3474  ( .IN0(n651), .IN1(\b/n3431 ), .SEL(\b/n3336 ), .F(\b/n3432 )
         );
  MUX \b/U3473  ( .IN0(\b/n673 ), .IN1(\b/n3303 ), .SEL(msg[50]), .F(\b/n3431 ) );
  MUX \b/U3472  ( .IN0(\b/n3429 ), .IN1(\b/n3421 ), .SEL(msg[48]), .F(
        \b/n3430 ) );
  MUX \b/U3471  ( .IN0(\b/n3428 ), .IN1(\b/n3425 ), .SEL(msg[53]), .F(
        \b/n3429 ) );
  MUX \b/U3470  ( .IN0(\b/n3427 ), .IN1(\b/n3426 ), .SEL(msg[50]), .F(
        \b/n3428 ) );
  MUX \b/U3469  ( .IN0(\b/n701 ), .IN1(msg[49]), .SEL(msg[55]), .F(\b/n3427 )
         );
  MUX \b/U3468  ( .IN0(n654), .IN1(\b/n3304 ), .SEL(msg[55]), .F(\b/n3426 ) );
  MUX \b/U3467  ( .IN0(\b/n3424 ), .IN1(\b/n3423 ), .SEL(msg[50]), .F(
        \b/n3425 ) );
  MUX \b/U3466  ( .IN0(\b/n706 ), .IN1(\b/n700 ), .SEL(msg[55]), .F(\b/n3424 )
         );
  MUX \b/U3465  ( .IN0(n654), .IN1(\b/n3422 ), .SEL(msg[55]), .F(\b/n3423 ) );
  MUX \b/U3464  ( .IN0(\b/n652 ), .IN1(\b/n689 ), .SEL(msg[49]), .F(\b/n3422 )
         );
  MUX \b/U3463  ( .IN0(\b/n3420 ), .IN1(\b/n3414 ), .SEL(msg[53]), .F(
        \b/n3421 ) );
  MUX \b/U3462  ( .IN0(\b/n3417 ), .IN1(\b/n3416 ), .SEL(msg[50]), .F(
        \b/n3420 ) );
  NAND \b/U3461  ( .A(\b/n3418 ), .B(\b/n3419 ), .Z(\b/n3417 ) );
  MUX \b/U3460  ( .IN0(\b/n3290 ), .IN1(\b/n3415 ), .SEL(n652), .F(\b/n3416 )
         );
  MUX \b/U3459  ( .IN0(msg[51]), .IN1(\b/n662 ), .SEL(msg[55]), .F(\b/n3415 )
         );
  MUX \b/U3458  ( .IN0(\b/n3413 ), .IN1(\b/n3412 ), .SEL(msg[50]), .F(
        \b/n3414 ) );
  MUX \b/U3457  ( .IN0(\b/n3335 ), .IN1(\b/n660 ), .SEL(msg[55]), .F(\b/n3413 ) );
  MUX \b/U3456  ( .IN0(\b/n3331 ), .IN1(\b/n3411 ), .SEL(msg[55]), .F(
        \b/n3412 ) );
  MUX \b/U3455  ( .IN0(\b/n3293 ), .IN1(\b/n3298 ), .SEL(msg[49]), .F(
        \b/n3411 ) );
  MUX \b/U3454  ( .IN0(\b/n3410 ), .IN1(\b/n3392 ), .SEL(msg[54]), .F(
        shift_row_out[113]) );
  MUX \b/U3453  ( .IN0(\b/n3409 ), .IN1(\b/n3400 ), .SEL(msg[48]), .F(
        \b/n3410 ) );
  MUX \b/U3452  ( .IN0(\b/n3408 ), .IN1(\b/n3404 ), .SEL(msg[53]), .F(
        \b/n3409 ) );
  MUX \b/U3451  ( .IN0(\b/n3407 ), .IN1(\b/n3406 ), .SEL(msg[50]), .F(
        \b/n3408 ) );
  MUX \b/U3450  ( .IN0(\b/n697 ), .IN1(n656), .SEL(msg[55]), .F(\b/n3407 ) );
  MUX \b/U3449  ( .IN0(\b/n3405 ), .IN1(n650), .SEL(msg[55]), .F(\b/n3406 ) );
  NAND \b/U3448  ( .A(\b/n709 ), .B(\b/n668 ), .Z(\b/n3405 ) );
  MUX \b/U3447  ( .IN0(\b/n3403 ), .IN1(\b/n3402 ), .SEL(msg[50]), .F(
        \b/n3404 ) );
  MUX \b/U3446  ( .IN0(\b/n645 ), .IN1(\b/n3305 ), .SEL(msg[55]), .F(\b/n3403 ) );
  MUX \b/U3445  ( .IN0(\b/n3295 ), .IN1(\b/n3401 ), .SEL(msg[55]), .F(
        \b/n3402 ) );
  AND \b/U3444  ( .A(msg[49]), .B(msg[52]), .Z(\b/n3401 ) );
  MUX \b/U3443  ( .IN0(\b/n3399 ), .IN1(\b/n3396 ), .SEL(msg[53]), .F(
        \b/n3400 ) );
  MUX \b/U3442  ( .IN0(\b/n3398 ), .IN1(\b/n3397 ), .SEL(msg[50]), .F(
        \b/n3399 ) );
  MUX \b/U3441  ( .IN0(\b/n3334 ), .IN1(\b/n706 ), .SEL(msg[55]), .F(\b/n3398 ) );
  MUX \b/U3440  ( .IN0(\b/n681 ), .IN1(\b/n3303 ), .SEL(msg[55]), .F(\b/n3397 ) );
  MUX \b/U3439  ( .IN0(\b/n3393 ), .IN1(\b/n3394 ), .SEL(msg[50]), .F(
        \b/n3396 ) );
  AND \b/U3438  ( .A(\b/n3395 ), .B(\b/n3350 ), .Z(\b/n3394 ) );
  MUX \b/U3437  ( .IN0(\b/n3309 ), .IN1(\b/n3298 ), .SEL(msg[55]), .F(
        \b/n3393 ) );
  MUX \b/U3436  ( .IN0(\b/n3391 ), .IN1(\b/n3383 ), .SEL(msg[48]), .F(
        \b/n3392 ) );
  MUX \b/U3435  ( .IN0(\b/n3390 ), .IN1(\b/n3386 ), .SEL(msg[53]), .F(
        \b/n3391 ) );
  MUX \b/U3434  ( .IN0(\b/n3389 ), .IN1(\b/n3388 ), .SEL(msg[50]), .F(
        \b/n3390 ) );
  MUX \b/U3433  ( .IN0(\b/n3297 ), .IN1(\b/n670 ), .SEL(msg[55]), .F(\b/n3389 ) );
  MUX \b/U3432  ( .IN0(\b/n3387 ), .IN1(\b/n654 ), .SEL(msg[55]), .F(\b/n3388 ) );
  MUX \b/U3431  ( .IN0(\b/n3295 ), .IN1(\b/n662 ), .SEL(msg[49]), .F(\b/n3387 ) );
  MUX \b/U3430  ( .IN0(\b/n3385 ), .IN1(\b/n3384 ), .SEL(msg[50]), .F(
        \b/n3386 ) );
  MUX \b/U3429  ( .IN0(\b/n701 ), .IN1(\b/n679 ), .SEL(msg[55]), .F(\b/n3385 )
         );
  MUX \b/U3428  ( .IN0(\b/n697 ), .IN1(\b/n657 ), .SEL(msg[55]), .F(\b/n3384 )
         );
  MUX \b/U3427  ( .IN0(\b/n3382 ), .IN1(\b/n3377 ), .SEL(msg[53]), .F(
        \b/n3383 ) );
  MUX \b/U3426  ( .IN0(\b/n3381 ), .IN1(\b/n3378 ), .SEL(msg[50]), .F(
        \b/n3382 ) );
  MUX \b/U3425  ( .IN0(\b/n3379 ), .IN1(\b/n3380 ), .SEL(msg[55]), .F(
        \b/n3381 ) );
  NAND \b/U3424  ( .A(\b/n3298 ), .B(\b/n3370 ), .Z(\b/n3380 ) );
  MUX \b/U3423  ( .IN0(\b/n3298 ), .IN1(\b/n662 ), .SEL(msg[49]), .F(\b/n3379 ) );
  MUX \b/U3422  ( .IN0(\b/n3315 ), .IN1(\b/n3313 ), .SEL(msg[55]), .F(
        \b/n3378 ) );
  MUX \b/U3421  ( .IN0(\b/n3333 ), .IN1(\b/n3376 ), .SEL(msg[50]), .F(
        \b/n3377 ) );
  MUX \b/U3420  ( .IN0(\b/n668 ), .IN1(\b/n700 ), .SEL(msg[55]), .F(\b/n3376 )
         );
  MUX \b/U3419  ( .IN0(\b/n3375 ), .IN1(\b/n3358 ), .SEL(msg[54]), .F(
        shift_row_out[112]) );
  MUX \b/U3418  ( .IN0(\b/n3374 ), .IN1(\b/n3366 ), .SEL(msg[48]), .F(
        \b/n3375 ) );
  MUX \b/U3417  ( .IN0(\b/n3373 ), .IN1(\b/n3371 ), .SEL(msg[50]), .F(
        \b/n3374 ) );
  MUX \b/U3416  ( .IN0(\b/n642 ), .IN1(\b/n3372 ), .SEL(msg[55]), .F(\b/n3373 ) );
  MUX \b/U3415  ( .IN0(\b/n695 ), .IN1(\b/n698 ), .SEL(msg[53]), .F(\b/n3372 )
         );
  MUX \b/U3414  ( .IN0(\b/n3368 ), .IN1(\b/n3367 ), .SEL(msg[55]), .F(
        \b/n3371 ) );
  NAND \b/U3413  ( .A(\b/n3369 ), .B(\b/n3370 ), .Z(\b/n3368 ) );
  MUX \b/U3412  ( .IN0(\b/n694 ), .IN1(\b/n709 ), .SEL(msg[53]), .F(\b/n3367 )
         );
  MUX \b/U3411  ( .IN0(\b/n3365 ), .IN1(\b/n3361 ), .SEL(msg[50]), .F(
        \b/n3366 ) );
  MUX \b/U3410  ( .IN0(\b/n3364 ), .IN1(\b/n3362 ), .SEL(msg[55]), .F(
        \b/n3365 ) );
  MUX \b/U3409  ( .IN0(\b/n3363 ), .IN1(\b/n647 ), .SEL(msg[53]), .F(\b/n3364 ) );
  NAND \b/U3408  ( .A(\b/n709 ), .B(\b/n3290 ), .Z(\b/n3363 ) );
  MUX \b/U3406  ( .IN0(\b/n3360 ), .IN1(\b/n3359 ), .SEL(msg[55]), .F(
        \b/n3361 ) );
  MUX \b/U3405  ( .IN0(n651), .IN1(\b/n644 ), .SEL(msg[53]), .F(\b/n3360 ) );
  MUX \b/U3404  ( .IN0(\b/n696 ), .IN1(\b/n652 ), .SEL(msg[53]), .F(\b/n3359 )
         );
  MUX \b/U3403  ( .IN0(\b/n3357 ), .IN1(\b/n3347 ), .SEL(msg[48]), .F(
        \b/n3358 ) );
  MUX \b/U3402  ( .IN0(\b/n3356 ), .IN1(\b/n3352 ), .SEL(msg[50]), .F(
        \b/n3357 ) );
  MUX \b/U3401  ( .IN0(\b/n3355 ), .IN1(\b/n3354 ), .SEL(msg[55]), .F(
        \b/n3356 ) );
  MUX \b/U3400  ( .IN0(n649), .IN1(\b/n648 ), .SEL(msg[53]), .F(\b/n3355 ) );
  MUX \b/U3399  ( .IN0(\b/n3353 ), .IN1(\b/n685 ), .SEL(msg[53]), .F(\b/n3354 ) );
  NAND \b/U3398  ( .A(\b/n3289 ), .B(\b/n3291 ), .Z(\b/n3353 ) );
  MUX \b/U3397  ( .IN0(\b/n3351 ), .IN1(\b/n3348 ), .SEL(msg[55]), .F(
        \b/n3352 ) );
  MUX \b/U3396  ( .IN0(\b/n655 ), .IN1(\b/n3349 ), .SEL(msg[53]), .F(\b/n3351 ) );
  NAND \b/U3395  ( .A(\b/n3293 ), .B(\b/n3350 ), .Z(\b/n3349 ) );
  MUX \b/U3394  ( .IN0(\b/n3308 ), .IN1(\b/n3299 ), .SEL(msg[53]), .F(
        \b/n3348 ) );
  MUX \b/U3393  ( .IN0(\b/n3346 ), .IN1(\b/n3342 ), .SEL(msg[50]), .F(
        \b/n3347 ) );
  MUX \b/U3392  ( .IN0(\b/n3344 ), .IN1(\b/n3343 ), .SEL(msg[55]), .F(
        \b/n3346 ) );
  NAND \b/U3391  ( .A(\b/n3345 ), .B(\b/n3332 ), .Z(\b/n3344 ) );
  MUX \b/U3390  ( .IN0(msg[51]), .IN1(\b/n3324 ), .SEL(msg[53]), .F(\b/n3343 )
         );
  MUX \b/U3389  ( .IN0(\b/n3341 ), .IN1(\b/n3340 ), .SEL(msg[55]), .F(
        \b/n3342 ) );
  MUX \b/U3388  ( .IN0(\b/n660 ), .IN1(\b/n676 ), .SEL(msg[53]), .F(\b/n3341 )
         );
  MUX \b/U3387  ( .IN0(\b/n693 ), .IN1(\b/n681 ), .SEL(msg[53]), .F(\b/n3340 )
         );
  XOR \b/U3386  ( .A(\b/n3290 ), .B(msg[49]), .Z(\b/n3339 ) );
  XOR \b/U3385  ( .A(msg[49]), .B(msg[50]), .Z(\b/n3338 ) );
  XOR \b/U3384  ( .A(msg[49]), .B(msg[51]), .Z(\b/n3337 ) );
  XOR \b/U3383  ( .A(msg[50]), .B(msg[55]), .Z(\b/n3336 ) );
  XOR \b/U3382  ( .A(\b/n709 ), .B(\b/n652 ), .Z(\b/n3335 ) );
  XOR \b/U3381  ( .A(msg[49]), .B(\b/n698 ), .Z(\b/n3334 ) );
  XOR \b/U3379  ( .A(msg[49]), .B(msg[53]), .Z(\b/n3332 ) );
  NAND \b/U3378  ( .A(msg[49]), .B(msg[51]), .Z(\b/n3331 ) );
  MUX \b/U3377  ( .IN0(\b/n3290 ), .IN1(\b/n652 ), .SEL(msg[49]), .F(\b/n3330 ) );
  MUX \b/U3375  ( .IN0(msg[51]), .IN1(\b/n689 ), .SEL(msg[49]), .F(\b/n3328 )
         );
  MUX \b/U3374  ( .IN0(\b/n668 ), .IN1(\b/n689 ), .SEL(msg[49]), .F(\b/n3327 )
         );
  MUX \b/U3373  ( .IN0(\b/n3293 ), .IN1(\b/n3295 ), .SEL(msg[49]), .F(
        \b/n3326 ) );
  MUX \b/U3372  ( .IN0(msg[52]), .IN1(\b/n668 ), .SEL(msg[49]), .F(\b/n3325 )
         );
  OR \b/U3371  ( .A(msg[49]), .B(msg[52]), .Z(\b/n3324 ) );
  NAND \b/U3369  ( .A(\b/n689 ), .B(\b/n709 ), .Z(\b/n3322 ) );
  MUX \b/U3368  ( .IN0(\b/n689 ), .IN1(msg[52]), .SEL(msg[49]), .F(\b/n3321 )
         );
  MUX \b/U3367  ( .IN0(\b/n3289 ), .IN1(\b/n3298 ), .SEL(msg[49]), .F(
        \b/n3320 ) );
  MUX \b/U3366  ( .IN0(\b/n704 ), .IN1(msg[52]), .SEL(msg[49]), .F(\b/n3319 )
         );
  MUX \b/U3365  ( .IN0(\b/n662 ), .IN1(\b/n689 ), .SEL(msg[49]), .F(\b/n3318 )
         );
  MUX \b/U3364  ( .IN0(\b/n3289 ), .IN1(msg[52]), .SEL(msg[49]), .F(\b/n3317 )
         );
  MUX \b/U3363  ( .IN0(\b/n679 ), .IN1(\b/n668 ), .SEL(msg[49]), .F(\b/n3316 )
         );
  XOR \b/U3362  ( .A(\b/n662 ), .B(msg[49]), .Z(\b/n3315 ) );
  MUX \b/U3361  ( .IN0(\b/n3295 ), .IN1(\b/n679 ), .SEL(msg[49]), .F(\b/n3314 ) );
  NANDN \b/U3360  ( .B(msg[49]), .A(msg[51]), .Z(\b/n3313 ) );
  MUX \b/U3359  ( .IN0(\b/n652 ), .IN1(msg[51]), .SEL(msg[49]), .F(\b/n3312 )
         );
  NAND \b/U3357  ( .A(\b/n3293 ), .B(\b/n709 ), .Z(\b/n3310 ) );
  MUX \b/U3356  ( .IN0(msg[52]), .IN1(\b/n3290 ), .SEL(msg[49]), .F(\b/n3309 )
         );
  MUX \b/U3355  ( .IN0(\b/n679 ), .IN1(msg[51]), .SEL(msg[49]), .F(\b/n3308 )
         );
  MUX \b/U3353  ( .IN0(msg[52]), .IN1(\b/n698 ), .SEL(msg[49]), .F(\b/n3306 )
         );
  MUX \b/U3352  ( .IN0(\b/n652 ), .IN1(\b/n704 ), .SEL(msg[49]), .F(\b/n3305 )
         );
  NAND \b/U3351  ( .A(\b/n3291 ), .B(\b/n652 ), .Z(\b/n3304 ) );
  MUX \b/U3350  ( .IN0(\b/n3290 ), .IN1(\b/n3298 ), .SEL(msg[49]), .F(
        \b/n3303 ) );
  NAND \b/U3349  ( .A(\b/n3302 ), .B(\b/n3289 ), .Z(\b/n3301 ) );
  MUX \b/U3348  ( .IN0(\b/n3293 ), .IN1(\b/n704 ), .SEL(msg[49]), .F(\b/n3300 ) );
  MUX \b/U3347  ( .IN0(\b/n704 ), .IN1(\b/n668 ), .SEL(msg[49]), .F(\b/n3299 )
         );
  NANDN \b/U3346  ( .B(msg[51]), .A(msg[52]), .Z(\b/n3298 ) );
  MUX \b/U3345  ( .IN0(\b/n3293 ), .IN1(msg[51]), .SEL(msg[49]), .F(\b/n3297 )
         );
  OR \b/U3344  ( .A(msg[51]), .B(msg[52]), .Z(\b/n3293 ) );
  MUX \b/U3343  ( .IN0(\b/n652 ), .IN1(\b/n668 ), .SEL(msg[49]), .F(\b/n3296 )
         );
  XOR \b/U3342  ( .A(\b/n662 ), .B(msg[51]), .Z(\b/n3295 ) );
  NANDN \b/U3341  ( .B(msg[51]), .A(msg[49]), .Z(\b/n3294 ) );
  NAND \b/U3340  ( .A(\b/n3293 ), .B(\b/n3291 ), .Z(\b/n3292 ) );
  NAND \b/U3339  ( .A(msg[49]), .B(\b/n3290 ), .Z(\b/n3291 ) );
  NANDN \b/U3338  ( .B(msg[52]), .A(msg[51]), .Z(\b/n3290 ) );
  NAND \b/U3337  ( .A(msg[51]), .B(msg[52]), .Z(\b/n3289 ) );
  MUX \b/U3336  ( .IN0(msg[44]), .IN1(\b/n2930 ), .SEL(msg[41]), .F(\b/n3288 )
         );
  MUX \b/U3335  ( .IN0(msg[44]), .IN1(\b/n2939 ), .SEL(msg[41]), .F(\b/n3287 )
         );
  MUX \b/U3334  ( .IN0(\b/n2931 ), .IN1(\b/n2934 ), .SEL(msg[41]), .F(
        \b/n3286 ) );
  MUX \b/U3333  ( .IN0(\b/n2936 ), .IN1(\b/n769 ), .SEL(msg[41]), .F(\b/n3285 ) );
  MUX \b/U3331  ( .IN0(\b/n2939 ), .IN1(\b/n2930 ), .SEL(msg[42]), .F(
        \b/n3112 ) );
  MUX \b/U3330  ( .IN0(\b/n2932 ), .IN1(\b/n780 ), .SEL(msg[42]), .F(\b/n3113 ) );
  MUX \b/U3329  ( .IN0(\b/n723 ), .IN1(\b/n733 ), .SEL(msg[41]), .F(\b/n3076 )
         );
  MUX \b/U3328  ( .IN0(\b/n2960 ), .IN1(\b/n3271 ), .SEL(msg[47]), .F(
        \b/n3283 ) );
  MUX \b/U3327  ( .IN0(\b/n2934 ), .IN1(\b/n2930 ), .SEL(msg[41]), .F(
        \b/n3274 ) );
  MUX \b/U3326  ( .IN0(\b/n775 ), .IN1(\b/n2936 ), .SEL(msg[41]), .F(\b/n3282 ) );
  MUX \b/U3325  ( .IN0(msg[43]), .IN1(\b/n769 ), .SEL(msg[41]), .F(\b/n3281 )
         );
  MUX \b/U3324  ( .IN0(\b/n2939 ), .IN1(\b/n775 ), .SEL(msg[41]), .F(\b/n3280 ) );
  MUX \b/U3323  ( .IN0(msg[44]), .IN1(\b/n2936 ), .SEL(msg[41]), .F(\b/n3279 )
         );
  MUX \b/U3322  ( .IN0(\b/n760 ), .IN1(\b/n739 ), .SEL(msg[45]), .F(\b/n2986 )
         );
  MUX \b/U3321  ( .IN0(\b/n2931 ), .IN1(\b/n733 ), .SEL(msg[41]), .F(\b/n3278 ) );
  NANDN \b/U3318  ( .B(\b/n2937 ), .A(msg[47]), .Z(\b/n3251 ) );
  NAND \b/U3317  ( .A(msg[47]), .B(\b/n736 ), .Z(\b/n3219 ) );
  NAND \b/U3316  ( .A(msg[47]), .B(\b/n748 ), .Z(\b/n3160 ) );
  NAND \b/U3315  ( .A(msg[47]), .B(\b/n3268 ), .Z(\b/n3193 ) );
  NAND \b/U3314  ( .A(msg[47]), .B(\b/n3188 ), .Z(\b/n3151 ) );
  NAND \b/U3312  ( .A(\b/n780 ), .B(\b/n769 ), .Z(\b/n3272 ) );
  NAND \b/U3311  ( .A(msg[47]), .B(\b/n3270 ), .Z(\b/n3265 ) );
  NAND \b/U3310  ( .A(n648), .B(msg[47]), .Z(\b/n3245 ) );
  NAND \b/U3308  ( .A(msg[42]), .B(\b/n2939 ), .Z(\b/n3105 ) );
  NAND \b/U3307  ( .A(\b/n769 ), .B(msg[41]), .Z(\b/n3060 ) );
  NAND \b/U3306  ( .A(msg[47]), .B(\b/n3274 ), .Z(\b/n3059 ) );
  NAND \b/U3304  ( .A(\b/n3272 ), .B(msg[47]), .Z(\b/n3075 ) );
  NAND \b/U3303  ( .A(\b/n3093 ), .B(\b/n2939 ), .Z(\b/n3271 ) );
  NANDN \b/U3302  ( .B(\b/n723 ), .A(\b/n780 ), .Z(\b/n3270 ) );
  NAND \b/U3300  ( .A(msg[41]), .B(\b/n2939 ), .Z(\b/n2991 ) );
  NAND \b/U3299  ( .A(\b/n723 ), .B(\b/n780 ), .Z(\b/n3268 ) );
  NAND \b/U3296  ( .A(msg[41]), .B(\b/n2934 ), .Z(\b/n3093 ) );
  ANDN \b/U3294  ( .A(msg[42]), .B(msg[41]), .Z(\b/n3121 ) );
  AND \b/U3293  ( .A(\b/n2931 ), .B(\b/n3265 ), .Z(\b/n3036 ) );
  MUX \b/U3292  ( .IN0(\b/n3264 ), .IN1(\b/n3248 ), .SEL(msg[46]), .F(
        shift_row_out[15]) );
  MUX \b/U3291  ( .IN0(\b/n3263 ), .IN1(\b/n3256 ), .SEL(msg[40]), .F(
        \b/n3264 ) );
  MUX \b/U3290  ( .IN0(\b/n3262 ), .IN1(\b/n3259 ), .SEL(msg[45]), .F(
        \b/n3263 ) );
  MUX \b/U3289  ( .IN0(\b/n3261 ), .IN1(\b/n3260 ), .SEL(msg[42]), .F(
        \b/n3262 ) );
  MUX \b/U3288  ( .IN0(msg[44]), .IN1(\b/n740 ), .SEL(msg[47]), .F(\b/n3261 )
         );
  MUX \b/U3287  ( .IN0(\b/n2932 ), .IN1(\b/n744 ), .SEL(msg[47]), .F(\b/n3260 ) );
  MUX \b/U3286  ( .IN0(\b/n3258 ), .IN1(\b/n3257 ), .SEL(msg[42]), .F(
        \b/n3259 ) );
  MUX \b/U3285  ( .IN0(\b/n2990 ), .IN1(\b/n736 ), .SEL(msg[47]), .F(\b/n3258 ) );
  MUX \b/U3284  ( .IN0(\b/n2942 ), .IN1(\b/n2953 ), .SEL(msg[47]), .F(
        \b/n3257 ) );
  MUX \b/U3283  ( .IN0(\b/n3255 ), .IN1(\b/n3252 ), .SEL(msg[45]), .F(
        \b/n3256 ) );
  MUX \b/U3282  ( .IN0(\b/n3254 ), .IN1(\b/n3253 ), .SEL(msg[42]), .F(
        \b/n3255 ) );
  MUX \b/U3281  ( .IN0(\b/n2966 ), .IN1(\b/n2941 ), .SEL(msg[47]), .F(
        \b/n3254 ) );
  MUX \b/U3280  ( .IN0(\b/n748 ), .IN1(\b/n2962 ), .SEL(msg[47]), .F(\b/n3253 ) );
  MUX \b/U3279  ( .IN0(\b/n3250 ), .IN1(\b/n3249 ), .SEL(msg[42]), .F(
        \b/n3252 ) );
  AND \b/U3278  ( .A(\b/n738 ), .B(\b/n3251 ), .Z(\b/n3250 ) );
  MUX \b/U3277  ( .IN0(\b/n2946 ), .IN1(n647), .SEL(msg[47]), .F(\b/n3249 ) );
  MUX \b/U3276  ( .IN0(\b/n3247 ), .IN1(\b/n3239 ), .SEL(msg[40]), .F(
        \b/n3248 ) );
  MUX \b/U3275  ( .IN0(\b/n3246 ), .IN1(\b/n3242 ), .SEL(msg[45]), .F(
        \b/n3247 ) );
  MUX \b/U3274  ( .IN0(\b/n3243 ), .IN1(\b/n3244 ), .SEL(msg[42]), .F(
        \b/n3246 ) );
  NAND \b/U3273  ( .A(\b/n3060 ), .B(\b/n3245 ), .Z(\b/n3244 ) );
  MUX \b/U3272  ( .IN0(\b/n778 ), .IN1(\b/n770 ), .SEL(msg[47]), .F(\b/n3243 )
         );
  MUX \b/U3271  ( .IN0(\b/n3241 ), .IN1(\b/n3240 ), .SEL(msg[42]), .F(
        \b/n3242 ) );
  MUX \b/U3270  ( .IN0(\b/n2936 ), .IN1(\b/n2930 ), .SEL(msg[47]), .F(
        \b/n3241 ) );
  MUX \b/U3269  ( .IN0(\b/n771 ), .IN1(\b/n2967 ), .SEL(msg[47]), .F(\b/n3240 ) );
  MUX \b/U3268  ( .IN0(\b/n3238 ), .IN1(\b/n3235 ), .SEL(msg[45]), .F(
        \b/n3239 ) );
  MUX \b/U3267  ( .IN0(\b/n3237 ), .IN1(\b/n3236 ), .SEL(msg[42]), .F(
        \b/n3238 ) );
  MUX \b/U3266  ( .IN0(\b/n2971 ), .IN1(\b/n2957 ), .SEL(msg[47]), .F(
        \b/n3237 ) );
  MUX \b/U3265  ( .IN0(\b/n724 ), .IN1(\b/n2939 ), .SEL(msg[47]), .F(\b/n3236 ) );
  MUX \b/U3264  ( .IN0(\b/n3234 ), .IN1(\b/n3233 ), .SEL(msg[42]), .F(
        \b/n3235 ) );
  MUX \b/U3263  ( .IN0(\b/n2972 ), .IN1(\b/n2980 ), .SEL(msg[47]), .F(
        \b/n3234 ) );
  MUX \b/U3262  ( .IN0(\b/n2965 ), .IN1(\b/n3232 ), .SEL(msg[47]), .F(
        \b/n3233 ) );
  MUX \b/U3261  ( .IN0(\b/n775 ), .IN1(\b/n733 ), .SEL(msg[41]), .F(\b/n3232 )
         );
  MUX \b/U3260  ( .IN0(\b/n3231 ), .IN1(\b/n3213 ), .SEL(msg[46]), .F(
        shift_row_out[14]) );
  MUX \b/U3259  ( .IN0(\b/n3230 ), .IN1(\b/n3221 ), .SEL(msg[40]), .F(
        \b/n3231 ) );
  MUX \b/U3258  ( .IN0(\b/n3229 ), .IN1(\b/n3224 ), .SEL(msg[45]), .F(
        \b/n3230 ) );
  MUX \b/U3257  ( .IN0(\b/n3228 ), .IN1(\b/n3226 ), .SEL(msg[42]), .F(
        \b/n3229 ) );
  MUX \b/U3256  ( .IN0(\b/n3227 ), .IN1(\b/n2943 ), .SEL(msg[47]), .F(
        \b/n3228 ) );
  MUX \b/U3255  ( .IN0(\b/n775 ), .IN1(\b/n2930 ), .SEL(msg[41]), .F(\b/n3227 ) );
  MUX \b/U3254  ( .IN0(\b/n3225 ), .IN1(\b/n763 ), .SEL(msg[47]), .F(\b/n3226 ) );
  MUX \b/U3253  ( .IN0(\b/n2930 ), .IN1(\b/n2931 ), .SEL(msg[41]), .F(
        \b/n3225 ) );
  MUX \b/U3252  ( .IN0(\b/n3223 ), .IN1(\b/n3222 ), .SEL(msg[42]), .F(
        \b/n3224 ) );
  MUX \b/U3251  ( .IN0(n646), .IN1(\b/n3011 ), .SEL(msg[47]), .F(\b/n3223 ) );
  MUX \b/U3250  ( .IN0(\b/n2969 ), .IN1(\b/n2976 ), .SEL(msg[47]), .F(
        \b/n3222 ) );
  MUX \b/U3249  ( .IN0(\b/n3220 ), .IN1(\b/n3216 ), .SEL(msg[45]), .F(
        \b/n3221 ) );
  MUX \b/U3248  ( .IN0(\b/n3218 ), .IN1(\b/n3217 ), .SEL(msg[42]), .F(
        \b/n3220 ) );
  AND \b/U3247  ( .A(\b/n716 ), .B(\b/n3219 ), .Z(\b/n3218 ) );
  MUX \b/U3246  ( .IN0(\b/n3046 ), .IN1(msg[43]), .SEL(msg[47]), .F(\b/n3217 )
         );
  MUX \b/U3245  ( .IN0(\b/n3215 ), .IN1(\b/n3214 ), .SEL(msg[42]), .F(
        \b/n3216 ) );
  MUX \b/U3244  ( .IN0(\b/n759 ), .IN1(\b/n2934 ), .SEL(msg[47]), .F(\b/n3215 ) );
  MUX \b/U3242  ( .IN0(\b/n3212 ), .IN1(\b/n3205 ), .SEL(msg[40]), .F(
        \b/n3213 ) );
  MUX \b/U3241  ( .IN0(\b/n3211 ), .IN1(\b/n3208 ), .SEL(msg[45]), .F(
        \b/n3212 ) );
  MUX \b/U3240  ( .IN0(\b/n3210 ), .IN1(\b/n3209 ), .SEL(msg[42]), .F(
        \b/n3211 ) );
  MUX \b/U3239  ( .IN0(\b/n755 ), .IN1(\b/n2938 ), .SEL(msg[47]), .F(\b/n3210 ) );
  MUX \b/U3238  ( .IN0(\b/n2942 ), .IN1(n647), .SEL(msg[47]), .F(\b/n3209 ) );
  MUX \b/U3237  ( .IN0(\b/n3207 ), .IN1(\b/n3206 ), .SEL(msg[42]), .F(
        \b/n3208 ) );
  MUX \b/U3236  ( .IN0(\b/n2958 ), .IN1(\b/n720 ), .SEL(msg[47]), .F(\b/n3207 ) );
  MUX \b/U3235  ( .IN0(\b/n740 ), .IN1(\b/n770 ), .SEL(msg[47]), .F(\b/n3206 )
         );
  MUX \b/U3234  ( .IN0(\b/n3204 ), .IN1(\b/n3200 ), .SEL(msg[45]), .F(
        \b/n3205 ) );
  MUX \b/U3233  ( .IN0(\b/n3203 ), .IN1(\b/n3202 ), .SEL(msg[42]), .F(
        \b/n3204 ) );
  MUX \b/U3232  ( .IN0(\b/n2947 ), .IN1(\b/n770 ), .SEL(msg[47]), .F(\b/n3203 ) );
  MUX \b/U3231  ( .IN0(\b/n3201 ), .IN1(\b/n2968 ), .SEL(msg[47]), .F(
        \b/n3202 ) );
  NANDN \b/U3230  ( .B(msg[44]), .A(msg[41]), .Z(\b/n3201 ) );
  MUX \b/U3229  ( .IN0(\b/n3199 ), .IN1(\b/n3197 ), .SEL(msg[42]), .F(
        \b/n3200 ) );
  MUX \b/U3228  ( .IN0(\b/n733 ), .IN1(\b/n3198 ), .SEL(msg[47]), .F(\b/n3199 ) );
  MUX \b/U3227  ( .IN0(\b/n760 ), .IN1(\b/n750 ), .SEL(msg[41]), .F(\b/n3198 )
         );
  MUX \b/U3226  ( .IN0(\b/n722 ), .IN1(\b/n2943 ), .SEL(msg[47]), .F(\b/n3197 ) );
  NANDN \b/U3225  ( .B(\b/n723 ), .A(msg[41]), .Z(\b/n2943 ) );
  MUX \b/U3224  ( .IN0(\b/n3196 ), .IN1(\b/n3175 ), .SEL(msg[46]), .F(
        shift_row_out[13]) );
  MUX \b/U3223  ( .IN0(\b/n3195 ), .IN1(\b/n3185 ), .SEL(msg[40]), .F(
        \b/n3196 ) );
  MUX \b/U3222  ( .IN0(\b/n3194 ), .IN1(\b/n3190 ), .SEL(msg[45]), .F(
        \b/n3195 ) );
  MUX \b/U3221  ( .IN0(\b/n3191 ), .IN1(\b/n3192 ), .SEL(msg[42]), .F(
        \b/n3194 ) );
  AND \b/U3220  ( .A(\b/n2961 ), .B(\b/n3193 ), .Z(\b/n3192 ) );
  MUX \b/U3219  ( .IN0(\b/n2939 ), .IN1(\b/n771 ), .SEL(msg[47]), .F(\b/n3191 ) );
  MUX \b/U3218  ( .IN0(\b/n3189 ), .IN1(\b/n3187 ), .SEL(msg[42]), .F(
        \b/n3190 ) );
  MUX \b/U3217  ( .IN0(\b/n726 ), .IN1(\b/n3188 ), .SEL(msg[47]), .F(\b/n3189 ) );
  NAND \b/U3216  ( .A(\b/n750 ), .B(\b/n780 ), .Z(\b/n3188 ) );
  MUX \b/U3215  ( .IN0(\b/n2939 ), .IN1(\b/n3186 ), .SEL(msg[47]), .F(
        \b/n3187 ) );
  NAND \b/U3214  ( .A(\b/n2930 ), .B(\b/n2991 ), .Z(\b/n3186 ) );
  MUX \b/U3213  ( .IN0(\b/n3184 ), .IN1(\b/n3180 ), .SEL(msg[45]), .F(
        \b/n3185 ) );
  MUX \b/U3212  ( .IN0(\b/n3183 ), .IN1(\b/n3182 ), .SEL(msg[42]), .F(
        \b/n3184 ) );
  MUX \b/U3211  ( .IN0(\b/n2951 ), .IN1(\b/n773 ), .SEL(msg[47]), .F(\b/n3183 ) );
  MUX \b/U3210  ( .IN0(\b/n2976 ), .IN1(\b/n3181 ), .SEL(msg[47]), .F(
        \b/n3182 ) );
  MUX \b/U3209  ( .IN0(\b/n769 ), .IN1(\b/n750 ), .SEL(msg[41]), .F(\b/n3181 )
         );
  MUX \b/U3208  ( .IN0(\b/n3179 ), .IN1(\b/n3178 ), .SEL(msg[42]), .F(
        \b/n3180 ) );
  MUX \b/U3207  ( .IN0(\b/n767 ), .IN1(n645), .SEL(msg[47]), .F(\b/n3179 ) );
  MUX \b/U3206  ( .IN0(\b/n3177 ), .IN1(\b/n3176 ), .SEL(msg[47]), .F(
        \b/n3178 ) );
  AND \b/U3205  ( .A(\b/n2936 ), .B(\b/n3011 ), .Z(\b/n3177 ) );
  MUX \b/U3204  ( .IN0(\b/n739 ), .IN1(\b/n723 ), .SEL(msg[41]), .F(\b/n3176 )
         );
  MUX \b/U3203  ( .IN0(\b/n3174 ), .IN1(\b/n3165 ), .SEL(msg[40]), .F(
        \b/n3175 ) );
  MUX \b/U3202  ( .IN0(\b/n3173 ), .IN1(\b/n3169 ), .SEL(msg[45]), .F(
        \b/n3174 ) );
  MUX \b/U3201  ( .IN0(\b/n3172 ), .IN1(\b/n3170 ), .SEL(msg[42]), .F(
        \b/n3173 ) );
  MUX \b/U3200  ( .IN0(\b/n2942 ), .IN1(\b/n3171 ), .SEL(msg[47]), .F(
        \b/n3172 ) );
  NAND \b/U3199  ( .A(msg[41]), .B(\b/n739 ), .Z(\b/n3171 ) );
  MUX \b/U3198  ( .IN0(\b/n723 ), .IN1(\b/n776 ), .SEL(msg[47]), .F(\b/n3170 )
         );
  MUX \b/U3197  ( .IN0(\b/n3168 ), .IN1(\b/n3167 ), .SEL(msg[42]), .F(
        \b/n3169 ) );
  MUX \b/U3196  ( .IN0(\b/n2968 ), .IN1(\b/n741 ), .SEL(msg[47]), .F(\b/n3168 ) );
  MUX \b/U3195  ( .IN0(\b/n3166 ), .IN1(\b/n2931 ), .SEL(n644), .F(\b/n3167 )
         );
  AND \b/U3194  ( .A(msg[47]), .B(msg[43]), .Z(\b/n3166 ) );
  MUX \b/U3193  ( .IN0(\b/n3164 ), .IN1(\b/n3161 ), .SEL(msg[45]), .F(
        \b/n3165 ) );
  MUX \b/U3192  ( .IN0(\b/n3163 ), .IN1(\b/n3162 ), .SEL(msg[42]), .F(
        \b/n3164 ) );
  MUX \b/U3191  ( .IN0(\b/n3092 ), .IN1(\b/n2931 ), .SEL(msg[47]), .F(
        \b/n3163 ) );
  MUX \b/U3190  ( .IN0(n643), .IN1(\b/n774 ), .SEL(msg[47]), .F(\b/n3162 ) );
  MUX \b/U3189  ( .IN0(\b/n3159 ), .IN1(\b/n3158 ), .SEL(msg[42]), .F(
        \b/n3161 ) );
  AND \b/U3188  ( .A(\b/n3160 ), .B(\b/n3060 ), .Z(\b/n3159 ) );
  MUX \b/U3187  ( .IN0(\b/n725 ), .IN1(\b/n769 ), .SEL(msg[47]), .F(\b/n3158 )
         );
  MUX \b/U3186  ( .IN0(\b/n3157 ), .IN1(\b/n3140 ), .SEL(msg[46]), .F(
        shift_row_out[12]) );
  MUX \b/U3185  ( .IN0(\b/n3156 ), .IN1(\b/n3148 ), .SEL(msg[40]), .F(
        \b/n3157 ) );
  MUX \b/U3184  ( .IN0(\b/n3155 ), .IN1(\b/n3152 ), .SEL(msg[45]), .F(
        \b/n3156 ) );
  MUX \b/U3183  ( .IN0(\b/n3154 ), .IN1(\b/n3153 ), .SEL(msg[42]), .F(
        \b/n3155 ) );
  MUX \b/U3182  ( .IN0(\b/n751 ), .IN1(\b/n772 ), .SEL(msg[47]), .F(\b/n3154 )
         );
  MUX \b/U3181  ( .IN0(\b/n3011 ), .IN1(\b/n2976 ), .SEL(msg[47]), .F(
        \b/n3153 ) );
  NAND \b/U3180  ( .A(msg[41]), .B(\b/n2930 ), .Z(\b/n3011 ) );
  MUX \b/U3179  ( .IN0(\b/n3149 ), .IN1(\b/n3150 ), .SEL(msg[42]), .F(
        \b/n3152 ) );
  AND \b/U3178  ( .A(\b/n2961 ), .B(\b/n3151 ), .Z(\b/n3150 ) );
  MUX \b/U3177  ( .IN0(\b/n2959 ), .IN1(\b/n754 ), .SEL(msg[47]), .F(\b/n3149 ) );
  MUX \b/U3176  ( .IN0(\b/n3147 ), .IN1(\b/n3144 ), .SEL(msg[45]), .F(
        \b/n3148 ) );
  MUX \b/U3175  ( .IN0(\b/n3146 ), .IN1(\b/n3145 ), .SEL(msg[42]), .F(
        \b/n3147 ) );
  MUX \b/U3174  ( .IN0(\b/n716 ), .IN1(\b/n762 ), .SEL(msg[47]), .F(\b/n3146 )
         );
  MUX \b/U3173  ( .IN0(\b/n723 ), .IN1(\b/n2939 ), .SEL(msg[47]), .F(\b/n3145 ) );
  MUX \b/U3172  ( .IN0(\b/n3143 ), .IN1(\b/n3141 ), .SEL(msg[42]), .F(
        \b/n3144 ) );
  MUX \b/U3171  ( .IN0(\b/n2955 ), .IN1(\b/n3142 ), .SEL(msg[47]), .F(
        \b/n3143 ) );
  AND \b/U3170  ( .A(\b/n2939 ), .B(\b/n780 ), .Z(\b/n3142 ) );
  MUX \b/U3169  ( .IN0(\b/n738 ), .IN1(\b/n757 ), .SEL(msg[47]), .F(\b/n3141 )
         );
  MUX \b/U3168  ( .IN0(\b/n3139 ), .IN1(\b/n3133 ), .SEL(msg[40]), .F(
        \b/n3140 ) );
  MUX \b/U3167  ( .IN0(\b/n3138 ), .IN1(\b/n3136 ), .SEL(msg[45]), .F(
        \b/n3139 ) );
  MUX \b/U3166  ( .IN0(\b/n3137 ), .IN1(\b/n2933 ), .SEL(msg[42]), .F(
        \b/n3138 ) );
  MUX \b/U3165  ( .IN0(\b/n2953 ), .IN1(\b/n759 ), .SEL(msg[47]), .F(\b/n3137 ) );
  MUX \b/U3164  ( .IN0(\b/n3135 ), .IN1(\b/n3134 ), .SEL(msg[42]), .F(
        \b/n3136 ) );
  MUX \b/U3163  ( .IN0(n642), .IN1(\b/n751 ), .SEL(msg[47]), .F(\b/n3135 ) );
  MUX \b/U3162  ( .IN0(\b/n2963 ), .IN1(\b/n2966 ), .SEL(msg[47]), .F(
        \b/n3134 ) );
  MUX \b/U3161  ( .IN0(\b/n3132 ), .IN1(\b/n3129 ), .SEL(msg[45]), .F(
        \b/n3133 ) );
  MUX \b/U3160  ( .IN0(\b/n3131 ), .IN1(\b/n3130 ), .SEL(msg[42]), .F(
        \b/n3132 ) );
  MUX \b/U3159  ( .IN0(\b/n724 ), .IN1(\b/n2935 ), .SEL(msg[47]), .F(\b/n3131 ) );
  MUX \b/U3158  ( .IN0(\b/n769 ), .IN1(\b/n2957 ), .SEL(msg[47]), .F(\b/n3130 ) );
  MUX \b/U3157  ( .IN0(\b/n712 ), .IN1(\b/n3128 ), .SEL(msg[42]), .F(\b/n3129 ) );
  MUX \b/U3156  ( .IN0(\b/n732 ), .IN1(\b/n2939 ), .SEL(msg[47]), .F(\b/n3128 ) );
  MUX \b/U3155  ( .IN0(\b/n3127 ), .IN1(\b/n3108 ), .SEL(msg[46]), .F(
        shift_row_out[11]) );
  MUX \b/U3154  ( .IN0(\b/n3126 ), .IN1(\b/n3118 ), .SEL(msg[40]), .F(
        \b/n3127 ) );
  MUX \b/U3153  ( .IN0(\b/n3125 ), .IN1(\b/n3122 ), .SEL(msg[45]), .F(
        \b/n3126 ) );
  MUX \b/U3152  ( .IN0(\b/n3124 ), .IN1(\b/n3123 ), .SEL(msg[47]), .F(
        \b/n3125 ) );
  MUX \b/U3151  ( .IN0(\b/n2947 ), .IN1(\b/n757 ), .SEL(msg[42]), .F(\b/n3124 ) );
  MUX \b/U3150  ( .IN0(n645), .IN1(\b/n715 ), .SEL(msg[42]), .F(\b/n3123 ) );
  MUX \b/U3149  ( .IN0(\b/n3120 ), .IN1(\b/n3119 ), .SEL(msg[47]), .F(
        \b/n3122 ) );
  AND \b/U3148  ( .A(\b/n3121 ), .B(msg[44]), .Z(\b/n3120 ) );
  MUX \b/U3147  ( .IN0(\b/n745 ), .IN1(\b/n2960 ), .SEL(msg[42]), .F(\b/n3119 ) );
  MUX \b/U3146  ( .IN0(\b/n3117 ), .IN1(\b/n3114 ), .SEL(msg[45]), .F(
        \b/n3118 ) );
  MUX \b/U3145  ( .IN0(\b/n3116 ), .IN1(\b/n3115 ), .SEL(msg[47]), .F(
        \b/n3117 ) );
  MUX \b/U3144  ( .IN0(\b/n2951 ), .IN1(n641), .SEL(msg[42]), .F(\b/n3116 ) );
  MUX \b/U3143  ( .IN0(\b/n713 ), .IN1(\b/n732 ), .SEL(msg[42]), .F(\b/n3115 )
         );
  MUX \b/U3142  ( .IN0(\b/n3110 ), .IN1(\b/n3111 ), .SEL(msg[47]), .F(
        \b/n3114 ) );
  NAND \b/U3141  ( .A(\b/n3112 ), .B(\b/n3113 ), .Z(\b/n3111 ) );
  MUX \b/U3140  ( .IN0(\b/n758 ), .IN1(\b/n3109 ), .SEL(msg[42]), .F(\b/n3110 ) );
  MUX \b/U3139  ( .IN0(\b/n733 ), .IN1(\b/n775 ), .SEL(msg[41]), .F(\b/n3109 )
         );
  MUX \b/U3138  ( .IN0(\b/n3107 ), .IN1(\b/n3098 ), .SEL(msg[40]), .F(
        \b/n3108 ) );
  MUX \b/U3137  ( .IN0(\b/n3106 ), .IN1(\b/n3102 ), .SEL(msg[45]), .F(
        \b/n3107 ) );
  MUX \b/U3136  ( .IN0(\b/n3104 ), .IN1(\b/n3103 ), .SEL(msg[47]), .F(
        \b/n3106 ) );
  NAND \b/U3135  ( .A(\b/n723 ), .B(\b/n3105 ), .Z(\b/n3104 ) );
  MUX \b/U3134  ( .IN0(\b/n774 ), .IN1(\b/n736 ), .SEL(msg[42]), .F(\b/n3103 )
         );
  MUX \b/U3133  ( .IN0(\b/n3101 ), .IN1(\b/n3099 ), .SEL(msg[47]), .F(
        \b/n3102 ) );
  MUX \b/U3132  ( .IN0(\b/n2942 ), .IN1(\b/n3100 ), .SEL(msg[42]), .F(
        \b/n3101 ) );
  AND \b/U3131  ( .A(msg[41]), .B(\b/n723 ), .Z(\b/n3100 ) );
  MUX \b/U3130  ( .IN0(\b/n728 ), .IN1(\b/n2961 ), .SEL(msg[42]), .F(\b/n3099 ) );
  MUX \b/U3129  ( .IN0(\b/n3097 ), .IN1(\b/n3091 ), .SEL(msg[45]), .F(
        \b/n3098 ) );
  MUX \b/U3128  ( .IN0(\b/n3096 ), .IN1(\b/n3094 ), .SEL(msg[47]), .F(
        \b/n3097 ) );
  MUX \b/U3127  ( .IN0(\b/n3095 ), .IN1(\b/n2931 ), .SEL(\b/n2979 ), .F(
        \b/n3096 ) );
  MUX \b/U3126  ( .IN0(msg[43]), .IN1(msg[44]), .SEL(msg[42]), .F(\b/n3095 )
         );
  MUX \b/U3125  ( .IN0(\b/n2961 ), .IN1(\b/n3092 ), .SEL(msg[42]), .F(
        \b/n3094 ) );
  NAND \b/U3124  ( .A(\b/n2931 ), .B(\b/n3093 ), .Z(\b/n3092 ) );
  MUX \b/U3123  ( .IN0(\b/n3088 ), .IN1(\b/n3089 ), .SEL(msg[47]), .F(
        \b/n3091 ) );
  AND \b/U3122  ( .A(\b/n756 ), .B(\b/n3090 ), .Z(\b/n3089 ) );
  MUX \b/U3121  ( .IN0(\b/n737 ), .IN1(\b/n2932 ), .SEL(msg[42]), .F(\b/n3088 ) );
  MUX \b/U3120  ( .IN0(\b/n3087 ), .IN1(\b/n3071 ), .SEL(msg[46]), .F(
        shift_row_out[10]) );
  MUX \b/U3119  ( .IN0(\b/n3086 ), .IN1(\b/n3078 ), .SEL(msg[40]), .F(
        \b/n3087 ) );
  MUX \b/U3118  ( .IN0(\b/n3085 ), .IN1(\b/n3081 ), .SEL(msg[45]), .F(
        \b/n3086 ) );
  MUX \b/U3117  ( .IN0(\b/n3084 ), .IN1(\b/n3082 ), .SEL(msg[42]), .F(
        \b/n3085 ) );
  MUX \b/U3116  ( .IN0(\b/n745 ), .IN1(\b/n3083 ), .SEL(msg[47]), .F(\b/n3084 ) );
  MUX \b/U3115  ( .IN0(\b/n2939 ), .IN1(\b/n723 ), .SEL(msg[41]), .F(\b/n3083 ) );
  MUX \b/U3114  ( .IN0(\b/n2978 ), .IN1(\b/n763 ), .SEL(msg[47]), .F(\b/n3082 ) );
  MUX \b/U3113  ( .IN0(\b/n3080 ), .IN1(\b/n3079 ), .SEL(msg[42]), .F(
        \b/n3081 ) );
  MUX \b/U3112  ( .IN0(\b/n2932 ), .IN1(\b/n730 ), .SEL(msg[47]), .F(\b/n3080 ) );
  MUX \b/U3111  ( .IN0(\b/n766 ), .IN1(\b/n2965 ), .SEL(msg[47]), .F(\b/n3079 ) );
  MUX \b/U3110  ( .IN0(\b/n3077 ), .IN1(\b/n3073 ), .SEL(msg[45]), .F(
        \b/n3078 ) );
  MUX \b/U3109  ( .IN0(\b/n3074 ), .IN1(\b/n712 ), .SEL(msg[42]), .F(\b/n3077 ) );
  NAND \b/U3108  ( .A(\b/n3075 ), .B(\b/n3076 ), .Z(\b/n3074 ) );
  MUX \b/U3107  ( .IN0(n643), .IN1(\b/n3072 ), .SEL(\b/n2977 ), .F(\b/n3073 )
         );
  MUX \b/U3106  ( .IN0(\b/n744 ), .IN1(\b/n2944 ), .SEL(msg[42]), .F(\b/n3072 ) );
  MUX \b/U3105  ( .IN0(\b/n3070 ), .IN1(\b/n3062 ), .SEL(msg[40]), .F(
        \b/n3071 ) );
  MUX \b/U3104  ( .IN0(\b/n3069 ), .IN1(\b/n3066 ), .SEL(msg[45]), .F(
        \b/n3070 ) );
  MUX \b/U3103  ( .IN0(\b/n3068 ), .IN1(\b/n3067 ), .SEL(msg[42]), .F(
        \b/n3069 ) );
  MUX \b/U3102  ( .IN0(\b/n772 ), .IN1(msg[41]), .SEL(msg[47]), .F(\b/n3068 )
         );
  MUX \b/U3101  ( .IN0(n646), .IN1(\b/n2945 ), .SEL(msg[47]), .F(\b/n3067 ) );
  MUX \b/U3100  ( .IN0(\b/n3065 ), .IN1(\b/n3064 ), .SEL(msg[42]), .F(
        \b/n3066 ) );
  MUX \b/U3099  ( .IN0(\b/n777 ), .IN1(\b/n771 ), .SEL(msg[47]), .F(\b/n3065 )
         );
  MUX \b/U3098  ( .IN0(n646), .IN1(\b/n3063 ), .SEL(msg[47]), .F(\b/n3064 ) );
  MUX \b/U3097  ( .IN0(\b/n723 ), .IN1(\b/n760 ), .SEL(msg[41]), .F(\b/n3063 )
         );
  MUX \b/U3096  ( .IN0(\b/n3061 ), .IN1(\b/n3055 ), .SEL(msg[45]), .F(
        \b/n3062 ) );
  MUX \b/U3095  ( .IN0(\b/n3058 ), .IN1(\b/n3057 ), .SEL(msg[42]), .F(
        \b/n3061 ) );
  NAND \b/U3094  ( .A(\b/n3059 ), .B(\b/n3060 ), .Z(\b/n3058 ) );
  MUX \b/U3093  ( .IN0(\b/n2931 ), .IN1(\b/n3056 ), .SEL(n644), .F(\b/n3057 )
         );
  MUX \b/U3092  ( .IN0(msg[43]), .IN1(\b/n733 ), .SEL(msg[47]), .F(\b/n3056 )
         );
  MUX \b/U3091  ( .IN0(\b/n3054 ), .IN1(\b/n3053 ), .SEL(msg[42]), .F(
        \b/n3055 ) );
  MUX \b/U3090  ( .IN0(\b/n2976 ), .IN1(\b/n731 ), .SEL(msg[47]), .F(\b/n3054 ) );
  MUX \b/U3089  ( .IN0(\b/n2972 ), .IN1(\b/n3052 ), .SEL(msg[47]), .F(
        \b/n3053 ) );
  MUX \b/U3088  ( .IN0(\b/n2934 ), .IN1(\b/n2939 ), .SEL(msg[41]), .F(
        \b/n3052 ) );
  MUX \b/U3087  ( .IN0(\b/n3051 ), .IN1(\b/n3033 ), .SEL(msg[46]), .F(
        shift_row_out[9]) );
  MUX \b/U3086  ( .IN0(\b/n3050 ), .IN1(\b/n3041 ), .SEL(msg[40]), .F(
        \b/n3051 ) );
  MUX \b/U3085  ( .IN0(\b/n3049 ), .IN1(\b/n3045 ), .SEL(msg[45]), .F(
        \b/n3050 ) );
  MUX \b/U3084  ( .IN0(\b/n3048 ), .IN1(\b/n3047 ), .SEL(msg[42]), .F(
        \b/n3049 ) );
  MUX \b/U3083  ( .IN0(\b/n768 ), .IN1(n648), .SEL(msg[47]), .F(\b/n3048 ) );
  MUX \b/U3082  ( .IN0(\b/n3046 ), .IN1(n642), .SEL(msg[47]), .F(\b/n3047 ) );
  NAND \b/U3081  ( .A(\b/n780 ), .B(\b/n739 ), .Z(\b/n3046 ) );
  MUX \b/U3080  ( .IN0(\b/n3044 ), .IN1(\b/n3043 ), .SEL(msg[42]), .F(
        \b/n3045 ) );
  MUX \b/U3079  ( .IN0(\b/n716 ), .IN1(\b/n2946 ), .SEL(msg[47]), .F(\b/n3044 ) );
  MUX \b/U3078  ( .IN0(\b/n2936 ), .IN1(\b/n3042 ), .SEL(msg[47]), .F(
        \b/n3043 ) );
  AND \b/U3077  ( .A(msg[41]), .B(msg[44]), .Z(\b/n3042 ) );
  MUX \b/U3076  ( .IN0(\b/n3040 ), .IN1(\b/n3037 ), .SEL(msg[45]), .F(
        \b/n3041 ) );
  MUX \b/U3075  ( .IN0(\b/n3039 ), .IN1(\b/n3038 ), .SEL(msg[42]), .F(
        \b/n3040 ) );
  MUX \b/U3074  ( .IN0(\b/n2975 ), .IN1(\b/n777 ), .SEL(msg[47]), .F(\b/n3039 ) );
  MUX \b/U3073  ( .IN0(\b/n752 ), .IN1(\b/n2944 ), .SEL(msg[47]), .F(\b/n3038 ) );
  MUX \b/U3072  ( .IN0(\b/n3034 ), .IN1(\b/n3035 ), .SEL(msg[42]), .F(
        \b/n3037 ) );
  AND \b/U3071  ( .A(\b/n3036 ), .B(\b/n2991 ), .Z(\b/n3035 ) );
  MUX \b/U3070  ( .IN0(\b/n2950 ), .IN1(\b/n2939 ), .SEL(msg[47]), .F(
        \b/n3034 ) );
  MUX \b/U3069  ( .IN0(\b/n3032 ), .IN1(\b/n3024 ), .SEL(msg[40]), .F(
        \b/n3033 ) );
  MUX \b/U3068  ( .IN0(\b/n3031 ), .IN1(\b/n3027 ), .SEL(msg[45]), .F(
        \b/n3032 ) );
  MUX \b/U3067  ( .IN0(\b/n3030 ), .IN1(\b/n3029 ), .SEL(msg[42]), .F(
        \b/n3031 ) );
  MUX \b/U3066  ( .IN0(\b/n2938 ), .IN1(\b/n741 ), .SEL(msg[47]), .F(\b/n3030 ) );
  MUX \b/U3065  ( .IN0(\b/n3028 ), .IN1(\b/n725 ), .SEL(msg[47]), .F(\b/n3029 ) );
  MUX \b/U3064  ( .IN0(\b/n2936 ), .IN1(\b/n733 ), .SEL(msg[41]), .F(\b/n3028 ) );
  MUX \b/U3063  ( .IN0(\b/n3026 ), .IN1(\b/n3025 ), .SEL(msg[42]), .F(
        \b/n3027 ) );
  MUX \b/U3062  ( .IN0(\b/n772 ), .IN1(\b/n750 ), .SEL(msg[47]), .F(\b/n3026 )
         );
  MUX \b/U3061  ( .IN0(\b/n768 ), .IN1(\b/n728 ), .SEL(msg[47]), .F(\b/n3025 )
         );
  MUX \b/U3060  ( .IN0(\b/n3023 ), .IN1(\b/n3018 ), .SEL(msg[45]), .F(
        \b/n3024 ) );
  MUX \b/U3059  ( .IN0(\b/n3022 ), .IN1(\b/n3019 ), .SEL(msg[42]), .F(
        \b/n3023 ) );
  MUX \b/U3058  ( .IN0(\b/n3020 ), .IN1(\b/n3021 ), .SEL(msg[47]), .F(
        \b/n3022 ) );
  NAND \b/U3057  ( .A(\b/n2939 ), .B(\b/n3011 ), .Z(\b/n3021 ) );
  MUX \b/U3056  ( .IN0(\b/n2939 ), .IN1(\b/n733 ), .SEL(msg[41]), .F(\b/n3020 ) );
  MUX \b/U3055  ( .IN0(\b/n2956 ), .IN1(\b/n2954 ), .SEL(msg[47]), .F(
        \b/n3019 ) );
  MUX \b/U3054  ( .IN0(\b/n2974 ), .IN1(\b/n3017 ), .SEL(msg[42]), .F(
        \b/n3018 ) );
  MUX \b/U3053  ( .IN0(\b/n739 ), .IN1(\b/n771 ), .SEL(msg[47]), .F(\b/n3017 )
         );
  MUX \b/U3052  ( .IN0(\b/n3016 ), .IN1(\b/n2999 ), .SEL(msg[46]), .F(
        shift_row_out[8]) );
  MUX \b/U3051  ( .IN0(\b/n3015 ), .IN1(\b/n3007 ), .SEL(msg[40]), .F(
        \b/n3016 ) );
  MUX \b/U3050  ( .IN0(\b/n3014 ), .IN1(\b/n3012 ), .SEL(msg[42]), .F(
        \b/n3015 ) );
  MUX \b/U3049  ( .IN0(\b/n713 ), .IN1(\b/n3013 ), .SEL(msg[47]), .F(\b/n3014 ) );
  MUX \b/U3048  ( .IN0(\b/n766 ), .IN1(\b/n769 ), .SEL(msg[45]), .F(\b/n3013 )
         );
  MUX \b/U3047  ( .IN0(\b/n3009 ), .IN1(\b/n3008 ), .SEL(msg[47]), .F(
        \b/n3012 ) );
  NAND \b/U3046  ( .A(\b/n3010 ), .B(\b/n3011 ), .Z(\b/n3009 ) );
  MUX \b/U3045  ( .IN0(\b/n765 ), .IN1(\b/n780 ), .SEL(msg[45]), .F(\b/n3008 )
         );
  MUX \b/U3044  ( .IN0(\b/n3006 ), .IN1(\b/n3002 ), .SEL(msg[42]), .F(
        \b/n3007 ) );
  MUX \b/U3043  ( .IN0(\b/n3005 ), .IN1(\b/n3003 ), .SEL(msg[47]), .F(
        \b/n3006 ) );
  MUX \b/U3042  ( .IN0(\b/n3004 ), .IN1(\b/n718 ), .SEL(msg[45]), .F(\b/n3005 ) );
  NAND \b/U3041  ( .A(\b/n780 ), .B(\b/n2931 ), .Z(\b/n3004 ) );
  MUX \b/U3039  ( .IN0(\b/n3001 ), .IN1(\b/n3000 ), .SEL(msg[47]), .F(
        \b/n3002 ) );
  MUX \b/U3038  ( .IN0(n643), .IN1(\b/n715 ), .SEL(msg[45]), .F(\b/n3001 ) );
  MUX \b/U3037  ( .IN0(\b/n767 ), .IN1(\b/n723 ), .SEL(msg[45]), .F(\b/n3000 )
         );
  MUX \b/U3036  ( .IN0(\b/n2998 ), .IN1(\b/n2988 ), .SEL(msg[40]), .F(
        \b/n2999 ) );
  MUX \b/U3035  ( .IN0(\b/n2997 ), .IN1(\b/n2993 ), .SEL(msg[42]), .F(
        \b/n2998 ) );
  MUX \b/U3034  ( .IN0(\b/n2996 ), .IN1(\b/n2995 ), .SEL(msg[47]), .F(
        \b/n2997 ) );
  MUX \b/U3033  ( .IN0(n641), .IN1(\b/n719 ), .SEL(msg[45]), .F(\b/n2996 ) );
  MUX \b/U3032  ( .IN0(\b/n2994 ), .IN1(\b/n756 ), .SEL(msg[45]), .F(\b/n2995 ) );
  NAND \b/U3031  ( .A(\b/n2930 ), .B(\b/n2932 ), .Z(\b/n2994 ) );
  MUX \b/U3030  ( .IN0(\b/n2992 ), .IN1(\b/n2989 ), .SEL(msg[47]), .F(
        \b/n2993 ) );
  MUX \b/U3029  ( .IN0(\b/n726 ), .IN1(\b/n2990 ), .SEL(msg[45]), .F(\b/n2992 ) );
  NAND \b/U3028  ( .A(\b/n2934 ), .B(\b/n2991 ), .Z(\b/n2990 ) );
  MUX \b/U3027  ( .IN0(\b/n2949 ), .IN1(\b/n2940 ), .SEL(msg[45]), .F(
        \b/n2989 ) );
  MUX \b/U3026  ( .IN0(\b/n2987 ), .IN1(\b/n2983 ), .SEL(msg[42]), .F(
        \b/n2988 ) );
  MUX \b/U3025  ( .IN0(\b/n2985 ), .IN1(\b/n2984 ), .SEL(msg[47]), .F(
        \b/n2987 ) );
  NAND \b/U3024  ( .A(\b/n2986 ), .B(\b/n2973 ), .Z(\b/n2985 ) );
  MUX \b/U3023  ( .IN0(msg[43]), .IN1(\b/n2965 ), .SEL(msg[45]), .F(\b/n2984 )
         );
  MUX \b/U3022  ( .IN0(\b/n2982 ), .IN1(\b/n2981 ), .SEL(msg[47]), .F(
        \b/n2983 ) );
  MUX \b/U3021  ( .IN0(\b/n731 ), .IN1(\b/n747 ), .SEL(msg[45]), .F(\b/n2982 )
         );
  MUX \b/U3020  ( .IN0(\b/n764 ), .IN1(\b/n752 ), .SEL(msg[45]), .F(\b/n2981 )
         );
  XOR \b/U3019  ( .A(\b/n2931 ), .B(msg[41]), .Z(\b/n2980 ) );
  XOR \b/U3018  ( .A(msg[41]), .B(msg[42]), .Z(\b/n2979 ) );
  XOR \b/U3017  ( .A(msg[41]), .B(msg[43]), .Z(\b/n2978 ) );
  XOR \b/U3016  ( .A(msg[42]), .B(msg[47]), .Z(\b/n2977 ) );
  XOR \b/U3015  ( .A(\b/n780 ), .B(\b/n723 ), .Z(\b/n2976 ) );
  XOR \b/U3014  ( .A(msg[41]), .B(\b/n769 ), .Z(\b/n2975 ) );
  XOR \b/U3012  ( .A(msg[41]), .B(msg[45]), .Z(\b/n2973 ) );
  NAND \b/U3011  ( .A(msg[41]), .B(msg[43]), .Z(\b/n2972 ) );
  MUX \b/U3010  ( .IN0(\b/n2931 ), .IN1(\b/n723 ), .SEL(msg[41]), .F(\b/n2971 ) );
  MUX \b/U3008  ( .IN0(msg[43]), .IN1(\b/n760 ), .SEL(msg[41]), .F(\b/n2969 )
         );
  MUX \b/U3007  ( .IN0(\b/n739 ), .IN1(\b/n760 ), .SEL(msg[41]), .F(\b/n2968 )
         );
  MUX \b/U3006  ( .IN0(\b/n2934 ), .IN1(\b/n2936 ), .SEL(msg[41]), .F(
        \b/n2967 ) );
  MUX \b/U3005  ( .IN0(msg[44]), .IN1(\b/n739 ), .SEL(msg[41]), .F(\b/n2966 )
         );
  OR \b/U3004  ( .A(msg[41]), .B(msg[44]), .Z(\b/n2965 ) );
  NAND \b/U3002  ( .A(\b/n760 ), .B(\b/n780 ), .Z(\b/n2963 ) );
  MUX \b/U3001  ( .IN0(\b/n760 ), .IN1(msg[44]), .SEL(msg[41]), .F(\b/n2962 )
         );
  MUX \b/U3000  ( .IN0(\b/n2930 ), .IN1(\b/n2939 ), .SEL(msg[41]), .F(
        \b/n2961 ) );
  MUX \b/U2999  ( .IN0(\b/n775 ), .IN1(msg[44]), .SEL(msg[41]), .F(\b/n2960 )
         );
  MUX \b/U2998  ( .IN0(\b/n733 ), .IN1(\b/n760 ), .SEL(msg[41]), .F(\b/n2959 )
         );
  MUX \b/U2997  ( .IN0(\b/n2930 ), .IN1(msg[44]), .SEL(msg[41]), .F(\b/n2958 )
         );
  MUX \b/U2996  ( .IN0(\b/n750 ), .IN1(\b/n739 ), .SEL(msg[41]), .F(\b/n2957 )
         );
  XOR \b/U2995  ( .A(\b/n733 ), .B(msg[41]), .Z(\b/n2956 ) );
  MUX \b/U2994  ( .IN0(\b/n2936 ), .IN1(\b/n750 ), .SEL(msg[41]), .F(\b/n2955 ) );
  NANDN \b/U2993  ( .B(msg[41]), .A(msg[43]), .Z(\b/n2954 ) );
  MUX \b/U2992  ( .IN0(\b/n723 ), .IN1(msg[43]), .SEL(msg[41]), .F(\b/n2953 )
         );
  NAND \b/U2990  ( .A(\b/n2934 ), .B(\b/n780 ), .Z(\b/n2951 ) );
  MUX \b/U2989  ( .IN0(msg[44]), .IN1(\b/n2931 ), .SEL(msg[41]), .F(\b/n2950 )
         );
  MUX \b/U2988  ( .IN0(\b/n750 ), .IN1(msg[43]), .SEL(msg[41]), .F(\b/n2949 )
         );
  MUX \b/U2986  ( .IN0(msg[44]), .IN1(\b/n769 ), .SEL(msg[41]), .F(\b/n2947 )
         );
  MUX \b/U2985  ( .IN0(\b/n723 ), .IN1(\b/n775 ), .SEL(msg[41]), .F(\b/n2946 )
         );
  NAND \b/U2984  ( .A(\b/n2932 ), .B(\b/n723 ), .Z(\b/n2945 ) );
  MUX \b/U2983  ( .IN0(\b/n2931 ), .IN1(\b/n2939 ), .SEL(msg[41]), .F(
        \b/n2944 ) );
  NAND \b/U2982  ( .A(\b/n2943 ), .B(\b/n2930 ), .Z(\b/n2942 ) );
  MUX \b/U2981  ( .IN0(\b/n2934 ), .IN1(\b/n775 ), .SEL(msg[41]), .F(\b/n2941 ) );
  MUX \b/U2980  ( .IN0(\b/n775 ), .IN1(\b/n739 ), .SEL(msg[41]), .F(\b/n2940 )
         );
  NANDN \b/U2979  ( .B(msg[43]), .A(msg[44]), .Z(\b/n2939 ) );
  MUX \b/U2978  ( .IN0(\b/n2934 ), .IN1(msg[43]), .SEL(msg[41]), .F(\b/n2938 )
         );
  OR \b/U2977  ( .A(msg[43]), .B(msg[44]), .Z(\b/n2934 ) );
  MUX \b/U2976  ( .IN0(\b/n723 ), .IN1(\b/n739 ), .SEL(msg[41]), .F(\b/n2937 )
         );
  XOR \b/U2975  ( .A(\b/n733 ), .B(msg[43]), .Z(\b/n2936 ) );
  NANDN \b/U2974  ( .B(msg[43]), .A(msg[41]), .Z(\b/n2935 ) );
  NAND \b/U2973  ( .A(\b/n2934 ), .B(\b/n2932 ), .Z(\b/n2933 ) );
  NAND \b/U2972  ( .A(msg[41]), .B(\b/n2931 ), .Z(\b/n2932 ) );
  NANDN \b/U2971  ( .B(msg[44]), .A(msg[43]), .Z(\b/n2931 ) );
  NAND \b/U2970  ( .A(msg[43]), .B(msg[44]), .Z(\b/n2930 ) );
  MUX \b/U2969  ( .IN0(msg[36]), .IN1(\b/n2571 ), .SEL(msg[33]), .F(\b/n2929 )
         );
  MUX \b/U2968  ( .IN0(msg[36]), .IN1(\b/n2580 ), .SEL(msg[33]), .F(\b/n2928 )
         );
  MUX \b/U2967  ( .IN0(\b/n2572 ), .IN1(\b/n2575 ), .SEL(msg[33]), .F(
        \b/n2927 ) );
  MUX \b/U2966  ( .IN0(\b/n2577 ), .IN1(\b/n840 ), .SEL(msg[33]), .F(\b/n2926 ) );
  MUX \b/U2964  ( .IN0(\b/n2580 ), .IN1(\b/n2571 ), .SEL(msg[34]), .F(
        \b/n2753 ) );
  MUX \b/U2963  ( .IN0(\b/n2573 ), .IN1(\b/n851 ), .SEL(msg[34]), .F(\b/n2754 ) );
  MUX \b/U2962  ( .IN0(\b/n794 ), .IN1(\b/n804 ), .SEL(msg[33]), .F(\b/n2717 )
         );
  MUX \b/U2961  ( .IN0(\b/n2601 ), .IN1(\b/n2912 ), .SEL(msg[39]), .F(
        \b/n2924 ) );
  MUX \b/U2960  ( .IN0(\b/n2575 ), .IN1(\b/n2571 ), .SEL(msg[33]), .F(
        \b/n2915 ) );
  MUX \b/U2959  ( .IN0(\b/n846 ), .IN1(\b/n2577 ), .SEL(msg[33]), .F(\b/n2923 ) );
  MUX \b/U2958  ( .IN0(msg[35]), .IN1(\b/n840 ), .SEL(msg[33]), .F(\b/n2922 )
         );
  MUX \b/U2957  ( .IN0(\b/n2580 ), .IN1(\b/n846 ), .SEL(msg[33]), .F(\b/n2921 ) );
  MUX \b/U2956  ( .IN0(msg[36]), .IN1(\b/n2577 ), .SEL(msg[33]), .F(\b/n2920 )
         );
  MUX \b/U2955  ( .IN0(\b/n831 ), .IN1(\b/n810 ), .SEL(msg[37]), .F(\b/n2627 )
         );
  MUX \b/U2954  ( .IN0(\b/n2572 ), .IN1(\b/n804 ), .SEL(msg[33]), .F(\b/n2919 ) );
  NANDN \b/U2951  ( .B(\b/n2578 ), .A(msg[39]), .Z(\b/n2892 ) );
  NAND \b/U2950  ( .A(msg[39]), .B(\b/n807 ), .Z(\b/n2860 ) );
  NAND \b/U2949  ( .A(msg[39]), .B(\b/n819 ), .Z(\b/n2801 ) );
  NAND \b/U2948  ( .A(msg[39]), .B(\b/n2909 ), .Z(\b/n2834 ) );
  NAND \b/U2947  ( .A(msg[39]), .B(\b/n2829 ), .Z(\b/n2792 ) );
  NAND \b/U2945  ( .A(\b/n851 ), .B(\b/n840 ), .Z(\b/n2913 ) );
  NAND \b/U2944  ( .A(msg[39]), .B(\b/n2911 ), .Z(\b/n2906 ) );
  NAND \b/U2943  ( .A(n640), .B(msg[39]), .Z(\b/n2886 ) );
  NAND \b/U2941  ( .A(msg[34]), .B(\b/n2580 ), .Z(\b/n2746 ) );
  NAND \b/U2940  ( .A(\b/n840 ), .B(msg[33]), .Z(\b/n2701 ) );
  NAND \b/U2939  ( .A(msg[39]), .B(\b/n2915 ), .Z(\b/n2700 ) );
  NAND \b/U2937  ( .A(\b/n2913 ), .B(msg[39]), .Z(\b/n2716 ) );
  NAND \b/U2936  ( .A(\b/n2734 ), .B(\b/n2580 ), .Z(\b/n2912 ) );
  NANDN \b/U2935  ( .B(\b/n794 ), .A(\b/n851 ), .Z(\b/n2911 ) );
  NAND \b/U2933  ( .A(msg[33]), .B(\b/n2580 ), .Z(\b/n2632 ) );
  NAND \b/U2932  ( .A(\b/n794 ), .B(\b/n851 ), .Z(\b/n2909 ) );
  NAND \b/U2929  ( .A(msg[33]), .B(\b/n2575 ), .Z(\b/n2734 ) );
  ANDN \b/U2927  ( .A(msg[34]), .B(msg[33]), .Z(\b/n2762 ) );
  AND \b/U2926  ( .A(\b/n2572 ), .B(\b/n2906 ), .Z(\b/n2677 ) );
  MUX \b/U2925  ( .IN0(\b/n2905 ), .IN1(\b/n2889 ), .SEL(msg[38]), .F(
        shift_row_out[39]) );
  MUX \b/U2924  ( .IN0(\b/n2904 ), .IN1(\b/n2897 ), .SEL(msg[32]), .F(
        \b/n2905 ) );
  MUX \b/U2923  ( .IN0(\b/n2903 ), .IN1(\b/n2900 ), .SEL(msg[37]), .F(
        \b/n2904 ) );
  MUX \b/U2922  ( .IN0(\b/n2902 ), .IN1(\b/n2901 ), .SEL(msg[34]), .F(
        \b/n2903 ) );
  MUX \b/U2921  ( .IN0(msg[36]), .IN1(\b/n811 ), .SEL(msg[39]), .F(\b/n2902 )
         );
  MUX \b/U2920  ( .IN0(\b/n2573 ), .IN1(\b/n815 ), .SEL(msg[39]), .F(\b/n2901 ) );
  MUX \b/U2919  ( .IN0(\b/n2899 ), .IN1(\b/n2898 ), .SEL(msg[34]), .F(
        \b/n2900 ) );
  MUX \b/U2918  ( .IN0(\b/n2631 ), .IN1(\b/n807 ), .SEL(msg[39]), .F(\b/n2899 ) );
  MUX \b/U2917  ( .IN0(\b/n2583 ), .IN1(\b/n2594 ), .SEL(msg[39]), .F(
        \b/n2898 ) );
  MUX \b/U2916  ( .IN0(\b/n2896 ), .IN1(\b/n2893 ), .SEL(msg[37]), .F(
        \b/n2897 ) );
  MUX \b/U2915  ( .IN0(\b/n2895 ), .IN1(\b/n2894 ), .SEL(msg[34]), .F(
        \b/n2896 ) );
  MUX \b/U2914  ( .IN0(\b/n2607 ), .IN1(\b/n2582 ), .SEL(msg[39]), .F(
        \b/n2895 ) );
  MUX \b/U2913  ( .IN0(\b/n819 ), .IN1(\b/n2603 ), .SEL(msg[39]), .F(\b/n2894 ) );
  MUX \b/U2912  ( .IN0(\b/n2891 ), .IN1(\b/n2890 ), .SEL(msg[34]), .F(
        \b/n2893 ) );
  AND \b/U2911  ( .A(\b/n809 ), .B(\b/n2892 ), .Z(\b/n2891 ) );
  MUX \b/U2910  ( .IN0(\b/n2587 ), .IN1(n639), .SEL(msg[39]), .F(\b/n2890 ) );
  MUX \b/U2909  ( .IN0(\b/n2888 ), .IN1(\b/n2880 ), .SEL(msg[32]), .F(
        \b/n2889 ) );
  MUX \b/U2908  ( .IN0(\b/n2887 ), .IN1(\b/n2883 ), .SEL(msg[37]), .F(
        \b/n2888 ) );
  MUX \b/U2907  ( .IN0(\b/n2884 ), .IN1(\b/n2885 ), .SEL(msg[34]), .F(
        \b/n2887 ) );
  NAND \b/U2906  ( .A(\b/n2701 ), .B(\b/n2886 ), .Z(\b/n2885 ) );
  MUX \b/U2905  ( .IN0(\b/n849 ), .IN1(\b/n841 ), .SEL(msg[39]), .F(\b/n2884 )
         );
  MUX \b/U2904  ( .IN0(\b/n2882 ), .IN1(\b/n2881 ), .SEL(msg[34]), .F(
        \b/n2883 ) );
  MUX \b/U2903  ( .IN0(\b/n2577 ), .IN1(\b/n2571 ), .SEL(msg[39]), .F(
        \b/n2882 ) );
  MUX \b/U2902  ( .IN0(\b/n842 ), .IN1(\b/n2608 ), .SEL(msg[39]), .F(\b/n2881 ) );
  MUX \b/U2901  ( .IN0(\b/n2879 ), .IN1(\b/n2876 ), .SEL(msg[37]), .F(
        \b/n2880 ) );
  MUX \b/U2900  ( .IN0(\b/n2878 ), .IN1(\b/n2877 ), .SEL(msg[34]), .F(
        \b/n2879 ) );
  MUX \b/U2899  ( .IN0(\b/n2612 ), .IN1(\b/n2598 ), .SEL(msg[39]), .F(
        \b/n2878 ) );
  MUX \b/U2898  ( .IN0(\b/n795 ), .IN1(\b/n2580 ), .SEL(msg[39]), .F(\b/n2877 ) );
  MUX \b/U2897  ( .IN0(\b/n2875 ), .IN1(\b/n2874 ), .SEL(msg[34]), .F(
        \b/n2876 ) );
  MUX \b/U2896  ( .IN0(\b/n2613 ), .IN1(\b/n2621 ), .SEL(msg[39]), .F(
        \b/n2875 ) );
  MUX \b/U2895  ( .IN0(\b/n2606 ), .IN1(\b/n2873 ), .SEL(msg[39]), .F(
        \b/n2874 ) );
  MUX \b/U2894  ( .IN0(\b/n846 ), .IN1(\b/n804 ), .SEL(msg[33]), .F(\b/n2873 )
         );
  MUX \b/U2893  ( .IN0(\b/n2872 ), .IN1(\b/n2854 ), .SEL(msg[38]), .F(
        shift_row_out[38]) );
  MUX \b/U2892  ( .IN0(\b/n2871 ), .IN1(\b/n2862 ), .SEL(msg[32]), .F(
        \b/n2872 ) );
  MUX \b/U2891  ( .IN0(\b/n2870 ), .IN1(\b/n2865 ), .SEL(msg[37]), .F(
        \b/n2871 ) );
  MUX \b/U2890  ( .IN0(\b/n2869 ), .IN1(\b/n2867 ), .SEL(msg[34]), .F(
        \b/n2870 ) );
  MUX \b/U2889  ( .IN0(\b/n2868 ), .IN1(\b/n2584 ), .SEL(msg[39]), .F(
        \b/n2869 ) );
  MUX \b/U2888  ( .IN0(\b/n846 ), .IN1(\b/n2571 ), .SEL(msg[33]), .F(\b/n2868 ) );
  MUX \b/U2887  ( .IN0(\b/n2866 ), .IN1(\b/n834 ), .SEL(msg[39]), .F(\b/n2867 ) );
  MUX \b/U2886  ( .IN0(\b/n2571 ), .IN1(\b/n2572 ), .SEL(msg[33]), .F(
        \b/n2866 ) );
  MUX \b/U2885  ( .IN0(\b/n2864 ), .IN1(\b/n2863 ), .SEL(msg[34]), .F(
        \b/n2865 ) );
  MUX \b/U2884  ( .IN0(n638), .IN1(\b/n2652 ), .SEL(msg[39]), .F(\b/n2864 ) );
  MUX \b/U2883  ( .IN0(\b/n2610 ), .IN1(\b/n2617 ), .SEL(msg[39]), .F(
        \b/n2863 ) );
  MUX \b/U2882  ( .IN0(\b/n2861 ), .IN1(\b/n2857 ), .SEL(msg[37]), .F(
        \b/n2862 ) );
  MUX \b/U2881  ( .IN0(\b/n2859 ), .IN1(\b/n2858 ), .SEL(msg[34]), .F(
        \b/n2861 ) );
  AND \b/U2880  ( .A(\b/n787 ), .B(\b/n2860 ), .Z(\b/n2859 ) );
  MUX \b/U2879  ( .IN0(\b/n2687 ), .IN1(msg[35]), .SEL(msg[39]), .F(\b/n2858 )
         );
  MUX \b/U2878  ( .IN0(\b/n2856 ), .IN1(\b/n2855 ), .SEL(msg[34]), .F(
        \b/n2857 ) );
  MUX \b/U2877  ( .IN0(\b/n830 ), .IN1(\b/n2575 ), .SEL(msg[39]), .F(\b/n2856 ) );
  MUX \b/U2875  ( .IN0(\b/n2853 ), .IN1(\b/n2846 ), .SEL(msg[32]), .F(
        \b/n2854 ) );
  MUX \b/U2874  ( .IN0(\b/n2852 ), .IN1(\b/n2849 ), .SEL(msg[37]), .F(
        \b/n2853 ) );
  MUX \b/U2873  ( .IN0(\b/n2851 ), .IN1(\b/n2850 ), .SEL(msg[34]), .F(
        \b/n2852 ) );
  MUX \b/U2872  ( .IN0(\b/n826 ), .IN1(\b/n2579 ), .SEL(msg[39]), .F(\b/n2851 ) );
  MUX \b/U2871  ( .IN0(\b/n2583 ), .IN1(n639), .SEL(msg[39]), .F(\b/n2850 ) );
  MUX \b/U2870  ( .IN0(\b/n2848 ), .IN1(\b/n2847 ), .SEL(msg[34]), .F(
        \b/n2849 ) );
  MUX \b/U2869  ( .IN0(\b/n2599 ), .IN1(\b/n791 ), .SEL(msg[39]), .F(\b/n2848 ) );
  MUX \b/U2868  ( .IN0(\b/n811 ), .IN1(\b/n841 ), .SEL(msg[39]), .F(\b/n2847 )
         );
  MUX \b/U2867  ( .IN0(\b/n2845 ), .IN1(\b/n2841 ), .SEL(msg[37]), .F(
        \b/n2846 ) );
  MUX \b/U2866  ( .IN0(\b/n2844 ), .IN1(\b/n2843 ), .SEL(msg[34]), .F(
        \b/n2845 ) );
  MUX \b/U2865  ( .IN0(\b/n2588 ), .IN1(\b/n841 ), .SEL(msg[39]), .F(\b/n2844 ) );
  MUX \b/U2864  ( .IN0(\b/n2842 ), .IN1(\b/n2609 ), .SEL(msg[39]), .F(
        \b/n2843 ) );
  NANDN \b/U2863  ( .B(msg[36]), .A(msg[33]), .Z(\b/n2842 ) );
  MUX \b/U2862  ( .IN0(\b/n2840 ), .IN1(\b/n2838 ), .SEL(msg[34]), .F(
        \b/n2841 ) );
  MUX \b/U2861  ( .IN0(\b/n804 ), .IN1(\b/n2839 ), .SEL(msg[39]), .F(\b/n2840 ) );
  MUX \b/U2860  ( .IN0(\b/n831 ), .IN1(\b/n821 ), .SEL(msg[33]), .F(\b/n2839 )
         );
  MUX \b/U2859  ( .IN0(\b/n793 ), .IN1(\b/n2584 ), .SEL(msg[39]), .F(\b/n2838 ) );
  NANDN \b/U2858  ( .B(\b/n794 ), .A(msg[33]), .Z(\b/n2584 ) );
  MUX \b/U2857  ( .IN0(\b/n2837 ), .IN1(\b/n2816 ), .SEL(msg[38]), .F(
        shift_row_out[37]) );
  MUX \b/U2856  ( .IN0(\b/n2836 ), .IN1(\b/n2826 ), .SEL(msg[32]), .F(
        \b/n2837 ) );
  MUX \b/U2855  ( .IN0(\b/n2835 ), .IN1(\b/n2831 ), .SEL(msg[37]), .F(
        \b/n2836 ) );
  MUX \b/U2854  ( .IN0(\b/n2832 ), .IN1(\b/n2833 ), .SEL(msg[34]), .F(
        \b/n2835 ) );
  AND \b/U2853  ( .A(\b/n2602 ), .B(\b/n2834 ), .Z(\b/n2833 ) );
  MUX \b/U2852  ( .IN0(\b/n2580 ), .IN1(\b/n842 ), .SEL(msg[39]), .F(\b/n2832 ) );
  MUX \b/U2851  ( .IN0(\b/n2830 ), .IN1(\b/n2828 ), .SEL(msg[34]), .F(
        \b/n2831 ) );
  MUX \b/U2850  ( .IN0(\b/n797 ), .IN1(\b/n2829 ), .SEL(msg[39]), .F(\b/n2830 ) );
  NAND \b/U2849  ( .A(\b/n821 ), .B(\b/n851 ), .Z(\b/n2829 ) );
  MUX \b/U2848  ( .IN0(\b/n2580 ), .IN1(\b/n2827 ), .SEL(msg[39]), .F(
        \b/n2828 ) );
  NAND \b/U2847  ( .A(\b/n2571 ), .B(\b/n2632 ), .Z(\b/n2827 ) );
  MUX \b/U2846  ( .IN0(\b/n2825 ), .IN1(\b/n2821 ), .SEL(msg[37]), .F(
        \b/n2826 ) );
  MUX \b/U2845  ( .IN0(\b/n2824 ), .IN1(\b/n2823 ), .SEL(msg[34]), .F(
        \b/n2825 ) );
  MUX \b/U2844  ( .IN0(\b/n2592 ), .IN1(\b/n844 ), .SEL(msg[39]), .F(\b/n2824 ) );
  MUX \b/U2843  ( .IN0(\b/n2617 ), .IN1(\b/n2822 ), .SEL(msg[39]), .F(
        \b/n2823 ) );
  MUX \b/U2842  ( .IN0(\b/n840 ), .IN1(\b/n821 ), .SEL(msg[33]), .F(\b/n2822 )
         );
  MUX \b/U2841  ( .IN0(\b/n2820 ), .IN1(\b/n2819 ), .SEL(msg[34]), .F(
        \b/n2821 ) );
  MUX \b/U2840  ( .IN0(\b/n838 ), .IN1(n637), .SEL(msg[39]), .F(\b/n2820 ) );
  MUX \b/U2839  ( .IN0(\b/n2818 ), .IN1(\b/n2817 ), .SEL(msg[39]), .F(
        \b/n2819 ) );
  AND \b/U2838  ( .A(\b/n2577 ), .B(\b/n2652 ), .Z(\b/n2818 ) );
  MUX \b/U2837  ( .IN0(\b/n810 ), .IN1(\b/n794 ), .SEL(msg[33]), .F(\b/n2817 )
         );
  MUX \b/U2836  ( .IN0(\b/n2815 ), .IN1(\b/n2806 ), .SEL(msg[32]), .F(
        \b/n2816 ) );
  MUX \b/U2835  ( .IN0(\b/n2814 ), .IN1(\b/n2810 ), .SEL(msg[37]), .F(
        \b/n2815 ) );
  MUX \b/U2834  ( .IN0(\b/n2813 ), .IN1(\b/n2811 ), .SEL(msg[34]), .F(
        \b/n2814 ) );
  MUX \b/U2833  ( .IN0(\b/n2583 ), .IN1(\b/n2812 ), .SEL(msg[39]), .F(
        \b/n2813 ) );
  NAND \b/U2832  ( .A(msg[33]), .B(\b/n810 ), .Z(\b/n2812 ) );
  MUX \b/U2831  ( .IN0(\b/n794 ), .IN1(\b/n847 ), .SEL(msg[39]), .F(\b/n2811 )
         );
  MUX \b/U2830  ( .IN0(\b/n2809 ), .IN1(\b/n2808 ), .SEL(msg[34]), .F(
        \b/n2810 ) );
  MUX \b/U2829  ( .IN0(\b/n2609 ), .IN1(\b/n812 ), .SEL(msg[39]), .F(\b/n2809 ) );
  MUX \b/U2828  ( .IN0(\b/n2807 ), .IN1(\b/n2572 ), .SEL(n636), .F(\b/n2808 )
         );
  AND \b/U2827  ( .A(msg[39]), .B(msg[35]), .Z(\b/n2807 ) );
  MUX \b/U2826  ( .IN0(\b/n2805 ), .IN1(\b/n2802 ), .SEL(msg[37]), .F(
        \b/n2806 ) );
  MUX \b/U2825  ( .IN0(\b/n2804 ), .IN1(\b/n2803 ), .SEL(msg[34]), .F(
        \b/n2805 ) );
  MUX \b/U2824  ( .IN0(\b/n2733 ), .IN1(\b/n2572 ), .SEL(msg[39]), .F(
        \b/n2804 ) );
  MUX \b/U2823  ( .IN0(n635), .IN1(\b/n845 ), .SEL(msg[39]), .F(\b/n2803 ) );
  MUX \b/U2822  ( .IN0(\b/n2800 ), .IN1(\b/n2799 ), .SEL(msg[34]), .F(
        \b/n2802 ) );
  AND \b/U2821  ( .A(\b/n2801 ), .B(\b/n2701 ), .Z(\b/n2800 ) );
  MUX \b/U2820  ( .IN0(\b/n796 ), .IN1(\b/n840 ), .SEL(msg[39]), .F(\b/n2799 )
         );
  MUX \b/U2819  ( .IN0(\b/n2798 ), .IN1(\b/n2781 ), .SEL(msg[38]), .F(
        shift_row_out[36]) );
  MUX \b/U2818  ( .IN0(\b/n2797 ), .IN1(\b/n2789 ), .SEL(msg[32]), .F(
        \b/n2798 ) );
  MUX \b/U2817  ( .IN0(\b/n2796 ), .IN1(\b/n2793 ), .SEL(msg[37]), .F(
        \b/n2797 ) );
  MUX \b/U2816  ( .IN0(\b/n2795 ), .IN1(\b/n2794 ), .SEL(msg[34]), .F(
        \b/n2796 ) );
  MUX \b/U2815  ( .IN0(\b/n822 ), .IN1(\b/n843 ), .SEL(msg[39]), .F(\b/n2795 )
         );
  MUX \b/U2814  ( .IN0(\b/n2652 ), .IN1(\b/n2617 ), .SEL(msg[39]), .F(
        \b/n2794 ) );
  NAND \b/U2813  ( .A(msg[33]), .B(\b/n2571 ), .Z(\b/n2652 ) );
  MUX \b/U2812  ( .IN0(\b/n2790 ), .IN1(\b/n2791 ), .SEL(msg[34]), .F(
        \b/n2793 ) );
  AND \b/U2811  ( .A(\b/n2602 ), .B(\b/n2792 ), .Z(\b/n2791 ) );
  MUX \b/U2810  ( .IN0(\b/n2600 ), .IN1(\b/n825 ), .SEL(msg[39]), .F(\b/n2790 ) );
  MUX \b/U2809  ( .IN0(\b/n2788 ), .IN1(\b/n2785 ), .SEL(msg[37]), .F(
        \b/n2789 ) );
  MUX \b/U2808  ( .IN0(\b/n2787 ), .IN1(\b/n2786 ), .SEL(msg[34]), .F(
        \b/n2788 ) );
  MUX \b/U2807  ( .IN0(\b/n787 ), .IN1(\b/n833 ), .SEL(msg[39]), .F(\b/n2787 )
         );
  MUX \b/U2806  ( .IN0(\b/n794 ), .IN1(\b/n2580 ), .SEL(msg[39]), .F(\b/n2786 ) );
  MUX \b/U2805  ( .IN0(\b/n2784 ), .IN1(\b/n2782 ), .SEL(msg[34]), .F(
        \b/n2785 ) );
  MUX \b/U2804  ( .IN0(\b/n2596 ), .IN1(\b/n2783 ), .SEL(msg[39]), .F(
        \b/n2784 ) );
  AND \b/U2803  ( .A(\b/n2580 ), .B(\b/n851 ), .Z(\b/n2783 ) );
  MUX \b/U2802  ( .IN0(\b/n809 ), .IN1(\b/n828 ), .SEL(msg[39]), .F(\b/n2782 )
         );
  MUX \b/U2801  ( .IN0(\b/n2780 ), .IN1(\b/n2774 ), .SEL(msg[32]), .F(
        \b/n2781 ) );
  MUX \b/U2800  ( .IN0(\b/n2779 ), .IN1(\b/n2777 ), .SEL(msg[37]), .F(
        \b/n2780 ) );
  MUX \b/U2799  ( .IN0(\b/n2778 ), .IN1(\b/n2574 ), .SEL(msg[34]), .F(
        \b/n2779 ) );
  MUX \b/U2798  ( .IN0(\b/n2594 ), .IN1(\b/n830 ), .SEL(msg[39]), .F(\b/n2778 ) );
  MUX \b/U2797  ( .IN0(\b/n2776 ), .IN1(\b/n2775 ), .SEL(msg[34]), .F(
        \b/n2777 ) );
  MUX \b/U2796  ( .IN0(n634), .IN1(\b/n822 ), .SEL(msg[39]), .F(\b/n2776 ) );
  MUX \b/U2795  ( .IN0(\b/n2604 ), .IN1(\b/n2607 ), .SEL(msg[39]), .F(
        \b/n2775 ) );
  MUX \b/U2794  ( .IN0(\b/n2773 ), .IN1(\b/n2770 ), .SEL(msg[37]), .F(
        \b/n2774 ) );
  MUX \b/U2793  ( .IN0(\b/n2772 ), .IN1(\b/n2771 ), .SEL(msg[34]), .F(
        \b/n2773 ) );
  MUX \b/U2792  ( .IN0(\b/n795 ), .IN1(\b/n2576 ), .SEL(msg[39]), .F(\b/n2772 ) );
  MUX \b/U2791  ( .IN0(\b/n840 ), .IN1(\b/n2598 ), .SEL(msg[39]), .F(\b/n2771 ) );
  MUX \b/U2790  ( .IN0(\b/n783 ), .IN1(\b/n2769 ), .SEL(msg[34]), .F(\b/n2770 ) );
  MUX \b/U2789  ( .IN0(\b/n803 ), .IN1(\b/n2580 ), .SEL(msg[39]), .F(\b/n2769 ) );
  MUX \b/U2788  ( .IN0(\b/n2768 ), .IN1(\b/n2749 ), .SEL(msg[38]), .F(
        shift_row_out[35]) );
  MUX \b/U2787  ( .IN0(\b/n2767 ), .IN1(\b/n2759 ), .SEL(msg[32]), .F(
        \b/n2768 ) );
  MUX \b/U2786  ( .IN0(\b/n2766 ), .IN1(\b/n2763 ), .SEL(msg[37]), .F(
        \b/n2767 ) );
  MUX \b/U2785  ( .IN0(\b/n2765 ), .IN1(\b/n2764 ), .SEL(msg[39]), .F(
        \b/n2766 ) );
  MUX \b/U2784  ( .IN0(\b/n2588 ), .IN1(\b/n828 ), .SEL(msg[34]), .F(\b/n2765 ) );
  MUX \b/U2783  ( .IN0(n637), .IN1(\b/n786 ), .SEL(msg[34]), .F(\b/n2764 ) );
  MUX \b/U2782  ( .IN0(\b/n2761 ), .IN1(\b/n2760 ), .SEL(msg[39]), .F(
        \b/n2763 ) );
  AND \b/U2781  ( .A(\b/n2762 ), .B(msg[36]), .Z(\b/n2761 ) );
  MUX \b/U2780  ( .IN0(\b/n816 ), .IN1(\b/n2601 ), .SEL(msg[34]), .F(\b/n2760 ) );
  MUX \b/U2779  ( .IN0(\b/n2758 ), .IN1(\b/n2755 ), .SEL(msg[37]), .F(
        \b/n2759 ) );
  MUX \b/U2778  ( .IN0(\b/n2757 ), .IN1(\b/n2756 ), .SEL(msg[39]), .F(
        \b/n2758 ) );
  MUX \b/U2777  ( .IN0(\b/n2592 ), .IN1(n633), .SEL(msg[34]), .F(\b/n2757 ) );
  MUX \b/U2776  ( .IN0(\b/n784 ), .IN1(\b/n803 ), .SEL(msg[34]), .F(\b/n2756 )
         );
  MUX \b/U2775  ( .IN0(\b/n2751 ), .IN1(\b/n2752 ), .SEL(msg[39]), .F(
        \b/n2755 ) );
  NAND \b/U2774  ( .A(\b/n2753 ), .B(\b/n2754 ), .Z(\b/n2752 ) );
  MUX \b/U2773  ( .IN0(\b/n829 ), .IN1(\b/n2750 ), .SEL(msg[34]), .F(\b/n2751 ) );
  MUX \b/U2772  ( .IN0(\b/n804 ), .IN1(\b/n846 ), .SEL(msg[33]), .F(\b/n2750 )
         );
  MUX \b/U2771  ( .IN0(\b/n2748 ), .IN1(\b/n2739 ), .SEL(msg[32]), .F(
        \b/n2749 ) );
  MUX \b/U2770  ( .IN0(\b/n2747 ), .IN1(\b/n2743 ), .SEL(msg[37]), .F(
        \b/n2748 ) );
  MUX \b/U2769  ( .IN0(\b/n2745 ), .IN1(\b/n2744 ), .SEL(msg[39]), .F(
        \b/n2747 ) );
  NAND \b/U2768  ( .A(\b/n794 ), .B(\b/n2746 ), .Z(\b/n2745 ) );
  MUX \b/U2767  ( .IN0(\b/n845 ), .IN1(\b/n807 ), .SEL(msg[34]), .F(\b/n2744 )
         );
  MUX \b/U2766  ( .IN0(\b/n2742 ), .IN1(\b/n2740 ), .SEL(msg[39]), .F(
        \b/n2743 ) );
  MUX \b/U2765  ( .IN0(\b/n2583 ), .IN1(\b/n2741 ), .SEL(msg[34]), .F(
        \b/n2742 ) );
  AND \b/U2764  ( .A(msg[33]), .B(\b/n794 ), .Z(\b/n2741 ) );
  MUX \b/U2763  ( .IN0(\b/n799 ), .IN1(\b/n2602 ), .SEL(msg[34]), .F(\b/n2740 ) );
  MUX \b/U2762  ( .IN0(\b/n2738 ), .IN1(\b/n2732 ), .SEL(msg[37]), .F(
        \b/n2739 ) );
  MUX \b/U2761  ( .IN0(\b/n2737 ), .IN1(\b/n2735 ), .SEL(msg[39]), .F(
        \b/n2738 ) );
  MUX \b/U2760  ( .IN0(\b/n2736 ), .IN1(\b/n2572 ), .SEL(\b/n2620 ), .F(
        \b/n2737 ) );
  MUX \b/U2759  ( .IN0(msg[35]), .IN1(msg[36]), .SEL(msg[34]), .F(\b/n2736 )
         );
  MUX \b/U2758  ( .IN0(\b/n2602 ), .IN1(\b/n2733 ), .SEL(msg[34]), .F(
        \b/n2735 ) );
  NAND \b/U2757  ( .A(\b/n2572 ), .B(\b/n2734 ), .Z(\b/n2733 ) );
  MUX \b/U2756  ( .IN0(\b/n2729 ), .IN1(\b/n2730 ), .SEL(msg[39]), .F(
        \b/n2732 ) );
  AND \b/U2755  ( .A(\b/n827 ), .B(\b/n2731 ), .Z(\b/n2730 ) );
  MUX \b/U2754  ( .IN0(\b/n808 ), .IN1(\b/n2573 ), .SEL(msg[34]), .F(\b/n2729 ) );
  MUX \b/U2753  ( .IN0(\b/n2728 ), .IN1(\b/n2712 ), .SEL(msg[38]), .F(
        shift_row_out[34]) );
  MUX \b/U2752  ( .IN0(\b/n2727 ), .IN1(\b/n2719 ), .SEL(msg[32]), .F(
        \b/n2728 ) );
  MUX \b/U2751  ( .IN0(\b/n2726 ), .IN1(\b/n2722 ), .SEL(msg[37]), .F(
        \b/n2727 ) );
  MUX \b/U2750  ( .IN0(\b/n2725 ), .IN1(\b/n2723 ), .SEL(msg[34]), .F(
        \b/n2726 ) );
  MUX \b/U2749  ( .IN0(\b/n816 ), .IN1(\b/n2724 ), .SEL(msg[39]), .F(\b/n2725 ) );
  MUX \b/U2748  ( .IN0(\b/n2580 ), .IN1(\b/n794 ), .SEL(msg[33]), .F(\b/n2724 ) );
  MUX \b/U2747  ( .IN0(\b/n2619 ), .IN1(\b/n834 ), .SEL(msg[39]), .F(\b/n2723 ) );
  MUX \b/U2746  ( .IN0(\b/n2721 ), .IN1(\b/n2720 ), .SEL(msg[34]), .F(
        \b/n2722 ) );
  MUX \b/U2745  ( .IN0(\b/n2573 ), .IN1(\b/n801 ), .SEL(msg[39]), .F(\b/n2721 ) );
  MUX \b/U2744  ( .IN0(\b/n837 ), .IN1(\b/n2606 ), .SEL(msg[39]), .F(\b/n2720 ) );
  MUX \b/U2743  ( .IN0(\b/n2718 ), .IN1(\b/n2714 ), .SEL(msg[37]), .F(
        \b/n2719 ) );
  MUX \b/U2742  ( .IN0(\b/n2715 ), .IN1(\b/n783 ), .SEL(msg[34]), .F(\b/n2718 ) );
  NAND \b/U2741  ( .A(\b/n2716 ), .B(\b/n2717 ), .Z(\b/n2715 ) );
  MUX \b/U2740  ( .IN0(n635), .IN1(\b/n2713 ), .SEL(\b/n2618 ), .F(\b/n2714 )
         );
  MUX \b/U2739  ( .IN0(\b/n815 ), .IN1(\b/n2585 ), .SEL(msg[34]), .F(\b/n2713 ) );
  MUX \b/U2738  ( .IN0(\b/n2711 ), .IN1(\b/n2703 ), .SEL(msg[32]), .F(
        \b/n2712 ) );
  MUX \b/U2737  ( .IN0(\b/n2710 ), .IN1(\b/n2707 ), .SEL(msg[37]), .F(
        \b/n2711 ) );
  MUX \b/U2736  ( .IN0(\b/n2709 ), .IN1(\b/n2708 ), .SEL(msg[34]), .F(
        \b/n2710 ) );
  MUX \b/U2735  ( .IN0(\b/n843 ), .IN1(msg[33]), .SEL(msg[39]), .F(\b/n2709 )
         );
  MUX \b/U2734  ( .IN0(n638), .IN1(\b/n2586 ), .SEL(msg[39]), .F(\b/n2708 ) );
  MUX \b/U2733  ( .IN0(\b/n2706 ), .IN1(\b/n2705 ), .SEL(msg[34]), .F(
        \b/n2707 ) );
  MUX \b/U2732  ( .IN0(\b/n848 ), .IN1(\b/n842 ), .SEL(msg[39]), .F(\b/n2706 )
         );
  MUX \b/U2731  ( .IN0(n638), .IN1(\b/n2704 ), .SEL(msg[39]), .F(\b/n2705 ) );
  MUX \b/U2730  ( .IN0(\b/n794 ), .IN1(\b/n831 ), .SEL(msg[33]), .F(\b/n2704 )
         );
  MUX \b/U2729  ( .IN0(\b/n2702 ), .IN1(\b/n2696 ), .SEL(msg[37]), .F(
        \b/n2703 ) );
  MUX \b/U2728  ( .IN0(\b/n2699 ), .IN1(\b/n2698 ), .SEL(msg[34]), .F(
        \b/n2702 ) );
  NAND \b/U2727  ( .A(\b/n2700 ), .B(\b/n2701 ), .Z(\b/n2699 ) );
  MUX \b/U2726  ( .IN0(\b/n2572 ), .IN1(\b/n2697 ), .SEL(n636), .F(\b/n2698 )
         );
  MUX \b/U2725  ( .IN0(msg[35]), .IN1(\b/n804 ), .SEL(msg[39]), .F(\b/n2697 )
         );
  MUX \b/U2724  ( .IN0(\b/n2695 ), .IN1(\b/n2694 ), .SEL(msg[34]), .F(
        \b/n2696 ) );
  MUX \b/U2723  ( .IN0(\b/n2617 ), .IN1(\b/n802 ), .SEL(msg[39]), .F(\b/n2695 ) );
  MUX \b/U2722  ( .IN0(\b/n2613 ), .IN1(\b/n2693 ), .SEL(msg[39]), .F(
        \b/n2694 ) );
  MUX \b/U2721  ( .IN0(\b/n2575 ), .IN1(\b/n2580 ), .SEL(msg[33]), .F(
        \b/n2693 ) );
  MUX \b/U2720  ( .IN0(\b/n2692 ), .IN1(\b/n2674 ), .SEL(msg[38]), .F(
        shift_row_out[33]) );
  MUX \b/U2719  ( .IN0(\b/n2691 ), .IN1(\b/n2682 ), .SEL(msg[32]), .F(
        \b/n2692 ) );
  MUX \b/U2718  ( .IN0(\b/n2690 ), .IN1(\b/n2686 ), .SEL(msg[37]), .F(
        \b/n2691 ) );
  MUX \b/U2717  ( .IN0(\b/n2689 ), .IN1(\b/n2688 ), .SEL(msg[34]), .F(
        \b/n2690 ) );
  MUX \b/U2716  ( .IN0(\b/n839 ), .IN1(n640), .SEL(msg[39]), .F(\b/n2689 ) );
  MUX \b/U2715  ( .IN0(\b/n2687 ), .IN1(n634), .SEL(msg[39]), .F(\b/n2688 ) );
  NAND \b/U2714  ( .A(\b/n851 ), .B(\b/n810 ), .Z(\b/n2687 ) );
  MUX \b/U2713  ( .IN0(\b/n2685 ), .IN1(\b/n2684 ), .SEL(msg[34]), .F(
        \b/n2686 ) );
  MUX \b/U2712  ( .IN0(\b/n787 ), .IN1(\b/n2587 ), .SEL(msg[39]), .F(\b/n2685 ) );
  MUX \b/U2711  ( .IN0(\b/n2577 ), .IN1(\b/n2683 ), .SEL(msg[39]), .F(
        \b/n2684 ) );
  AND \b/U2710  ( .A(msg[33]), .B(msg[36]), .Z(\b/n2683 ) );
  MUX \b/U2709  ( .IN0(\b/n2681 ), .IN1(\b/n2678 ), .SEL(msg[37]), .F(
        \b/n2682 ) );
  MUX \b/U2708  ( .IN0(\b/n2680 ), .IN1(\b/n2679 ), .SEL(msg[34]), .F(
        \b/n2681 ) );
  MUX \b/U2707  ( .IN0(\b/n2616 ), .IN1(\b/n848 ), .SEL(msg[39]), .F(\b/n2680 ) );
  MUX \b/U2706  ( .IN0(\b/n823 ), .IN1(\b/n2585 ), .SEL(msg[39]), .F(\b/n2679 ) );
  MUX \b/U2705  ( .IN0(\b/n2675 ), .IN1(\b/n2676 ), .SEL(msg[34]), .F(
        \b/n2678 ) );
  AND \b/U2704  ( .A(\b/n2677 ), .B(\b/n2632 ), .Z(\b/n2676 ) );
  MUX \b/U2703  ( .IN0(\b/n2591 ), .IN1(\b/n2580 ), .SEL(msg[39]), .F(
        \b/n2675 ) );
  MUX \b/U2702  ( .IN0(\b/n2673 ), .IN1(\b/n2665 ), .SEL(msg[32]), .F(
        \b/n2674 ) );
  MUX \b/U2701  ( .IN0(\b/n2672 ), .IN1(\b/n2668 ), .SEL(msg[37]), .F(
        \b/n2673 ) );
  MUX \b/U2700  ( .IN0(\b/n2671 ), .IN1(\b/n2670 ), .SEL(msg[34]), .F(
        \b/n2672 ) );
  MUX \b/U2699  ( .IN0(\b/n2579 ), .IN1(\b/n812 ), .SEL(msg[39]), .F(\b/n2671 ) );
  MUX \b/U2698  ( .IN0(\b/n2669 ), .IN1(\b/n796 ), .SEL(msg[39]), .F(\b/n2670 ) );
  MUX \b/U2697  ( .IN0(\b/n2577 ), .IN1(\b/n804 ), .SEL(msg[33]), .F(\b/n2669 ) );
  MUX \b/U2696  ( .IN0(\b/n2667 ), .IN1(\b/n2666 ), .SEL(msg[34]), .F(
        \b/n2668 ) );
  MUX \b/U2695  ( .IN0(\b/n843 ), .IN1(\b/n821 ), .SEL(msg[39]), .F(\b/n2667 )
         );
  MUX \b/U2694  ( .IN0(\b/n839 ), .IN1(\b/n799 ), .SEL(msg[39]), .F(\b/n2666 )
         );
  MUX \b/U2693  ( .IN0(\b/n2664 ), .IN1(\b/n2659 ), .SEL(msg[37]), .F(
        \b/n2665 ) );
  MUX \b/U2692  ( .IN0(\b/n2663 ), .IN1(\b/n2660 ), .SEL(msg[34]), .F(
        \b/n2664 ) );
  MUX \b/U2691  ( .IN0(\b/n2661 ), .IN1(\b/n2662 ), .SEL(msg[39]), .F(
        \b/n2663 ) );
  NAND \b/U2690  ( .A(\b/n2580 ), .B(\b/n2652 ), .Z(\b/n2662 ) );
  MUX \b/U2689  ( .IN0(\b/n2580 ), .IN1(\b/n804 ), .SEL(msg[33]), .F(\b/n2661 ) );
  MUX \b/U2688  ( .IN0(\b/n2597 ), .IN1(\b/n2595 ), .SEL(msg[39]), .F(
        \b/n2660 ) );
  MUX \b/U2687  ( .IN0(\b/n2615 ), .IN1(\b/n2658 ), .SEL(msg[34]), .F(
        \b/n2659 ) );
  MUX \b/U2686  ( .IN0(\b/n810 ), .IN1(\b/n842 ), .SEL(msg[39]), .F(\b/n2658 )
         );
  MUX \b/U2685  ( .IN0(\b/n2657 ), .IN1(\b/n2640 ), .SEL(msg[38]), .F(
        shift_row_out[32]) );
  MUX \b/U2684  ( .IN0(\b/n2656 ), .IN1(\b/n2648 ), .SEL(msg[32]), .F(
        \b/n2657 ) );
  MUX \b/U2683  ( .IN0(\b/n2655 ), .IN1(\b/n2653 ), .SEL(msg[34]), .F(
        \b/n2656 ) );
  MUX \b/U2682  ( .IN0(\b/n784 ), .IN1(\b/n2654 ), .SEL(msg[39]), .F(\b/n2655 ) );
  MUX \b/U2681  ( .IN0(\b/n837 ), .IN1(\b/n840 ), .SEL(msg[37]), .F(\b/n2654 )
         );
  MUX \b/U2680  ( .IN0(\b/n2650 ), .IN1(\b/n2649 ), .SEL(msg[39]), .F(
        \b/n2653 ) );
  NAND \b/U2679  ( .A(\b/n2651 ), .B(\b/n2652 ), .Z(\b/n2650 ) );
  MUX \b/U2678  ( .IN0(\b/n836 ), .IN1(\b/n851 ), .SEL(msg[37]), .F(\b/n2649 )
         );
  MUX \b/U2677  ( .IN0(\b/n2647 ), .IN1(\b/n2643 ), .SEL(msg[34]), .F(
        \b/n2648 ) );
  MUX \b/U2676  ( .IN0(\b/n2646 ), .IN1(\b/n2644 ), .SEL(msg[39]), .F(
        \b/n2647 ) );
  MUX \b/U2675  ( .IN0(\b/n2645 ), .IN1(\b/n789 ), .SEL(msg[37]), .F(\b/n2646 ) );
  NAND \b/U2674  ( .A(\b/n851 ), .B(\b/n2572 ), .Z(\b/n2645 ) );
  MUX \b/U2672  ( .IN0(\b/n2642 ), .IN1(\b/n2641 ), .SEL(msg[39]), .F(
        \b/n2643 ) );
  MUX \b/U2671  ( .IN0(n635), .IN1(\b/n786 ), .SEL(msg[37]), .F(\b/n2642 ) );
  MUX \b/U2670  ( .IN0(\b/n838 ), .IN1(\b/n794 ), .SEL(msg[37]), .F(\b/n2641 )
         );
  MUX \b/U2669  ( .IN0(\b/n2639 ), .IN1(\b/n2629 ), .SEL(msg[32]), .F(
        \b/n2640 ) );
  MUX \b/U2668  ( .IN0(\b/n2638 ), .IN1(\b/n2634 ), .SEL(msg[34]), .F(
        \b/n2639 ) );
  MUX \b/U2667  ( .IN0(\b/n2637 ), .IN1(\b/n2636 ), .SEL(msg[39]), .F(
        \b/n2638 ) );
  MUX \b/U2666  ( .IN0(n633), .IN1(\b/n790 ), .SEL(msg[37]), .F(\b/n2637 ) );
  MUX \b/U2665  ( .IN0(\b/n2635 ), .IN1(\b/n827 ), .SEL(msg[37]), .F(\b/n2636 ) );
  NAND \b/U2664  ( .A(\b/n2571 ), .B(\b/n2573 ), .Z(\b/n2635 ) );
  MUX \b/U2663  ( .IN0(\b/n2633 ), .IN1(\b/n2630 ), .SEL(msg[39]), .F(
        \b/n2634 ) );
  MUX \b/U2662  ( .IN0(\b/n797 ), .IN1(\b/n2631 ), .SEL(msg[37]), .F(\b/n2633 ) );
  NAND \b/U2661  ( .A(\b/n2575 ), .B(\b/n2632 ), .Z(\b/n2631 ) );
  MUX \b/U2660  ( .IN0(\b/n2590 ), .IN1(\b/n2581 ), .SEL(msg[37]), .F(
        \b/n2630 ) );
  MUX \b/U2659  ( .IN0(\b/n2628 ), .IN1(\b/n2624 ), .SEL(msg[34]), .F(
        \b/n2629 ) );
  MUX \b/U2658  ( .IN0(\b/n2626 ), .IN1(\b/n2625 ), .SEL(msg[39]), .F(
        \b/n2628 ) );
  NAND \b/U2657  ( .A(\b/n2627 ), .B(\b/n2614 ), .Z(\b/n2626 ) );
  MUX \b/U2656  ( .IN0(msg[35]), .IN1(\b/n2606 ), .SEL(msg[37]), .F(\b/n2625 )
         );
  MUX \b/U2655  ( .IN0(\b/n2623 ), .IN1(\b/n2622 ), .SEL(msg[39]), .F(
        \b/n2624 ) );
  MUX \b/U2654  ( .IN0(\b/n802 ), .IN1(\b/n818 ), .SEL(msg[37]), .F(\b/n2623 )
         );
  MUX \b/U2653  ( .IN0(\b/n835 ), .IN1(\b/n823 ), .SEL(msg[37]), .F(\b/n2622 )
         );
  XOR \b/U2652  ( .A(\b/n2572 ), .B(msg[33]), .Z(\b/n2621 ) );
  XOR \b/U2651  ( .A(msg[33]), .B(msg[34]), .Z(\b/n2620 ) );
  XOR \b/U2650  ( .A(msg[33]), .B(msg[35]), .Z(\b/n2619 ) );
  XOR \b/U2649  ( .A(msg[34]), .B(msg[39]), .Z(\b/n2618 ) );
  XOR \b/U2648  ( .A(\b/n851 ), .B(\b/n794 ), .Z(\b/n2617 ) );
  XOR \b/U2647  ( .A(msg[33]), .B(\b/n840 ), .Z(\b/n2616 ) );
  XOR \b/U2645  ( .A(msg[33]), .B(msg[37]), .Z(\b/n2614 ) );
  NAND \b/U2644  ( .A(msg[33]), .B(msg[35]), .Z(\b/n2613 ) );
  MUX \b/U2643  ( .IN0(\b/n2572 ), .IN1(\b/n794 ), .SEL(msg[33]), .F(\b/n2612 ) );
  MUX \b/U2641  ( .IN0(msg[35]), .IN1(\b/n831 ), .SEL(msg[33]), .F(\b/n2610 )
         );
  MUX \b/U2640  ( .IN0(\b/n810 ), .IN1(\b/n831 ), .SEL(msg[33]), .F(\b/n2609 )
         );
  MUX \b/U2639  ( .IN0(\b/n2575 ), .IN1(\b/n2577 ), .SEL(msg[33]), .F(
        \b/n2608 ) );
  MUX \b/U2638  ( .IN0(msg[36]), .IN1(\b/n810 ), .SEL(msg[33]), .F(\b/n2607 )
         );
  OR \b/U2637  ( .A(msg[33]), .B(msg[36]), .Z(\b/n2606 ) );
  NAND \b/U2635  ( .A(\b/n831 ), .B(\b/n851 ), .Z(\b/n2604 ) );
  MUX \b/U2634  ( .IN0(\b/n831 ), .IN1(msg[36]), .SEL(msg[33]), .F(\b/n2603 )
         );
  MUX \b/U2633  ( .IN0(\b/n2571 ), .IN1(\b/n2580 ), .SEL(msg[33]), .F(
        \b/n2602 ) );
  MUX \b/U2632  ( .IN0(\b/n846 ), .IN1(msg[36]), .SEL(msg[33]), .F(\b/n2601 )
         );
  MUX \b/U2631  ( .IN0(\b/n804 ), .IN1(\b/n831 ), .SEL(msg[33]), .F(\b/n2600 )
         );
  MUX \b/U2630  ( .IN0(\b/n2571 ), .IN1(msg[36]), .SEL(msg[33]), .F(\b/n2599 )
         );
  MUX \b/U2629  ( .IN0(\b/n821 ), .IN1(\b/n810 ), .SEL(msg[33]), .F(\b/n2598 )
         );
  XOR \b/U2628  ( .A(\b/n804 ), .B(msg[33]), .Z(\b/n2597 ) );
  MUX \b/U2627  ( .IN0(\b/n2577 ), .IN1(\b/n821 ), .SEL(msg[33]), .F(\b/n2596 ) );
  NANDN \b/U2626  ( .B(msg[33]), .A(msg[35]), .Z(\b/n2595 ) );
  MUX \b/U2625  ( .IN0(\b/n794 ), .IN1(msg[35]), .SEL(msg[33]), .F(\b/n2594 )
         );
  NAND \b/U2623  ( .A(\b/n2575 ), .B(\b/n851 ), .Z(\b/n2592 ) );
  MUX \b/U2622  ( .IN0(msg[36]), .IN1(\b/n2572 ), .SEL(msg[33]), .F(\b/n2591 )
         );
  MUX \b/U2621  ( .IN0(\b/n821 ), .IN1(msg[35]), .SEL(msg[33]), .F(\b/n2590 )
         );
  MUX \b/U2619  ( .IN0(msg[36]), .IN1(\b/n840 ), .SEL(msg[33]), .F(\b/n2588 )
         );
  MUX \b/U2618  ( .IN0(\b/n794 ), .IN1(\b/n846 ), .SEL(msg[33]), .F(\b/n2587 )
         );
  NAND \b/U2617  ( .A(\b/n2573 ), .B(\b/n794 ), .Z(\b/n2586 ) );
  MUX \b/U2616  ( .IN0(\b/n2572 ), .IN1(\b/n2580 ), .SEL(msg[33]), .F(
        \b/n2585 ) );
  NAND \b/U2615  ( .A(\b/n2584 ), .B(\b/n2571 ), .Z(\b/n2583 ) );
  MUX \b/U2614  ( .IN0(\b/n2575 ), .IN1(\b/n846 ), .SEL(msg[33]), .F(\b/n2582 ) );
  MUX \b/U2613  ( .IN0(\b/n846 ), .IN1(\b/n810 ), .SEL(msg[33]), .F(\b/n2581 )
         );
  NANDN \b/U2612  ( .B(msg[35]), .A(msg[36]), .Z(\b/n2580 ) );
  MUX \b/U2611  ( .IN0(\b/n2575 ), .IN1(msg[35]), .SEL(msg[33]), .F(\b/n2579 )
         );
  OR \b/U2610  ( .A(msg[35]), .B(msg[36]), .Z(\b/n2575 ) );
  MUX \b/U2609  ( .IN0(\b/n794 ), .IN1(\b/n810 ), .SEL(msg[33]), .F(\b/n2578 )
         );
  XOR \b/U2608  ( .A(\b/n804 ), .B(msg[35]), .Z(\b/n2577 ) );
  NANDN \b/U2607  ( .B(msg[35]), .A(msg[33]), .Z(\b/n2576 ) );
  NAND \b/U2606  ( .A(\b/n2575 ), .B(\b/n2573 ), .Z(\b/n2574 ) );
  NAND \b/U2605  ( .A(msg[33]), .B(\b/n2572 ), .Z(\b/n2573 ) );
  NANDN \b/U2604  ( .B(msg[36]), .A(msg[35]), .Z(\b/n2572 ) );
  NAND \b/U2603  ( .A(msg[35]), .B(msg[36]), .Z(\b/n2571 ) );
  MUX \b/U2602  ( .IN0(msg[28]), .IN1(\b/n2212 ), .SEL(msg[25]), .F(\b/n2570 )
         );
  MUX \b/U2601  ( .IN0(msg[28]), .IN1(\b/n2221 ), .SEL(msg[25]), .F(\b/n2569 )
         );
  MUX \b/U2600  ( .IN0(\b/n2213 ), .IN1(\b/n2216 ), .SEL(msg[25]), .F(
        \b/n2568 ) );
  MUX \b/U2599  ( .IN0(\b/n2218 ), .IN1(\b/n911 ), .SEL(msg[25]), .F(\b/n2567 ) );
  MUX \b/U2597  ( .IN0(\b/n2221 ), .IN1(\b/n2212 ), .SEL(msg[26]), .F(
        \b/n2394 ) );
  MUX \b/U2596  ( .IN0(\b/n2214 ), .IN1(\b/n922 ), .SEL(msg[26]), .F(\b/n2395 ) );
  MUX \b/U2595  ( .IN0(\b/n865 ), .IN1(\b/n875 ), .SEL(msg[25]), .F(\b/n2358 )
         );
  MUX \b/U2594  ( .IN0(\b/n2242 ), .IN1(\b/n2553 ), .SEL(msg[31]), .F(
        \b/n2565 ) );
  MUX \b/U2593  ( .IN0(\b/n2216 ), .IN1(\b/n2212 ), .SEL(msg[25]), .F(
        \b/n2556 ) );
  MUX \b/U2592  ( .IN0(\b/n917 ), .IN1(\b/n2218 ), .SEL(msg[25]), .F(\b/n2564 ) );
  MUX \b/U2591  ( .IN0(msg[27]), .IN1(\b/n911 ), .SEL(msg[25]), .F(\b/n2563 )
         );
  MUX \b/U2590  ( .IN0(\b/n2221 ), .IN1(\b/n917 ), .SEL(msg[25]), .F(\b/n2562 ) );
  MUX \b/U2589  ( .IN0(msg[28]), .IN1(\b/n2218 ), .SEL(msg[25]), .F(\b/n2561 )
         );
  MUX \b/U2588  ( .IN0(\b/n902 ), .IN1(\b/n881 ), .SEL(msg[29]), .F(\b/n2268 )
         );
  MUX \b/U2587  ( .IN0(\b/n2213 ), .IN1(\b/n875 ), .SEL(msg[25]), .F(\b/n2560 ) );
  NANDN \b/U2584  ( .B(\b/n2219 ), .A(msg[31]), .Z(\b/n2533 ) );
  NAND \b/U2583  ( .A(msg[31]), .B(\b/n878 ), .Z(\b/n2501 ) );
  NAND \b/U2582  ( .A(msg[31]), .B(\b/n890 ), .Z(\b/n2442 ) );
  NAND \b/U2581  ( .A(msg[31]), .B(\b/n2550 ), .Z(\b/n2475 ) );
  NAND \b/U2580  ( .A(msg[31]), .B(\b/n2470 ), .Z(\b/n2433 ) );
  NAND \b/U2578  ( .A(\b/n922 ), .B(\b/n911 ), .Z(\b/n2554 ) );
  NAND \b/U2577  ( .A(msg[31]), .B(\b/n2552 ), .Z(\b/n2547 ) );
  NAND \b/U2576  ( .A(n632), .B(msg[31]), .Z(\b/n2527 ) );
  NAND \b/U2574  ( .A(msg[26]), .B(\b/n2221 ), .Z(\b/n2387 ) );
  NAND \b/U2573  ( .A(\b/n911 ), .B(msg[25]), .Z(\b/n2342 ) );
  NAND \b/U2572  ( .A(msg[31]), .B(\b/n2556 ), .Z(\b/n2341 ) );
  NAND \b/U2570  ( .A(\b/n2554 ), .B(msg[31]), .Z(\b/n2357 ) );
  NAND \b/U2569  ( .A(\b/n2375 ), .B(\b/n2221 ), .Z(\b/n2553 ) );
  NANDN \b/U2568  ( .B(\b/n865 ), .A(\b/n922 ), .Z(\b/n2552 ) );
  NAND \b/U2566  ( .A(msg[25]), .B(\b/n2221 ), .Z(\b/n2273 ) );
  NAND \b/U2565  ( .A(\b/n865 ), .B(\b/n922 ), .Z(\b/n2550 ) );
  NAND \b/U2562  ( .A(msg[25]), .B(\b/n2216 ), .Z(\b/n2375 ) );
  ANDN \b/U2560  ( .A(msg[26]), .B(msg[25]), .Z(\b/n2403 ) );
  AND \b/U2559  ( .A(\b/n2213 ), .B(\b/n2547 ), .Z(\b/n2318 ) );
  MUX \b/U2558  ( .IN0(\b/n2546 ), .IN1(\b/n2530 ), .SEL(msg[30]), .F(
        shift_row_out[63]) );
  MUX \b/U2557  ( .IN0(\b/n2545 ), .IN1(\b/n2538 ), .SEL(msg[24]), .F(
        \b/n2546 ) );
  MUX \b/U2556  ( .IN0(\b/n2544 ), .IN1(\b/n2541 ), .SEL(msg[29]), .F(
        \b/n2545 ) );
  MUX \b/U2555  ( .IN0(\b/n2543 ), .IN1(\b/n2542 ), .SEL(msg[26]), .F(
        \b/n2544 ) );
  MUX \b/U2554  ( .IN0(msg[28]), .IN1(\b/n882 ), .SEL(msg[31]), .F(\b/n2543 )
         );
  MUX \b/U2553  ( .IN0(\b/n2214 ), .IN1(\b/n886 ), .SEL(msg[31]), .F(\b/n2542 ) );
  MUX \b/U2552  ( .IN0(\b/n2540 ), .IN1(\b/n2539 ), .SEL(msg[26]), .F(
        \b/n2541 ) );
  MUX \b/U2551  ( .IN0(\b/n2272 ), .IN1(\b/n878 ), .SEL(msg[31]), .F(\b/n2540 ) );
  MUX \b/U2550  ( .IN0(\b/n2224 ), .IN1(\b/n2235 ), .SEL(msg[31]), .F(
        \b/n2539 ) );
  MUX \b/U2549  ( .IN0(\b/n2537 ), .IN1(\b/n2534 ), .SEL(msg[29]), .F(
        \b/n2538 ) );
  MUX \b/U2548  ( .IN0(\b/n2536 ), .IN1(\b/n2535 ), .SEL(msg[26]), .F(
        \b/n2537 ) );
  MUX \b/U2547  ( .IN0(\b/n2248 ), .IN1(\b/n2223 ), .SEL(msg[31]), .F(
        \b/n2536 ) );
  MUX \b/U2546  ( .IN0(\b/n890 ), .IN1(\b/n2244 ), .SEL(msg[31]), .F(\b/n2535 ) );
  MUX \b/U2545  ( .IN0(\b/n2532 ), .IN1(\b/n2531 ), .SEL(msg[26]), .F(
        \b/n2534 ) );
  AND \b/U2544  ( .A(\b/n880 ), .B(\b/n2533 ), .Z(\b/n2532 ) );
  MUX \b/U2543  ( .IN0(\b/n2228 ), .IN1(n631), .SEL(msg[31]), .F(\b/n2531 ) );
  MUX \b/U2542  ( .IN0(\b/n2529 ), .IN1(\b/n2521 ), .SEL(msg[24]), .F(
        \b/n2530 ) );
  MUX \b/U2541  ( .IN0(\b/n2528 ), .IN1(\b/n2524 ), .SEL(msg[29]), .F(
        \b/n2529 ) );
  MUX \b/U2540  ( .IN0(\b/n2525 ), .IN1(\b/n2526 ), .SEL(msg[26]), .F(
        \b/n2528 ) );
  NAND \b/U2539  ( .A(\b/n2342 ), .B(\b/n2527 ), .Z(\b/n2526 ) );
  MUX \b/U2538  ( .IN0(\b/n920 ), .IN1(\b/n912 ), .SEL(msg[31]), .F(\b/n2525 )
         );
  MUX \b/U2537  ( .IN0(\b/n2523 ), .IN1(\b/n2522 ), .SEL(msg[26]), .F(
        \b/n2524 ) );
  MUX \b/U2536  ( .IN0(\b/n2218 ), .IN1(\b/n2212 ), .SEL(msg[31]), .F(
        \b/n2523 ) );
  MUX \b/U2535  ( .IN0(\b/n913 ), .IN1(\b/n2249 ), .SEL(msg[31]), .F(\b/n2522 ) );
  MUX \b/U2534  ( .IN0(\b/n2520 ), .IN1(\b/n2517 ), .SEL(msg[29]), .F(
        \b/n2521 ) );
  MUX \b/U2533  ( .IN0(\b/n2519 ), .IN1(\b/n2518 ), .SEL(msg[26]), .F(
        \b/n2520 ) );
  MUX \b/U2532  ( .IN0(\b/n2253 ), .IN1(\b/n2239 ), .SEL(msg[31]), .F(
        \b/n2519 ) );
  MUX \b/U2531  ( .IN0(\b/n866 ), .IN1(\b/n2221 ), .SEL(msg[31]), .F(\b/n2518 ) );
  MUX \b/U2530  ( .IN0(\b/n2516 ), .IN1(\b/n2515 ), .SEL(msg[26]), .F(
        \b/n2517 ) );
  MUX \b/U2529  ( .IN0(\b/n2254 ), .IN1(\b/n2262 ), .SEL(msg[31]), .F(
        \b/n2516 ) );
  MUX \b/U2528  ( .IN0(\b/n2247 ), .IN1(\b/n2514 ), .SEL(msg[31]), .F(
        \b/n2515 ) );
  MUX \b/U2527  ( .IN0(\b/n917 ), .IN1(\b/n875 ), .SEL(msg[25]), .F(\b/n2514 )
         );
  MUX \b/U2526  ( .IN0(\b/n2513 ), .IN1(\b/n2495 ), .SEL(msg[30]), .F(
        shift_row_out[62]) );
  MUX \b/U2525  ( .IN0(\b/n2512 ), .IN1(\b/n2503 ), .SEL(msg[24]), .F(
        \b/n2513 ) );
  MUX \b/U2524  ( .IN0(\b/n2511 ), .IN1(\b/n2506 ), .SEL(msg[29]), .F(
        \b/n2512 ) );
  MUX \b/U2523  ( .IN0(\b/n2510 ), .IN1(\b/n2508 ), .SEL(msg[26]), .F(
        \b/n2511 ) );
  MUX \b/U2522  ( .IN0(\b/n2509 ), .IN1(\b/n2225 ), .SEL(msg[31]), .F(
        \b/n2510 ) );
  MUX \b/U2521  ( .IN0(\b/n917 ), .IN1(\b/n2212 ), .SEL(msg[25]), .F(\b/n2509 ) );
  MUX \b/U2520  ( .IN0(\b/n2507 ), .IN1(\b/n905 ), .SEL(msg[31]), .F(\b/n2508 ) );
  MUX \b/U2519  ( .IN0(\b/n2212 ), .IN1(\b/n2213 ), .SEL(msg[25]), .F(
        \b/n2507 ) );
  MUX \b/U2518  ( .IN0(\b/n2505 ), .IN1(\b/n2504 ), .SEL(msg[26]), .F(
        \b/n2506 ) );
  MUX \b/U2517  ( .IN0(n630), .IN1(\b/n2293 ), .SEL(msg[31]), .F(\b/n2505 ) );
  MUX \b/U2516  ( .IN0(\b/n2251 ), .IN1(\b/n2258 ), .SEL(msg[31]), .F(
        \b/n2504 ) );
  MUX \b/U2515  ( .IN0(\b/n2502 ), .IN1(\b/n2498 ), .SEL(msg[29]), .F(
        \b/n2503 ) );
  MUX \b/U2514  ( .IN0(\b/n2500 ), .IN1(\b/n2499 ), .SEL(msg[26]), .F(
        \b/n2502 ) );
  AND \b/U2513  ( .A(\b/n858 ), .B(\b/n2501 ), .Z(\b/n2500 ) );
  MUX \b/U2512  ( .IN0(\b/n2328 ), .IN1(msg[27]), .SEL(msg[31]), .F(\b/n2499 )
         );
  MUX \b/U2511  ( .IN0(\b/n2497 ), .IN1(\b/n2496 ), .SEL(msg[26]), .F(
        \b/n2498 ) );
  MUX \b/U2510  ( .IN0(\b/n901 ), .IN1(\b/n2216 ), .SEL(msg[31]), .F(\b/n2497 ) );
  MUX \b/U2508  ( .IN0(\b/n2494 ), .IN1(\b/n2487 ), .SEL(msg[24]), .F(
        \b/n2495 ) );
  MUX \b/U2507  ( .IN0(\b/n2493 ), .IN1(\b/n2490 ), .SEL(msg[29]), .F(
        \b/n2494 ) );
  MUX \b/U2506  ( .IN0(\b/n2492 ), .IN1(\b/n2491 ), .SEL(msg[26]), .F(
        \b/n2493 ) );
  MUX \b/U2505  ( .IN0(\b/n897 ), .IN1(\b/n2220 ), .SEL(msg[31]), .F(\b/n2492 ) );
  MUX \b/U2504  ( .IN0(\b/n2224 ), .IN1(n631), .SEL(msg[31]), .F(\b/n2491 ) );
  MUX \b/U2503  ( .IN0(\b/n2489 ), .IN1(\b/n2488 ), .SEL(msg[26]), .F(
        \b/n2490 ) );
  MUX \b/U2502  ( .IN0(\b/n2240 ), .IN1(\b/n862 ), .SEL(msg[31]), .F(\b/n2489 ) );
  MUX \b/U2501  ( .IN0(\b/n882 ), .IN1(\b/n912 ), .SEL(msg[31]), .F(\b/n2488 )
         );
  MUX \b/U2500  ( .IN0(\b/n2486 ), .IN1(\b/n2482 ), .SEL(msg[29]), .F(
        \b/n2487 ) );
  MUX \b/U2499  ( .IN0(\b/n2485 ), .IN1(\b/n2484 ), .SEL(msg[26]), .F(
        \b/n2486 ) );
  MUX \b/U2498  ( .IN0(\b/n2229 ), .IN1(\b/n912 ), .SEL(msg[31]), .F(\b/n2485 ) );
  MUX \b/U2497  ( .IN0(\b/n2483 ), .IN1(\b/n2250 ), .SEL(msg[31]), .F(
        \b/n2484 ) );
  NANDN \b/U2496  ( .B(msg[28]), .A(msg[25]), .Z(\b/n2483 ) );
  MUX \b/U2495  ( .IN0(\b/n2481 ), .IN1(\b/n2479 ), .SEL(msg[26]), .F(
        \b/n2482 ) );
  MUX \b/U2494  ( .IN0(\b/n875 ), .IN1(\b/n2480 ), .SEL(msg[31]), .F(\b/n2481 ) );
  MUX \b/U2493  ( .IN0(\b/n902 ), .IN1(\b/n892 ), .SEL(msg[25]), .F(\b/n2480 )
         );
  MUX \b/U2492  ( .IN0(\b/n864 ), .IN1(\b/n2225 ), .SEL(msg[31]), .F(\b/n2479 ) );
  NANDN \b/U2491  ( .B(\b/n865 ), .A(msg[25]), .Z(\b/n2225 ) );
  MUX \b/U2490  ( .IN0(\b/n2478 ), .IN1(\b/n2457 ), .SEL(msg[30]), .F(
        shift_row_out[61]) );
  MUX \b/U2489  ( .IN0(\b/n2477 ), .IN1(\b/n2467 ), .SEL(msg[24]), .F(
        \b/n2478 ) );
  MUX \b/U2488  ( .IN0(\b/n2476 ), .IN1(\b/n2472 ), .SEL(msg[29]), .F(
        \b/n2477 ) );
  MUX \b/U2487  ( .IN0(\b/n2473 ), .IN1(\b/n2474 ), .SEL(msg[26]), .F(
        \b/n2476 ) );
  AND \b/U2486  ( .A(\b/n2243 ), .B(\b/n2475 ), .Z(\b/n2474 ) );
  MUX \b/U2485  ( .IN0(\b/n2221 ), .IN1(\b/n913 ), .SEL(msg[31]), .F(\b/n2473 ) );
  MUX \b/U2484  ( .IN0(\b/n2471 ), .IN1(\b/n2469 ), .SEL(msg[26]), .F(
        \b/n2472 ) );
  MUX \b/U2483  ( .IN0(\b/n868 ), .IN1(\b/n2470 ), .SEL(msg[31]), .F(\b/n2471 ) );
  NAND \b/U2482  ( .A(\b/n892 ), .B(\b/n922 ), .Z(\b/n2470 ) );
  MUX \b/U2481  ( .IN0(\b/n2221 ), .IN1(\b/n2468 ), .SEL(msg[31]), .F(
        \b/n2469 ) );
  NAND \b/U2480  ( .A(\b/n2212 ), .B(\b/n2273 ), .Z(\b/n2468 ) );
  MUX \b/U2479  ( .IN0(\b/n2466 ), .IN1(\b/n2462 ), .SEL(msg[29]), .F(
        \b/n2467 ) );
  MUX \b/U2478  ( .IN0(\b/n2465 ), .IN1(\b/n2464 ), .SEL(msg[26]), .F(
        \b/n2466 ) );
  MUX \b/U2477  ( .IN0(\b/n2233 ), .IN1(\b/n915 ), .SEL(msg[31]), .F(\b/n2465 ) );
  MUX \b/U2476  ( .IN0(\b/n2258 ), .IN1(\b/n2463 ), .SEL(msg[31]), .F(
        \b/n2464 ) );
  MUX \b/U2475  ( .IN0(\b/n911 ), .IN1(\b/n892 ), .SEL(msg[25]), .F(\b/n2463 )
         );
  MUX \b/U2474  ( .IN0(\b/n2461 ), .IN1(\b/n2460 ), .SEL(msg[26]), .F(
        \b/n2462 ) );
  MUX \b/U2473  ( .IN0(\b/n909 ), .IN1(n629), .SEL(msg[31]), .F(\b/n2461 ) );
  MUX \b/U2472  ( .IN0(\b/n2459 ), .IN1(\b/n2458 ), .SEL(msg[31]), .F(
        \b/n2460 ) );
  AND \b/U2471  ( .A(\b/n2218 ), .B(\b/n2293 ), .Z(\b/n2459 ) );
  MUX \b/U2470  ( .IN0(\b/n881 ), .IN1(\b/n865 ), .SEL(msg[25]), .F(\b/n2458 )
         );
  MUX \b/U2469  ( .IN0(\b/n2456 ), .IN1(\b/n2447 ), .SEL(msg[24]), .F(
        \b/n2457 ) );
  MUX \b/U2468  ( .IN0(\b/n2455 ), .IN1(\b/n2451 ), .SEL(msg[29]), .F(
        \b/n2456 ) );
  MUX \b/U2467  ( .IN0(\b/n2454 ), .IN1(\b/n2452 ), .SEL(msg[26]), .F(
        \b/n2455 ) );
  MUX \b/U2466  ( .IN0(\b/n2224 ), .IN1(\b/n2453 ), .SEL(msg[31]), .F(
        \b/n2454 ) );
  NAND \b/U2465  ( .A(msg[25]), .B(\b/n881 ), .Z(\b/n2453 ) );
  MUX \b/U2464  ( .IN0(\b/n865 ), .IN1(\b/n918 ), .SEL(msg[31]), .F(\b/n2452 )
         );
  MUX \b/U2463  ( .IN0(\b/n2450 ), .IN1(\b/n2449 ), .SEL(msg[26]), .F(
        \b/n2451 ) );
  MUX \b/U2462  ( .IN0(\b/n2250 ), .IN1(\b/n883 ), .SEL(msg[31]), .F(\b/n2450 ) );
  MUX \b/U2461  ( .IN0(\b/n2448 ), .IN1(\b/n2213 ), .SEL(n628), .F(\b/n2449 )
         );
  AND \b/U2460  ( .A(msg[31]), .B(msg[27]), .Z(\b/n2448 ) );
  MUX \b/U2459  ( .IN0(\b/n2446 ), .IN1(\b/n2443 ), .SEL(msg[29]), .F(
        \b/n2447 ) );
  MUX \b/U2458  ( .IN0(\b/n2445 ), .IN1(\b/n2444 ), .SEL(msg[26]), .F(
        \b/n2446 ) );
  MUX \b/U2457  ( .IN0(\b/n2374 ), .IN1(\b/n2213 ), .SEL(msg[31]), .F(
        \b/n2445 ) );
  MUX \b/U2456  ( .IN0(n627), .IN1(\b/n916 ), .SEL(msg[31]), .F(\b/n2444 ) );
  MUX \b/U2455  ( .IN0(\b/n2441 ), .IN1(\b/n2440 ), .SEL(msg[26]), .F(
        \b/n2443 ) );
  AND \b/U2454  ( .A(\b/n2442 ), .B(\b/n2342 ), .Z(\b/n2441 ) );
  MUX \b/U2453  ( .IN0(\b/n867 ), .IN1(\b/n911 ), .SEL(msg[31]), .F(\b/n2440 )
         );
  MUX \b/U2452  ( .IN0(\b/n2439 ), .IN1(\b/n2422 ), .SEL(msg[30]), .F(
        shift_row_out[60]) );
  MUX \b/U2451  ( .IN0(\b/n2438 ), .IN1(\b/n2430 ), .SEL(msg[24]), .F(
        \b/n2439 ) );
  MUX \b/U2450  ( .IN0(\b/n2437 ), .IN1(\b/n2434 ), .SEL(msg[29]), .F(
        \b/n2438 ) );
  MUX \b/U2449  ( .IN0(\b/n2436 ), .IN1(\b/n2435 ), .SEL(msg[26]), .F(
        \b/n2437 ) );
  MUX \b/U2448  ( .IN0(\b/n893 ), .IN1(\b/n914 ), .SEL(msg[31]), .F(\b/n2436 )
         );
  MUX \b/U2447  ( .IN0(\b/n2293 ), .IN1(\b/n2258 ), .SEL(msg[31]), .F(
        \b/n2435 ) );
  NAND \b/U2446  ( .A(msg[25]), .B(\b/n2212 ), .Z(\b/n2293 ) );
  MUX \b/U2445  ( .IN0(\b/n2431 ), .IN1(\b/n2432 ), .SEL(msg[26]), .F(
        \b/n2434 ) );
  AND \b/U2444  ( .A(\b/n2243 ), .B(\b/n2433 ), .Z(\b/n2432 ) );
  MUX \b/U2443  ( .IN0(\b/n2241 ), .IN1(\b/n896 ), .SEL(msg[31]), .F(\b/n2431 ) );
  MUX \b/U2442  ( .IN0(\b/n2429 ), .IN1(\b/n2426 ), .SEL(msg[29]), .F(
        \b/n2430 ) );
  MUX \b/U2441  ( .IN0(\b/n2428 ), .IN1(\b/n2427 ), .SEL(msg[26]), .F(
        \b/n2429 ) );
  MUX \b/U2440  ( .IN0(\b/n858 ), .IN1(\b/n904 ), .SEL(msg[31]), .F(\b/n2428 )
         );
  MUX \b/U2439  ( .IN0(\b/n865 ), .IN1(\b/n2221 ), .SEL(msg[31]), .F(\b/n2427 ) );
  MUX \b/U2438  ( .IN0(\b/n2425 ), .IN1(\b/n2423 ), .SEL(msg[26]), .F(
        \b/n2426 ) );
  MUX \b/U2437  ( .IN0(\b/n2237 ), .IN1(\b/n2424 ), .SEL(msg[31]), .F(
        \b/n2425 ) );
  AND \b/U2436  ( .A(\b/n2221 ), .B(\b/n922 ), .Z(\b/n2424 ) );
  MUX \b/U2435  ( .IN0(\b/n880 ), .IN1(\b/n899 ), .SEL(msg[31]), .F(\b/n2423 )
         );
  MUX \b/U2434  ( .IN0(\b/n2421 ), .IN1(\b/n2415 ), .SEL(msg[24]), .F(
        \b/n2422 ) );
  MUX \b/U2433  ( .IN0(\b/n2420 ), .IN1(\b/n2418 ), .SEL(msg[29]), .F(
        \b/n2421 ) );
  MUX \b/U2432  ( .IN0(\b/n2419 ), .IN1(\b/n2215 ), .SEL(msg[26]), .F(
        \b/n2420 ) );
  MUX \b/U2431  ( .IN0(\b/n2235 ), .IN1(\b/n901 ), .SEL(msg[31]), .F(\b/n2419 ) );
  MUX \b/U2430  ( .IN0(\b/n2417 ), .IN1(\b/n2416 ), .SEL(msg[26]), .F(
        \b/n2418 ) );
  MUX \b/U2429  ( .IN0(n626), .IN1(\b/n893 ), .SEL(msg[31]), .F(\b/n2417 ) );
  MUX \b/U2428  ( .IN0(\b/n2245 ), .IN1(\b/n2248 ), .SEL(msg[31]), .F(
        \b/n2416 ) );
  MUX \b/U2427  ( .IN0(\b/n2414 ), .IN1(\b/n2411 ), .SEL(msg[29]), .F(
        \b/n2415 ) );
  MUX \b/U2426  ( .IN0(\b/n2413 ), .IN1(\b/n2412 ), .SEL(msg[26]), .F(
        \b/n2414 ) );
  MUX \b/U2425  ( .IN0(\b/n866 ), .IN1(\b/n2217 ), .SEL(msg[31]), .F(\b/n2413 ) );
  MUX \b/U2424  ( .IN0(\b/n911 ), .IN1(\b/n2239 ), .SEL(msg[31]), .F(\b/n2412 ) );
  MUX \b/U2423  ( .IN0(\b/n854 ), .IN1(\b/n2410 ), .SEL(msg[26]), .F(\b/n2411 ) );
  MUX \b/U2422  ( .IN0(\b/n874 ), .IN1(\b/n2221 ), .SEL(msg[31]), .F(\b/n2410 ) );
  MUX \b/U2421  ( .IN0(\b/n2409 ), .IN1(\b/n2390 ), .SEL(msg[30]), .F(
        shift_row_out[59]) );
  MUX \b/U2420  ( .IN0(\b/n2408 ), .IN1(\b/n2400 ), .SEL(msg[24]), .F(
        \b/n2409 ) );
  MUX \b/U2419  ( .IN0(\b/n2407 ), .IN1(\b/n2404 ), .SEL(msg[29]), .F(
        \b/n2408 ) );
  MUX \b/U2418  ( .IN0(\b/n2406 ), .IN1(\b/n2405 ), .SEL(msg[31]), .F(
        \b/n2407 ) );
  MUX \b/U2417  ( .IN0(\b/n2229 ), .IN1(\b/n899 ), .SEL(msg[26]), .F(\b/n2406 ) );
  MUX \b/U2416  ( .IN0(n629), .IN1(\b/n857 ), .SEL(msg[26]), .F(\b/n2405 ) );
  MUX \b/U2415  ( .IN0(\b/n2402 ), .IN1(\b/n2401 ), .SEL(msg[31]), .F(
        \b/n2404 ) );
  AND \b/U2414  ( .A(\b/n2403 ), .B(msg[28]), .Z(\b/n2402 ) );
  MUX \b/U2413  ( .IN0(\b/n887 ), .IN1(\b/n2242 ), .SEL(msg[26]), .F(\b/n2401 ) );
  MUX \b/U2412  ( .IN0(\b/n2399 ), .IN1(\b/n2396 ), .SEL(msg[29]), .F(
        \b/n2400 ) );
  MUX \b/U2411  ( .IN0(\b/n2398 ), .IN1(\b/n2397 ), .SEL(msg[31]), .F(
        \b/n2399 ) );
  MUX \b/U2410  ( .IN0(\b/n2233 ), .IN1(n625), .SEL(msg[26]), .F(\b/n2398 ) );
  MUX \b/U2409  ( .IN0(\b/n855 ), .IN1(\b/n874 ), .SEL(msg[26]), .F(\b/n2397 )
         );
  MUX \b/U2408  ( .IN0(\b/n2392 ), .IN1(\b/n2393 ), .SEL(msg[31]), .F(
        \b/n2396 ) );
  NAND \b/U2407  ( .A(\b/n2394 ), .B(\b/n2395 ), .Z(\b/n2393 ) );
  MUX \b/U2406  ( .IN0(\b/n900 ), .IN1(\b/n2391 ), .SEL(msg[26]), .F(\b/n2392 ) );
  MUX \b/U2405  ( .IN0(\b/n875 ), .IN1(\b/n917 ), .SEL(msg[25]), .F(\b/n2391 )
         );
  MUX \b/U2404  ( .IN0(\b/n2389 ), .IN1(\b/n2380 ), .SEL(msg[24]), .F(
        \b/n2390 ) );
  MUX \b/U2403  ( .IN0(\b/n2388 ), .IN1(\b/n2384 ), .SEL(msg[29]), .F(
        \b/n2389 ) );
  MUX \b/U2402  ( .IN0(\b/n2386 ), .IN1(\b/n2385 ), .SEL(msg[31]), .F(
        \b/n2388 ) );
  NAND \b/U2401  ( .A(\b/n865 ), .B(\b/n2387 ), .Z(\b/n2386 ) );
  MUX \b/U2400  ( .IN0(\b/n916 ), .IN1(\b/n878 ), .SEL(msg[26]), .F(\b/n2385 )
         );
  MUX \b/U2399  ( .IN0(\b/n2383 ), .IN1(\b/n2381 ), .SEL(msg[31]), .F(
        \b/n2384 ) );
  MUX \b/U2398  ( .IN0(\b/n2224 ), .IN1(\b/n2382 ), .SEL(msg[26]), .F(
        \b/n2383 ) );
  AND \b/U2397  ( .A(msg[25]), .B(\b/n865 ), .Z(\b/n2382 ) );
  MUX \b/U2396  ( .IN0(\b/n870 ), .IN1(\b/n2243 ), .SEL(msg[26]), .F(\b/n2381 ) );
  MUX \b/U2395  ( .IN0(\b/n2379 ), .IN1(\b/n2373 ), .SEL(msg[29]), .F(
        \b/n2380 ) );
  MUX \b/U2394  ( .IN0(\b/n2378 ), .IN1(\b/n2376 ), .SEL(msg[31]), .F(
        \b/n2379 ) );
  MUX \b/U2393  ( .IN0(\b/n2377 ), .IN1(\b/n2213 ), .SEL(\b/n2261 ), .F(
        \b/n2378 ) );
  MUX \b/U2392  ( .IN0(msg[27]), .IN1(msg[28]), .SEL(msg[26]), .F(\b/n2377 )
         );
  MUX \b/U2391  ( .IN0(\b/n2243 ), .IN1(\b/n2374 ), .SEL(msg[26]), .F(
        \b/n2376 ) );
  NAND \b/U2390  ( .A(\b/n2213 ), .B(\b/n2375 ), .Z(\b/n2374 ) );
  MUX \b/U2389  ( .IN0(\b/n2370 ), .IN1(\b/n2371 ), .SEL(msg[31]), .F(
        \b/n2373 ) );
  AND \b/U2388  ( .A(\b/n898 ), .B(\b/n2372 ), .Z(\b/n2371 ) );
  MUX \b/U2387  ( .IN0(\b/n879 ), .IN1(\b/n2214 ), .SEL(msg[26]), .F(\b/n2370 ) );
  MUX \b/U2386  ( .IN0(\b/n2369 ), .IN1(\b/n2353 ), .SEL(msg[30]), .F(
        shift_row_out[58]) );
  MUX \b/U2385  ( .IN0(\b/n2368 ), .IN1(\b/n2360 ), .SEL(msg[24]), .F(
        \b/n2369 ) );
  MUX \b/U2384  ( .IN0(\b/n2367 ), .IN1(\b/n2363 ), .SEL(msg[29]), .F(
        \b/n2368 ) );
  MUX \b/U2383  ( .IN0(\b/n2366 ), .IN1(\b/n2364 ), .SEL(msg[26]), .F(
        \b/n2367 ) );
  MUX \b/U2382  ( .IN0(\b/n887 ), .IN1(\b/n2365 ), .SEL(msg[31]), .F(\b/n2366 ) );
  MUX \b/U2381  ( .IN0(\b/n2221 ), .IN1(\b/n865 ), .SEL(msg[25]), .F(\b/n2365 ) );
  MUX \b/U2380  ( .IN0(\b/n2260 ), .IN1(\b/n905 ), .SEL(msg[31]), .F(\b/n2364 ) );
  MUX \b/U2379  ( .IN0(\b/n2362 ), .IN1(\b/n2361 ), .SEL(msg[26]), .F(
        \b/n2363 ) );
  MUX \b/U2378  ( .IN0(\b/n2214 ), .IN1(\b/n872 ), .SEL(msg[31]), .F(\b/n2362 ) );
  MUX \b/U2377  ( .IN0(\b/n908 ), .IN1(\b/n2247 ), .SEL(msg[31]), .F(\b/n2361 ) );
  MUX \b/U2376  ( .IN0(\b/n2359 ), .IN1(\b/n2355 ), .SEL(msg[29]), .F(
        \b/n2360 ) );
  MUX \b/U2375  ( .IN0(\b/n2356 ), .IN1(\b/n854 ), .SEL(msg[26]), .F(\b/n2359 ) );
  NAND \b/U2374  ( .A(\b/n2357 ), .B(\b/n2358 ), .Z(\b/n2356 ) );
  MUX \b/U2373  ( .IN0(n627), .IN1(\b/n2354 ), .SEL(\b/n2259 ), .F(\b/n2355 )
         );
  MUX \b/U2372  ( .IN0(\b/n886 ), .IN1(\b/n2226 ), .SEL(msg[26]), .F(\b/n2354 ) );
  MUX \b/U2371  ( .IN0(\b/n2352 ), .IN1(\b/n2344 ), .SEL(msg[24]), .F(
        \b/n2353 ) );
  MUX \b/U2370  ( .IN0(\b/n2351 ), .IN1(\b/n2348 ), .SEL(msg[29]), .F(
        \b/n2352 ) );
  MUX \b/U2369  ( .IN0(\b/n2350 ), .IN1(\b/n2349 ), .SEL(msg[26]), .F(
        \b/n2351 ) );
  MUX \b/U2368  ( .IN0(\b/n914 ), .IN1(msg[25]), .SEL(msg[31]), .F(\b/n2350 )
         );
  MUX \b/U2367  ( .IN0(n630), .IN1(\b/n2227 ), .SEL(msg[31]), .F(\b/n2349 ) );
  MUX \b/U2366  ( .IN0(\b/n2347 ), .IN1(\b/n2346 ), .SEL(msg[26]), .F(
        \b/n2348 ) );
  MUX \b/U2365  ( .IN0(\b/n919 ), .IN1(\b/n913 ), .SEL(msg[31]), .F(\b/n2347 )
         );
  MUX \b/U2364  ( .IN0(n630), .IN1(\b/n2345 ), .SEL(msg[31]), .F(\b/n2346 ) );
  MUX \b/U2363  ( .IN0(\b/n865 ), .IN1(\b/n902 ), .SEL(msg[25]), .F(\b/n2345 )
         );
  MUX \b/U2362  ( .IN0(\b/n2343 ), .IN1(\b/n2337 ), .SEL(msg[29]), .F(
        \b/n2344 ) );
  MUX \b/U2361  ( .IN0(\b/n2340 ), .IN1(\b/n2339 ), .SEL(msg[26]), .F(
        \b/n2343 ) );
  NAND \b/U2360  ( .A(\b/n2341 ), .B(\b/n2342 ), .Z(\b/n2340 ) );
  MUX \b/U2359  ( .IN0(\b/n2213 ), .IN1(\b/n2338 ), .SEL(n628), .F(\b/n2339 )
         );
  MUX \b/U2358  ( .IN0(msg[27]), .IN1(\b/n875 ), .SEL(msg[31]), .F(\b/n2338 )
         );
  MUX \b/U2357  ( .IN0(\b/n2336 ), .IN1(\b/n2335 ), .SEL(msg[26]), .F(
        \b/n2337 ) );
  MUX \b/U2356  ( .IN0(\b/n2258 ), .IN1(\b/n873 ), .SEL(msg[31]), .F(\b/n2336 ) );
  MUX \b/U2355  ( .IN0(\b/n2254 ), .IN1(\b/n2334 ), .SEL(msg[31]), .F(
        \b/n2335 ) );
  MUX \b/U2354  ( .IN0(\b/n2216 ), .IN1(\b/n2221 ), .SEL(msg[25]), .F(
        \b/n2334 ) );
  MUX \b/U2353  ( .IN0(\b/n2333 ), .IN1(\b/n2315 ), .SEL(msg[30]), .F(
        shift_row_out[57]) );
  MUX \b/U2352  ( .IN0(\b/n2332 ), .IN1(\b/n2323 ), .SEL(msg[24]), .F(
        \b/n2333 ) );
  MUX \b/U2351  ( .IN0(\b/n2331 ), .IN1(\b/n2327 ), .SEL(msg[29]), .F(
        \b/n2332 ) );
  MUX \b/U2350  ( .IN0(\b/n2330 ), .IN1(\b/n2329 ), .SEL(msg[26]), .F(
        \b/n2331 ) );
  MUX \b/U2349  ( .IN0(\b/n910 ), .IN1(n632), .SEL(msg[31]), .F(\b/n2330 ) );
  MUX \b/U2348  ( .IN0(\b/n2328 ), .IN1(n626), .SEL(msg[31]), .F(\b/n2329 ) );
  NAND \b/U2347  ( .A(\b/n922 ), .B(\b/n881 ), .Z(\b/n2328 ) );
  MUX \b/U2346  ( .IN0(\b/n2326 ), .IN1(\b/n2325 ), .SEL(msg[26]), .F(
        \b/n2327 ) );
  MUX \b/U2345  ( .IN0(\b/n858 ), .IN1(\b/n2228 ), .SEL(msg[31]), .F(\b/n2326 ) );
  MUX \b/U2344  ( .IN0(\b/n2218 ), .IN1(\b/n2324 ), .SEL(msg[31]), .F(
        \b/n2325 ) );
  AND \b/U2343  ( .A(msg[25]), .B(msg[28]), .Z(\b/n2324 ) );
  MUX \b/U2342  ( .IN0(\b/n2322 ), .IN1(\b/n2319 ), .SEL(msg[29]), .F(
        \b/n2323 ) );
  MUX \b/U2341  ( .IN0(\b/n2321 ), .IN1(\b/n2320 ), .SEL(msg[26]), .F(
        \b/n2322 ) );
  MUX \b/U2340  ( .IN0(\b/n2257 ), .IN1(\b/n919 ), .SEL(msg[31]), .F(\b/n2321 ) );
  MUX \b/U2339  ( .IN0(\b/n894 ), .IN1(\b/n2226 ), .SEL(msg[31]), .F(\b/n2320 ) );
  MUX \b/U2338  ( .IN0(\b/n2316 ), .IN1(\b/n2317 ), .SEL(msg[26]), .F(
        \b/n2319 ) );
  AND \b/U2337  ( .A(\b/n2318 ), .B(\b/n2273 ), .Z(\b/n2317 ) );
  MUX \b/U2336  ( .IN0(\b/n2232 ), .IN1(\b/n2221 ), .SEL(msg[31]), .F(
        \b/n2316 ) );
  MUX \b/U2335  ( .IN0(\b/n2314 ), .IN1(\b/n2306 ), .SEL(msg[24]), .F(
        \b/n2315 ) );
  MUX \b/U2334  ( .IN0(\b/n2313 ), .IN1(\b/n2309 ), .SEL(msg[29]), .F(
        \b/n2314 ) );
  MUX \b/U2333  ( .IN0(\b/n2312 ), .IN1(\b/n2311 ), .SEL(msg[26]), .F(
        \b/n2313 ) );
  MUX \b/U2332  ( .IN0(\b/n2220 ), .IN1(\b/n883 ), .SEL(msg[31]), .F(\b/n2312 ) );
  MUX \b/U2331  ( .IN0(\b/n2310 ), .IN1(\b/n867 ), .SEL(msg[31]), .F(\b/n2311 ) );
  MUX \b/U2330  ( .IN0(\b/n2218 ), .IN1(\b/n875 ), .SEL(msg[25]), .F(\b/n2310 ) );
  MUX \b/U2329  ( .IN0(\b/n2308 ), .IN1(\b/n2307 ), .SEL(msg[26]), .F(
        \b/n2309 ) );
  MUX \b/U2328  ( .IN0(\b/n914 ), .IN1(\b/n892 ), .SEL(msg[31]), .F(\b/n2308 )
         );
  MUX \b/U2327  ( .IN0(\b/n910 ), .IN1(\b/n870 ), .SEL(msg[31]), .F(\b/n2307 )
         );
  MUX \b/U2326  ( .IN0(\b/n2305 ), .IN1(\b/n2300 ), .SEL(msg[29]), .F(
        \b/n2306 ) );
  MUX \b/U2325  ( .IN0(\b/n2304 ), .IN1(\b/n2301 ), .SEL(msg[26]), .F(
        \b/n2305 ) );
  MUX \b/U2324  ( .IN0(\b/n2302 ), .IN1(\b/n2303 ), .SEL(msg[31]), .F(
        \b/n2304 ) );
  NAND \b/U2323  ( .A(\b/n2221 ), .B(\b/n2293 ), .Z(\b/n2303 ) );
  MUX \b/U2322  ( .IN0(\b/n2221 ), .IN1(\b/n875 ), .SEL(msg[25]), .F(\b/n2302 ) );
  MUX \b/U2321  ( .IN0(\b/n2238 ), .IN1(\b/n2236 ), .SEL(msg[31]), .F(
        \b/n2301 ) );
  MUX \b/U2320  ( .IN0(\b/n2256 ), .IN1(\b/n2299 ), .SEL(msg[26]), .F(
        \b/n2300 ) );
  MUX \b/U2319  ( .IN0(\b/n881 ), .IN1(\b/n913 ), .SEL(msg[31]), .F(\b/n2299 )
         );
  MUX \b/U2318  ( .IN0(\b/n2298 ), .IN1(\b/n2281 ), .SEL(msg[30]), .F(
        shift_row_out[56]) );
  MUX \b/U2317  ( .IN0(\b/n2297 ), .IN1(\b/n2289 ), .SEL(msg[24]), .F(
        \b/n2298 ) );
  MUX \b/U2316  ( .IN0(\b/n2296 ), .IN1(\b/n2294 ), .SEL(msg[26]), .F(
        \b/n2297 ) );
  MUX \b/U2315  ( .IN0(\b/n855 ), .IN1(\b/n2295 ), .SEL(msg[31]), .F(\b/n2296 ) );
  MUX \b/U2314  ( .IN0(\b/n908 ), .IN1(\b/n911 ), .SEL(msg[29]), .F(\b/n2295 )
         );
  MUX \b/U2313  ( .IN0(\b/n2291 ), .IN1(\b/n2290 ), .SEL(msg[31]), .F(
        \b/n2294 ) );
  NAND \b/U2312  ( .A(\b/n2292 ), .B(\b/n2293 ), .Z(\b/n2291 ) );
  MUX \b/U2311  ( .IN0(\b/n907 ), .IN1(\b/n922 ), .SEL(msg[29]), .F(\b/n2290 )
         );
  MUX \b/U2310  ( .IN0(\b/n2288 ), .IN1(\b/n2284 ), .SEL(msg[26]), .F(
        \b/n2289 ) );
  MUX \b/U2309  ( .IN0(\b/n2287 ), .IN1(\b/n2285 ), .SEL(msg[31]), .F(
        \b/n2288 ) );
  MUX \b/U2308  ( .IN0(\b/n2286 ), .IN1(\b/n860 ), .SEL(msg[29]), .F(\b/n2287 ) );
  NAND \b/U2307  ( .A(\b/n922 ), .B(\b/n2213 ), .Z(\b/n2286 ) );
  MUX \b/U2305  ( .IN0(\b/n2283 ), .IN1(\b/n2282 ), .SEL(msg[31]), .F(
        \b/n2284 ) );
  MUX \b/U2304  ( .IN0(n627), .IN1(\b/n857 ), .SEL(msg[29]), .F(\b/n2283 ) );
  MUX \b/U2303  ( .IN0(\b/n909 ), .IN1(\b/n865 ), .SEL(msg[29]), .F(\b/n2282 )
         );
  MUX \b/U2302  ( .IN0(\b/n2280 ), .IN1(\b/n2270 ), .SEL(msg[24]), .F(
        \b/n2281 ) );
  MUX \b/U2301  ( .IN0(\b/n2279 ), .IN1(\b/n2275 ), .SEL(msg[26]), .F(
        \b/n2280 ) );
  MUX \b/U2300  ( .IN0(\b/n2278 ), .IN1(\b/n2277 ), .SEL(msg[31]), .F(
        \b/n2279 ) );
  MUX \b/U2299  ( .IN0(n625), .IN1(\b/n861 ), .SEL(msg[29]), .F(\b/n2278 ) );
  MUX \b/U2298  ( .IN0(\b/n2276 ), .IN1(\b/n898 ), .SEL(msg[29]), .F(\b/n2277 ) );
  NAND \b/U2297  ( .A(\b/n2212 ), .B(\b/n2214 ), .Z(\b/n2276 ) );
  MUX \b/U2296  ( .IN0(\b/n2274 ), .IN1(\b/n2271 ), .SEL(msg[31]), .F(
        \b/n2275 ) );
  MUX \b/U2295  ( .IN0(\b/n868 ), .IN1(\b/n2272 ), .SEL(msg[29]), .F(\b/n2274 ) );
  NAND \b/U2294  ( .A(\b/n2216 ), .B(\b/n2273 ), .Z(\b/n2272 ) );
  MUX \b/U2293  ( .IN0(\b/n2231 ), .IN1(\b/n2222 ), .SEL(msg[29]), .F(
        \b/n2271 ) );
  MUX \b/U2292  ( .IN0(\b/n2269 ), .IN1(\b/n2265 ), .SEL(msg[26]), .F(
        \b/n2270 ) );
  MUX \b/U2291  ( .IN0(\b/n2267 ), .IN1(\b/n2266 ), .SEL(msg[31]), .F(
        \b/n2269 ) );
  NAND \b/U2290  ( .A(\b/n2268 ), .B(\b/n2255 ), .Z(\b/n2267 ) );
  MUX \b/U2289  ( .IN0(msg[27]), .IN1(\b/n2247 ), .SEL(msg[29]), .F(\b/n2266 )
         );
  MUX \b/U2288  ( .IN0(\b/n2264 ), .IN1(\b/n2263 ), .SEL(msg[31]), .F(
        \b/n2265 ) );
  MUX \b/U2287  ( .IN0(\b/n873 ), .IN1(\b/n889 ), .SEL(msg[29]), .F(\b/n2264 )
         );
  MUX \b/U2286  ( .IN0(\b/n906 ), .IN1(\b/n894 ), .SEL(msg[29]), .F(\b/n2263 )
         );
  XOR \b/U2285  ( .A(\b/n2213 ), .B(msg[25]), .Z(\b/n2262 ) );
  XOR \b/U2284  ( .A(msg[25]), .B(msg[26]), .Z(\b/n2261 ) );
  XOR \b/U2283  ( .A(msg[25]), .B(msg[27]), .Z(\b/n2260 ) );
  XOR \b/U2282  ( .A(msg[26]), .B(msg[31]), .Z(\b/n2259 ) );
  XOR \b/U2281  ( .A(\b/n922 ), .B(\b/n865 ), .Z(\b/n2258 ) );
  XOR \b/U2280  ( .A(msg[25]), .B(\b/n911 ), .Z(\b/n2257 ) );
  XOR \b/U2278  ( .A(msg[25]), .B(msg[29]), .Z(\b/n2255 ) );
  NAND \b/U2277  ( .A(msg[25]), .B(msg[27]), .Z(\b/n2254 ) );
  MUX \b/U2276  ( .IN0(\b/n2213 ), .IN1(\b/n865 ), .SEL(msg[25]), .F(\b/n2253 ) );
  MUX \b/U2274  ( .IN0(msg[27]), .IN1(\b/n902 ), .SEL(msg[25]), .F(\b/n2251 )
         );
  MUX \b/U2273  ( .IN0(\b/n881 ), .IN1(\b/n902 ), .SEL(msg[25]), .F(\b/n2250 )
         );
  MUX \b/U2272  ( .IN0(\b/n2216 ), .IN1(\b/n2218 ), .SEL(msg[25]), .F(
        \b/n2249 ) );
  MUX \b/U2271  ( .IN0(msg[28]), .IN1(\b/n881 ), .SEL(msg[25]), .F(\b/n2248 )
         );
  OR \b/U2270  ( .A(msg[25]), .B(msg[28]), .Z(\b/n2247 ) );
  NAND \b/U2268  ( .A(\b/n902 ), .B(\b/n922 ), .Z(\b/n2245 ) );
  MUX \b/U2267  ( .IN0(\b/n902 ), .IN1(msg[28]), .SEL(msg[25]), .F(\b/n2244 )
         );
  MUX \b/U2266  ( .IN0(\b/n2212 ), .IN1(\b/n2221 ), .SEL(msg[25]), .F(
        \b/n2243 ) );
  MUX \b/U2265  ( .IN0(\b/n917 ), .IN1(msg[28]), .SEL(msg[25]), .F(\b/n2242 )
         );
  MUX \b/U2264  ( .IN0(\b/n875 ), .IN1(\b/n902 ), .SEL(msg[25]), .F(\b/n2241 )
         );
  MUX \b/U2263  ( .IN0(\b/n2212 ), .IN1(msg[28]), .SEL(msg[25]), .F(\b/n2240 )
         );
  MUX \b/U2262  ( .IN0(\b/n892 ), .IN1(\b/n881 ), .SEL(msg[25]), .F(\b/n2239 )
         );
  XOR \b/U2261  ( .A(\b/n875 ), .B(msg[25]), .Z(\b/n2238 ) );
  MUX \b/U2260  ( .IN0(\b/n2218 ), .IN1(\b/n892 ), .SEL(msg[25]), .F(\b/n2237 ) );
  NANDN \b/U2259  ( .B(msg[25]), .A(msg[27]), .Z(\b/n2236 ) );
  MUX \b/U2258  ( .IN0(\b/n865 ), .IN1(msg[27]), .SEL(msg[25]), .F(\b/n2235 )
         );
  NAND \b/U2256  ( .A(\b/n2216 ), .B(\b/n922 ), .Z(\b/n2233 ) );
  MUX \b/U2255  ( .IN0(msg[28]), .IN1(\b/n2213 ), .SEL(msg[25]), .F(\b/n2232 )
         );
  MUX \b/U2254  ( .IN0(\b/n892 ), .IN1(msg[27]), .SEL(msg[25]), .F(\b/n2231 )
         );
  MUX \b/U2252  ( .IN0(msg[28]), .IN1(\b/n911 ), .SEL(msg[25]), .F(\b/n2229 )
         );
  MUX \b/U2251  ( .IN0(\b/n865 ), .IN1(\b/n917 ), .SEL(msg[25]), .F(\b/n2228 )
         );
  NAND \b/U2250  ( .A(\b/n2214 ), .B(\b/n865 ), .Z(\b/n2227 ) );
  MUX \b/U2249  ( .IN0(\b/n2213 ), .IN1(\b/n2221 ), .SEL(msg[25]), .F(
        \b/n2226 ) );
  NAND \b/U2248  ( .A(\b/n2225 ), .B(\b/n2212 ), .Z(\b/n2224 ) );
  MUX \b/U2247  ( .IN0(\b/n2216 ), .IN1(\b/n917 ), .SEL(msg[25]), .F(\b/n2223 ) );
  MUX \b/U2246  ( .IN0(\b/n917 ), .IN1(\b/n881 ), .SEL(msg[25]), .F(\b/n2222 )
         );
  NANDN \b/U2245  ( .B(msg[27]), .A(msg[28]), .Z(\b/n2221 ) );
  MUX \b/U2244  ( .IN0(\b/n2216 ), .IN1(msg[27]), .SEL(msg[25]), .F(\b/n2220 )
         );
  OR \b/U2243  ( .A(msg[27]), .B(msg[28]), .Z(\b/n2216 ) );
  MUX \b/U2242  ( .IN0(\b/n865 ), .IN1(\b/n881 ), .SEL(msg[25]), .F(\b/n2219 )
         );
  XOR \b/U2241  ( .A(\b/n875 ), .B(msg[27]), .Z(\b/n2218 ) );
  NANDN \b/U2240  ( .B(msg[27]), .A(msg[25]), .Z(\b/n2217 ) );
  NAND \b/U2239  ( .A(\b/n2216 ), .B(\b/n2214 ), .Z(\b/n2215 ) );
  NAND \b/U2238  ( .A(msg[25]), .B(\b/n2213 ), .Z(\b/n2214 ) );
  NANDN \b/U2237  ( .B(msg[28]), .A(msg[27]), .Z(\b/n2213 ) );
  NAND \b/U2236  ( .A(msg[27]), .B(msg[28]), .Z(\b/n2212 ) );
  MUX \b/U2235  ( .IN0(msg[20]), .IN1(\b/n1853 ), .SEL(msg[17]), .F(\b/n2211 )
         );
  MUX \b/U2234  ( .IN0(msg[20]), .IN1(\b/n1862 ), .SEL(msg[17]), .F(\b/n2210 )
         );
  MUX \b/U2233  ( .IN0(\b/n1854 ), .IN1(\b/n1857 ), .SEL(msg[17]), .F(
        \b/n2209 ) );
  MUX \b/U2232  ( .IN0(\b/n1859 ), .IN1(\b/n982 ), .SEL(msg[17]), .F(\b/n2208 ) );
  MUX \b/U2230  ( .IN0(\b/n1862 ), .IN1(\b/n1853 ), .SEL(msg[18]), .F(
        \b/n2035 ) );
  MUX \b/U2229  ( .IN0(\b/n1855 ), .IN1(\b/n993 ), .SEL(msg[18]), .F(\b/n2036 ) );
  MUX \b/U2228  ( .IN0(\b/n936 ), .IN1(\b/n946 ), .SEL(msg[17]), .F(\b/n1999 )
         );
  MUX \b/U2227  ( .IN0(\b/n1883 ), .IN1(\b/n2194 ), .SEL(msg[23]), .F(
        \b/n2206 ) );
  MUX \b/U2226  ( .IN0(\b/n1857 ), .IN1(\b/n1853 ), .SEL(msg[17]), .F(
        \b/n2197 ) );
  MUX \b/U2225  ( .IN0(\b/n988 ), .IN1(\b/n1859 ), .SEL(msg[17]), .F(\b/n2205 ) );
  MUX \b/U2224  ( .IN0(msg[19]), .IN1(\b/n982 ), .SEL(msg[17]), .F(\b/n2204 )
         );
  MUX \b/U2223  ( .IN0(\b/n1862 ), .IN1(\b/n988 ), .SEL(msg[17]), .F(\b/n2203 ) );
  MUX \b/U2222  ( .IN0(msg[20]), .IN1(\b/n1859 ), .SEL(msg[17]), .F(\b/n2202 )
         );
  MUX \b/U2221  ( .IN0(\b/n973 ), .IN1(\b/n952 ), .SEL(msg[21]), .F(\b/n1909 )
         );
  MUX \b/U2220  ( .IN0(\b/n1854 ), .IN1(\b/n946 ), .SEL(msg[17]), .F(\b/n2201 ) );
  NANDN \b/U2217  ( .B(\b/n1860 ), .A(msg[23]), .Z(\b/n2174 ) );
  NAND \b/U2216  ( .A(msg[23]), .B(\b/n949 ), .Z(\b/n2142 ) );
  NAND \b/U2215  ( .A(msg[23]), .B(\b/n961 ), .Z(\b/n2083 ) );
  NAND \b/U2214  ( .A(msg[23]), .B(\b/n2191 ), .Z(\b/n2116 ) );
  NAND \b/U2213  ( .A(msg[23]), .B(\b/n2111 ), .Z(\b/n2074 ) );
  NAND \b/U2211  ( .A(\b/n993 ), .B(\b/n982 ), .Z(\b/n2195 ) );
  NAND \b/U2210  ( .A(msg[23]), .B(\b/n2193 ), .Z(\b/n2188 ) );
  NAND \b/U2209  ( .A(n624), .B(msg[23]), .Z(\b/n2168 ) );
  NAND \b/U2207  ( .A(msg[18]), .B(\b/n1862 ), .Z(\b/n2028 ) );
  NAND \b/U2206  ( .A(\b/n982 ), .B(msg[17]), .Z(\b/n1983 ) );
  NAND \b/U2205  ( .A(msg[23]), .B(\b/n2197 ), .Z(\b/n1982 ) );
  NAND \b/U2203  ( .A(\b/n2195 ), .B(msg[23]), .Z(\b/n1998 ) );
  NAND \b/U2202  ( .A(\b/n2016 ), .B(\b/n1862 ), .Z(\b/n2194 ) );
  NANDN \b/U2201  ( .B(\b/n936 ), .A(\b/n993 ), .Z(\b/n2193 ) );
  NAND \b/U2199  ( .A(msg[17]), .B(\b/n1862 ), .Z(\b/n1914 ) );
  NAND \b/U2198  ( .A(\b/n936 ), .B(\b/n993 ), .Z(\b/n2191 ) );
  NAND \b/U2195  ( .A(msg[17]), .B(\b/n1857 ), .Z(\b/n2016 ) );
  ANDN \b/U2193  ( .A(msg[18]), .B(msg[17]), .Z(\b/n2044 ) );
  AND \b/U2192  ( .A(\b/n1854 ), .B(\b/n2188 ), .Z(\b/n1959 ) );
  MUX \b/U2191  ( .IN0(\b/n2187 ), .IN1(\b/n2171 ), .SEL(msg[22]), .F(
        shift_row_out[87]) );
  MUX \b/U2190  ( .IN0(\b/n2186 ), .IN1(\b/n2179 ), .SEL(msg[16]), .F(
        \b/n2187 ) );
  MUX \b/U2189  ( .IN0(\b/n2185 ), .IN1(\b/n2182 ), .SEL(msg[21]), .F(
        \b/n2186 ) );
  MUX \b/U2188  ( .IN0(\b/n2184 ), .IN1(\b/n2183 ), .SEL(msg[18]), .F(
        \b/n2185 ) );
  MUX \b/U2187  ( .IN0(msg[20]), .IN1(\b/n953 ), .SEL(msg[23]), .F(\b/n2184 )
         );
  MUX \b/U2186  ( .IN0(\b/n1855 ), .IN1(\b/n957 ), .SEL(msg[23]), .F(\b/n2183 ) );
  MUX \b/U2185  ( .IN0(\b/n2181 ), .IN1(\b/n2180 ), .SEL(msg[18]), .F(
        \b/n2182 ) );
  MUX \b/U2184  ( .IN0(\b/n1913 ), .IN1(\b/n949 ), .SEL(msg[23]), .F(\b/n2181 ) );
  MUX \b/U2183  ( .IN0(\b/n1865 ), .IN1(\b/n1876 ), .SEL(msg[23]), .F(
        \b/n2180 ) );
  MUX \b/U2182  ( .IN0(\b/n2178 ), .IN1(\b/n2175 ), .SEL(msg[21]), .F(
        \b/n2179 ) );
  MUX \b/U2181  ( .IN0(\b/n2177 ), .IN1(\b/n2176 ), .SEL(msg[18]), .F(
        \b/n2178 ) );
  MUX \b/U2180  ( .IN0(\b/n1889 ), .IN1(\b/n1864 ), .SEL(msg[23]), .F(
        \b/n2177 ) );
  MUX \b/U2179  ( .IN0(\b/n961 ), .IN1(\b/n1885 ), .SEL(msg[23]), .F(\b/n2176 ) );
  MUX \b/U2178  ( .IN0(\b/n2173 ), .IN1(\b/n2172 ), .SEL(msg[18]), .F(
        \b/n2175 ) );
  AND \b/U2177  ( .A(\b/n951 ), .B(\b/n2174 ), .Z(\b/n2173 ) );
  MUX \b/U2176  ( .IN0(\b/n1869 ), .IN1(n623), .SEL(msg[23]), .F(\b/n2172 ) );
  MUX \b/U2175  ( .IN0(\b/n2170 ), .IN1(\b/n2162 ), .SEL(msg[16]), .F(
        \b/n2171 ) );
  MUX \b/U2174  ( .IN0(\b/n2169 ), .IN1(\b/n2165 ), .SEL(msg[21]), .F(
        \b/n2170 ) );
  MUX \b/U2173  ( .IN0(\b/n2166 ), .IN1(\b/n2167 ), .SEL(msg[18]), .F(
        \b/n2169 ) );
  NAND \b/U2172  ( .A(\b/n1983 ), .B(\b/n2168 ), .Z(\b/n2167 ) );
  MUX \b/U2171  ( .IN0(\b/n991 ), .IN1(\b/n983 ), .SEL(msg[23]), .F(\b/n2166 )
         );
  MUX \b/U2170  ( .IN0(\b/n2164 ), .IN1(\b/n2163 ), .SEL(msg[18]), .F(
        \b/n2165 ) );
  MUX \b/U2169  ( .IN0(\b/n1859 ), .IN1(\b/n1853 ), .SEL(msg[23]), .F(
        \b/n2164 ) );
  MUX \b/U2168  ( .IN0(\b/n984 ), .IN1(\b/n1890 ), .SEL(msg[23]), .F(\b/n2163 ) );
  MUX \b/U2167  ( .IN0(\b/n2161 ), .IN1(\b/n2158 ), .SEL(msg[21]), .F(
        \b/n2162 ) );
  MUX \b/U2166  ( .IN0(\b/n2160 ), .IN1(\b/n2159 ), .SEL(msg[18]), .F(
        \b/n2161 ) );
  MUX \b/U2165  ( .IN0(\b/n1894 ), .IN1(\b/n1880 ), .SEL(msg[23]), .F(
        \b/n2160 ) );
  MUX \b/U2164  ( .IN0(\b/n937 ), .IN1(\b/n1862 ), .SEL(msg[23]), .F(\b/n2159 ) );
  MUX \b/U2163  ( .IN0(\b/n2157 ), .IN1(\b/n2156 ), .SEL(msg[18]), .F(
        \b/n2158 ) );
  MUX \b/U2162  ( .IN0(\b/n1895 ), .IN1(\b/n1903 ), .SEL(msg[23]), .F(
        \b/n2157 ) );
  MUX \b/U2161  ( .IN0(\b/n1888 ), .IN1(\b/n2155 ), .SEL(msg[23]), .F(
        \b/n2156 ) );
  MUX \b/U2160  ( .IN0(\b/n988 ), .IN1(\b/n946 ), .SEL(msg[17]), .F(\b/n2155 )
         );
  MUX \b/U2159  ( .IN0(\b/n2154 ), .IN1(\b/n2136 ), .SEL(msg[22]), .F(
        shift_row_out[86]) );
  MUX \b/U2158  ( .IN0(\b/n2153 ), .IN1(\b/n2144 ), .SEL(msg[16]), .F(
        \b/n2154 ) );
  MUX \b/U2157  ( .IN0(\b/n2152 ), .IN1(\b/n2147 ), .SEL(msg[21]), .F(
        \b/n2153 ) );
  MUX \b/U2156  ( .IN0(\b/n2151 ), .IN1(\b/n2149 ), .SEL(msg[18]), .F(
        \b/n2152 ) );
  MUX \b/U2155  ( .IN0(\b/n2150 ), .IN1(\b/n1866 ), .SEL(msg[23]), .F(
        \b/n2151 ) );
  MUX \b/U2154  ( .IN0(\b/n988 ), .IN1(\b/n1853 ), .SEL(msg[17]), .F(\b/n2150 ) );
  MUX \b/U2153  ( .IN0(\b/n2148 ), .IN1(\b/n976 ), .SEL(msg[23]), .F(\b/n2149 ) );
  MUX \b/U2152  ( .IN0(\b/n1853 ), .IN1(\b/n1854 ), .SEL(msg[17]), .F(
        \b/n2148 ) );
  MUX \b/U2151  ( .IN0(\b/n2146 ), .IN1(\b/n2145 ), .SEL(msg[18]), .F(
        \b/n2147 ) );
  MUX \b/U2150  ( .IN0(n622), .IN1(\b/n1934 ), .SEL(msg[23]), .F(\b/n2146 ) );
  MUX \b/U2149  ( .IN0(\b/n1892 ), .IN1(\b/n1899 ), .SEL(msg[23]), .F(
        \b/n2145 ) );
  MUX \b/U2148  ( .IN0(\b/n2143 ), .IN1(\b/n2139 ), .SEL(msg[21]), .F(
        \b/n2144 ) );
  MUX \b/U2147  ( .IN0(\b/n2141 ), .IN1(\b/n2140 ), .SEL(msg[18]), .F(
        \b/n2143 ) );
  AND \b/U2146  ( .A(\b/n929 ), .B(\b/n2142 ), .Z(\b/n2141 ) );
  MUX \b/U2145  ( .IN0(\b/n1969 ), .IN1(msg[19]), .SEL(msg[23]), .F(\b/n2140 )
         );
  MUX \b/U2144  ( .IN0(\b/n2138 ), .IN1(\b/n2137 ), .SEL(msg[18]), .F(
        \b/n2139 ) );
  MUX \b/U2143  ( .IN0(\b/n972 ), .IN1(\b/n1857 ), .SEL(msg[23]), .F(\b/n2138 ) );
  MUX \b/U2141  ( .IN0(\b/n2135 ), .IN1(\b/n2128 ), .SEL(msg[16]), .F(
        \b/n2136 ) );
  MUX \b/U2140  ( .IN0(\b/n2134 ), .IN1(\b/n2131 ), .SEL(msg[21]), .F(
        \b/n2135 ) );
  MUX \b/U2139  ( .IN0(\b/n2133 ), .IN1(\b/n2132 ), .SEL(msg[18]), .F(
        \b/n2134 ) );
  MUX \b/U2138  ( .IN0(\b/n968 ), .IN1(\b/n1861 ), .SEL(msg[23]), .F(\b/n2133 ) );
  MUX \b/U2137  ( .IN0(\b/n1865 ), .IN1(n623), .SEL(msg[23]), .F(\b/n2132 ) );
  MUX \b/U2136  ( .IN0(\b/n2130 ), .IN1(\b/n2129 ), .SEL(msg[18]), .F(
        \b/n2131 ) );
  MUX \b/U2135  ( .IN0(\b/n1881 ), .IN1(\b/n933 ), .SEL(msg[23]), .F(\b/n2130 ) );
  MUX \b/U2134  ( .IN0(\b/n953 ), .IN1(\b/n983 ), .SEL(msg[23]), .F(\b/n2129 )
         );
  MUX \b/U2133  ( .IN0(\b/n2127 ), .IN1(\b/n2123 ), .SEL(msg[21]), .F(
        \b/n2128 ) );
  MUX \b/U2132  ( .IN0(\b/n2126 ), .IN1(\b/n2125 ), .SEL(msg[18]), .F(
        \b/n2127 ) );
  MUX \b/U2131  ( .IN0(\b/n1870 ), .IN1(\b/n983 ), .SEL(msg[23]), .F(\b/n2126 ) );
  MUX \b/U2130  ( .IN0(\b/n2124 ), .IN1(\b/n1891 ), .SEL(msg[23]), .F(
        \b/n2125 ) );
  NANDN \b/U2129  ( .B(msg[20]), .A(msg[17]), .Z(\b/n2124 ) );
  MUX \b/U2128  ( .IN0(\b/n2122 ), .IN1(\b/n2120 ), .SEL(msg[18]), .F(
        \b/n2123 ) );
  MUX \b/U2127  ( .IN0(\b/n946 ), .IN1(\b/n2121 ), .SEL(msg[23]), .F(\b/n2122 ) );
  MUX \b/U2126  ( .IN0(\b/n973 ), .IN1(\b/n963 ), .SEL(msg[17]), .F(\b/n2121 )
         );
  MUX \b/U2125  ( .IN0(\b/n935 ), .IN1(\b/n1866 ), .SEL(msg[23]), .F(\b/n2120 ) );
  NANDN \b/U2124  ( .B(\b/n936 ), .A(msg[17]), .Z(\b/n1866 ) );
  MUX \b/U2123  ( .IN0(\b/n2119 ), .IN1(\b/n2098 ), .SEL(msg[22]), .F(
        shift_row_out[85]) );
  MUX \b/U2122  ( .IN0(\b/n2118 ), .IN1(\b/n2108 ), .SEL(msg[16]), .F(
        \b/n2119 ) );
  MUX \b/U2121  ( .IN0(\b/n2117 ), .IN1(\b/n2113 ), .SEL(msg[21]), .F(
        \b/n2118 ) );
  MUX \b/U2120  ( .IN0(\b/n2114 ), .IN1(\b/n2115 ), .SEL(msg[18]), .F(
        \b/n2117 ) );
  AND \b/U2119  ( .A(\b/n1884 ), .B(\b/n2116 ), .Z(\b/n2115 ) );
  MUX \b/U2118  ( .IN0(\b/n1862 ), .IN1(\b/n984 ), .SEL(msg[23]), .F(\b/n2114 ) );
  MUX \b/U2117  ( .IN0(\b/n2112 ), .IN1(\b/n2110 ), .SEL(msg[18]), .F(
        \b/n2113 ) );
  MUX \b/U2116  ( .IN0(\b/n939 ), .IN1(\b/n2111 ), .SEL(msg[23]), .F(\b/n2112 ) );
  NAND \b/U2115  ( .A(\b/n963 ), .B(\b/n993 ), .Z(\b/n2111 ) );
  MUX \b/U2114  ( .IN0(\b/n1862 ), .IN1(\b/n2109 ), .SEL(msg[23]), .F(
        \b/n2110 ) );
  NAND \b/U2113  ( .A(\b/n1853 ), .B(\b/n1914 ), .Z(\b/n2109 ) );
  MUX \b/U2112  ( .IN0(\b/n2107 ), .IN1(\b/n2103 ), .SEL(msg[21]), .F(
        \b/n2108 ) );
  MUX \b/U2111  ( .IN0(\b/n2106 ), .IN1(\b/n2105 ), .SEL(msg[18]), .F(
        \b/n2107 ) );
  MUX \b/U2110  ( .IN0(\b/n1874 ), .IN1(\b/n986 ), .SEL(msg[23]), .F(\b/n2106 ) );
  MUX \b/U2109  ( .IN0(\b/n1899 ), .IN1(\b/n2104 ), .SEL(msg[23]), .F(
        \b/n2105 ) );
  MUX \b/U2108  ( .IN0(\b/n982 ), .IN1(\b/n963 ), .SEL(msg[17]), .F(\b/n2104 )
         );
  MUX \b/U2107  ( .IN0(\b/n2102 ), .IN1(\b/n2101 ), .SEL(msg[18]), .F(
        \b/n2103 ) );
  MUX \b/U2106  ( .IN0(\b/n980 ), .IN1(n621), .SEL(msg[23]), .F(\b/n2102 ) );
  MUX \b/U2105  ( .IN0(\b/n2100 ), .IN1(\b/n2099 ), .SEL(msg[23]), .F(
        \b/n2101 ) );
  AND \b/U2104  ( .A(\b/n1859 ), .B(\b/n1934 ), .Z(\b/n2100 ) );
  MUX \b/U2103  ( .IN0(\b/n952 ), .IN1(\b/n936 ), .SEL(msg[17]), .F(\b/n2099 )
         );
  MUX \b/U2102  ( .IN0(\b/n2097 ), .IN1(\b/n2088 ), .SEL(msg[16]), .F(
        \b/n2098 ) );
  MUX \b/U2101  ( .IN0(\b/n2096 ), .IN1(\b/n2092 ), .SEL(msg[21]), .F(
        \b/n2097 ) );
  MUX \b/U2100  ( .IN0(\b/n2095 ), .IN1(\b/n2093 ), .SEL(msg[18]), .F(
        \b/n2096 ) );
  MUX \b/U2099  ( .IN0(\b/n1865 ), .IN1(\b/n2094 ), .SEL(msg[23]), .F(
        \b/n2095 ) );
  NAND \b/U2098  ( .A(msg[17]), .B(\b/n952 ), .Z(\b/n2094 ) );
  MUX \b/U2097  ( .IN0(\b/n936 ), .IN1(\b/n989 ), .SEL(msg[23]), .F(\b/n2093 )
         );
  MUX \b/U2096  ( .IN0(\b/n2091 ), .IN1(\b/n2090 ), .SEL(msg[18]), .F(
        \b/n2092 ) );
  MUX \b/U2095  ( .IN0(\b/n1891 ), .IN1(\b/n954 ), .SEL(msg[23]), .F(\b/n2091 ) );
  MUX \b/U2094  ( .IN0(\b/n2089 ), .IN1(\b/n1854 ), .SEL(n620), .F(\b/n2090 )
         );
  AND \b/U2093  ( .A(msg[23]), .B(msg[19]), .Z(\b/n2089 ) );
  MUX \b/U2092  ( .IN0(\b/n2087 ), .IN1(\b/n2084 ), .SEL(msg[21]), .F(
        \b/n2088 ) );
  MUX \b/U2091  ( .IN0(\b/n2086 ), .IN1(\b/n2085 ), .SEL(msg[18]), .F(
        \b/n2087 ) );
  MUX \b/U2090  ( .IN0(\b/n2015 ), .IN1(\b/n1854 ), .SEL(msg[23]), .F(
        \b/n2086 ) );
  MUX \b/U2089  ( .IN0(n619), .IN1(\b/n987 ), .SEL(msg[23]), .F(\b/n2085 ) );
  MUX \b/U2088  ( .IN0(\b/n2082 ), .IN1(\b/n2081 ), .SEL(msg[18]), .F(
        \b/n2084 ) );
  AND \b/U2087  ( .A(\b/n2083 ), .B(\b/n1983 ), .Z(\b/n2082 ) );
  MUX \b/U2086  ( .IN0(\b/n938 ), .IN1(\b/n982 ), .SEL(msg[23]), .F(\b/n2081 )
         );
  MUX \b/U2085  ( .IN0(\b/n2080 ), .IN1(\b/n2063 ), .SEL(msg[22]), .F(
        shift_row_out[84]) );
  MUX \b/U2084  ( .IN0(\b/n2079 ), .IN1(\b/n2071 ), .SEL(msg[16]), .F(
        \b/n2080 ) );
  MUX \b/U2083  ( .IN0(\b/n2078 ), .IN1(\b/n2075 ), .SEL(msg[21]), .F(
        \b/n2079 ) );
  MUX \b/U2082  ( .IN0(\b/n2077 ), .IN1(\b/n2076 ), .SEL(msg[18]), .F(
        \b/n2078 ) );
  MUX \b/U2081  ( .IN0(\b/n964 ), .IN1(\b/n985 ), .SEL(msg[23]), .F(\b/n2077 )
         );
  MUX \b/U2080  ( .IN0(\b/n1934 ), .IN1(\b/n1899 ), .SEL(msg[23]), .F(
        \b/n2076 ) );
  NAND \b/U2079  ( .A(msg[17]), .B(\b/n1853 ), .Z(\b/n1934 ) );
  MUX \b/U2078  ( .IN0(\b/n2072 ), .IN1(\b/n2073 ), .SEL(msg[18]), .F(
        \b/n2075 ) );
  AND \b/U2077  ( .A(\b/n1884 ), .B(\b/n2074 ), .Z(\b/n2073 ) );
  MUX \b/U2076  ( .IN0(\b/n1882 ), .IN1(\b/n967 ), .SEL(msg[23]), .F(\b/n2072 ) );
  MUX \b/U2075  ( .IN0(\b/n2070 ), .IN1(\b/n2067 ), .SEL(msg[21]), .F(
        \b/n2071 ) );
  MUX \b/U2074  ( .IN0(\b/n2069 ), .IN1(\b/n2068 ), .SEL(msg[18]), .F(
        \b/n2070 ) );
  MUX \b/U2073  ( .IN0(\b/n929 ), .IN1(\b/n975 ), .SEL(msg[23]), .F(\b/n2069 )
         );
  MUX \b/U2072  ( .IN0(\b/n936 ), .IN1(\b/n1862 ), .SEL(msg[23]), .F(\b/n2068 ) );
  MUX \b/U2071  ( .IN0(\b/n2066 ), .IN1(\b/n2064 ), .SEL(msg[18]), .F(
        \b/n2067 ) );
  MUX \b/U2070  ( .IN0(\b/n1878 ), .IN1(\b/n2065 ), .SEL(msg[23]), .F(
        \b/n2066 ) );
  AND \b/U2069  ( .A(\b/n1862 ), .B(\b/n993 ), .Z(\b/n2065 ) );
  MUX \b/U2068  ( .IN0(\b/n951 ), .IN1(\b/n970 ), .SEL(msg[23]), .F(\b/n2064 )
         );
  MUX \b/U2067  ( .IN0(\b/n2062 ), .IN1(\b/n2056 ), .SEL(msg[16]), .F(
        \b/n2063 ) );
  MUX \b/U2066  ( .IN0(\b/n2061 ), .IN1(\b/n2059 ), .SEL(msg[21]), .F(
        \b/n2062 ) );
  MUX \b/U2065  ( .IN0(\b/n2060 ), .IN1(\b/n1856 ), .SEL(msg[18]), .F(
        \b/n2061 ) );
  MUX \b/U2064  ( .IN0(\b/n1876 ), .IN1(\b/n972 ), .SEL(msg[23]), .F(\b/n2060 ) );
  MUX \b/U2063  ( .IN0(\b/n2058 ), .IN1(\b/n2057 ), .SEL(msg[18]), .F(
        \b/n2059 ) );
  MUX \b/U2062  ( .IN0(n618), .IN1(\b/n964 ), .SEL(msg[23]), .F(\b/n2058 ) );
  MUX \b/U2061  ( .IN0(\b/n1886 ), .IN1(\b/n1889 ), .SEL(msg[23]), .F(
        \b/n2057 ) );
  MUX \b/U2060  ( .IN0(\b/n2055 ), .IN1(\b/n2052 ), .SEL(msg[21]), .F(
        \b/n2056 ) );
  MUX \b/U2059  ( .IN0(\b/n2054 ), .IN1(\b/n2053 ), .SEL(msg[18]), .F(
        \b/n2055 ) );
  MUX \b/U2058  ( .IN0(\b/n937 ), .IN1(\b/n1858 ), .SEL(msg[23]), .F(\b/n2054 ) );
  MUX \b/U2057  ( .IN0(\b/n982 ), .IN1(\b/n1880 ), .SEL(msg[23]), .F(\b/n2053 ) );
  MUX \b/U2056  ( .IN0(\b/n925 ), .IN1(\b/n2051 ), .SEL(msg[18]), .F(\b/n2052 ) );
  MUX \b/U2055  ( .IN0(\b/n945 ), .IN1(\b/n1862 ), .SEL(msg[23]), .F(\b/n2051 ) );
  MUX \b/U2054  ( .IN0(\b/n2050 ), .IN1(\b/n2031 ), .SEL(msg[22]), .F(
        shift_row_out[83]) );
  MUX \b/U2053  ( .IN0(\b/n2049 ), .IN1(\b/n2041 ), .SEL(msg[16]), .F(
        \b/n2050 ) );
  MUX \b/U2052  ( .IN0(\b/n2048 ), .IN1(\b/n2045 ), .SEL(msg[21]), .F(
        \b/n2049 ) );
  MUX \b/U2051  ( .IN0(\b/n2047 ), .IN1(\b/n2046 ), .SEL(msg[23]), .F(
        \b/n2048 ) );
  MUX \b/U2050  ( .IN0(\b/n1870 ), .IN1(\b/n970 ), .SEL(msg[18]), .F(\b/n2047 ) );
  MUX \b/U2049  ( .IN0(n621), .IN1(\b/n928 ), .SEL(msg[18]), .F(\b/n2046 ) );
  MUX \b/U2048  ( .IN0(\b/n2043 ), .IN1(\b/n2042 ), .SEL(msg[23]), .F(
        \b/n2045 ) );
  AND \b/U2047  ( .A(\b/n2044 ), .B(msg[20]), .Z(\b/n2043 ) );
  MUX \b/U2046  ( .IN0(\b/n958 ), .IN1(\b/n1883 ), .SEL(msg[18]), .F(\b/n2042 ) );
  MUX \b/U2045  ( .IN0(\b/n2040 ), .IN1(\b/n2037 ), .SEL(msg[21]), .F(
        \b/n2041 ) );
  MUX \b/U2044  ( .IN0(\b/n2039 ), .IN1(\b/n2038 ), .SEL(msg[23]), .F(
        \b/n2040 ) );
  MUX \b/U2043  ( .IN0(\b/n1874 ), .IN1(n617), .SEL(msg[18]), .F(\b/n2039 ) );
  MUX \b/U2042  ( .IN0(\b/n926 ), .IN1(\b/n945 ), .SEL(msg[18]), .F(\b/n2038 )
         );
  MUX \b/U2041  ( .IN0(\b/n2033 ), .IN1(\b/n2034 ), .SEL(msg[23]), .F(
        \b/n2037 ) );
  NAND \b/U2040  ( .A(\b/n2035 ), .B(\b/n2036 ), .Z(\b/n2034 ) );
  MUX \b/U2039  ( .IN0(\b/n971 ), .IN1(\b/n2032 ), .SEL(msg[18]), .F(\b/n2033 ) );
  MUX \b/U2038  ( .IN0(\b/n946 ), .IN1(\b/n988 ), .SEL(msg[17]), .F(\b/n2032 )
         );
  MUX \b/U2037  ( .IN0(\b/n2030 ), .IN1(\b/n2021 ), .SEL(msg[16]), .F(
        \b/n2031 ) );
  MUX \b/U2036  ( .IN0(\b/n2029 ), .IN1(\b/n2025 ), .SEL(msg[21]), .F(
        \b/n2030 ) );
  MUX \b/U2035  ( .IN0(\b/n2027 ), .IN1(\b/n2026 ), .SEL(msg[23]), .F(
        \b/n2029 ) );
  NAND \b/U2034  ( .A(\b/n936 ), .B(\b/n2028 ), .Z(\b/n2027 ) );
  MUX \b/U2033  ( .IN0(\b/n987 ), .IN1(\b/n949 ), .SEL(msg[18]), .F(\b/n2026 )
         );
  MUX \b/U2032  ( .IN0(\b/n2024 ), .IN1(\b/n2022 ), .SEL(msg[23]), .F(
        \b/n2025 ) );
  MUX \b/U2031  ( .IN0(\b/n1865 ), .IN1(\b/n2023 ), .SEL(msg[18]), .F(
        \b/n2024 ) );
  AND \b/U2030  ( .A(msg[17]), .B(\b/n936 ), .Z(\b/n2023 ) );
  MUX \b/U2029  ( .IN0(\b/n941 ), .IN1(\b/n1884 ), .SEL(msg[18]), .F(\b/n2022 ) );
  MUX \b/U2028  ( .IN0(\b/n2020 ), .IN1(\b/n2014 ), .SEL(msg[21]), .F(
        \b/n2021 ) );
  MUX \b/U2027  ( .IN0(\b/n2019 ), .IN1(\b/n2017 ), .SEL(msg[23]), .F(
        \b/n2020 ) );
  MUX \b/U2026  ( .IN0(\b/n2018 ), .IN1(\b/n1854 ), .SEL(\b/n1902 ), .F(
        \b/n2019 ) );
  MUX \b/U2025  ( .IN0(msg[19]), .IN1(msg[20]), .SEL(msg[18]), .F(\b/n2018 )
         );
  MUX \b/U2024  ( .IN0(\b/n1884 ), .IN1(\b/n2015 ), .SEL(msg[18]), .F(
        \b/n2017 ) );
  NAND \b/U2023  ( .A(\b/n1854 ), .B(\b/n2016 ), .Z(\b/n2015 ) );
  MUX \b/U2022  ( .IN0(\b/n2011 ), .IN1(\b/n2012 ), .SEL(msg[23]), .F(
        \b/n2014 ) );
  AND \b/U2021  ( .A(\b/n969 ), .B(\b/n2013 ), .Z(\b/n2012 ) );
  MUX \b/U2020  ( .IN0(\b/n950 ), .IN1(\b/n1855 ), .SEL(msg[18]), .F(\b/n2011 ) );
  MUX \b/U2019  ( .IN0(\b/n2010 ), .IN1(\b/n1994 ), .SEL(msg[22]), .F(
        shift_row_out[82]) );
  MUX \b/U2018  ( .IN0(\b/n2009 ), .IN1(\b/n2001 ), .SEL(msg[16]), .F(
        \b/n2010 ) );
  MUX \b/U2017  ( .IN0(\b/n2008 ), .IN1(\b/n2004 ), .SEL(msg[21]), .F(
        \b/n2009 ) );
  MUX \b/U2016  ( .IN0(\b/n2007 ), .IN1(\b/n2005 ), .SEL(msg[18]), .F(
        \b/n2008 ) );
  MUX \b/U2015  ( .IN0(\b/n958 ), .IN1(\b/n2006 ), .SEL(msg[23]), .F(\b/n2007 ) );
  MUX \b/U2014  ( .IN0(\b/n1862 ), .IN1(\b/n936 ), .SEL(msg[17]), .F(\b/n2006 ) );
  MUX \b/U2013  ( .IN0(\b/n1901 ), .IN1(\b/n976 ), .SEL(msg[23]), .F(\b/n2005 ) );
  MUX \b/U2012  ( .IN0(\b/n2003 ), .IN1(\b/n2002 ), .SEL(msg[18]), .F(
        \b/n2004 ) );
  MUX \b/U2011  ( .IN0(\b/n1855 ), .IN1(\b/n943 ), .SEL(msg[23]), .F(\b/n2003 ) );
  MUX \b/U2010  ( .IN0(\b/n979 ), .IN1(\b/n1888 ), .SEL(msg[23]), .F(\b/n2002 ) );
  MUX \b/U2009  ( .IN0(\b/n2000 ), .IN1(\b/n1996 ), .SEL(msg[21]), .F(
        \b/n2001 ) );
  MUX \b/U2008  ( .IN0(\b/n1997 ), .IN1(\b/n925 ), .SEL(msg[18]), .F(\b/n2000 ) );
  NAND \b/U2007  ( .A(\b/n1998 ), .B(\b/n1999 ), .Z(\b/n1997 ) );
  MUX \b/U2006  ( .IN0(n619), .IN1(\b/n1995 ), .SEL(\b/n1900 ), .F(\b/n1996 )
         );
  MUX \b/U2005  ( .IN0(\b/n957 ), .IN1(\b/n1867 ), .SEL(msg[18]), .F(\b/n1995 ) );
  MUX \b/U2004  ( .IN0(\b/n1993 ), .IN1(\b/n1985 ), .SEL(msg[16]), .F(
        \b/n1994 ) );
  MUX \b/U2003  ( .IN0(\b/n1992 ), .IN1(\b/n1989 ), .SEL(msg[21]), .F(
        \b/n1993 ) );
  MUX \b/U2002  ( .IN0(\b/n1991 ), .IN1(\b/n1990 ), .SEL(msg[18]), .F(
        \b/n1992 ) );
  MUX \b/U2001  ( .IN0(\b/n985 ), .IN1(msg[17]), .SEL(msg[23]), .F(\b/n1991 )
         );
  MUX \b/U2000  ( .IN0(n622), .IN1(\b/n1868 ), .SEL(msg[23]), .F(\b/n1990 ) );
  MUX \b/U1999  ( .IN0(\b/n1988 ), .IN1(\b/n1987 ), .SEL(msg[18]), .F(
        \b/n1989 ) );
  MUX \b/U1998  ( .IN0(\b/n990 ), .IN1(\b/n984 ), .SEL(msg[23]), .F(\b/n1988 )
         );
  MUX \b/U1997  ( .IN0(n622), .IN1(\b/n1986 ), .SEL(msg[23]), .F(\b/n1987 ) );
  MUX \b/U1996  ( .IN0(\b/n936 ), .IN1(\b/n973 ), .SEL(msg[17]), .F(\b/n1986 )
         );
  MUX \b/U1995  ( .IN0(\b/n1984 ), .IN1(\b/n1978 ), .SEL(msg[21]), .F(
        \b/n1985 ) );
  MUX \b/U1994  ( .IN0(\b/n1981 ), .IN1(\b/n1980 ), .SEL(msg[18]), .F(
        \b/n1984 ) );
  NAND \b/U1993  ( .A(\b/n1982 ), .B(\b/n1983 ), .Z(\b/n1981 ) );
  MUX \b/U1992  ( .IN0(\b/n1854 ), .IN1(\b/n1979 ), .SEL(n620), .F(\b/n1980 )
         );
  MUX \b/U1991  ( .IN0(msg[19]), .IN1(\b/n946 ), .SEL(msg[23]), .F(\b/n1979 )
         );
  MUX \b/U1990  ( .IN0(\b/n1977 ), .IN1(\b/n1976 ), .SEL(msg[18]), .F(
        \b/n1978 ) );
  MUX \b/U1989  ( .IN0(\b/n1899 ), .IN1(\b/n944 ), .SEL(msg[23]), .F(\b/n1977 ) );
  MUX \b/U1988  ( .IN0(\b/n1895 ), .IN1(\b/n1975 ), .SEL(msg[23]), .F(
        \b/n1976 ) );
  MUX \b/U1987  ( .IN0(\b/n1857 ), .IN1(\b/n1862 ), .SEL(msg[17]), .F(
        \b/n1975 ) );
  MUX \b/U1986  ( .IN0(\b/n1974 ), .IN1(\b/n1956 ), .SEL(msg[22]), .F(
        shift_row_out[81]) );
  MUX \b/U1985  ( .IN0(\b/n1973 ), .IN1(\b/n1964 ), .SEL(msg[16]), .F(
        \b/n1974 ) );
  MUX \b/U1984  ( .IN0(\b/n1972 ), .IN1(\b/n1968 ), .SEL(msg[21]), .F(
        \b/n1973 ) );
  MUX \b/U1983  ( .IN0(\b/n1971 ), .IN1(\b/n1970 ), .SEL(msg[18]), .F(
        \b/n1972 ) );
  MUX \b/U1982  ( .IN0(\b/n981 ), .IN1(n624), .SEL(msg[23]), .F(\b/n1971 ) );
  MUX \b/U1981  ( .IN0(\b/n1969 ), .IN1(n618), .SEL(msg[23]), .F(\b/n1970 ) );
  NAND \b/U1980  ( .A(\b/n993 ), .B(\b/n952 ), .Z(\b/n1969 ) );
  MUX \b/U1979  ( .IN0(\b/n1967 ), .IN1(\b/n1966 ), .SEL(msg[18]), .F(
        \b/n1968 ) );
  MUX \b/U1978  ( .IN0(\b/n929 ), .IN1(\b/n1869 ), .SEL(msg[23]), .F(\b/n1967 ) );
  MUX \b/U1977  ( .IN0(\b/n1859 ), .IN1(\b/n1965 ), .SEL(msg[23]), .F(
        \b/n1966 ) );
  AND \b/U1976  ( .A(msg[17]), .B(msg[20]), .Z(\b/n1965 ) );
  MUX \b/U1975  ( .IN0(\b/n1963 ), .IN1(\b/n1960 ), .SEL(msg[21]), .F(
        \b/n1964 ) );
  MUX \b/U1974  ( .IN0(\b/n1962 ), .IN1(\b/n1961 ), .SEL(msg[18]), .F(
        \b/n1963 ) );
  MUX \b/U1973  ( .IN0(\b/n1898 ), .IN1(\b/n990 ), .SEL(msg[23]), .F(\b/n1962 ) );
  MUX \b/U1972  ( .IN0(\b/n965 ), .IN1(\b/n1867 ), .SEL(msg[23]), .F(\b/n1961 ) );
  MUX \b/U1971  ( .IN0(\b/n1957 ), .IN1(\b/n1958 ), .SEL(msg[18]), .F(
        \b/n1960 ) );
  AND \b/U1970  ( .A(\b/n1959 ), .B(\b/n1914 ), .Z(\b/n1958 ) );
  MUX \b/U1969  ( .IN0(\b/n1873 ), .IN1(\b/n1862 ), .SEL(msg[23]), .F(
        \b/n1957 ) );
  MUX \b/U1968  ( .IN0(\b/n1955 ), .IN1(\b/n1947 ), .SEL(msg[16]), .F(
        \b/n1956 ) );
  MUX \b/U1967  ( .IN0(\b/n1954 ), .IN1(\b/n1950 ), .SEL(msg[21]), .F(
        \b/n1955 ) );
  MUX \b/U1966  ( .IN0(\b/n1953 ), .IN1(\b/n1952 ), .SEL(msg[18]), .F(
        \b/n1954 ) );
  MUX \b/U1965  ( .IN0(\b/n1861 ), .IN1(\b/n954 ), .SEL(msg[23]), .F(\b/n1953 ) );
  MUX \b/U1964  ( .IN0(\b/n1951 ), .IN1(\b/n938 ), .SEL(msg[23]), .F(\b/n1952 ) );
  MUX \b/U1963  ( .IN0(\b/n1859 ), .IN1(\b/n946 ), .SEL(msg[17]), .F(\b/n1951 ) );
  MUX \b/U1962  ( .IN0(\b/n1949 ), .IN1(\b/n1948 ), .SEL(msg[18]), .F(
        \b/n1950 ) );
  MUX \b/U1961  ( .IN0(\b/n985 ), .IN1(\b/n963 ), .SEL(msg[23]), .F(\b/n1949 )
         );
  MUX \b/U1960  ( .IN0(\b/n981 ), .IN1(\b/n941 ), .SEL(msg[23]), .F(\b/n1948 )
         );
  MUX \b/U1959  ( .IN0(\b/n1946 ), .IN1(\b/n1941 ), .SEL(msg[21]), .F(
        \b/n1947 ) );
  MUX \b/U1958  ( .IN0(\b/n1945 ), .IN1(\b/n1942 ), .SEL(msg[18]), .F(
        \b/n1946 ) );
  MUX \b/U1957  ( .IN0(\b/n1943 ), .IN1(\b/n1944 ), .SEL(msg[23]), .F(
        \b/n1945 ) );
  NAND \b/U1956  ( .A(\b/n1862 ), .B(\b/n1934 ), .Z(\b/n1944 ) );
  MUX \b/U1955  ( .IN0(\b/n1862 ), .IN1(\b/n946 ), .SEL(msg[17]), .F(\b/n1943 ) );
  MUX \b/U1954  ( .IN0(\b/n1879 ), .IN1(\b/n1877 ), .SEL(msg[23]), .F(
        \b/n1942 ) );
  MUX \b/U1953  ( .IN0(\b/n1897 ), .IN1(\b/n1940 ), .SEL(msg[18]), .F(
        \b/n1941 ) );
  MUX \b/U1952  ( .IN0(\b/n952 ), .IN1(\b/n984 ), .SEL(msg[23]), .F(\b/n1940 )
         );
  MUX \b/U1951  ( .IN0(\b/n1939 ), .IN1(\b/n1922 ), .SEL(msg[22]), .F(
        shift_row_out[80]) );
  MUX \b/U1950  ( .IN0(\b/n1938 ), .IN1(\b/n1930 ), .SEL(msg[16]), .F(
        \b/n1939 ) );
  MUX \b/U1949  ( .IN0(\b/n1937 ), .IN1(\b/n1935 ), .SEL(msg[18]), .F(
        \b/n1938 ) );
  MUX \b/U1948  ( .IN0(\b/n926 ), .IN1(\b/n1936 ), .SEL(msg[23]), .F(\b/n1937 ) );
  MUX \b/U1947  ( .IN0(\b/n979 ), .IN1(\b/n982 ), .SEL(msg[21]), .F(\b/n1936 )
         );
  MUX \b/U1946  ( .IN0(\b/n1932 ), .IN1(\b/n1931 ), .SEL(msg[23]), .F(
        \b/n1935 ) );
  NAND \b/U1945  ( .A(\b/n1933 ), .B(\b/n1934 ), .Z(\b/n1932 ) );
  MUX \b/U1944  ( .IN0(\b/n978 ), .IN1(\b/n993 ), .SEL(msg[21]), .F(\b/n1931 )
         );
  MUX \b/U1943  ( .IN0(\b/n1929 ), .IN1(\b/n1925 ), .SEL(msg[18]), .F(
        \b/n1930 ) );
  MUX \b/U1942  ( .IN0(\b/n1928 ), .IN1(\b/n1926 ), .SEL(msg[23]), .F(
        \b/n1929 ) );
  MUX \b/U1941  ( .IN0(\b/n1927 ), .IN1(\b/n931 ), .SEL(msg[21]), .F(\b/n1928 ) );
  NAND \b/U1940  ( .A(\b/n993 ), .B(\b/n1854 ), .Z(\b/n1927 ) );
  MUX \b/U1938  ( .IN0(\b/n1924 ), .IN1(\b/n1923 ), .SEL(msg[23]), .F(
        \b/n1925 ) );
  MUX \b/U1937  ( .IN0(n619), .IN1(\b/n928 ), .SEL(msg[21]), .F(\b/n1924 ) );
  MUX \b/U1936  ( .IN0(\b/n980 ), .IN1(\b/n936 ), .SEL(msg[21]), .F(\b/n1923 )
         );
  MUX \b/U1935  ( .IN0(\b/n1921 ), .IN1(\b/n1911 ), .SEL(msg[16]), .F(
        \b/n1922 ) );
  MUX \b/U1934  ( .IN0(\b/n1920 ), .IN1(\b/n1916 ), .SEL(msg[18]), .F(
        \b/n1921 ) );
  MUX \b/U1933  ( .IN0(\b/n1919 ), .IN1(\b/n1918 ), .SEL(msg[23]), .F(
        \b/n1920 ) );
  MUX \b/U1932  ( .IN0(n617), .IN1(\b/n932 ), .SEL(msg[21]), .F(\b/n1919 ) );
  MUX \b/U1931  ( .IN0(\b/n1917 ), .IN1(\b/n969 ), .SEL(msg[21]), .F(\b/n1918 ) );
  NAND \b/U1930  ( .A(\b/n1853 ), .B(\b/n1855 ), .Z(\b/n1917 ) );
  MUX \b/U1929  ( .IN0(\b/n1915 ), .IN1(\b/n1912 ), .SEL(msg[23]), .F(
        \b/n1916 ) );
  MUX \b/U1928  ( .IN0(\b/n939 ), .IN1(\b/n1913 ), .SEL(msg[21]), .F(\b/n1915 ) );
  NAND \b/U1927  ( .A(\b/n1857 ), .B(\b/n1914 ), .Z(\b/n1913 ) );
  MUX \b/U1926  ( .IN0(\b/n1872 ), .IN1(\b/n1863 ), .SEL(msg[21]), .F(
        \b/n1912 ) );
  MUX \b/U1925  ( .IN0(\b/n1910 ), .IN1(\b/n1906 ), .SEL(msg[18]), .F(
        \b/n1911 ) );
  MUX \b/U1924  ( .IN0(\b/n1908 ), .IN1(\b/n1907 ), .SEL(msg[23]), .F(
        \b/n1910 ) );
  NAND \b/U1923  ( .A(\b/n1909 ), .B(\b/n1896 ), .Z(\b/n1908 ) );
  MUX \b/U1922  ( .IN0(msg[19]), .IN1(\b/n1888 ), .SEL(msg[21]), .F(\b/n1907 )
         );
  MUX \b/U1921  ( .IN0(\b/n1905 ), .IN1(\b/n1904 ), .SEL(msg[23]), .F(
        \b/n1906 ) );
  MUX \b/U1920  ( .IN0(\b/n944 ), .IN1(\b/n960 ), .SEL(msg[21]), .F(\b/n1905 )
         );
  MUX \b/U1919  ( .IN0(\b/n977 ), .IN1(\b/n965 ), .SEL(msg[21]), .F(\b/n1904 )
         );
  XOR \b/U1918  ( .A(\b/n1854 ), .B(msg[17]), .Z(\b/n1903 ) );
  XOR \b/U1917  ( .A(msg[17]), .B(msg[18]), .Z(\b/n1902 ) );
  XOR \b/U1916  ( .A(msg[17]), .B(msg[19]), .Z(\b/n1901 ) );
  XOR \b/U1915  ( .A(msg[18]), .B(msg[23]), .Z(\b/n1900 ) );
  XOR \b/U1914  ( .A(\b/n993 ), .B(\b/n936 ), .Z(\b/n1899 ) );
  XOR \b/U1913  ( .A(msg[17]), .B(\b/n982 ), .Z(\b/n1898 ) );
  XOR \b/U1911  ( .A(msg[17]), .B(msg[21]), .Z(\b/n1896 ) );
  NAND \b/U1910  ( .A(msg[17]), .B(msg[19]), .Z(\b/n1895 ) );
  MUX \b/U1909  ( .IN0(\b/n1854 ), .IN1(\b/n936 ), .SEL(msg[17]), .F(\b/n1894 ) );
  MUX \b/U1907  ( .IN0(msg[19]), .IN1(\b/n973 ), .SEL(msg[17]), .F(\b/n1892 )
         );
  MUX \b/U1906  ( .IN0(\b/n952 ), .IN1(\b/n973 ), .SEL(msg[17]), .F(\b/n1891 )
         );
  MUX \b/U1905  ( .IN0(\b/n1857 ), .IN1(\b/n1859 ), .SEL(msg[17]), .F(
        \b/n1890 ) );
  MUX \b/U1904  ( .IN0(msg[20]), .IN1(\b/n952 ), .SEL(msg[17]), .F(\b/n1889 )
         );
  OR \b/U1903  ( .A(msg[17]), .B(msg[20]), .Z(\b/n1888 ) );
  NAND \b/U1901  ( .A(\b/n973 ), .B(\b/n993 ), .Z(\b/n1886 ) );
  MUX \b/U1900  ( .IN0(\b/n973 ), .IN1(msg[20]), .SEL(msg[17]), .F(\b/n1885 )
         );
  MUX \b/U1899  ( .IN0(\b/n1853 ), .IN1(\b/n1862 ), .SEL(msg[17]), .F(
        \b/n1884 ) );
  MUX \b/U1898  ( .IN0(\b/n988 ), .IN1(msg[20]), .SEL(msg[17]), .F(\b/n1883 )
         );
  MUX \b/U1897  ( .IN0(\b/n946 ), .IN1(\b/n973 ), .SEL(msg[17]), .F(\b/n1882 )
         );
  MUX \b/U1896  ( .IN0(\b/n1853 ), .IN1(msg[20]), .SEL(msg[17]), .F(\b/n1881 )
         );
  MUX \b/U1895  ( .IN0(\b/n963 ), .IN1(\b/n952 ), .SEL(msg[17]), .F(\b/n1880 )
         );
  XOR \b/U1894  ( .A(\b/n946 ), .B(msg[17]), .Z(\b/n1879 ) );
  MUX \b/U1893  ( .IN0(\b/n1859 ), .IN1(\b/n963 ), .SEL(msg[17]), .F(\b/n1878 ) );
  NANDN \b/U1892  ( .B(msg[17]), .A(msg[19]), .Z(\b/n1877 ) );
  MUX \b/U1891  ( .IN0(\b/n936 ), .IN1(msg[19]), .SEL(msg[17]), .F(\b/n1876 )
         );
  NAND \b/U1889  ( .A(\b/n1857 ), .B(\b/n993 ), .Z(\b/n1874 ) );
  MUX \b/U1888  ( .IN0(msg[20]), .IN1(\b/n1854 ), .SEL(msg[17]), .F(\b/n1873 )
         );
  MUX \b/U1887  ( .IN0(\b/n963 ), .IN1(msg[19]), .SEL(msg[17]), .F(\b/n1872 )
         );
  MUX \b/U1885  ( .IN0(msg[20]), .IN1(\b/n982 ), .SEL(msg[17]), .F(\b/n1870 )
         );
  MUX \b/U1884  ( .IN0(\b/n936 ), .IN1(\b/n988 ), .SEL(msg[17]), .F(\b/n1869 )
         );
  NAND \b/U1883  ( .A(\b/n1855 ), .B(\b/n936 ), .Z(\b/n1868 ) );
  MUX \b/U1882  ( .IN0(\b/n1854 ), .IN1(\b/n1862 ), .SEL(msg[17]), .F(
        \b/n1867 ) );
  NAND \b/U1881  ( .A(\b/n1866 ), .B(\b/n1853 ), .Z(\b/n1865 ) );
  MUX \b/U1880  ( .IN0(\b/n1857 ), .IN1(\b/n988 ), .SEL(msg[17]), .F(\b/n1864 ) );
  MUX \b/U1879  ( .IN0(\b/n988 ), .IN1(\b/n952 ), .SEL(msg[17]), .F(\b/n1863 )
         );
  NANDN \b/U1878  ( .B(msg[19]), .A(msg[20]), .Z(\b/n1862 ) );
  MUX \b/U1877  ( .IN0(\b/n1857 ), .IN1(msg[19]), .SEL(msg[17]), .F(\b/n1861 )
         );
  OR \b/U1876  ( .A(msg[19]), .B(msg[20]), .Z(\b/n1857 ) );
  MUX \b/U1875  ( .IN0(\b/n936 ), .IN1(\b/n952 ), .SEL(msg[17]), .F(\b/n1860 )
         );
  XOR \b/U1874  ( .A(\b/n946 ), .B(msg[19]), .Z(\b/n1859 ) );
  NANDN \b/U1873  ( .B(msg[19]), .A(msg[17]), .Z(\b/n1858 ) );
  NAND \b/U1872  ( .A(\b/n1857 ), .B(\b/n1855 ), .Z(\b/n1856 ) );
  NAND \b/U1871  ( .A(msg[17]), .B(\b/n1854 ), .Z(\b/n1855 ) );
  NANDN \b/U1870  ( .B(msg[20]), .A(msg[19]), .Z(\b/n1854 ) );
  NAND \b/U1869  ( .A(msg[19]), .B(msg[20]), .Z(\b/n1853 ) );
  MUX \b/U1868  ( .IN0(msg[12]), .IN1(\b/n1494 ), .SEL(msg[9]), .F(\b/n1852 )
         );
  MUX \b/U1867  ( .IN0(msg[12]), .IN1(\b/n1495 ), .SEL(msg[9]), .F(\b/n1851 )
         );
  MUX \b/U1866  ( .IN0(\b/n1497 ), .IN1(\b/n1501 ), .SEL(msg[9]), .F(\b/n1850 ) );
  MUX \b/U1865  ( .IN0(\b/n1519 ), .IN1(\b/n1032 ), .SEL(msg[9]), .F(\b/n1849 ) );
  MUX \b/U1863  ( .IN0(\b/n1495 ), .IN1(\b/n1494 ), .SEL(msg[10]), .F(
        \b/n1666 ) );
  MUX \b/U1862  ( .IN0(\b/n1496 ), .IN1(\b/n1063 ), .SEL(msg[10]), .F(
        \b/n1667 ) );
  MUX \b/U1861  ( .IN0(\b/n1007 ), .IN1(\b/n1015 ), .SEL(msg[9]), .F(\b/n1631 ) );
  MUX \b/U1860  ( .IN0(\b/n1524 ), .IN1(\b/n1835 ), .SEL(msg[15]), .F(
        \b/n1847 ) );
  MUX \b/U1859  ( .IN0(\b/n1501 ), .IN1(\b/n1494 ), .SEL(msg[9]), .F(\b/n1838 ) );
  MUX \b/U1858  ( .IN0(\b/n1058 ), .IN1(\b/n1519 ), .SEL(msg[9]), .F(\b/n1846 ) );
  MUX \b/U1857  ( .IN0(msg[11]), .IN1(\b/n1032 ), .SEL(msg[9]), .F(\b/n1845 )
         );
  MUX \b/U1856  ( .IN0(\b/n1495 ), .IN1(\b/n1058 ), .SEL(msg[9]), .F(\b/n1844 ) );
  MUX \b/U1855  ( .IN0(msg[12]), .IN1(\b/n1519 ), .SEL(msg[9]), .F(\b/n1843 )
         );
  MUX \b/U1854  ( .IN0(\b/n1042 ), .IN1(\b/n1021 ), .SEL(msg[13]), .F(
        \b/n1550 ) );
  MUX \b/U1853  ( .IN0(\b/n1497 ), .IN1(\b/n1015 ), .SEL(msg[9]), .F(\b/n1842 ) );
  NANDN \b/U1850  ( .B(\b/n1502 ), .A(msg[15]), .Z(\b/n1806 ) );
  NAND \b/U1849  ( .A(msg[15]), .B(\b/n1018 ), .Z(\b/n1775 ) );
  NAND \b/U1848  ( .A(msg[15]), .B(\b/n1050 ), .Z(\b/n1724 ) );
  NAND \b/U1847  ( .A(msg[15]), .B(\b/n1831 ), .Z(\b/n1757 ) );
  NAND \b/U1846  ( .A(msg[15]), .B(\b/n1752 ), .Z(\b/n1715 ) );
  NAND \b/U1844  ( .A(\b/n1063 ), .B(\b/n1032 ), .Z(\b/n1837 ) );
  NAND \b/U1843  ( .A(msg[15]), .B(\b/n1834 ), .Z(\b/n1829 ) );
  NAND \b/U1842  ( .A(n616), .B(msg[15]), .Z(\b/n1818 ) );
  NAND \b/U1840  ( .A(msg[10]), .B(\b/n1495 ), .Z(\b/n1680 ) );
  NAND \b/U1839  ( .A(msg[9]), .B(\b/n1032 ), .Z(\b/n1624 ) );
  NAND \b/U1838  ( .A(msg[15]), .B(\b/n1838 ), .Z(\b/n1623 ) );
  NAND \b/U1837  ( .A(\b/n1837 ), .B(msg[15]), .Z(\b/n1630 ) );
  NAND \b/U1835  ( .A(\b/n1495 ), .B(\b/n1657 ), .Z(\b/n1835 ) );
  NANDN \b/U1834  ( .B(\b/n1007 ), .A(\b/n1063 ), .Z(\b/n1834 ) );
  NAND \b/U1831  ( .A(msg[9]), .B(\b/n1501 ), .Z(\b/n1657 ) );
  NAND \b/U1830  ( .A(\b/n1495 ), .B(msg[9]), .Z(\b/n1564 ) );
  NAND \b/U1829  ( .A(\b/n1007 ), .B(\b/n1063 ), .Z(\b/n1831 ) );
  ANDN \b/U1826  ( .A(msg[10]), .B(msg[9]), .Z(\b/n1685 ) );
  AND \b/U1825  ( .A(\b/n1829 ), .B(\b/n1497 ), .Z(\b/n1591 ) );
  MUX \b/U1824  ( .IN0(\b/n1828 ), .IN1(\b/n1812 ), .SEL(msg[8]), .F(
        shift_row_out[111]) );
  MUX \b/U1823  ( .IN0(\b/n1827 ), .IN1(\b/n1820 ), .SEL(msg[14]), .F(
        \b/n1828 ) );
  MUX \b/U1822  ( .IN0(\b/n1826 ), .IN1(\b/n1823 ), .SEL(msg[13]), .F(
        \b/n1827 ) );
  MUX \b/U1821  ( .IN0(\b/n1825 ), .IN1(\b/n1824 ), .SEL(msg[10]), .F(
        \b/n1826 ) );
  MUX \b/U1820  ( .IN0(msg[12]), .IN1(\b/n1022 ), .SEL(msg[15]), .F(\b/n1825 )
         );
  MUX \b/U1819  ( .IN0(\b/n1496 ), .IN1(\b/n1026 ), .SEL(msg[15]), .F(
        \b/n1824 ) );
  MUX \b/U1818  ( .IN0(\b/n1822 ), .IN1(\b/n1821 ), .SEL(msg[10]), .F(
        \b/n1823 ) );
  MUX \b/U1817  ( .IN0(\b/n1563 ), .IN1(\b/n1018 ), .SEL(msg[15]), .F(
        \b/n1822 ) );
  MUX \b/U1816  ( .IN0(\b/n1508 ), .IN1(\b/n1517 ), .SEL(msg[15]), .F(
        \b/n1821 ) );
  MUX \b/U1815  ( .IN0(\b/n1819 ), .IN1(\b/n1815 ), .SEL(msg[13]), .F(
        \b/n1820 ) );
  MUX \b/U1814  ( .IN0(\b/n1816 ), .IN1(\b/n1817 ), .SEL(msg[10]), .F(
        \b/n1819 ) );
  NAND \b/U1813  ( .A(\b/n1624 ), .B(\b/n1818 ), .Z(\b/n1817 ) );
  MUX \b/U1812  ( .IN0(\b/n1059 ), .IN1(\b/n1033 ), .SEL(msg[15]), .F(
        \b/n1816 ) );
  MUX \b/U1811  ( .IN0(\b/n1814 ), .IN1(\b/n1813 ), .SEL(msg[10]), .F(
        \b/n1815 ) );
  MUX \b/U1810  ( .IN0(\b/n1519 ), .IN1(\b/n1494 ), .SEL(msg[15]), .F(
        \b/n1814 ) );
  MUX \b/U1809  ( .IN0(\b/n1034 ), .IN1(\b/n1530 ), .SEL(msg[15]), .F(
        \b/n1813 ) );
  MUX \b/U1808  ( .IN0(\b/n1811 ), .IN1(\b/n1803 ), .SEL(msg[14]), .F(
        \b/n1812 ) );
  MUX \b/U1807  ( .IN0(\b/n1810 ), .IN1(\b/n1807 ), .SEL(msg[13]), .F(
        \b/n1811 ) );
  MUX \b/U1806  ( .IN0(\b/n1809 ), .IN1(\b/n1808 ), .SEL(msg[10]), .F(
        \b/n1810 ) );
  MUX \b/U1805  ( .IN0(\b/n1529 ), .IN1(\b/n1505 ), .SEL(msg[15]), .F(
        \b/n1809 ) );
  MUX \b/U1804  ( .IN0(\b/n1050 ), .IN1(\b/n1526 ), .SEL(msg[15]), .F(
        \b/n1808 ) );
  MUX \b/U1803  ( .IN0(\b/n1805 ), .IN1(\b/n1804 ), .SEL(msg[10]), .F(
        \b/n1807 ) );
  AND \b/U1802  ( .A(\b/n1020 ), .B(\b/n1806 ), .Z(\b/n1805 ) );
  MUX \b/U1801  ( .IN0(\b/n1512 ), .IN1(n615), .SEL(msg[15]), .F(\b/n1804 ) );
  MUX \b/U1800  ( .IN0(\b/n1802 ), .IN1(\b/n1799 ), .SEL(msg[13]), .F(
        \b/n1803 ) );
  MUX \b/U1799  ( .IN0(\b/n1801 ), .IN1(\b/n1800 ), .SEL(msg[10]), .F(
        \b/n1802 ) );
  MUX \b/U1798  ( .IN0(\b/n1535 ), .IN1(\b/n1521 ), .SEL(msg[15]), .F(
        \b/n1801 ) );
  MUX \b/U1797  ( .IN0(\b/n1008 ), .IN1(\b/n1495 ), .SEL(msg[15]), .F(
        \b/n1800 ) );
  MUX \b/U1796  ( .IN0(\b/n1798 ), .IN1(\b/n1797 ), .SEL(msg[10]), .F(
        \b/n1799 ) );
  MUX \b/U1795  ( .IN0(\b/n1499 ), .IN1(\b/n1544 ), .SEL(msg[15]), .F(
        \b/n1798 ) );
  MUX \b/U1794  ( .IN0(\b/n1498 ), .IN1(\b/n1796 ), .SEL(msg[15]), .F(
        \b/n1797 ) );
  MUX \b/U1793  ( .IN0(\b/n1058 ), .IN1(\b/n1015 ), .SEL(msg[9]), .F(\b/n1796 ) );
  MUX \b/U1792  ( .IN0(\b/n1795 ), .IN1(\b/n1778 ), .SEL(msg[8]), .F(
        shift_row_out[110]) );
  MUX \b/U1791  ( .IN0(\b/n1794 ), .IN1(\b/n1785 ), .SEL(msg[14]), .F(
        \b/n1795 ) );
  MUX \b/U1790  ( .IN0(\b/n1793 ), .IN1(\b/n1788 ), .SEL(msg[13]), .F(
        \b/n1794 ) );
  MUX \b/U1789  ( .IN0(\b/n1792 ), .IN1(\b/n1790 ), .SEL(msg[10]), .F(
        \b/n1793 ) );
  MUX \b/U1788  ( .IN0(\b/n1791 ), .IN1(\b/n1509 ), .SEL(msg[15]), .F(
        \b/n1792 ) );
  MUX \b/U1787  ( .IN0(\b/n1058 ), .IN1(\b/n1494 ), .SEL(msg[9]), .F(\b/n1791 ) );
  MUX \b/U1786  ( .IN0(\b/n1789 ), .IN1(\b/n1035 ), .SEL(msg[15]), .F(
        \b/n1790 ) );
  MUX \b/U1785  ( .IN0(\b/n1494 ), .IN1(\b/n1497 ), .SEL(msg[9]), .F(\b/n1789 ) );
  MUX \b/U1784  ( .IN0(\b/n1787 ), .IN1(\b/n1786 ), .SEL(msg[10]), .F(
        \b/n1788 ) );
  MUX \b/U1783  ( .IN0(n614), .IN1(\b/n1575 ), .SEL(msg[15]), .F(\b/n1787 ) );
  MUX \b/U1782  ( .IN0(\b/n1531 ), .IN1(\b/n1540 ), .SEL(msg[15]), .F(
        \b/n1786 ) );
  MUX \b/U1781  ( .IN0(\b/n1784 ), .IN1(\b/n1781 ), .SEL(msg[13]), .F(
        \b/n1785 ) );
  MUX \b/U1780  ( .IN0(\b/n1783 ), .IN1(\b/n1782 ), .SEL(msg[10]), .F(
        \b/n1784 ) );
  MUX \b/U1779  ( .IN0(\b/n1049 ), .IN1(\b/n1503 ), .SEL(msg[15]), .F(
        \b/n1783 ) );
  MUX \b/U1778  ( .IN0(\b/n1508 ), .IN1(n615), .SEL(msg[15]), .F(\b/n1782 ) );
  MUX \b/U1777  ( .IN0(\b/n1780 ), .IN1(\b/n1779 ), .SEL(msg[10]), .F(
        \b/n1781 ) );
  MUX \b/U1776  ( .IN0(\b/n1522 ), .IN1(\b/n1004 ), .SEL(msg[15]), .F(
        \b/n1780 ) );
  MUX \b/U1775  ( .IN0(\b/n1022 ), .IN1(\b/n1033 ), .SEL(msg[15]), .F(
        \b/n1779 ) );
  MUX \b/U1774  ( .IN0(\b/n1777 ), .IN1(\b/n1769 ), .SEL(msg[14]), .F(
        \b/n1778 ) );
  MUX \b/U1773  ( .IN0(\b/n1776 ), .IN1(\b/n1772 ), .SEL(msg[13]), .F(
        \b/n1777 ) );
  MUX \b/U1772  ( .IN0(\b/n1774 ), .IN1(\b/n1773 ), .SEL(msg[10]), .F(
        \b/n1776 ) );
  AND \b/U1771  ( .A(\b/n1000 ), .B(\b/n1775 ), .Z(\b/n1774 ) );
  MUX \b/U1770  ( .IN0(\b/n1610 ), .IN1(msg[11]), .SEL(msg[15]), .F(\b/n1773 )
         );
  MUX \b/U1769  ( .IN0(\b/n1771 ), .IN1(\b/n1770 ), .SEL(msg[10]), .F(
        \b/n1772 ) );
  MUX \b/U1768  ( .IN0(\b/n1041 ), .IN1(\b/n1501 ), .SEL(msg[15]), .F(
        \b/n1771 ) );
  MUX \b/U1766  ( .IN0(\b/n1768 ), .IN1(\b/n1764 ), .SEL(msg[13]), .F(
        \b/n1769 ) );
  MUX \b/U1765  ( .IN0(\b/n1767 ), .IN1(\b/n1766 ), .SEL(msg[10]), .F(
        \b/n1768 ) );
  MUX \b/U1764  ( .IN0(\b/n1513 ), .IN1(\b/n1033 ), .SEL(msg[15]), .F(
        \b/n1767 ) );
  MUX \b/U1763  ( .IN0(\b/n1765 ), .IN1(\b/n1532 ), .SEL(msg[15]), .F(
        \b/n1766 ) );
  NANDN \b/U1762  ( .B(msg[12]), .A(msg[9]), .Z(\b/n1765 ) );
  MUX \b/U1761  ( .IN0(\b/n1763 ), .IN1(\b/n1761 ), .SEL(msg[10]), .F(
        \b/n1764 ) );
  MUX \b/U1760  ( .IN0(\b/n1015 ), .IN1(\b/n1762 ), .SEL(msg[15]), .F(
        \b/n1763 ) );
  MUX \b/U1759  ( .IN0(\b/n1042 ), .IN1(\b/n1052 ), .SEL(msg[9]), .F(\b/n1762 ) );
  MUX \b/U1758  ( .IN0(\b/n1006 ), .IN1(\b/n1509 ), .SEL(msg[15]), .F(
        \b/n1761 ) );
  NANDN \b/U1757  ( .B(\b/n1007 ), .A(msg[9]), .Z(\b/n1509 ) );
  MUX \b/U1756  ( .IN0(\b/n1760 ), .IN1(\b/n1740 ), .SEL(msg[8]), .F(
        shift_row_out[109]) );
  MUX \b/U1755  ( .IN0(\b/n1759 ), .IN1(\b/n1749 ), .SEL(msg[14]), .F(
        \b/n1760 ) );
  MUX \b/U1754  ( .IN0(\b/n1758 ), .IN1(\b/n1754 ), .SEL(msg[13]), .F(
        \b/n1759 ) );
  MUX \b/U1753  ( .IN0(\b/n1755 ), .IN1(\b/n1756 ), .SEL(msg[10]), .F(
        \b/n1758 ) );
  AND \b/U1752  ( .A(\b/n1525 ), .B(\b/n1757 ), .Z(\b/n1756 ) );
  MUX \b/U1751  ( .IN0(\b/n1495 ), .IN1(\b/n1034 ), .SEL(msg[15]), .F(
        \b/n1755 ) );
  MUX \b/U1750  ( .IN0(\b/n1753 ), .IN1(\b/n1751 ), .SEL(msg[10]), .F(
        \b/n1754 ) );
  MUX \b/U1749  ( .IN0(\b/n1010 ), .IN1(\b/n1752 ), .SEL(msg[15]), .F(
        \b/n1753 ) );
  NAND \b/U1748  ( .A(\b/n1052 ), .B(\b/n1063 ), .Z(\b/n1752 ) );
  MUX \b/U1747  ( .IN0(\b/n1495 ), .IN1(\b/n1750 ), .SEL(msg[15]), .F(
        \b/n1751 ) );
  NAND \b/U1746  ( .A(\b/n1494 ), .B(\b/n1564 ), .Z(\b/n1750 ) );
  MUX \b/U1745  ( .IN0(\b/n1748 ), .IN1(\b/n1744 ), .SEL(msg[13]), .F(
        \b/n1749 ) );
  MUX \b/U1744  ( .IN0(\b/n1747 ), .IN1(\b/n1745 ), .SEL(msg[10]), .F(
        \b/n1748 ) );
  MUX \b/U1743  ( .IN0(\b/n1508 ), .IN1(\b/n1746 ), .SEL(msg[15]), .F(
        \b/n1747 ) );
  NAND \b/U1742  ( .A(msg[9]), .B(\b/n1021 ), .Z(\b/n1746 ) );
  MUX \b/U1741  ( .IN0(\b/n1007 ), .IN1(\b/n1061 ), .SEL(msg[15]), .F(
        \b/n1745 ) );
  MUX \b/U1740  ( .IN0(\b/n1743 ), .IN1(\b/n1742 ), .SEL(msg[10]), .F(
        \b/n1744 ) );
  MUX \b/U1739  ( .IN0(\b/n1532 ), .IN1(\b/n1023 ), .SEL(msg[15]), .F(
        \b/n1743 ) );
  MUX \b/U1738  ( .IN0(\b/n1741 ), .IN1(\b/n1497 ), .SEL(n613), .F(\b/n1742 )
         );
  AND \b/U1737  ( .A(msg[15]), .B(msg[11]), .Z(\b/n1741 ) );
  MUX \b/U1736  ( .IN0(\b/n1739 ), .IN1(\b/n1729 ), .SEL(msg[14]), .F(
        \b/n1740 ) );
  MUX \b/U1735  ( .IN0(\b/n1738 ), .IN1(\b/n1734 ), .SEL(msg[13]), .F(
        \b/n1739 ) );
  MUX \b/U1734  ( .IN0(\b/n1737 ), .IN1(\b/n1736 ), .SEL(msg[10]), .F(
        \b/n1738 ) );
  MUX \b/U1733  ( .IN0(\b/n1515 ), .IN1(\b/n1056 ), .SEL(msg[15]), .F(
        \b/n1737 ) );
  MUX \b/U1732  ( .IN0(\b/n1540 ), .IN1(\b/n1735 ), .SEL(msg[15]), .F(
        \b/n1736 ) );
  MUX \b/U1731  ( .IN0(\b/n1032 ), .IN1(\b/n1052 ), .SEL(msg[9]), .F(\b/n1735 ) );
  MUX \b/U1730  ( .IN0(\b/n1733 ), .IN1(\b/n1732 ), .SEL(msg[10]), .F(
        \b/n1734 ) );
  MUX \b/U1729  ( .IN0(\b/n1030 ), .IN1(n612), .SEL(msg[15]), .F(\b/n1733 ) );
  MUX \b/U1728  ( .IN0(\b/n1731 ), .IN1(\b/n1730 ), .SEL(msg[15]), .F(
        \b/n1732 ) );
  AND \b/U1727  ( .A(\b/n1519 ), .B(\b/n1575 ), .Z(\b/n1731 ) );
  MUX \b/U1726  ( .IN0(\b/n1021 ), .IN1(\b/n1007 ), .SEL(msg[9]), .F(\b/n1730 ) );
  MUX \b/U1725  ( .IN0(\b/n1728 ), .IN1(\b/n1725 ), .SEL(msg[13]), .F(
        \b/n1729 ) );
  MUX \b/U1724  ( .IN0(\b/n1727 ), .IN1(\b/n1726 ), .SEL(msg[10]), .F(
        \b/n1728 ) );
  MUX \b/U1723  ( .IN0(\b/n1656 ), .IN1(\b/n1497 ), .SEL(msg[15]), .F(
        \b/n1727 ) );
  MUX \b/U1722  ( .IN0(n611), .IN1(\b/n1038 ), .SEL(msg[15]), .F(\b/n1726 ) );
  MUX \b/U1721  ( .IN0(\b/n1723 ), .IN1(\b/n1722 ), .SEL(msg[10]), .F(
        \b/n1725 ) );
  AND \b/U1720  ( .A(\b/n1724 ), .B(\b/n1624 ), .Z(\b/n1723 ) );
  MUX \b/U1719  ( .IN0(\b/n1009 ), .IN1(\b/n1032 ), .SEL(msg[15]), .F(
        \b/n1722 ) );
  MUX \b/U1718  ( .IN0(\b/n1721 ), .IN1(\b/n1706 ), .SEL(msg[8]), .F(
        shift_row_out[108]) );
  MUX \b/U1717  ( .IN0(\b/n1720 ), .IN1(\b/n1712 ), .SEL(msg[14]), .F(
        \b/n1721 ) );
  MUX \b/U1716  ( .IN0(\b/n1719 ), .IN1(\b/n1716 ), .SEL(msg[13]), .F(
        \b/n1720 ) );
  MUX \b/U1715  ( .IN0(\b/n1718 ), .IN1(\b/n1717 ), .SEL(msg[10]), .F(
        \b/n1719 ) );
  MUX \b/U1714  ( .IN0(\b/n1043 ), .IN1(\b/n1036 ), .SEL(msg[15]), .F(
        \b/n1718 ) );
  MUX \b/U1713  ( .IN0(\b/n1575 ), .IN1(\b/n1540 ), .SEL(msg[15]), .F(
        \b/n1717 ) );
  NAND \b/U1712  ( .A(msg[9]), .B(\b/n1494 ), .Z(\b/n1575 ) );
  MUX \b/U1711  ( .IN0(\b/n1713 ), .IN1(\b/n1714 ), .SEL(msg[10]), .F(
        \b/n1716 ) );
  AND \b/U1710  ( .A(\b/n1525 ), .B(\b/n1715 ), .Z(\b/n1714 ) );
  MUX \b/U1709  ( .IN0(\b/n1523 ), .IN1(\b/n1055 ), .SEL(msg[15]), .F(
        \b/n1713 ) );
  MUX \b/U1708  ( .IN0(\b/n1711 ), .IN1(\b/n1709 ), .SEL(msg[13]), .F(
        \b/n1712 ) );
  MUX \b/U1707  ( .IN0(\b/n1710 ), .IN1(\b/n1500 ), .SEL(msg[10]), .F(
        \b/n1711 ) );
  MUX \b/U1706  ( .IN0(\b/n1517 ), .IN1(\b/n1041 ), .SEL(msg[15]), .F(
        \b/n1710 ) );
  MUX \b/U1705  ( .IN0(\b/n1708 ), .IN1(\b/n1707 ), .SEL(msg[10]), .F(
        \b/n1709 ) );
  MUX \b/U1704  ( .IN0(n610), .IN1(\b/n1043 ), .SEL(msg[15]), .F(\b/n1708 ) );
  MUX \b/U1703  ( .IN0(\b/n1528 ), .IN1(\b/n1529 ), .SEL(msg[15]), .F(
        \b/n1707 ) );
  MUX \b/U1702  ( .IN0(\b/n1705 ), .IN1(\b/n1697 ), .SEL(msg[14]), .F(
        \b/n1706 ) );
  MUX \b/U1701  ( .IN0(\b/n1704 ), .IN1(\b/n1701 ), .SEL(msg[13]), .F(
        \b/n1705 ) );
  MUX \b/U1700  ( .IN0(\b/n1703 ), .IN1(\b/n1702 ), .SEL(msg[10]), .F(
        \b/n1704 ) );
  MUX \b/U1699  ( .IN0(\b/n1000 ), .IN1(\b/n1045 ), .SEL(msg[15]), .F(
        \b/n1703 ) );
  MUX \b/U1698  ( .IN0(\b/n1007 ), .IN1(\b/n1495 ), .SEL(msg[15]), .F(
        \b/n1702 ) );
  MUX \b/U1697  ( .IN0(\b/n1700 ), .IN1(\b/n1698 ), .SEL(msg[10]), .F(
        \b/n1701 ) );
  MUX \b/U1696  ( .IN0(\b/n1518 ), .IN1(\b/n1699 ), .SEL(msg[15]), .F(
        \b/n1700 ) );
  AND \b/U1695  ( .A(\b/n1495 ), .B(\b/n1063 ), .Z(\b/n1699 ) );
  MUX \b/U1694  ( .IN0(\b/n1020 ), .IN1(\b/n1039 ), .SEL(msg[15]), .F(
        \b/n1698 ) );
  MUX \b/U1693  ( .IN0(\b/n1696 ), .IN1(\b/n1693 ), .SEL(msg[13]), .F(
        \b/n1697 ) );
  MUX \b/U1692  ( .IN0(\b/n1695 ), .IN1(\b/n1694 ), .SEL(msg[10]), .F(
        \b/n1696 ) );
  MUX \b/U1691  ( .IN0(\b/n1008 ), .IN1(\b/n1533 ), .SEL(msg[15]), .F(
        \b/n1695 ) );
  MUX \b/U1690  ( .IN0(\b/n1032 ), .IN1(\b/n1521 ), .SEL(msg[15]), .F(
        \b/n1694 ) );
  MUX \b/U1689  ( .IN0(\b/n995 ), .IN1(\b/n1692 ), .SEL(msg[10]), .F(\b/n1693 ) );
  MUX \b/U1688  ( .IN0(\b/n1014 ), .IN1(\b/n1495 ), .SEL(msg[15]), .F(
        \b/n1692 ) );
  MUX \b/U1687  ( .IN0(\b/n1691 ), .IN1(\b/n1673 ), .SEL(msg[8]), .F(
        shift_row_out[107]) );
  MUX \b/U1686  ( .IN0(\b/n1690 ), .IN1(\b/n1682 ), .SEL(msg[14]), .F(
        \b/n1691 ) );
  MUX \b/U1685  ( .IN0(\b/n1689 ), .IN1(\b/n1686 ), .SEL(msg[13]), .F(
        \b/n1690 ) );
  MUX \b/U1684  ( .IN0(\b/n1688 ), .IN1(\b/n1687 ), .SEL(msg[15]), .F(
        \b/n1689 ) );
  MUX \b/U1683  ( .IN0(\b/n1513 ), .IN1(\b/n1039 ), .SEL(msg[10]), .F(
        \b/n1688 ) );
  MUX \b/U1682  ( .IN0(n612), .IN1(\b/n999 ), .SEL(msg[10]), .F(\b/n1687 ) );
  MUX \b/U1681  ( .IN0(\b/n1684 ), .IN1(\b/n1683 ), .SEL(msg[15]), .F(
        \b/n1686 ) );
  AND \b/U1680  ( .A(\b/n1685 ), .B(msg[12]), .Z(\b/n1684 ) );
  MUX \b/U1679  ( .IN0(\b/n1027 ), .IN1(\b/n1524 ), .SEL(msg[10]), .F(
        \b/n1683 ) );
  MUX \b/U1678  ( .IN0(\b/n1681 ), .IN1(\b/n1677 ), .SEL(msg[13]), .F(
        \b/n1682 ) );
  MUX \b/U1677  ( .IN0(\b/n1679 ), .IN1(\b/n1678 ), .SEL(msg[15]), .F(
        \b/n1681 ) );
  NAND \b/U1676  ( .A(\b/n1007 ), .B(\b/n1680 ), .Z(\b/n1679 ) );
  MUX \b/U1675  ( .IN0(\b/n1038 ), .IN1(\b/n1018 ), .SEL(msg[10]), .F(
        \b/n1678 ) );
  MUX \b/U1674  ( .IN0(\b/n1676 ), .IN1(\b/n1674 ), .SEL(msg[15]), .F(
        \b/n1677 ) );
  MUX \b/U1673  ( .IN0(\b/n1508 ), .IN1(\b/n1675 ), .SEL(msg[10]), .F(
        \b/n1676 ) );
  AND \b/U1672  ( .A(msg[9]), .B(\b/n1007 ), .Z(\b/n1675 ) );
  MUX \b/U1671  ( .IN0(\b/n1012 ), .IN1(\b/n1525 ), .SEL(msg[10]), .F(
        \b/n1674 ) );
  MUX \b/U1670  ( .IN0(\b/n1672 ), .IN1(\b/n1662 ), .SEL(msg[14]), .F(
        \b/n1673 ) );
  MUX \b/U1669  ( .IN0(\b/n1671 ), .IN1(\b/n1668 ), .SEL(msg[13]), .F(
        \b/n1672 ) );
  MUX \b/U1668  ( .IN0(\b/n1670 ), .IN1(\b/n1669 ), .SEL(msg[15]), .F(
        \b/n1671 ) );
  MUX \b/U1667  ( .IN0(\b/n1515 ), .IN1(n609), .SEL(msg[10]), .F(\b/n1670 ) );
  MUX \b/U1666  ( .IN0(\b/n997 ), .IN1(\b/n1014 ), .SEL(msg[10]), .F(\b/n1669 ) );
  MUX \b/U1665  ( .IN0(\b/n1664 ), .IN1(\b/n1665 ), .SEL(msg[15]), .F(
        \b/n1668 ) );
  NAND \b/U1664  ( .A(\b/n1666 ), .B(\b/n1667 ), .Z(\b/n1665 ) );
  MUX \b/U1663  ( .IN0(\b/n1040 ), .IN1(\b/n1663 ), .SEL(msg[10]), .F(
        \b/n1664 ) );
  MUX \b/U1662  ( .IN0(\b/n1015 ), .IN1(\b/n1058 ), .SEL(msg[9]), .F(\b/n1663 ) );
  MUX \b/U1661  ( .IN0(\b/n1661 ), .IN1(\b/n1655 ), .SEL(msg[13]), .F(
        \b/n1662 ) );
  MUX \b/U1660  ( .IN0(\b/n1660 ), .IN1(\b/n1658 ), .SEL(msg[15]), .F(
        \b/n1661 ) );
  MUX \b/U1659  ( .IN0(\b/n1659 ), .IN1(\b/n1497 ), .SEL(\b/n1543 ), .F(
        \b/n1660 ) );
  MUX \b/U1658  ( .IN0(msg[11]), .IN1(msg[12]), .SEL(msg[10]), .F(\b/n1659 )
         );
  MUX \b/U1657  ( .IN0(\b/n1525 ), .IN1(\b/n1656 ), .SEL(msg[10]), .F(
        \b/n1658 ) );
  NAND \b/U1656  ( .A(\b/n1497 ), .B(\b/n1657 ), .Z(\b/n1656 ) );
  MUX \b/U1655  ( .IN0(\b/n1652 ), .IN1(\b/n1653 ), .SEL(msg[15]), .F(
        \b/n1655 ) );
  AND \b/U1654  ( .A(\b/n1029 ), .B(\b/n1654 ), .Z(\b/n1653 ) );
  MUX \b/U1653  ( .IN0(\b/n1019 ), .IN1(\b/n1496 ), .SEL(msg[10]), .F(
        \b/n1652 ) );
  MUX \b/U1652  ( .IN0(\b/n1651 ), .IN1(\b/n1634 ), .SEL(msg[8]), .F(
        shift_row_out[106]) );
  MUX \b/U1651  ( .IN0(\b/n1650 ), .IN1(\b/n1642 ), .SEL(msg[14]), .F(
        \b/n1651 ) );
  MUX \b/U1650  ( .IN0(\b/n1649 ), .IN1(\b/n1645 ), .SEL(msg[13]), .F(
        \b/n1650 ) );
  MUX \b/U1649  ( .IN0(\b/n1648 ), .IN1(\b/n1646 ), .SEL(msg[10]), .F(
        \b/n1649 ) );
  MUX \b/U1648  ( .IN0(\b/n1027 ), .IN1(\b/n1647 ), .SEL(msg[15]), .F(
        \b/n1648 ) );
  MUX \b/U1647  ( .IN0(\b/n1495 ), .IN1(\b/n1007 ), .SEL(msg[9]), .F(\b/n1647 ) );
  MUX \b/U1646  ( .IN0(\b/n1542 ), .IN1(\b/n1035 ), .SEL(msg[15]), .F(
        \b/n1646 ) );
  MUX \b/U1645  ( .IN0(\b/n1644 ), .IN1(\b/n1643 ), .SEL(msg[10]), .F(
        \b/n1645 ) );
  MUX \b/U1644  ( .IN0(\b/n1496 ), .IN1(\b/n996 ), .SEL(msg[15]), .F(\b/n1644 ) );
  MUX \b/U1643  ( .IN0(\b/n1048 ), .IN1(\b/n1498 ), .SEL(msg[15]), .F(
        \b/n1643 ) );
  MUX \b/U1642  ( .IN0(\b/n1641 ), .IN1(\b/n1638 ), .SEL(msg[13]), .F(
        \b/n1642 ) );
  MUX \b/U1641  ( .IN0(\b/n1640 ), .IN1(\b/n1639 ), .SEL(msg[10]), .F(
        \b/n1641 ) );
  MUX \b/U1640  ( .IN0(\b/n1036 ), .IN1(msg[9]), .SEL(msg[15]), .F(\b/n1640 )
         );
  MUX \b/U1639  ( .IN0(n614), .IN1(\b/n1511 ), .SEL(msg[15]), .F(\b/n1639 ) );
  MUX \b/U1638  ( .IN0(\b/n1637 ), .IN1(\b/n1636 ), .SEL(msg[10]), .F(
        \b/n1638 ) );
  MUX \b/U1637  ( .IN0(\b/n1060 ), .IN1(\b/n1034 ), .SEL(msg[15]), .F(
        \b/n1637 ) );
  MUX \b/U1636  ( .IN0(n614), .IN1(\b/n1635 ), .SEL(msg[15]), .F(\b/n1636 ) );
  MUX \b/U1635  ( .IN0(\b/n1007 ), .IN1(\b/n1042 ), .SEL(msg[9]), .F(\b/n1635 ) );
  MUX \b/U1634  ( .IN0(\b/n1633 ), .IN1(\b/n1626 ), .SEL(msg[14]), .F(
        \b/n1634 ) );
  MUX \b/U1633  ( .IN0(\b/n1632 ), .IN1(\b/n1628 ), .SEL(msg[13]), .F(
        \b/n1633 ) );
  MUX \b/U1632  ( .IN0(\b/n1629 ), .IN1(\b/n995 ), .SEL(msg[10]), .F(\b/n1632 ) );
  NAND \b/U1631  ( .A(\b/n1630 ), .B(\b/n1631 ), .Z(\b/n1629 ) );
  MUX \b/U1630  ( .IN0(n611), .IN1(\b/n1627 ), .SEL(\b/n1541 ), .F(\b/n1628 )
         );
  MUX \b/U1629  ( .IN0(\b/n1026 ), .IN1(\b/n1510 ), .SEL(msg[10]), .F(
        \b/n1627 ) );
  MUX \b/U1628  ( .IN0(\b/n1625 ), .IN1(\b/n1619 ), .SEL(msg[13]), .F(
        \b/n1626 ) );
  MUX \b/U1627  ( .IN0(\b/n1622 ), .IN1(\b/n1621 ), .SEL(msg[10]), .F(
        \b/n1625 ) );
  NAND \b/U1626  ( .A(\b/n1623 ), .B(\b/n1624 ), .Z(\b/n1622 ) );
  MUX \b/U1625  ( .IN0(\b/n1497 ), .IN1(\b/n1620 ), .SEL(n613), .F(\b/n1621 )
         );
  MUX \b/U1624  ( .IN0(msg[11]), .IN1(\b/n1015 ), .SEL(msg[15]), .F(\b/n1620 )
         );
  MUX \b/U1623  ( .IN0(\b/n1618 ), .IN1(\b/n1617 ), .SEL(msg[10]), .F(
        \b/n1619 ) );
  MUX \b/U1622  ( .IN0(\b/n1540 ), .IN1(\b/n1013 ), .SEL(msg[15]), .F(
        \b/n1618 ) );
  MUX \b/U1621  ( .IN0(\b/n1499 ), .IN1(\b/n1616 ), .SEL(msg[15]), .F(
        \b/n1617 ) );
  MUX \b/U1620  ( .IN0(\b/n1501 ), .IN1(\b/n1495 ), .SEL(msg[9]), .F(\b/n1616 ) );
  MUX \b/U1619  ( .IN0(\b/n1615 ), .IN1(\b/n1597 ), .SEL(msg[8]), .F(
        shift_row_out[105]) );
  MUX \b/U1618  ( .IN0(\b/n1614 ), .IN1(\b/n1605 ), .SEL(msg[14]), .F(
        \b/n1615 ) );
  MUX \b/U1617  ( .IN0(\b/n1613 ), .IN1(\b/n1609 ), .SEL(msg[13]), .F(
        \b/n1614 ) );
  MUX \b/U1616  ( .IN0(\b/n1612 ), .IN1(\b/n1611 ), .SEL(msg[10]), .F(
        \b/n1613 ) );
  MUX \b/U1615  ( .IN0(\b/n1031 ), .IN1(n616), .SEL(msg[15]), .F(\b/n1612 ) );
  MUX \b/U1614  ( .IN0(\b/n1610 ), .IN1(n610), .SEL(msg[15]), .F(\b/n1611 ) );
  NAND \b/U1613  ( .A(\b/n1063 ), .B(\b/n1021 ), .Z(\b/n1610 ) );
  MUX \b/U1612  ( .IN0(\b/n1608 ), .IN1(\b/n1607 ), .SEL(msg[10]), .F(
        \b/n1609 ) );
  MUX \b/U1611  ( .IN0(\b/n1000 ), .IN1(\b/n1512 ), .SEL(msg[15]), .F(
        \b/n1608 ) );
  MUX \b/U1610  ( .IN0(\b/n1519 ), .IN1(\b/n1606 ), .SEL(msg[15]), .F(
        \b/n1607 ) );
  AND \b/U1609  ( .A(msg[9]), .B(msg[12]), .Z(\b/n1606 ) );
  MUX \b/U1608  ( .IN0(\b/n1604 ), .IN1(\b/n1600 ), .SEL(msg[13]), .F(
        \b/n1605 ) );
  MUX \b/U1607  ( .IN0(\b/n1603 ), .IN1(\b/n1602 ), .SEL(msg[10]), .F(
        \b/n1604 ) );
  MUX \b/U1606  ( .IN0(\b/n1503 ), .IN1(\b/n1023 ), .SEL(msg[15]), .F(
        \b/n1603 ) );
  MUX \b/U1605  ( .IN0(\b/n1601 ), .IN1(\b/n1009 ), .SEL(msg[15]), .F(
        \b/n1602 ) );
  MUX \b/U1604  ( .IN0(\b/n1519 ), .IN1(\b/n1015 ), .SEL(msg[9]), .F(\b/n1601 ) );
  MUX \b/U1603  ( .IN0(\b/n1599 ), .IN1(\b/n1598 ), .SEL(msg[10]), .F(
        \b/n1600 ) );
  MUX \b/U1602  ( .IN0(\b/n1036 ), .IN1(\b/n1052 ), .SEL(msg[15]), .F(
        \b/n1599 ) );
  MUX \b/U1601  ( .IN0(\b/n1031 ), .IN1(\b/n1012 ), .SEL(msg[15]), .F(
        \b/n1598 ) );
  MUX \b/U1600  ( .IN0(\b/n1596 ), .IN1(\b/n1588 ), .SEL(msg[14]), .F(
        \b/n1597 ) );
  MUX \b/U1599  ( .IN0(\b/n1595 ), .IN1(\b/n1592 ), .SEL(msg[13]), .F(
        \b/n1596 ) );
  MUX \b/U1598  ( .IN0(\b/n1594 ), .IN1(\b/n1593 ), .SEL(msg[10]), .F(
        \b/n1595 ) );
  MUX \b/U1597  ( .IN0(\b/n1539 ), .IN1(\b/n1060 ), .SEL(msg[15]), .F(
        \b/n1594 ) );
  MUX \b/U1596  ( .IN0(\b/n1053 ), .IN1(\b/n1510 ), .SEL(msg[15]), .F(
        \b/n1593 ) );
  MUX \b/U1595  ( .IN0(\b/n1589 ), .IN1(\b/n1590 ), .SEL(msg[10]), .F(
        \b/n1592 ) );
  AND \b/U1594  ( .A(\b/n1591 ), .B(\b/n1564 ), .Z(\b/n1590 ) );
  MUX \b/U1593  ( .IN0(\b/n1514 ), .IN1(\b/n1495 ), .SEL(msg[15]), .F(
        \b/n1589 ) );
  MUX \b/U1592  ( .IN0(\b/n1587 ), .IN1(\b/n1582 ), .SEL(msg[13]), .F(
        \b/n1588 ) );
  MUX \b/U1591  ( .IN0(\b/n1586 ), .IN1(\b/n1583 ), .SEL(msg[10]), .F(
        \b/n1587 ) );
  MUX \b/U1590  ( .IN0(\b/n1584 ), .IN1(\b/n1585 ), .SEL(msg[15]), .F(
        \b/n1586 ) );
  NAND \b/U1589  ( .A(\b/n1495 ), .B(\b/n1575 ), .Z(\b/n1585 ) );
  MUX \b/U1588  ( .IN0(\b/n1495 ), .IN1(\b/n1015 ), .SEL(msg[9]), .F(\b/n1584 ) );
  MUX \b/U1587  ( .IN0(\b/n1538 ), .IN1(\b/n1520 ), .SEL(msg[15]), .F(
        \b/n1583 ) );
  MUX \b/U1586  ( .IN0(\b/n1537 ), .IN1(\b/n1581 ), .SEL(msg[10]), .F(
        \b/n1582 ) );
  MUX \b/U1585  ( .IN0(\b/n1021 ), .IN1(\b/n1034 ), .SEL(msg[15]), .F(
        \b/n1581 ) );
  MUX \b/U1584  ( .IN0(\b/n1580 ), .IN1(\b/n1561 ), .SEL(msg[8]), .F(
        shift_row_out[104]) );
  MUX \b/U1583  ( .IN0(\b/n1579 ), .IN1(\b/n1571 ), .SEL(msg[14]), .F(
        \b/n1580 ) );
  MUX \b/U1582  ( .IN0(\b/n1578 ), .IN1(\b/n1576 ), .SEL(msg[10]), .F(
        \b/n1579 ) );
  MUX \b/U1581  ( .IN0(\b/n997 ), .IN1(\b/n1577 ), .SEL(msg[15]), .F(\b/n1578 ) );
  MUX \b/U1580  ( .IN0(\b/n1048 ), .IN1(\b/n1032 ), .SEL(msg[13]), .F(
        \b/n1577 ) );
  MUX \b/U1579  ( .IN0(\b/n1573 ), .IN1(\b/n1572 ), .SEL(msg[15]), .F(
        \b/n1576 ) );
  NAND \b/U1578  ( .A(\b/n1574 ), .B(\b/n1575 ), .Z(\b/n1573 ) );
  MUX \b/U1577  ( .IN0(\b/n1047 ), .IN1(\b/n1063 ), .SEL(msg[13]), .F(
        \b/n1572 ) );
  MUX \b/U1576  ( .IN0(\b/n1570 ), .IN1(\b/n1566 ), .SEL(msg[10]), .F(
        \b/n1571 ) );
  MUX \b/U1575  ( .IN0(\b/n1569 ), .IN1(\b/n1568 ), .SEL(msg[15]), .F(
        \b/n1570 ) );
  MUX \b/U1574  ( .IN0(n609), .IN1(\b/n1003 ), .SEL(msg[13]), .F(\b/n1569 ) );
  MUX \b/U1573  ( .IN0(\b/n1567 ), .IN1(\b/n1029 ), .SEL(msg[13]), .F(
        \b/n1568 ) );
  NAND \b/U1572  ( .A(\b/n1494 ), .B(\b/n1496 ), .Z(\b/n1567 ) );
  MUX \b/U1571  ( .IN0(\b/n1565 ), .IN1(\b/n1562 ), .SEL(msg[15]), .F(
        \b/n1566 ) );
  MUX \b/U1570  ( .IN0(\b/n1010 ), .IN1(\b/n1563 ), .SEL(msg[13]), .F(
        \b/n1565 ) );
  NAND \b/U1569  ( .A(\b/n1501 ), .B(\b/n1564 ), .Z(\b/n1563 ) );
  MUX \b/U1568  ( .IN0(\b/n1054 ), .IN1(\b/n1504 ), .SEL(msg[13]), .F(
        \b/n1562 ) );
  MUX \b/U1567  ( .IN0(\b/n1560 ), .IN1(\b/n1552 ), .SEL(msg[14]), .F(
        \b/n1561 ) );
  MUX \b/U1566  ( .IN0(\b/n1559 ), .IN1(\b/n1555 ), .SEL(msg[10]), .F(
        \b/n1560 ) );
  MUX \b/U1565  ( .IN0(\b/n1558 ), .IN1(\b/n1556 ), .SEL(msg[15]), .F(
        \b/n1559 ) );
  MUX \b/U1564  ( .IN0(\b/n1557 ), .IN1(\b/n1002 ), .SEL(msg[13]), .F(
        \b/n1558 ) );
  NAND \b/U1563  ( .A(\b/n1063 ), .B(\b/n1497 ), .Z(\b/n1557 ) );
  MUX \b/U1561  ( .IN0(\b/n1554 ), .IN1(\b/n1553 ), .SEL(msg[15]), .F(
        \b/n1555 ) );
  MUX \b/U1560  ( .IN0(n611), .IN1(\b/n999 ), .SEL(msg[13]), .F(\b/n1554 ) );
  MUX \b/U1559  ( .IN0(\b/n1030 ), .IN1(\b/n1007 ), .SEL(msg[13]), .F(
        \b/n1553 ) );
  MUX \b/U1558  ( .IN0(\b/n1551 ), .IN1(\b/n1547 ), .SEL(msg[10]), .F(
        \b/n1552 ) );
  MUX \b/U1557  ( .IN0(\b/n1549 ), .IN1(\b/n1548 ), .SEL(msg[15]), .F(
        \b/n1551 ) );
  NAND \b/U1556  ( .A(\b/n1550 ), .B(\b/n1536 ), .Z(\b/n1549 ) );
  MUX \b/U1555  ( .IN0(msg[11]), .IN1(\b/n1498 ), .SEL(msg[13]), .F(\b/n1548 )
         );
  MUX \b/U1554  ( .IN0(\b/n1546 ), .IN1(\b/n1545 ), .SEL(msg[15]), .F(
        \b/n1547 ) );
  MUX \b/U1553  ( .IN0(\b/n1013 ), .IN1(\b/n1507 ), .SEL(msg[13]), .F(
        \b/n1546 ) );
  MUX \b/U1552  ( .IN0(\b/n1046 ), .IN1(\b/n1053 ), .SEL(msg[13]), .F(
        \b/n1545 ) );
  XOR \b/U1551  ( .A(\b/n1497 ), .B(msg[9]), .Z(\b/n1544 ) );
  XOR \b/U1550  ( .A(msg[10]), .B(msg[9]), .Z(\b/n1543 ) );
  XOR \b/U1549  ( .A(msg[11]), .B(msg[9]), .Z(\b/n1542 ) );
  XOR \b/U1548  ( .A(msg[10]), .B(msg[15]), .Z(\b/n1541 ) );
  XOR \b/U1547  ( .A(\b/n1063 ), .B(\b/n1007 ), .Z(\b/n1540 ) );
  XOR \b/U1546  ( .A(msg[9]), .B(\b/n1032 ), .Z(\b/n1539 ) );
  XOR \b/U1545  ( .A(\b/n1063 ), .B(msg[12]), .Z(\b/n1538 ) );
  XOR \b/U1543  ( .A(\b/n1015 ), .B(msg[11]), .Z(\b/n1519 ) );
  XOR \b/U1542  ( .A(msg[13]), .B(msg[9]), .Z(\b/n1536 ) );
  MUX \b/U1541  ( .IN0(\b/n1497 ), .IN1(\b/n1007 ), .SEL(msg[9]), .F(\b/n1535 ) );
  NANDN \b/U1539  ( .B(msg[11]), .A(msg[9]), .Z(\b/n1533 ) );
  MUX \b/U1538  ( .IN0(\b/n1021 ), .IN1(\b/n1042 ), .SEL(msg[9]), .F(\b/n1532 ) );
  MUX \b/U1537  ( .IN0(msg[11]), .IN1(\b/n1042 ), .SEL(msg[9]), .F(\b/n1531 )
         );
  MUX \b/U1536  ( .IN0(\b/n1501 ), .IN1(\b/n1519 ), .SEL(msg[9]), .F(\b/n1530 ) );
  MUX \b/U1535  ( .IN0(msg[12]), .IN1(\b/n1021 ), .SEL(msg[9]), .F(\b/n1529 )
         );
  NAND \b/U1534  ( .A(\b/n1042 ), .B(\b/n1063 ), .Z(\b/n1528 ) );
  MUX \b/U1532  ( .IN0(\b/n1042 ), .IN1(msg[12]), .SEL(msg[9]), .F(\b/n1526 )
         );
  MUX \b/U1531  ( .IN0(\b/n1494 ), .IN1(\b/n1495 ), .SEL(msg[9]), .F(\b/n1525 ) );
  MUX \b/U1530  ( .IN0(\b/n1058 ), .IN1(msg[12]), .SEL(msg[9]), .F(\b/n1524 )
         );
  MUX \b/U1529  ( .IN0(\b/n1015 ), .IN1(\b/n1042 ), .SEL(msg[9]), .F(\b/n1523 ) );
  MUX \b/U1528  ( .IN0(\b/n1494 ), .IN1(msg[12]), .SEL(msg[9]), .F(\b/n1522 )
         );
  MUX \b/U1527  ( .IN0(\b/n1052 ), .IN1(\b/n1021 ), .SEL(msg[9]), .F(\b/n1521 ) );
  NANDN \b/U1526  ( .B(msg[9]), .A(msg[11]), .Z(\b/n1520 ) );
  MUX \b/U1525  ( .IN0(\b/n1519 ), .IN1(\b/n1052 ), .SEL(msg[9]), .F(\b/n1518 ) );
  MUX \b/U1524  ( .IN0(\b/n1007 ), .IN1(msg[11]), .SEL(msg[9]), .F(\b/n1517 )
         );
  NAND \b/U1522  ( .A(\b/n1501 ), .B(\b/n1063 ), .Z(\b/n1515 ) );
  MUX \b/U1521  ( .IN0(msg[12]), .IN1(\b/n1497 ), .SEL(msg[9]), .F(\b/n1514 )
         );
  MUX \b/U1520  ( .IN0(msg[12]), .IN1(\b/n1032 ), .SEL(msg[9]), .F(\b/n1513 )
         );
  MUX \b/U1519  ( .IN0(\b/n1007 ), .IN1(\b/n1058 ), .SEL(msg[9]), .F(\b/n1512 ) );
  NAND \b/U1518  ( .A(\b/n1496 ), .B(\b/n1007 ), .Z(\b/n1511 ) );
  MUX \b/U1517  ( .IN0(\b/n1497 ), .IN1(\b/n1495 ), .SEL(msg[9]), .F(\b/n1510 ) );
  NAND \b/U1516  ( .A(\b/n1509 ), .B(\b/n1494 ), .Z(\b/n1508 ) );
  MUX \b/U1515  ( .IN0(\b/n1497 ), .IN1(\b/n1058 ), .SEL(msg[9]), .F(\b/n1507 ) );
  NANDN \b/U1513  ( .B(msg[12]), .A(msg[11]), .Z(\b/n1497 ) );
  MUX \b/U1512  ( .IN0(\b/n1501 ), .IN1(\b/n1058 ), .SEL(msg[9]), .F(\b/n1505 ) );
  MUX \b/U1511  ( .IN0(\b/n1058 ), .IN1(\b/n1021 ), .SEL(msg[9]), .F(\b/n1504 ) );
  MUX \b/U1510  ( .IN0(\b/n1501 ), .IN1(msg[11]), .SEL(msg[9]), .F(\b/n1503 )
         );
  OR \b/U1509  ( .A(msg[11]), .B(msg[12]), .Z(\b/n1501 ) );
  MUX \b/U1508  ( .IN0(\b/n1007 ), .IN1(\b/n1021 ), .SEL(msg[9]), .F(\b/n1502 ) );
  NAND \b/U1507  ( .A(\b/n1501 ), .B(\b/n1496 ), .Z(\b/n1500 ) );
  NAND \b/U1506  ( .A(msg[11]), .B(msg[9]), .Z(\b/n1499 ) );
  OR \b/U1505  ( .A(msg[9]), .B(msg[12]), .Z(\b/n1498 ) );
  NAND \b/U1504  ( .A(msg[9]), .B(\b/n1497 ), .Z(\b/n1496 ) );
  NANDN \b/U1503  ( .B(msg[11]), .A(msg[12]), .Z(\b/n1495 ) );
  NAND \b/U1502  ( .A(msg[11]), .B(msg[12]), .Z(\b/n1494 ) );
  MUX \b/U1501  ( .IN0(msg[4]), .IN1(\b/n1135 ), .SEL(msg[1]), .F(\b/n1493 )
         );
  MUX \b/U1500  ( .IN0(msg[4]), .IN1(\b/n1144 ), .SEL(msg[1]), .F(\b/n1492 )
         );
  MUX \b/U1499  ( .IN0(\b/n1136 ), .IN1(\b/n1139 ), .SEL(msg[1]), .F(\b/n1491 ) );
  MUX \b/U1498  ( .IN0(\b/n1141 ), .IN1(\b/n1123 ), .SEL(msg[1]), .F(\b/n1490 ) );
  MUX \b/U1496  ( .IN0(\b/n1144 ), .IN1(\b/n1135 ), .SEL(msg[2]), .F(\b/n1317 ) );
  MUX \b/U1495  ( .IN0(\b/n1137 ), .IN1(\b/n1134 ), .SEL(msg[2]), .F(\b/n1318 ) );
  MUX \b/U1494  ( .IN0(\b/n1077 ), .IN1(\b/n1087 ), .SEL(msg[1]), .F(\b/n1281 ) );
  MUX \b/U1493  ( .IN0(\b/n1165 ), .IN1(\b/n1476 ), .SEL(msg[7]), .F(\b/n1488 ) );
  MUX \b/U1492  ( .IN0(\b/n1139 ), .IN1(\b/n1135 ), .SEL(msg[1]), .F(\b/n1479 ) );
  MUX \b/U1491  ( .IN0(\b/n1129 ), .IN1(\b/n1141 ), .SEL(msg[1]), .F(\b/n1487 ) );
  MUX \b/U1490  ( .IN0(msg[3]), .IN1(\b/n1123 ), .SEL(msg[1]), .F(\b/n1486 )
         );
  MUX \b/U1489  ( .IN0(\b/n1144 ), .IN1(\b/n1129 ), .SEL(msg[1]), .F(\b/n1485 ) );
  MUX \b/U1488  ( .IN0(msg[4]), .IN1(\b/n1141 ), .SEL(msg[1]), .F(\b/n1484 )
         );
  MUX \b/U1487  ( .IN0(\b/n1114 ), .IN1(\b/n1093 ), .SEL(msg[5]), .F(\b/n1191 ) );
  MUX \b/U1486  ( .IN0(\b/n1136 ), .IN1(\b/n1087 ), .SEL(msg[1]), .F(\b/n1483 ) );
  NANDN \b/U1483  ( .B(\b/n1142 ), .A(msg[7]), .Z(\b/n1456 ) );
  NAND \b/U1482  ( .A(msg[7]), .B(\b/n1090 ), .Z(\b/n1424 ) );
  NAND \b/U1481  ( .A(msg[7]), .B(\b/n1102 ), .Z(\b/n1365 ) );
  NAND \b/U1480  ( .A(msg[7]), .B(\b/n1473 ), .Z(\b/n1398 ) );
  NAND \b/U1479  ( .A(msg[7]), .B(\b/n1393 ), .Z(\b/n1356 ) );
  NAND \b/U1477  ( .A(\b/n1134 ), .B(\b/n1123 ), .Z(\b/n1477 ) );
  NAND \b/U1476  ( .A(msg[7]), .B(\b/n1475 ), .Z(\b/n1470 ) );
  NAND \b/U1475  ( .A(n608), .B(msg[7]), .Z(\b/n1450 ) );
  NAND \b/U1473  ( .A(msg[2]), .B(\b/n1144 ), .Z(\b/n1310 ) );
  NAND \b/U1472  ( .A(\b/n1123 ), .B(msg[1]), .Z(\b/n1265 ) );
  NAND \b/U1471  ( .A(msg[7]), .B(\b/n1479 ), .Z(\b/n1264 ) );
  NAND \b/U1469  ( .A(\b/n1477 ), .B(msg[7]), .Z(\b/n1280 ) );
  NAND \b/U1468  ( .A(\b/n1298 ), .B(\b/n1144 ), .Z(\b/n1476 ) );
  NANDN \b/U1467  ( .B(\b/n1077 ), .A(\b/n1134 ), .Z(\b/n1475 ) );
  NAND \b/U1465  ( .A(msg[1]), .B(\b/n1144 ), .Z(\b/n1196 ) );
  NAND \b/U1464  ( .A(\b/n1077 ), .B(\b/n1134 ), .Z(\b/n1473 ) );
  NAND \b/U1461  ( .A(msg[1]), .B(\b/n1139 ), .Z(\b/n1298 ) );
  ANDN \b/U1459  ( .A(msg[2]), .B(msg[1]), .Z(\b/n1326 ) );
  AND \b/U1458  ( .A(\b/n1136 ), .B(\b/n1470 ), .Z(\b/n1241 ) );
  MUX \b/U1457  ( .IN0(\b/n1469 ), .IN1(\b/n1453 ), .SEL(msg[6]), .F(
        shift_row_out[7]) );
  MUX \b/U1456  ( .IN0(\b/n1468 ), .IN1(\b/n1461 ), .SEL(msg[0]), .F(\b/n1469 ) );
  MUX \b/U1455  ( .IN0(\b/n1467 ), .IN1(\b/n1464 ), .SEL(msg[5]), .F(\b/n1468 ) );
  MUX \b/U1454  ( .IN0(\b/n1466 ), .IN1(\b/n1465 ), .SEL(msg[2]), .F(\b/n1467 ) );
  MUX \b/U1453  ( .IN0(msg[4]), .IN1(\b/n1094 ), .SEL(msg[7]), .F(\b/n1466 )
         );
  MUX \b/U1452  ( .IN0(\b/n1137 ), .IN1(\b/n1098 ), .SEL(msg[7]), .F(\b/n1465 ) );
  MUX \b/U1451  ( .IN0(\b/n1463 ), .IN1(\b/n1462 ), .SEL(msg[2]), .F(\b/n1464 ) );
  MUX \b/U1450  ( .IN0(\b/n1195 ), .IN1(\b/n1090 ), .SEL(msg[7]), .F(\b/n1463 ) );
  MUX \b/U1449  ( .IN0(\b/n1147 ), .IN1(\b/n1158 ), .SEL(msg[7]), .F(\b/n1462 ) );
  MUX \b/U1448  ( .IN0(\b/n1460 ), .IN1(\b/n1457 ), .SEL(msg[5]), .F(\b/n1461 ) );
  MUX \b/U1447  ( .IN0(\b/n1459 ), .IN1(\b/n1458 ), .SEL(msg[2]), .F(\b/n1460 ) );
  MUX \b/U1446  ( .IN0(\b/n1171 ), .IN1(\b/n1146 ), .SEL(msg[7]), .F(\b/n1459 ) );
  MUX \b/U1445  ( .IN0(\b/n1102 ), .IN1(\b/n1167 ), .SEL(msg[7]), .F(\b/n1458 ) );
  MUX \b/U1444  ( .IN0(\b/n1455 ), .IN1(\b/n1454 ), .SEL(msg[2]), .F(\b/n1457 ) );
  AND \b/U1443  ( .A(\b/n1092 ), .B(\b/n1456 ), .Z(\b/n1455 ) );
  MUX \b/U1442  ( .IN0(\b/n1151 ), .IN1(n607), .SEL(msg[7]), .F(\b/n1454 ) );
  MUX \b/U1441  ( .IN0(\b/n1452 ), .IN1(\b/n1444 ), .SEL(msg[0]), .F(\b/n1453 ) );
  MUX \b/U1440  ( .IN0(\b/n1451 ), .IN1(\b/n1447 ), .SEL(msg[5]), .F(\b/n1452 ) );
  MUX \b/U1439  ( .IN0(\b/n1448 ), .IN1(\b/n1449 ), .SEL(msg[2]), .F(\b/n1451 ) );
  NAND \b/U1438  ( .A(\b/n1265 ), .B(\b/n1450 ), .Z(\b/n1449 ) );
  MUX \b/U1437  ( .IN0(\b/n1132 ), .IN1(\b/n1124 ), .SEL(msg[7]), .F(\b/n1448 ) );
  MUX \b/U1436  ( .IN0(\b/n1446 ), .IN1(\b/n1445 ), .SEL(msg[2]), .F(\b/n1447 ) );
  MUX \b/U1435  ( .IN0(\b/n1141 ), .IN1(\b/n1135 ), .SEL(msg[7]), .F(\b/n1446 ) );
  MUX \b/U1434  ( .IN0(\b/n1125 ), .IN1(\b/n1172 ), .SEL(msg[7]), .F(\b/n1445 ) );
  MUX \b/U1433  ( .IN0(\b/n1443 ), .IN1(\b/n1440 ), .SEL(msg[5]), .F(\b/n1444 ) );
  MUX \b/U1432  ( .IN0(\b/n1442 ), .IN1(\b/n1441 ), .SEL(msg[2]), .F(\b/n1443 ) );
  MUX \b/U1431  ( .IN0(\b/n1176 ), .IN1(\b/n1162 ), .SEL(msg[7]), .F(\b/n1442 ) );
  MUX \b/U1430  ( .IN0(\b/n1078 ), .IN1(\b/n1144 ), .SEL(msg[7]), .F(\b/n1441 ) );
  MUX \b/U1429  ( .IN0(\b/n1439 ), .IN1(\b/n1438 ), .SEL(msg[2]), .F(\b/n1440 ) );
  MUX \b/U1428  ( .IN0(\b/n1177 ), .IN1(\b/n1185 ), .SEL(msg[7]), .F(\b/n1439 ) );
  MUX \b/U1427  ( .IN0(\b/n1170 ), .IN1(\b/n1437 ), .SEL(msg[7]), .F(\b/n1438 ) );
  MUX \b/U1426  ( .IN0(\b/n1129 ), .IN1(\b/n1087 ), .SEL(msg[1]), .F(\b/n1437 ) );
  MUX \b/U1425  ( .IN0(\b/n1436 ), .IN1(\b/n1418 ), .SEL(msg[6]), .F(
        shift_row_out[6]) );
  MUX \b/U1424  ( .IN0(\b/n1435 ), .IN1(\b/n1426 ), .SEL(msg[0]), .F(\b/n1436 ) );
  MUX \b/U1423  ( .IN0(\b/n1434 ), .IN1(\b/n1429 ), .SEL(msg[5]), .F(\b/n1435 ) );
  MUX \b/U1422  ( .IN0(\b/n1433 ), .IN1(\b/n1431 ), .SEL(msg[2]), .F(\b/n1434 ) );
  MUX \b/U1421  ( .IN0(\b/n1432 ), .IN1(\b/n1148 ), .SEL(msg[7]), .F(\b/n1433 ) );
  MUX \b/U1420  ( .IN0(\b/n1129 ), .IN1(\b/n1135 ), .SEL(msg[1]), .F(\b/n1432 ) );
  MUX \b/U1419  ( .IN0(\b/n1430 ), .IN1(\b/n1117 ), .SEL(msg[7]), .F(\b/n1431 ) );
  MUX \b/U1418  ( .IN0(\b/n1135 ), .IN1(\b/n1136 ), .SEL(msg[1]), .F(\b/n1430 ) );
  MUX \b/U1417  ( .IN0(\b/n1428 ), .IN1(\b/n1427 ), .SEL(msg[2]), .F(\b/n1429 ) );
  MUX \b/U1416  ( .IN0(n606), .IN1(\b/n1216 ), .SEL(msg[7]), .F(\b/n1428 ) );
  MUX \b/U1415  ( .IN0(\b/n1174 ), .IN1(\b/n1181 ), .SEL(msg[7]), .F(\b/n1427 ) );
  MUX \b/U1414  ( .IN0(\b/n1425 ), .IN1(\b/n1421 ), .SEL(msg[5]), .F(\b/n1426 ) );
  MUX \b/U1413  ( .IN0(\b/n1423 ), .IN1(\b/n1422 ), .SEL(msg[2]), .F(\b/n1425 ) );
  AND \b/U1412  ( .A(\b/n1070 ), .B(\b/n1424 ), .Z(\b/n1423 ) );
  MUX \b/U1411  ( .IN0(\b/n1251 ), .IN1(msg[3]), .SEL(msg[7]), .F(\b/n1422 )
         );
  MUX \b/U1410  ( .IN0(\b/n1420 ), .IN1(\b/n1419 ), .SEL(msg[2]), .F(\b/n1421 ) );
  MUX \b/U1409  ( .IN0(\b/n1113 ), .IN1(\b/n1139 ), .SEL(msg[7]), .F(\b/n1420 ) );
  MUX \b/U1407  ( .IN0(\b/n1417 ), .IN1(\b/n1410 ), .SEL(msg[0]), .F(\b/n1418 ) );
  MUX \b/U1406  ( .IN0(\b/n1416 ), .IN1(\b/n1413 ), .SEL(msg[5]), .F(\b/n1417 ) );
  MUX \b/U1405  ( .IN0(\b/n1415 ), .IN1(\b/n1414 ), .SEL(msg[2]), .F(\b/n1416 ) );
  MUX \b/U1404  ( .IN0(\b/n1109 ), .IN1(\b/n1143 ), .SEL(msg[7]), .F(\b/n1415 ) );
  MUX \b/U1403  ( .IN0(\b/n1147 ), .IN1(n607), .SEL(msg[7]), .F(\b/n1414 ) );
  MUX \b/U1402  ( .IN0(\b/n1412 ), .IN1(\b/n1411 ), .SEL(msg[2]), .F(\b/n1413 ) );
  MUX \b/U1401  ( .IN0(\b/n1163 ), .IN1(\b/n1074 ), .SEL(msg[7]), .F(\b/n1412 ) );
  MUX \b/U1400  ( .IN0(\b/n1094 ), .IN1(\b/n1124 ), .SEL(msg[7]), .F(\b/n1411 ) );
  MUX \b/U1399  ( .IN0(\b/n1409 ), .IN1(\b/n1405 ), .SEL(msg[5]), .F(\b/n1410 ) );
  MUX \b/U1398  ( .IN0(\b/n1408 ), .IN1(\b/n1407 ), .SEL(msg[2]), .F(\b/n1409 ) );
  MUX \b/U1397  ( .IN0(\b/n1152 ), .IN1(\b/n1124 ), .SEL(msg[7]), .F(\b/n1408 ) );
  MUX \b/U1396  ( .IN0(\b/n1406 ), .IN1(\b/n1173 ), .SEL(msg[7]), .F(\b/n1407 ) );
  NANDN \b/U1395  ( .B(msg[4]), .A(msg[1]), .Z(\b/n1406 ) );
  MUX \b/U1394  ( .IN0(\b/n1404 ), .IN1(\b/n1402 ), .SEL(msg[2]), .F(\b/n1405 ) );
  MUX \b/U1393  ( .IN0(\b/n1087 ), .IN1(\b/n1403 ), .SEL(msg[7]), .F(\b/n1404 ) );
  MUX \b/U1392  ( .IN0(\b/n1114 ), .IN1(\b/n1104 ), .SEL(msg[1]), .F(\b/n1403 ) );
  MUX \b/U1391  ( .IN0(\b/n1076 ), .IN1(\b/n1148 ), .SEL(msg[7]), .F(\b/n1402 ) );
  NANDN \b/U1390  ( .B(\b/n1077 ), .A(msg[1]), .Z(\b/n1148 ) );
  MUX \b/U1389  ( .IN0(\b/n1401 ), .IN1(\b/n1380 ), .SEL(msg[6]), .F(
        shift_row_out[5]) );
  MUX \b/U1388  ( .IN0(\b/n1400 ), .IN1(\b/n1390 ), .SEL(msg[0]), .F(\b/n1401 ) );
  MUX \b/U1387  ( .IN0(\b/n1399 ), .IN1(\b/n1395 ), .SEL(msg[5]), .F(\b/n1400 ) );
  MUX \b/U1386  ( .IN0(\b/n1396 ), .IN1(\b/n1397 ), .SEL(msg[2]), .F(\b/n1399 ) );
  AND \b/U1385  ( .A(\b/n1166 ), .B(\b/n1398 ), .Z(\b/n1397 ) );
  MUX \b/U1384  ( .IN0(\b/n1144 ), .IN1(\b/n1125 ), .SEL(msg[7]), .F(\b/n1396 ) );
  MUX \b/U1383  ( .IN0(\b/n1394 ), .IN1(\b/n1392 ), .SEL(msg[2]), .F(\b/n1395 ) );
  MUX \b/U1382  ( .IN0(\b/n1080 ), .IN1(\b/n1393 ), .SEL(msg[7]), .F(\b/n1394 ) );
  NAND \b/U1381  ( .A(\b/n1104 ), .B(\b/n1134 ), .Z(\b/n1393 ) );
  MUX \b/U1380  ( .IN0(\b/n1144 ), .IN1(\b/n1391 ), .SEL(msg[7]), .F(\b/n1392 ) );
  NAND \b/U1379  ( .A(\b/n1135 ), .B(\b/n1196 ), .Z(\b/n1391 ) );
  MUX \b/U1378  ( .IN0(\b/n1389 ), .IN1(\b/n1385 ), .SEL(msg[5]), .F(\b/n1390 ) );
  MUX \b/U1377  ( .IN0(\b/n1388 ), .IN1(\b/n1387 ), .SEL(msg[2]), .F(\b/n1389 ) );
  MUX \b/U1376  ( .IN0(\b/n1156 ), .IN1(\b/n1127 ), .SEL(msg[7]), .F(\b/n1388 ) );
  MUX \b/U1375  ( .IN0(\b/n1181 ), .IN1(\b/n1386 ), .SEL(msg[7]), .F(\b/n1387 ) );
  MUX \b/U1374  ( .IN0(\b/n1123 ), .IN1(\b/n1104 ), .SEL(msg[1]), .F(\b/n1386 ) );
  MUX \b/U1373  ( .IN0(\b/n1384 ), .IN1(\b/n1383 ), .SEL(msg[2]), .F(\b/n1385 ) );
  MUX \b/U1372  ( .IN0(\b/n1121 ), .IN1(n605), .SEL(msg[7]), .F(\b/n1384 ) );
  MUX \b/U1371  ( .IN0(\b/n1382 ), .IN1(\b/n1381 ), .SEL(msg[7]), .F(\b/n1383 ) );
  AND \b/U1370  ( .A(\b/n1141 ), .B(\b/n1216 ), .Z(\b/n1382 ) );
  MUX \b/U1369  ( .IN0(\b/n1093 ), .IN1(\b/n1077 ), .SEL(msg[1]), .F(\b/n1381 ) );
  MUX \b/U1368  ( .IN0(\b/n1379 ), .IN1(\b/n1370 ), .SEL(msg[0]), .F(\b/n1380 ) );
  MUX \b/U1367  ( .IN0(\b/n1378 ), .IN1(\b/n1374 ), .SEL(msg[5]), .F(\b/n1379 ) );
  MUX \b/U1366  ( .IN0(\b/n1377 ), .IN1(\b/n1375 ), .SEL(msg[2]), .F(\b/n1378 ) );
  MUX \b/U1365  ( .IN0(\b/n1147 ), .IN1(\b/n1376 ), .SEL(msg[7]), .F(\b/n1377 ) );
  NAND \b/U1364  ( .A(msg[1]), .B(\b/n1093 ), .Z(\b/n1376 ) );
  MUX \b/U1363  ( .IN0(\b/n1077 ), .IN1(\b/n1130 ), .SEL(msg[7]), .F(\b/n1375 ) );
  MUX \b/U1362  ( .IN0(\b/n1373 ), .IN1(\b/n1372 ), .SEL(msg[2]), .F(\b/n1374 ) );
  MUX \b/U1361  ( .IN0(\b/n1173 ), .IN1(\b/n1095 ), .SEL(msg[7]), .F(\b/n1373 ) );
  MUX \b/U1360  ( .IN0(\b/n1371 ), .IN1(\b/n1136 ), .SEL(n604), .F(\b/n1372 )
         );
  AND \b/U1359  ( .A(msg[7]), .B(msg[3]), .Z(\b/n1371 ) );
  MUX \b/U1358  ( .IN0(\b/n1369 ), .IN1(\b/n1366 ), .SEL(msg[5]), .F(\b/n1370 ) );
  MUX \b/U1357  ( .IN0(\b/n1368 ), .IN1(\b/n1367 ), .SEL(msg[2]), .F(\b/n1369 ) );
  MUX \b/U1356  ( .IN0(\b/n1297 ), .IN1(\b/n1136 ), .SEL(msg[7]), .F(\b/n1368 ) );
  MUX \b/U1355  ( .IN0(n603), .IN1(\b/n1128 ), .SEL(msg[7]), .F(\b/n1367 ) );
  MUX \b/U1354  ( .IN0(\b/n1364 ), .IN1(\b/n1363 ), .SEL(msg[2]), .F(\b/n1366 ) );
  AND \b/U1353  ( .A(\b/n1365 ), .B(\b/n1265 ), .Z(\b/n1364 ) );
  MUX \b/U1352  ( .IN0(\b/n1079 ), .IN1(\b/n1123 ), .SEL(msg[7]), .F(\b/n1363 ) );
  MUX \b/U1351  ( .IN0(\b/n1362 ), .IN1(\b/n1345 ), .SEL(msg[6]), .F(
        shift_row_out[4]) );
  MUX \b/U1350  ( .IN0(\b/n1361 ), .IN1(\b/n1353 ), .SEL(msg[0]), .F(\b/n1362 ) );
  MUX \b/U1349  ( .IN0(\b/n1360 ), .IN1(\b/n1357 ), .SEL(msg[5]), .F(\b/n1361 ) );
  MUX \b/U1348  ( .IN0(\b/n1359 ), .IN1(\b/n1358 ), .SEL(msg[2]), .F(\b/n1360 ) );
  MUX \b/U1347  ( .IN0(\b/n1105 ), .IN1(\b/n1126 ), .SEL(msg[7]), .F(\b/n1359 ) );
  MUX \b/U1346  ( .IN0(\b/n1216 ), .IN1(\b/n1181 ), .SEL(msg[7]), .F(\b/n1358 ) );
  NAND \b/U1345  ( .A(msg[1]), .B(\b/n1135 ), .Z(\b/n1216 ) );
  MUX \b/U1344  ( .IN0(\b/n1354 ), .IN1(\b/n1355 ), .SEL(msg[2]), .F(\b/n1357 ) );
  AND \b/U1343  ( .A(\b/n1166 ), .B(\b/n1356 ), .Z(\b/n1355 ) );
  MUX \b/U1342  ( .IN0(\b/n1164 ), .IN1(\b/n1108 ), .SEL(msg[7]), .F(\b/n1354 ) );
  MUX \b/U1341  ( .IN0(\b/n1352 ), .IN1(\b/n1349 ), .SEL(msg[5]), .F(\b/n1353 ) );
  MUX \b/U1340  ( .IN0(\b/n1351 ), .IN1(\b/n1350 ), .SEL(msg[2]), .F(\b/n1352 ) );
  MUX \b/U1339  ( .IN0(\b/n1070 ), .IN1(\b/n1116 ), .SEL(msg[7]), .F(\b/n1351 ) );
  MUX \b/U1338  ( .IN0(\b/n1077 ), .IN1(\b/n1144 ), .SEL(msg[7]), .F(\b/n1350 ) );
  MUX \b/U1337  ( .IN0(\b/n1348 ), .IN1(\b/n1346 ), .SEL(msg[2]), .F(\b/n1349 ) );
  MUX \b/U1336  ( .IN0(\b/n1160 ), .IN1(\b/n1347 ), .SEL(msg[7]), .F(\b/n1348 ) );
  AND \b/U1335  ( .A(\b/n1144 ), .B(\b/n1134 ), .Z(\b/n1347 ) );
  MUX \b/U1334  ( .IN0(\b/n1092 ), .IN1(\b/n1111 ), .SEL(msg[7]), .F(\b/n1346 ) );
  MUX \b/U1333  ( .IN0(\b/n1344 ), .IN1(\b/n1338 ), .SEL(msg[0]), .F(\b/n1345 ) );
  MUX \b/U1332  ( .IN0(\b/n1343 ), .IN1(\b/n1341 ), .SEL(msg[5]), .F(\b/n1344 ) );
  MUX \b/U1331  ( .IN0(\b/n1342 ), .IN1(\b/n1138 ), .SEL(msg[2]), .F(\b/n1343 ) );
  MUX \b/U1330  ( .IN0(\b/n1158 ), .IN1(\b/n1113 ), .SEL(msg[7]), .F(\b/n1342 ) );
  MUX \b/U1329  ( .IN0(\b/n1340 ), .IN1(\b/n1339 ), .SEL(msg[2]), .F(\b/n1341 ) );
  MUX \b/U1328  ( .IN0(n602), .IN1(\b/n1105 ), .SEL(msg[7]), .F(\b/n1340 ) );
  MUX \b/U1327  ( .IN0(\b/n1168 ), .IN1(\b/n1171 ), .SEL(msg[7]), .F(\b/n1339 ) );
  MUX \b/U1326  ( .IN0(\b/n1337 ), .IN1(\b/n1334 ), .SEL(msg[5]), .F(\b/n1338 ) );
  MUX \b/U1325  ( .IN0(\b/n1336 ), .IN1(\b/n1335 ), .SEL(msg[2]), .F(\b/n1337 ) );
  MUX \b/U1324  ( .IN0(\b/n1078 ), .IN1(\b/n1140 ), .SEL(msg[7]), .F(\b/n1336 ) );
  MUX \b/U1323  ( .IN0(\b/n1123 ), .IN1(\b/n1162 ), .SEL(msg[7]), .F(\b/n1335 ) );
  MUX \b/U1322  ( .IN0(\b/n1066 ), .IN1(\b/n1333 ), .SEL(msg[2]), .F(\b/n1334 ) );
  MUX \b/U1321  ( .IN0(\b/n1086 ), .IN1(\b/n1144 ), .SEL(msg[7]), .F(\b/n1333 ) );
  MUX \b/U1320  ( .IN0(\b/n1332 ), .IN1(\b/n1313 ), .SEL(msg[6]), .F(
        shift_row_out[3]) );
  MUX \b/U1319  ( .IN0(\b/n1331 ), .IN1(\b/n1323 ), .SEL(msg[0]), .F(\b/n1332 ) );
  MUX \b/U1318  ( .IN0(\b/n1330 ), .IN1(\b/n1327 ), .SEL(msg[5]), .F(\b/n1331 ) );
  MUX \b/U1317  ( .IN0(\b/n1329 ), .IN1(\b/n1328 ), .SEL(msg[7]), .F(\b/n1330 ) );
  MUX \b/U1316  ( .IN0(\b/n1152 ), .IN1(\b/n1111 ), .SEL(msg[2]), .F(\b/n1329 ) );
  MUX \b/U1315  ( .IN0(n605), .IN1(\b/n1069 ), .SEL(msg[2]), .F(\b/n1328 ) );
  MUX \b/U1314  ( .IN0(\b/n1325 ), .IN1(\b/n1324 ), .SEL(msg[7]), .F(\b/n1327 ) );
  AND \b/U1313  ( .A(\b/n1326 ), .B(msg[4]), .Z(\b/n1325 ) );
  MUX \b/U1312  ( .IN0(\b/n1099 ), .IN1(\b/n1165 ), .SEL(msg[2]), .F(\b/n1324 ) );
  MUX \b/U1311  ( .IN0(\b/n1322 ), .IN1(\b/n1319 ), .SEL(msg[5]), .F(\b/n1323 ) );
  MUX \b/U1310  ( .IN0(\b/n1321 ), .IN1(\b/n1320 ), .SEL(msg[7]), .F(\b/n1322 ) );
  MUX \b/U1309  ( .IN0(\b/n1156 ), .IN1(n601), .SEL(msg[2]), .F(\b/n1321 ) );
  MUX \b/U1308  ( .IN0(\b/n1067 ), .IN1(\b/n1086 ), .SEL(msg[2]), .F(\b/n1320 ) );
  MUX \b/U1307  ( .IN0(\b/n1315 ), .IN1(\b/n1316 ), .SEL(msg[7]), .F(\b/n1319 ) );
  NAND \b/U1306  ( .A(\b/n1317 ), .B(\b/n1318 ), .Z(\b/n1316 ) );
  MUX \b/U1305  ( .IN0(\b/n1112 ), .IN1(\b/n1314 ), .SEL(msg[2]), .F(\b/n1315 ) );
  MUX \b/U1304  ( .IN0(\b/n1087 ), .IN1(\b/n1129 ), .SEL(msg[1]), .F(\b/n1314 ) );
  MUX \b/U1303  ( .IN0(\b/n1312 ), .IN1(\b/n1303 ), .SEL(msg[0]), .F(\b/n1313 ) );
  MUX \b/U1302  ( .IN0(\b/n1311 ), .IN1(\b/n1307 ), .SEL(msg[5]), .F(\b/n1312 ) );
  MUX \b/U1301  ( .IN0(\b/n1309 ), .IN1(\b/n1308 ), .SEL(msg[7]), .F(\b/n1311 ) );
  NAND \b/U1300  ( .A(\b/n1077 ), .B(\b/n1310 ), .Z(\b/n1309 ) );
  MUX \b/U1299  ( .IN0(\b/n1128 ), .IN1(\b/n1090 ), .SEL(msg[2]), .F(\b/n1308 ) );
  MUX \b/U1298  ( .IN0(\b/n1306 ), .IN1(\b/n1304 ), .SEL(msg[7]), .F(\b/n1307 ) );
  MUX \b/U1297  ( .IN0(\b/n1147 ), .IN1(\b/n1305 ), .SEL(msg[2]), .F(\b/n1306 ) );
  AND \b/U1296  ( .A(msg[1]), .B(\b/n1077 ), .Z(\b/n1305 ) );
  MUX \b/U1295  ( .IN0(\b/n1082 ), .IN1(\b/n1166 ), .SEL(msg[2]), .F(\b/n1304 ) );
  MUX \b/U1294  ( .IN0(\b/n1302 ), .IN1(\b/n1296 ), .SEL(msg[5]), .F(\b/n1303 ) );
  MUX \b/U1293  ( .IN0(\b/n1301 ), .IN1(\b/n1299 ), .SEL(msg[7]), .F(\b/n1302 ) );
  MUX \b/U1292  ( .IN0(\b/n1300 ), .IN1(\b/n1136 ), .SEL(\b/n1184 ), .F(
        \b/n1301 ) );
  MUX \b/U1291  ( .IN0(msg[3]), .IN1(msg[4]), .SEL(msg[2]), .F(\b/n1300 ) );
  MUX \b/U1290  ( .IN0(\b/n1166 ), .IN1(\b/n1297 ), .SEL(msg[2]), .F(\b/n1299 ) );
  NAND \b/U1289  ( .A(\b/n1136 ), .B(\b/n1298 ), .Z(\b/n1297 ) );
  MUX \b/U1288  ( .IN0(\b/n1293 ), .IN1(\b/n1294 ), .SEL(msg[7]), .F(\b/n1296 ) );
  AND \b/U1287  ( .A(\b/n1110 ), .B(\b/n1295 ), .Z(\b/n1294 ) );
  MUX \b/U1286  ( .IN0(\b/n1091 ), .IN1(\b/n1137 ), .SEL(msg[2]), .F(\b/n1293 ) );
  MUX \b/U1285  ( .IN0(\b/n1292 ), .IN1(\b/n1276 ), .SEL(msg[6]), .F(
        shift_row_out[2]) );
  MUX \b/U1284  ( .IN0(\b/n1291 ), .IN1(\b/n1283 ), .SEL(msg[0]), .F(\b/n1292 ) );
  MUX \b/U1283  ( .IN0(\b/n1290 ), .IN1(\b/n1286 ), .SEL(msg[5]), .F(\b/n1291 ) );
  MUX \b/U1282  ( .IN0(\b/n1289 ), .IN1(\b/n1287 ), .SEL(msg[2]), .F(\b/n1290 ) );
  MUX \b/U1281  ( .IN0(\b/n1099 ), .IN1(\b/n1288 ), .SEL(msg[7]), .F(\b/n1289 ) );
  MUX \b/U1280  ( .IN0(\b/n1144 ), .IN1(\b/n1077 ), .SEL(msg[1]), .F(\b/n1288 ) );
  MUX \b/U1279  ( .IN0(\b/n1183 ), .IN1(\b/n1117 ), .SEL(msg[7]), .F(\b/n1287 ) );
  MUX \b/U1278  ( .IN0(\b/n1285 ), .IN1(\b/n1284 ), .SEL(msg[2]), .F(\b/n1286 ) );
  MUX \b/U1277  ( .IN0(\b/n1137 ), .IN1(\b/n1084 ), .SEL(msg[7]), .F(\b/n1285 ) );
  MUX \b/U1276  ( .IN0(\b/n1120 ), .IN1(\b/n1170 ), .SEL(msg[7]), .F(\b/n1284 ) );
  MUX \b/U1275  ( .IN0(\b/n1282 ), .IN1(\b/n1278 ), .SEL(msg[5]), .F(\b/n1283 ) );
  MUX \b/U1274  ( .IN0(\b/n1279 ), .IN1(\b/n1066 ), .SEL(msg[2]), .F(\b/n1282 ) );
  NAND \b/U1273  ( .A(\b/n1280 ), .B(\b/n1281 ), .Z(\b/n1279 ) );
  MUX \b/U1272  ( .IN0(n603), .IN1(\b/n1277 ), .SEL(\b/n1182 ), .F(\b/n1278 )
         );
  MUX \b/U1271  ( .IN0(\b/n1098 ), .IN1(\b/n1149 ), .SEL(msg[2]), .F(\b/n1277 ) );
  MUX \b/U1270  ( .IN0(\b/n1275 ), .IN1(\b/n1267 ), .SEL(msg[0]), .F(\b/n1276 ) );
  MUX \b/U1269  ( .IN0(\b/n1274 ), .IN1(\b/n1271 ), .SEL(msg[5]), .F(\b/n1275 ) );
  MUX \b/U1268  ( .IN0(\b/n1273 ), .IN1(\b/n1272 ), .SEL(msg[2]), .F(\b/n1274 ) );
  MUX \b/U1267  ( .IN0(\b/n1126 ), .IN1(msg[1]), .SEL(msg[7]), .F(\b/n1273 )
         );
  MUX \b/U1266  ( .IN0(n606), .IN1(\b/n1150 ), .SEL(msg[7]), .F(\b/n1272 ) );
  MUX \b/U1265  ( .IN0(\b/n1270 ), .IN1(\b/n1269 ), .SEL(msg[2]), .F(\b/n1271 ) );
  MUX \b/U1264  ( .IN0(\b/n1131 ), .IN1(\b/n1125 ), .SEL(msg[7]), .F(\b/n1270 ) );
  MUX \b/U1263  ( .IN0(n606), .IN1(\b/n1268 ), .SEL(msg[7]), .F(\b/n1269 ) );
  MUX \b/U1262  ( .IN0(\b/n1077 ), .IN1(\b/n1114 ), .SEL(msg[1]), .F(\b/n1268 ) );
  MUX \b/U1261  ( .IN0(\b/n1266 ), .IN1(\b/n1260 ), .SEL(msg[5]), .F(\b/n1267 ) );
  MUX \b/U1260  ( .IN0(\b/n1263 ), .IN1(\b/n1262 ), .SEL(msg[2]), .F(\b/n1266 ) );
  NAND \b/U1259  ( .A(\b/n1264 ), .B(\b/n1265 ), .Z(\b/n1263 ) );
  MUX \b/U1258  ( .IN0(\b/n1136 ), .IN1(\b/n1261 ), .SEL(n604), .F(\b/n1262 )
         );
  MUX \b/U1257  ( .IN0(msg[3]), .IN1(\b/n1087 ), .SEL(msg[7]), .F(\b/n1261 )
         );
  MUX \b/U1256  ( .IN0(\b/n1259 ), .IN1(\b/n1258 ), .SEL(msg[2]), .F(\b/n1260 ) );
  MUX \b/U1255  ( .IN0(\b/n1181 ), .IN1(\b/n1085 ), .SEL(msg[7]), .F(\b/n1259 ) );
  MUX \b/U1254  ( .IN0(\b/n1177 ), .IN1(\b/n1257 ), .SEL(msg[7]), .F(\b/n1258 ) );
  MUX \b/U1253  ( .IN0(\b/n1139 ), .IN1(\b/n1144 ), .SEL(msg[1]), .F(\b/n1257 ) );
  MUX \b/U1252  ( .IN0(\b/n1256 ), .IN1(\b/n1238 ), .SEL(msg[6]), .F(
        shift_row_out[1]) );
  MUX \b/U1251  ( .IN0(\b/n1255 ), .IN1(\b/n1246 ), .SEL(msg[0]), .F(\b/n1256 ) );
  MUX \b/U1250  ( .IN0(\b/n1254 ), .IN1(\b/n1250 ), .SEL(msg[5]), .F(\b/n1255 ) );
  MUX \b/U1249  ( .IN0(\b/n1253 ), .IN1(\b/n1252 ), .SEL(msg[2]), .F(\b/n1254 ) );
  MUX \b/U1248  ( .IN0(\b/n1122 ), .IN1(n608), .SEL(msg[7]), .F(\b/n1253 ) );
  MUX \b/U1247  ( .IN0(\b/n1251 ), .IN1(n602), .SEL(msg[7]), .F(\b/n1252 ) );
  NAND \b/U1246  ( .A(\b/n1134 ), .B(\b/n1093 ), .Z(\b/n1251 ) );
  MUX \b/U1245  ( .IN0(\b/n1249 ), .IN1(\b/n1248 ), .SEL(msg[2]), .F(\b/n1250 ) );
  MUX \b/U1244  ( .IN0(\b/n1070 ), .IN1(\b/n1151 ), .SEL(msg[7]), .F(\b/n1249 ) );
  MUX \b/U1243  ( .IN0(\b/n1141 ), .IN1(\b/n1247 ), .SEL(msg[7]), .F(\b/n1248 ) );
  AND \b/U1242  ( .A(msg[1]), .B(msg[4]), .Z(\b/n1247 ) );
  MUX \b/U1241  ( .IN0(\b/n1245 ), .IN1(\b/n1242 ), .SEL(msg[5]), .F(\b/n1246 ) );
  MUX \b/U1240  ( .IN0(\b/n1244 ), .IN1(\b/n1243 ), .SEL(msg[2]), .F(\b/n1245 ) );
  MUX \b/U1239  ( .IN0(\b/n1180 ), .IN1(\b/n1131 ), .SEL(msg[7]), .F(\b/n1244 ) );
  MUX \b/U1238  ( .IN0(\b/n1106 ), .IN1(\b/n1149 ), .SEL(msg[7]), .F(\b/n1243 ) );
  MUX \b/U1237  ( .IN0(\b/n1239 ), .IN1(\b/n1240 ), .SEL(msg[2]), .F(\b/n1242 ) );
  AND \b/U1236  ( .A(\b/n1241 ), .B(\b/n1196 ), .Z(\b/n1240 ) );
  MUX \b/U1235  ( .IN0(\b/n1155 ), .IN1(\b/n1144 ), .SEL(msg[7]), .F(\b/n1239 ) );
  MUX \b/U1234  ( .IN0(\b/n1237 ), .IN1(\b/n1229 ), .SEL(msg[0]), .F(\b/n1238 ) );
  MUX \b/U1233  ( .IN0(\b/n1236 ), .IN1(\b/n1232 ), .SEL(msg[5]), .F(\b/n1237 ) );
  MUX \b/U1232  ( .IN0(\b/n1235 ), .IN1(\b/n1234 ), .SEL(msg[2]), .F(\b/n1236 ) );
  MUX \b/U1231  ( .IN0(\b/n1143 ), .IN1(\b/n1095 ), .SEL(msg[7]), .F(\b/n1235 ) );
  MUX \b/U1230  ( .IN0(\b/n1233 ), .IN1(\b/n1079 ), .SEL(msg[7]), .F(\b/n1234 ) );
  MUX \b/U1229  ( .IN0(\b/n1141 ), .IN1(\b/n1087 ), .SEL(msg[1]), .F(\b/n1233 ) );
  MUX \b/U1228  ( .IN0(\b/n1231 ), .IN1(\b/n1230 ), .SEL(msg[2]), .F(\b/n1232 ) );
  MUX \b/U1227  ( .IN0(\b/n1126 ), .IN1(\b/n1104 ), .SEL(msg[7]), .F(\b/n1231 ) );
  MUX \b/U1226  ( .IN0(\b/n1122 ), .IN1(\b/n1082 ), .SEL(msg[7]), .F(\b/n1230 ) );
  MUX \b/U1225  ( .IN0(\b/n1228 ), .IN1(\b/n1223 ), .SEL(msg[5]), .F(\b/n1229 ) );
  MUX \b/U1224  ( .IN0(\b/n1227 ), .IN1(\b/n1224 ), .SEL(msg[2]), .F(\b/n1228 ) );
  MUX \b/U1223  ( .IN0(\b/n1225 ), .IN1(\b/n1226 ), .SEL(msg[7]), .F(\b/n1227 ) );
  NAND \b/U1222  ( .A(\b/n1144 ), .B(\b/n1216 ), .Z(\b/n1226 ) );
  MUX \b/U1221  ( .IN0(\b/n1144 ), .IN1(\b/n1087 ), .SEL(msg[1]), .F(\b/n1225 ) );
  MUX \b/U1220  ( .IN0(\b/n1161 ), .IN1(\b/n1159 ), .SEL(msg[7]), .F(\b/n1224 ) );
  MUX \b/U1219  ( .IN0(\b/n1179 ), .IN1(\b/n1222 ), .SEL(msg[2]), .F(\b/n1223 ) );
  MUX \b/U1218  ( .IN0(\b/n1093 ), .IN1(\b/n1125 ), .SEL(msg[7]), .F(\b/n1222 ) );
  MUX \b/U1217  ( .IN0(\b/n1221 ), .IN1(\b/n1204 ), .SEL(msg[6]), .F(
        shift_row_out[0]) );
  MUX \b/U1216  ( .IN0(\b/n1220 ), .IN1(\b/n1212 ), .SEL(msg[0]), .F(\b/n1221 ) );
  MUX \b/U1215  ( .IN0(\b/n1219 ), .IN1(\b/n1217 ), .SEL(msg[2]), .F(\b/n1220 ) );
  MUX \b/U1214  ( .IN0(\b/n1067 ), .IN1(\b/n1218 ), .SEL(msg[7]), .F(\b/n1219 ) );
  MUX \b/U1213  ( .IN0(\b/n1120 ), .IN1(\b/n1123 ), .SEL(msg[5]), .F(\b/n1218 ) );
  MUX \b/U1212  ( .IN0(\b/n1214 ), .IN1(\b/n1213 ), .SEL(msg[7]), .F(\b/n1217 ) );
  NAND \b/U1211  ( .A(\b/n1215 ), .B(\b/n1216 ), .Z(\b/n1214 ) );
  MUX \b/U1210  ( .IN0(\b/n1119 ), .IN1(\b/n1134 ), .SEL(msg[5]), .F(\b/n1213 ) );
  MUX \b/U1209  ( .IN0(\b/n1211 ), .IN1(\b/n1207 ), .SEL(msg[2]), .F(\b/n1212 ) );
  MUX \b/U1208  ( .IN0(\b/n1210 ), .IN1(\b/n1208 ), .SEL(msg[7]), .F(\b/n1211 ) );
  MUX \b/U1207  ( .IN0(\b/n1209 ), .IN1(\b/n1072 ), .SEL(msg[5]), .F(\b/n1210 ) );
  NAND \b/U1206  ( .A(\b/n1134 ), .B(\b/n1136 ), .Z(\b/n1209 ) );
  MUX \b/U1204  ( .IN0(\b/n1206 ), .IN1(\b/n1205 ), .SEL(msg[7]), .F(\b/n1207 ) );
  MUX \b/U1203  ( .IN0(n603), .IN1(\b/n1069 ), .SEL(msg[5]), .F(\b/n1206 ) );
  MUX \b/U1202  ( .IN0(\b/n1121 ), .IN1(\b/n1077 ), .SEL(msg[5]), .F(\b/n1205 ) );
  MUX \b/U1201  ( .IN0(\b/n1203 ), .IN1(\b/n1193 ), .SEL(msg[0]), .F(\b/n1204 ) );
  MUX \b/U1200  ( .IN0(\b/n1202 ), .IN1(\b/n1198 ), .SEL(msg[2]), .F(\b/n1203 ) );
  MUX \b/U1199  ( .IN0(\b/n1201 ), .IN1(\b/n1200 ), .SEL(msg[7]), .F(\b/n1202 ) );
  MUX \b/U1198  ( .IN0(n601), .IN1(\b/n1073 ), .SEL(msg[5]), .F(\b/n1201 ) );
  MUX \b/U1197  ( .IN0(\b/n1199 ), .IN1(\b/n1110 ), .SEL(msg[5]), .F(\b/n1200 ) );
  NAND \b/U1196  ( .A(\b/n1135 ), .B(\b/n1137 ), .Z(\b/n1199 ) );
  MUX \b/U1195  ( .IN0(\b/n1197 ), .IN1(\b/n1194 ), .SEL(msg[7]), .F(\b/n1198 ) );
  MUX \b/U1194  ( .IN0(\b/n1080 ), .IN1(\b/n1195 ), .SEL(msg[5]), .F(\b/n1197 ) );
  NAND \b/U1193  ( .A(\b/n1139 ), .B(\b/n1196 ), .Z(\b/n1195 ) );
  MUX \b/U1192  ( .IN0(\b/n1154 ), .IN1(\b/n1145 ), .SEL(msg[5]), .F(\b/n1194 ) );
  MUX \b/U1191  ( .IN0(\b/n1192 ), .IN1(\b/n1188 ), .SEL(msg[2]), .F(\b/n1193 ) );
  MUX \b/U1190  ( .IN0(\b/n1190 ), .IN1(\b/n1189 ), .SEL(msg[7]), .F(\b/n1192 ) );
  NAND \b/U1189  ( .A(\b/n1191 ), .B(\b/n1178 ), .Z(\b/n1190 ) );
  MUX \b/U1188  ( .IN0(msg[3]), .IN1(\b/n1170 ), .SEL(msg[5]), .F(\b/n1189 )
         );
  MUX \b/U1187  ( .IN0(\b/n1187 ), .IN1(\b/n1186 ), .SEL(msg[7]), .F(\b/n1188 ) );
  MUX \b/U1186  ( .IN0(\b/n1085 ), .IN1(\b/n1101 ), .SEL(msg[5]), .F(\b/n1187 ) );
  MUX \b/U1185  ( .IN0(\b/n1118 ), .IN1(\b/n1106 ), .SEL(msg[5]), .F(\b/n1186 ) );
  XOR \b/U1184  ( .A(\b/n1136 ), .B(msg[1]), .Z(\b/n1185 ) );
  XOR \b/U1183  ( .A(msg[1]), .B(msg[2]), .Z(\b/n1184 ) );
  XOR \b/U1182  ( .A(msg[1]), .B(msg[3]), .Z(\b/n1183 ) );
  XOR \b/U1181  ( .A(msg[2]), .B(msg[7]), .Z(\b/n1182 ) );
  XOR \b/U1180  ( .A(\b/n1134 ), .B(\b/n1077 ), .Z(\b/n1181 ) );
  XOR \b/U1179  ( .A(msg[1]), .B(\b/n1123 ), .Z(\b/n1180 ) );
  XOR \b/U1177  ( .A(msg[1]), .B(msg[5]), .Z(\b/n1178 ) );
  NAND \b/U1176  ( .A(msg[1]), .B(msg[3]), .Z(\b/n1177 ) );
  MUX \b/U1175  ( .IN0(\b/n1136 ), .IN1(\b/n1077 ), .SEL(msg[1]), .F(\b/n1176 ) );
  MUX \b/U1173  ( .IN0(msg[3]), .IN1(\b/n1114 ), .SEL(msg[1]), .F(\b/n1174 )
         );
  MUX \b/U1172  ( .IN0(\b/n1093 ), .IN1(\b/n1114 ), .SEL(msg[1]), .F(\b/n1173 ) );
  MUX \b/U1171  ( .IN0(\b/n1139 ), .IN1(\b/n1141 ), .SEL(msg[1]), .F(\b/n1172 ) );
  MUX \b/U1170  ( .IN0(msg[4]), .IN1(\b/n1093 ), .SEL(msg[1]), .F(\b/n1171 )
         );
  OR \b/U1169  ( .A(msg[1]), .B(msg[4]), .Z(\b/n1170 ) );
  NAND \b/U1167  ( .A(\b/n1114 ), .B(\b/n1134 ), .Z(\b/n1168 ) );
  MUX \b/U1166  ( .IN0(\b/n1114 ), .IN1(msg[4]), .SEL(msg[1]), .F(\b/n1167 )
         );
  MUX \b/U1165  ( .IN0(\b/n1135 ), .IN1(\b/n1144 ), .SEL(msg[1]), .F(\b/n1166 ) );
  MUX \b/U1164  ( .IN0(\b/n1129 ), .IN1(msg[4]), .SEL(msg[1]), .F(\b/n1165 )
         );
  MUX \b/U1163  ( .IN0(\b/n1087 ), .IN1(\b/n1114 ), .SEL(msg[1]), .F(\b/n1164 ) );
  MUX \b/U1162  ( .IN0(\b/n1135 ), .IN1(msg[4]), .SEL(msg[1]), .F(\b/n1163 )
         );
  MUX \b/U1161  ( .IN0(\b/n1104 ), .IN1(\b/n1093 ), .SEL(msg[1]), .F(\b/n1162 ) );
  XOR \b/U1160  ( .A(\b/n1087 ), .B(msg[1]), .Z(\b/n1161 ) );
  MUX \b/U1159  ( .IN0(\b/n1141 ), .IN1(\b/n1104 ), .SEL(msg[1]), .F(\b/n1160 ) );
  NANDN \b/U1158  ( .B(msg[1]), .A(msg[3]), .Z(\b/n1159 ) );
  MUX \b/U1157  ( .IN0(\b/n1077 ), .IN1(msg[3]), .SEL(msg[1]), .F(\b/n1158 )
         );
  NAND \b/U1155  ( .A(\b/n1139 ), .B(\b/n1134 ), .Z(\b/n1156 ) );
  MUX \b/U1154  ( .IN0(msg[4]), .IN1(\b/n1136 ), .SEL(msg[1]), .F(\b/n1155 )
         );
  MUX \b/U1153  ( .IN0(\b/n1104 ), .IN1(msg[3]), .SEL(msg[1]), .F(\b/n1154 )
         );
  MUX \b/U1151  ( .IN0(msg[4]), .IN1(\b/n1123 ), .SEL(msg[1]), .F(\b/n1152 )
         );
  MUX \b/U1150  ( .IN0(\b/n1077 ), .IN1(\b/n1129 ), .SEL(msg[1]), .F(\b/n1151 ) );
  NAND \b/U1149  ( .A(\b/n1137 ), .B(\b/n1077 ), .Z(\b/n1150 ) );
  MUX \b/U1148  ( .IN0(\b/n1136 ), .IN1(\b/n1144 ), .SEL(msg[1]), .F(\b/n1149 ) );
  NAND \b/U1147  ( .A(\b/n1148 ), .B(\b/n1135 ), .Z(\b/n1147 ) );
  MUX \b/U1146  ( .IN0(\b/n1139 ), .IN1(\b/n1129 ), .SEL(msg[1]), .F(\b/n1146 ) );
  MUX \b/U1145  ( .IN0(\b/n1129 ), .IN1(\b/n1093 ), .SEL(msg[1]), .F(\b/n1145 ) );
  NANDN \b/U1144  ( .B(msg[3]), .A(msg[4]), .Z(\b/n1144 ) );
  MUX \b/U1143  ( .IN0(\b/n1139 ), .IN1(msg[3]), .SEL(msg[1]), .F(\b/n1143 )
         );
  OR \b/U1142  ( .A(msg[3]), .B(msg[4]), .Z(\b/n1139 ) );
  MUX \b/U1141  ( .IN0(\b/n1077 ), .IN1(\b/n1093 ), .SEL(msg[1]), .F(\b/n1142 ) );
  XOR \b/U1140  ( .A(\b/n1087 ), .B(msg[3]), .Z(\b/n1141 ) );
  NANDN \b/U1139  ( .B(msg[3]), .A(msg[1]), .Z(\b/n1140 ) );
  NAND \b/U1138  ( .A(\b/n1139 ), .B(\b/n1137 ), .Z(\b/n1138 ) );
  NAND \b/U1137  ( .A(msg[1]), .B(\b/n1136 ), .Z(\b/n1137 ) );
  NANDN \b/U1136  ( .B(msg[4]), .A(msg[3]), .Z(\b/n1136 ) );
  NAND \b/U1135  ( .A(msg[3]), .B(msg[4]), .Z(\b/n1135 ) );
  XOR \d/U548  ( .A(shift_row_out[25]), .B(shift_row_out[17]), .Z(\d/n337 ) );
  XOR \d/U547  ( .A(\d/n337 ), .B(\d/n117 ), .Z(\d/n421 ) );
  XOR \d/U546  ( .A(shift_row_out[9]), .B(\d/n420 ), .Z(\d/n117 ) );
  XOR \d/U545  ( .A(\d/n119 ), .B(\d/n118 ), .Z(\d/n422 ) );
  XOR \d/U544  ( .A(shift_row_out[11]), .B(\d/n419 ), .Z(\d/n118 ) );
  XOR \d/U543  ( .A(shift_row_out[27]), .B(shift_row_out[19]), .Z(\d/n119 ) );
  XOR \d/U542  ( .A(shift_row_out[28]), .B(shift_row_out[20]), .Z(\d/n338 ) );
  XOR \d/U541  ( .A(\d/n338 ), .B(\d/n120 ), .Z(\d/n423 ) );
  XOR \d/U540  ( .A(shift_row_out[12]), .B(\d/n418 ), .Z(\d/n120 ) );
  XOR \d/U539  ( .A(\d/n337 ), .B(\d/n121 ), .Z(\d/n424 ) );
  XOR \d/U538  ( .A(shift_row_out[1]), .B(\d/n417 ), .Z(\d/n121 ) );
  XOR \d/U537  ( .A(\d/n123 ), .B(\d/n122 ), .Z(\d/n425 ) );
  XOR \d/U536  ( .A(shift_row_out[3]), .B(\d/n416 ), .Z(\d/n122 ) );
  XOR \d/U535  ( .A(shift_row_out[27]), .B(shift_row_out[19]), .Z(\d/n123 ) );
  XOR \d/U534  ( .A(\d/n338 ), .B(\d/n124 ), .Z(\d/n426 ) );
  XOR \d/U533  ( .A(shift_row_out[4]), .B(\d/n415 ), .Z(\d/n124 ) );
  XOR \d/U532  ( .A(\d/n126 ), .B(\d/n125 ), .Z(\d/n427 ) );
  XOR \d/U531  ( .A(shift_row_out[1]), .B(\d/n414 ), .Z(\d/n125 ) );
  XOR \d/U530  ( .A(shift_row_out[25]), .B(shift_row_out[9]), .Z(\d/n126 ) );
  XOR \d/U529  ( .A(\d/n128 ), .B(\d/n127 ), .Z(\d/n428 ) );
  XOR \d/U528  ( .A(shift_row_out[3]), .B(\d/n413 ), .Z(\d/n127 ) );
  XOR \d/U527  ( .A(shift_row_out[27]), .B(shift_row_out[11]), .Z(\d/n128 ) );
  XOR \d/U526  ( .A(shift_row_out[12]), .B(shift_row_out[4]), .Z(\d/n333 ) );
  XOR \d/U525  ( .A(\d/n333 ), .B(\d/n129 ), .Z(\d/n429 ) );
  XOR \d/U524  ( .A(shift_row_out[28]), .B(\d/n412 ), .Z(\d/n129 ) );
  XOR \d/U523  ( .A(\d/n131 ), .B(\d/n130 ), .Z(\d/n430 ) );
  XOR \d/U522  ( .A(shift_row_out[1]), .B(\d/n411 ), .Z(\d/n130 ) );
  XOR \d/U521  ( .A(shift_row_out[17]), .B(shift_row_out[9]), .Z(\d/n131 ) );
  XOR \d/U520  ( .A(\d/n133 ), .B(\d/n132 ), .Z(\d/n431 ) );
  XOR \d/U519  ( .A(shift_row_out[3]), .B(\d/n410 ), .Z(\d/n132 ) );
  XOR \d/U518  ( .A(shift_row_out[19]), .B(shift_row_out[11]), .Z(\d/n133 ) );
  XOR \d/U517  ( .A(\d/n333 ), .B(\d/n134 ), .Z(\d/n432 ) );
  XOR \d/U516  ( .A(shift_row_out[20]), .B(\d/n409 ), .Z(\d/n134 ) );
  XOR \d/U515  ( .A(shift_row_out[57]), .B(shift_row_out[49]), .Z(\d/n347 ) );
  XOR \d/U514  ( .A(\d/n347 ), .B(\d/n135 ), .Z(\d/n433 ) );
  XOR \d/U513  ( .A(shift_row_out[41]), .B(\d/n408 ), .Z(\d/n135 ) );
  XOR \d/U512  ( .A(\d/n137 ), .B(\d/n136 ), .Z(\d/n434 ) );
  XOR \d/U511  ( .A(shift_row_out[43]), .B(\d/n407 ), .Z(\d/n136 ) );
  XOR \d/U510  ( .A(shift_row_out[59]), .B(shift_row_out[51]), .Z(\d/n137 ) );
  XOR \d/U509  ( .A(shift_row_out[60]), .B(shift_row_out[52]), .Z(\d/n348 ) );
  XOR \d/U508  ( .A(\d/n348 ), .B(\d/n138 ), .Z(\d/n435 ) );
  XOR \d/U507  ( .A(shift_row_out[44]), .B(\d/n406 ), .Z(\d/n138 ) );
  XOR \d/U506  ( .A(\d/n347 ), .B(\d/n139 ), .Z(\d/n436 ) );
  XOR \d/U505  ( .A(shift_row_out[33]), .B(\d/n405 ), .Z(\d/n139 ) );
  XOR \d/U504  ( .A(\d/n141 ), .B(\d/n140 ), .Z(\d/n437 ) );
  XOR \d/U503  ( .A(shift_row_out[35]), .B(\d/n404 ), .Z(\d/n140 ) );
  XOR \d/U502  ( .A(shift_row_out[59]), .B(shift_row_out[51]), .Z(\d/n141 ) );
  XOR \d/U501  ( .A(\d/n348 ), .B(\d/n142 ), .Z(\d/n438 ) );
  XOR \d/U500  ( .A(shift_row_out[36]), .B(\d/n403 ), .Z(\d/n142 ) );
  XOR \d/U499  ( .A(\d/n144 ), .B(\d/n143 ), .Z(\d/n439 ) );
  XOR \d/U498  ( .A(shift_row_out[33]), .B(\d/n402 ), .Z(\d/n143 ) );
  XOR \d/U497  ( .A(shift_row_out[57]), .B(shift_row_out[41]), .Z(\d/n144 ) );
  XOR \d/U496  ( .A(\d/n146 ), .B(\d/n145 ), .Z(\d/n440 ) );
  XOR \d/U495  ( .A(shift_row_out[35]), .B(\d/n401 ), .Z(\d/n145 ) );
  XOR \d/U494  ( .A(shift_row_out[59]), .B(shift_row_out[43]), .Z(\d/n146 ) );
  XOR \d/U493  ( .A(shift_row_out[44]), .B(shift_row_out[36]), .Z(\d/n343 ) );
  XOR \d/U492  ( .A(\d/n343 ), .B(\d/n147 ), .Z(\d/n441 ) );
  XOR \d/U491  ( .A(shift_row_out[60]), .B(\d/n400 ), .Z(\d/n147 ) );
  XOR \d/U490  ( .A(\d/n149 ), .B(\d/n148 ), .Z(\d/n442 ) );
  XOR \d/U489  ( .A(shift_row_out[33]), .B(\d/n399 ), .Z(\d/n148 ) );
  XOR \d/U488  ( .A(shift_row_out[49]), .B(shift_row_out[41]), .Z(\d/n149 ) );
  XOR \d/U487  ( .A(\d/n151 ), .B(\d/n150 ), .Z(\d/n443 ) );
  XOR \d/U486  ( .A(shift_row_out[35]), .B(\d/n398 ), .Z(\d/n150 ) );
  XOR \d/U485  ( .A(shift_row_out[51]), .B(shift_row_out[43]), .Z(\d/n151 ) );
  XOR \d/U484  ( .A(\d/n343 ), .B(\d/n152 ), .Z(\d/n444 ) );
  XOR \d/U483  ( .A(shift_row_out[52]), .B(\d/n397 ), .Z(\d/n152 ) );
  XOR \d/U482  ( .A(shift_row_out[89]), .B(shift_row_out[81]), .Z(\d/n357 ) );
  XOR \d/U481  ( .A(\d/n357 ), .B(\d/n153 ), .Z(\d/n445 ) );
  XOR \d/U480  ( .A(shift_row_out[73]), .B(\d/n396 ), .Z(\d/n153 ) );
  XOR \d/U479  ( .A(\d/n155 ), .B(\d/n154 ), .Z(\d/n446 ) );
  XOR \d/U478  ( .A(shift_row_out[75]), .B(\d/n395 ), .Z(\d/n154 ) );
  XOR \d/U477  ( .A(shift_row_out[91]), .B(shift_row_out[83]), .Z(\d/n155 ) );
  XOR \d/U476  ( .A(shift_row_out[92]), .B(shift_row_out[84]), .Z(\d/n358 ) );
  XOR \d/U475  ( .A(\d/n358 ), .B(\d/n156 ), .Z(\d/n447 ) );
  XOR \d/U474  ( .A(shift_row_out[76]), .B(\d/n394 ), .Z(\d/n156 ) );
  XOR \d/U473  ( .A(\d/n357 ), .B(\d/n157 ), .Z(\d/n448 ) );
  XOR \d/U472  ( .A(shift_row_out[65]), .B(\d/n393 ), .Z(\d/n157 ) );
  XOR \d/U471  ( .A(\d/n159 ), .B(\d/n158 ), .Z(\d/n449 ) );
  XOR \d/U470  ( .A(shift_row_out[67]), .B(\d/n392 ), .Z(\d/n158 ) );
  XOR \d/U469  ( .A(shift_row_out[91]), .B(shift_row_out[83]), .Z(\d/n159 ) );
  XOR \d/U468  ( .A(\d/n358 ), .B(\d/n160 ), .Z(\d/n450 ) );
  XOR \d/U467  ( .A(shift_row_out[68]), .B(\d/n391 ), .Z(\d/n160 ) );
  XOR \d/U466  ( .A(\d/n162 ), .B(\d/n161 ), .Z(\d/n451 ) );
  XOR \d/U465  ( .A(shift_row_out[65]), .B(\d/n390 ), .Z(\d/n161 ) );
  XOR \d/U464  ( .A(shift_row_out[89]), .B(shift_row_out[73]), .Z(\d/n162 ) );
  XOR \d/U463  ( .A(\d/n164 ), .B(\d/n163 ), .Z(\d/n452 ) );
  XOR \d/U462  ( .A(shift_row_out[67]), .B(\d/n389 ), .Z(\d/n163 ) );
  XOR \d/U461  ( .A(shift_row_out[91]), .B(shift_row_out[75]), .Z(\d/n164 ) );
  XOR \d/U460  ( .A(shift_row_out[76]), .B(shift_row_out[68]), .Z(\d/n353 ) );
  XOR \d/U459  ( .A(\d/n353 ), .B(\d/n165 ), .Z(\d/n453 ) );
  XOR \d/U458  ( .A(shift_row_out[92]), .B(\d/n388 ), .Z(\d/n165 ) );
  XOR \d/U457  ( .A(\d/n167 ), .B(\d/n166 ), .Z(\d/n454 ) );
  XOR \d/U456  ( .A(shift_row_out[65]), .B(\d/n387 ), .Z(\d/n166 ) );
  XOR \d/U455  ( .A(shift_row_out[81]), .B(shift_row_out[73]), .Z(\d/n167 ) );
  XOR \d/U454  ( .A(\d/n169 ), .B(\d/n168 ), .Z(\d/n455 ) );
  XOR \d/U453  ( .A(shift_row_out[67]), .B(\d/n386 ), .Z(\d/n168 ) );
  XOR \d/U452  ( .A(shift_row_out[83]), .B(shift_row_out[75]), .Z(\d/n169 ) );
  XOR \d/U451  ( .A(\d/n353 ), .B(\d/n170 ), .Z(\d/n456 ) );
  XOR \d/U450  ( .A(shift_row_out[84]), .B(\d/n385 ), .Z(\d/n170 ) );
  XOR \d/U449  ( .A(shift_row_out[121]), .B(shift_row_out[113]), .Z(\d/n367 )
         );
  XOR \d/U448  ( .A(\d/n367 ), .B(\d/n171 ), .Z(\d/n457 ) );
  XOR \d/U447  ( .A(shift_row_out[105]), .B(\d/n384 ), .Z(\d/n171 ) );
  XOR \d/U446  ( .A(\d/n173 ), .B(\d/n172 ), .Z(\d/n458 ) );
  XOR \d/U445  ( .A(shift_row_out[107]), .B(\d/n383 ), .Z(\d/n172 ) );
  XOR \d/U444  ( .A(shift_row_out[123]), .B(shift_row_out[115]), .Z(\d/n173 )
         );
  XOR \d/U443  ( .A(shift_row_out[124]), .B(shift_row_out[116]), .Z(\d/n368 )
         );
  XOR \d/U442  ( .A(\d/n368 ), .B(\d/n174 ), .Z(\d/n459 ) );
  XOR \d/U441  ( .A(shift_row_out[108]), .B(\d/n382 ), .Z(\d/n174 ) );
  XOR \d/U440  ( .A(\d/n367 ), .B(\d/n175 ), .Z(\d/n460 ) );
  XOR \d/U439  ( .A(shift_row_out[97]), .B(\d/n381 ), .Z(\d/n175 ) );
  XOR \d/U438  ( .A(\d/n177 ), .B(\d/n176 ), .Z(\d/n461 ) );
  XOR \d/U437  ( .A(shift_row_out[99]), .B(\d/n380 ), .Z(\d/n176 ) );
  XOR \d/U436  ( .A(shift_row_out[123]), .B(shift_row_out[115]), .Z(\d/n177 )
         );
  XOR \d/U435  ( .A(\d/n368 ), .B(\d/n178 ), .Z(\d/n462 ) );
  XOR \d/U434  ( .A(shift_row_out[100]), .B(\d/n379 ), .Z(\d/n178 ) );
  XOR \d/U433  ( .A(\d/n180 ), .B(\d/n179 ), .Z(\d/n463 ) );
  XOR \d/U432  ( .A(shift_row_out[97]), .B(\d/n378 ), .Z(\d/n179 ) );
  XOR \d/U431  ( .A(shift_row_out[121]), .B(shift_row_out[105]), .Z(\d/n180 )
         );
  XOR \d/U430  ( .A(\d/n182 ), .B(\d/n181 ), .Z(\d/n464 ) );
  XOR \d/U429  ( .A(shift_row_out[99]), .B(\d/n377 ), .Z(\d/n181 ) );
  XOR \d/U428  ( .A(shift_row_out[123]), .B(shift_row_out[107]), .Z(\d/n182 )
         );
  XOR \d/U427  ( .A(shift_row_out[108]), .B(shift_row_out[100]), .Z(\d/n363 )
         );
  XOR \d/U426  ( .A(\d/n363 ), .B(\d/n183 ), .Z(\d/n465 ) );
  XOR \d/U425  ( .A(shift_row_out[124]), .B(\d/n376 ), .Z(\d/n183 ) );
  XOR \d/U424  ( .A(\d/n185 ), .B(\d/n184 ), .Z(\d/n466 ) );
  XOR \d/U423  ( .A(shift_row_out[97]), .B(\d/n375 ), .Z(\d/n184 ) );
  XOR \d/U422  ( .A(shift_row_out[113]), .B(shift_row_out[105]), .Z(\d/n185 )
         );
  XOR \d/U421  ( .A(\d/n187 ), .B(\d/n186 ), .Z(\d/n467 ) );
  XOR \d/U420  ( .A(shift_row_out[99]), .B(\d/n374 ), .Z(\d/n186 ) );
  XOR \d/U419  ( .A(shift_row_out[115]), .B(shift_row_out[107]), .Z(\d/n187 )
         );
  XOR \d/U418  ( .A(\d/n363 ), .B(\d/n188 ), .Z(\d/n468 ) );
  XOR \d/U417  ( .A(shift_row_out[116]), .B(\d/n373 ), .Z(\d/n188 ) );
  XOR \d/U416  ( .A(shift_row_out[15]), .B(\d/n189 ), .Z(\d/n334 ) );
  XOR \d/U415  ( .A(shift_row_out[24]), .B(shift_row_out[16]), .Z(\d/n189 ) );
  XOR \d/U414  ( .A(\d/n334 ), .B(\d/n190 ), .Z(mix_col_out[0]) );
  XOR \d/U413  ( .A(shift_row_out[8]), .B(shift_row_out[7]), .Z(\d/n190 ) );
  XOR \d/U412  ( .A(shift_row_out[9]), .B(\d/n191 ), .Z(\d/n335 ) );
  XOR \d/U411  ( .A(shift_row_out[26]), .B(shift_row_out[18]), .Z(\d/n191 ) );
  XOR \d/U410  ( .A(\d/n335 ), .B(\d/n192 ), .Z(mix_col_out[2]) );
  XOR \d/U409  ( .A(shift_row_out[10]), .B(shift_row_out[1]), .Z(\d/n192 ) );
  XOR \d/U408  ( .A(shift_row_out[29]), .B(shift_row_out[21]), .Z(\d/n339 ) );
  XOR \d/U407  ( .A(\d/n333 ), .B(\d/n193 ), .Z(mix_col_out[5]) );
  XOR \d/U406  ( .A(shift_row_out[13]), .B(\d/n339 ), .Z(\d/n193 ) );
  XOR \d/U405  ( .A(shift_row_out[30]), .B(shift_row_out[22]), .Z(\d/n340 ) );
  XOR \d/U404  ( .A(shift_row_out[13]), .B(shift_row_out[5]), .Z(\d/n341 ) );
  XOR \d/U403  ( .A(\d/n341 ), .B(\d/n194 ), .Z(mix_col_out[6]) );
  XOR \d/U402  ( .A(shift_row_out[14]), .B(\d/n340 ), .Z(\d/n194 ) );
  XOR \d/U401  ( .A(shift_row_out[31]), .B(shift_row_out[23]), .Z(\d/n336 ) );
  XOR \d/U400  ( .A(shift_row_out[14]), .B(shift_row_out[6]), .Z(\d/n342 ) );
  XOR \d/U399  ( .A(\d/n342 ), .B(\d/n195 ), .Z(mix_col_out[7]) );
  XOR \d/U398  ( .A(shift_row_out[15]), .B(\d/n336 ), .Z(\d/n195 ) );
  XOR \d/U397  ( .A(\d/n334 ), .B(\d/n196 ), .Z(mix_col_out[8]) );
  XOR \d/U396  ( .A(shift_row_out[23]), .B(shift_row_out[0]), .Z(\d/n196 ) );
  XOR \d/U395  ( .A(\d/n335 ), .B(\d/n197 ), .Z(mix_col_out[10]) );
  XOR \d/U394  ( .A(shift_row_out[17]), .B(shift_row_out[2]), .Z(\d/n197 ) );
  XOR \d/U393  ( .A(\d/n199 ), .B(\d/n198 ), .Z(mix_col_out[13]) );
  XOR \d/U392  ( .A(shift_row_out[5]), .B(\d/n339 ), .Z(\d/n198 ) );
  XOR \d/U391  ( .A(shift_row_out[20]), .B(shift_row_out[12]), .Z(\d/n199 ) );
  XOR \d/U390  ( .A(\d/n201 ), .B(\d/n200 ), .Z(mix_col_out[14]) );
  XOR \d/U389  ( .A(shift_row_out[6]), .B(\d/n340 ), .Z(\d/n200 ) );
  XOR \d/U388  ( .A(shift_row_out[21]), .B(shift_row_out[13]), .Z(\d/n201 ) );
  XOR \d/U387  ( .A(\d/n203 ), .B(\d/n202 ), .Z(mix_col_out[15]) );
  XOR \d/U386  ( .A(shift_row_out[7]), .B(\d/n336 ), .Z(\d/n202 ) );
  XOR \d/U385  ( .A(shift_row_out[22]), .B(shift_row_out[14]), .Z(\d/n203 ) );
  XOR \d/U384  ( .A(\d/n205 ), .B(\d/n204 ), .Z(mix_col_out[16]) );
  XOR \d/U383  ( .A(shift_row_out[0]), .B(\d/n336 ), .Z(\d/n204 ) );
  XOR \d/U382  ( .A(shift_row_out[24]), .B(shift_row_out[8]), .Z(\d/n205 ) );
  XOR \d/U381  ( .A(\d/n207 ), .B(\d/n206 ), .Z(mix_col_out[18]) );
  XOR \d/U380  ( .A(shift_row_out[2]), .B(\d/n337 ), .Z(\d/n206 ) );
  XOR \d/U379  ( .A(shift_row_out[26]), .B(shift_row_out[10]), .Z(\d/n207 ) );
  XOR \d/U378  ( .A(\d/n341 ), .B(\d/n208 ), .Z(mix_col_out[21]) );
  XOR \d/U377  ( .A(shift_row_out[29]), .B(\d/n338 ), .Z(\d/n208 ) );
  XOR \d/U376  ( .A(\d/n342 ), .B(\d/n209 ), .Z(mix_col_out[22]) );
  XOR \d/U375  ( .A(shift_row_out[30]), .B(\d/n339 ), .Z(\d/n209 ) );
  XOR \d/U374  ( .A(\d/n211 ), .B(\d/n210 ), .Z(mix_col_out[23]) );
  XOR \d/U373  ( .A(shift_row_out[7]), .B(\d/n340 ), .Z(\d/n210 ) );
  XOR \d/U372  ( .A(shift_row_out[31]), .B(shift_row_out[15]), .Z(\d/n211 ) );
  XOR \d/U371  ( .A(\d/n213 ), .B(\d/n212 ), .Z(mix_col_out[24]) );
  XOR \d/U370  ( .A(shift_row_out[0]), .B(\d/n214 ), .Z(\d/n212 ) );
  XOR \d/U369  ( .A(shift_row_out[8]), .B(shift_row_out[7]), .Z(\d/n213 ) );
  XOR \d/U368  ( .A(shift_row_out[31]), .B(shift_row_out[16]), .Z(\d/n214 ) );
  XOR \d/U367  ( .A(\d/n216 ), .B(\d/n215 ), .Z(mix_col_out[26]) );
  XOR \d/U366  ( .A(shift_row_out[1]), .B(\d/n217 ), .Z(\d/n215 ) );
  XOR \d/U365  ( .A(shift_row_out[10]), .B(shift_row_out[2]), .Z(\d/n216 ) );
  XOR \d/U364  ( .A(shift_row_out[25]), .B(shift_row_out[18]), .Z(\d/n217 ) );
  XOR \d/U363  ( .A(\d/n219 ), .B(\d/n218 ), .Z(mix_col_out[29]) );
  XOR \d/U362  ( .A(shift_row_out[4]), .B(\d/n341 ), .Z(\d/n218 ) );
  XOR \d/U361  ( .A(shift_row_out[28]), .B(shift_row_out[21]), .Z(\d/n219 ) );
  XOR \d/U360  ( .A(\d/n221 ), .B(\d/n220 ), .Z(mix_col_out[30]) );
  XOR \d/U359  ( .A(shift_row_out[5]), .B(\d/n342 ), .Z(\d/n220 ) );
  XOR \d/U358  ( .A(shift_row_out[29]), .B(shift_row_out[22]), .Z(\d/n221 ) );
  XOR \d/U357  ( .A(\d/n223 ), .B(\d/n222 ), .Z(mix_col_out[31]) );
  XOR \d/U356  ( .A(shift_row_out[6]), .B(\d/n224 ), .Z(\d/n222 ) );
  XOR \d/U355  ( .A(shift_row_out[15]), .B(shift_row_out[7]), .Z(\d/n223 ) );
  XOR \d/U354  ( .A(shift_row_out[30]), .B(shift_row_out[23]), .Z(\d/n224 ) );
  XOR \d/U353  ( .A(shift_row_out[47]), .B(\d/n225 ), .Z(\d/n344 ) );
  XOR \d/U352  ( .A(shift_row_out[56]), .B(shift_row_out[48]), .Z(\d/n225 ) );
  XOR \d/U351  ( .A(\d/n344 ), .B(\d/n226 ), .Z(mix_col_out[32]) );
  XOR \d/U350  ( .A(shift_row_out[40]), .B(shift_row_out[39]), .Z(\d/n226 ) );
  XOR \d/U349  ( .A(shift_row_out[41]), .B(\d/n227 ), .Z(\d/n345 ) );
  XOR \d/U348  ( .A(shift_row_out[58]), .B(shift_row_out[50]), .Z(\d/n227 ) );
  XOR \d/U347  ( .A(\d/n345 ), .B(\d/n228 ), .Z(mix_col_out[34]) );
  XOR \d/U346  ( .A(shift_row_out[42]), .B(shift_row_out[33]), .Z(\d/n228 ) );
  XOR \d/U345  ( .A(shift_row_out[61]), .B(shift_row_out[53]), .Z(\d/n349 ) );
  XOR \d/U344  ( .A(\d/n343 ), .B(\d/n229 ), .Z(mix_col_out[37]) );
  XOR \d/U343  ( .A(shift_row_out[45]), .B(\d/n349 ), .Z(\d/n229 ) );
  XOR \d/U342  ( .A(shift_row_out[62]), .B(shift_row_out[54]), .Z(\d/n350 ) );
  XOR \d/U341  ( .A(shift_row_out[45]), .B(shift_row_out[37]), .Z(\d/n351 ) );
  XOR \d/U340  ( .A(\d/n351 ), .B(\d/n230 ), .Z(mix_col_out[38]) );
  XOR \d/U339  ( .A(shift_row_out[46]), .B(\d/n350 ), .Z(\d/n230 ) );
  XOR \d/U338  ( .A(shift_row_out[63]), .B(shift_row_out[55]), .Z(\d/n346 ) );
  XOR \d/U337  ( .A(shift_row_out[46]), .B(shift_row_out[38]), .Z(\d/n352 ) );
  XOR \d/U336  ( .A(\d/n352 ), .B(\d/n231 ), .Z(mix_col_out[39]) );
  XOR \d/U335  ( .A(shift_row_out[47]), .B(\d/n346 ), .Z(\d/n231 ) );
  XOR \d/U334  ( .A(\d/n344 ), .B(\d/n232 ), .Z(mix_col_out[40]) );
  XOR \d/U333  ( .A(shift_row_out[55]), .B(shift_row_out[32]), .Z(\d/n232 ) );
  XOR \d/U332  ( .A(\d/n345 ), .B(\d/n233 ), .Z(mix_col_out[42]) );
  XOR \d/U331  ( .A(shift_row_out[49]), .B(shift_row_out[34]), .Z(\d/n233 ) );
  XOR \d/U330  ( .A(\d/n235 ), .B(\d/n234 ), .Z(mix_col_out[45]) );
  XOR \d/U329  ( .A(shift_row_out[37]), .B(\d/n349 ), .Z(\d/n234 ) );
  XOR \d/U328  ( .A(shift_row_out[52]), .B(shift_row_out[44]), .Z(\d/n235 ) );
  XOR \d/U327  ( .A(\d/n237 ), .B(\d/n236 ), .Z(mix_col_out[46]) );
  XOR \d/U326  ( .A(shift_row_out[38]), .B(\d/n350 ), .Z(\d/n236 ) );
  XOR \d/U325  ( .A(shift_row_out[53]), .B(shift_row_out[45]), .Z(\d/n237 ) );
  XOR \d/U324  ( .A(\d/n239 ), .B(\d/n238 ), .Z(mix_col_out[47]) );
  XOR \d/U323  ( .A(shift_row_out[39]), .B(\d/n346 ), .Z(\d/n238 ) );
  XOR \d/U322  ( .A(shift_row_out[54]), .B(shift_row_out[46]), .Z(\d/n239 ) );
  XOR \d/U321  ( .A(\d/n241 ), .B(\d/n240 ), .Z(mix_col_out[48]) );
  XOR \d/U320  ( .A(shift_row_out[32]), .B(\d/n346 ), .Z(\d/n240 ) );
  XOR \d/U319  ( .A(shift_row_out[56]), .B(shift_row_out[40]), .Z(\d/n241 ) );
  XOR \d/U318  ( .A(\d/n243 ), .B(\d/n242 ), .Z(mix_col_out[50]) );
  XOR \d/U317  ( .A(shift_row_out[34]), .B(\d/n347 ), .Z(\d/n242 ) );
  XOR \d/U316  ( .A(shift_row_out[58]), .B(shift_row_out[42]), .Z(\d/n243 ) );
  XOR \d/U315  ( .A(\d/n351 ), .B(\d/n244 ), .Z(mix_col_out[53]) );
  XOR \d/U314  ( .A(shift_row_out[61]), .B(\d/n348 ), .Z(\d/n244 ) );
  XOR \d/U313  ( .A(\d/n352 ), .B(\d/n245 ), .Z(mix_col_out[54]) );
  XOR \d/U312  ( .A(shift_row_out[62]), .B(\d/n349 ), .Z(\d/n245 ) );
  XOR \d/U311  ( .A(\d/n247 ), .B(\d/n246 ), .Z(mix_col_out[55]) );
  XOR \d/U310  ( .A(shift_row_out[39]), .B(\d/n350 ), .Z(\d/n246 ) );
  XOR \d/U309  ( .A(shift_row_out[63]), .B(shift_row_out[47]), .Z(\d/n247 ) );
  XOR \d/U308  ( .A(\d/n249 ), .B(\d/n248 ), .Z(mix_col_out[56]) );
  XOR \d/U307  ( .A(shift_row_out[32]), .B(\d/n250 ), .Z(\d/n248 ) );
  XOR \d/U306  ( .A(shift_row_out[40]), .B(shift_row_out[39]), .Z(\d/n249 ) );
  XOR \d/U305  ( .A(shift_row_out[63]), .B(shift_row_out[48]), .Z(\d/n250 ) );
  XOR \d/U304  ( .A(\d/n252 ), .B(\d/n251 ), .Z(mix_col_out[58]) );
  XOR \d/U303  ( .A(shift_row_out[33]), .B(\d/n253 ), .Z(\d/n251 ) );
  XOR \d/U302  ( .A(shift_row_out[42]), .B(shift_row_out[34]), .Z(\d/n252 ) );
  XOR \d/U301  ( .A(shift_row_out[57]), .B(shift_row_out[50]), .Z(\d/n253 ) );
  XOR \d/U300  ( .A(\d/n255 ), .B(\d/n254 ), .Z(mix_col_out[61]) );
  XOR \d/U299  ( .A(shift_row_out[36]), .B(\d/n351 ), .Z(\d/n254 ) );
  XOR \d/U298  ( .A(shift_row_out[60]), .B(shift_row_out[53]), .Z(\d/n255 ) );
  XOR \d/U297  ( .A(\d/n257 ), .B(\d/n256 ), .Z(mix_col_out[62]) );
  XOR \d/U296  ( .A(shift_row_out[37]), .B(\d/n352 ), .Z(\d/n256 ) );
  XOR \d/U295  ( .A(shift_row_out[61]), .B(shift_row_out[54]), .Z(\d/n257 ) );
  XOR \d/U294  ( .A(\d/n259 ), .B(\d/n258 ), .Z(mix_col_out[63]) );
  XOR \d/U293  ( .A(shift_row_out[38]), .B(\d/n260 ), .Z(\d/n258 ) );
  XOR \d/U292  ( .A(shift_row_out[47]), .B(shift_row_out[39]), .Z(\d/n259 ) );
  XOR \d/U291  ( .A(shift_row_out[62]), .B(shift_row_out[55]), .Z(\d/n260 ) );
  XOR \d/U290  ( .A(shift_row_out[79]), .B(\d/n261 ), .Z(\d/n354 ) );
  XOR \d/U289  ( .A(shift_row_out[88]), .B(shift_row_out[80]), .Z(\d/n261 ) );
  XOR \d/U288  ( .A(\d/n354 ), .B(\d/n262 ), .Z(mix_col_out[64]) );
  XOR \d/U287  ( .A(shift_row_out[72]), .B(shift_row_out[71]), .Z(\d/n262 ) );
  XOR \d/U286  ( .A(shift_row_out[73]), .B(\d/n263 ), .Z(\d/n355 ) );
  XOR \d/U285  ( .A(shift_row_out[90]), .B(shift_row_out[82]), .Z(\d/n263 ) );
  XOR \d/U284  ( .A(\d/n355 ), .B(\d/n264 ), .Z(mix_col_out[66]) );
  XOR \d/U283  ( .A(shift_row_out[74]), .B(shift_row_out[65]), .Z(\d/n264 ) );
  XOR \d/U282  ( .A(shift_row_out[93]), .B(shift_row_out[85]), .Z(\d/n359 ) );
  XOR \d/U281  ( .A(\d/n353 ), .B(\d/n265 ), .Z(mix_col_out[69]) );
  XOR \d/U280  ( .A(shift_row_out[77]), .B(\d/n359 ), .Z(\d/n265 ) );
  XOR \d/U279  ( .A(shift_row_out[94]), .B(shift_row_out[86]), .Z(\d/n360 ) );
  XOR \d/U278  ( .A(shift_row_out[77]), .B(shift_row_out[69]), .Z(\d/n361 ) );
  XOR \d/U277  ( .A(\d/n361 ), .B(\d/n266 ), .Z(mix_col_out[70]) );
  XOR \d/U276  ( .A(shift_row_out[78]), .B(\d/n360 ), .Z(\d/n266 ) );
  XOR \d/U275  ( .A(shift_row_out[95]), .B(shift_row_out[87]), .Z(\d/n356 ) );
  XOR \d/U274  ( .A(shift_row_out[78]), .B(shift_row_out[70]), .Z(\d/n362 ) );
  XOR \d/U273  ( .A(\d/n362 ), .B(\d/n267 ), .Z(mix_col_out[71]) );
  XOR \d/U272  ( .A(shift_row_out[79]), .B(\d/n356 ), .Z(\d/n267 ) );
  XOR \d/U271  ( .A(\d/n354 ), .B(\d/n268 ), .Z(mix_col_out[72]) );
  XOR \d/U270  ( .A(shift_row_out[87]), .B(shift_row_out[64]), .Z(\d/n268 ) );
  XOR \d/U269  ( .A(\d/n355 ), .B(\d/n269 ), .Z(mix_col_out[74]) );
  XOR \d/U268  ( .A(shift_row_out[81]), .B(shift_row_out[66]), .Z(\d/n269 ) );
  XOR \d/U267  ( .A(\d/n271 ), .B(\d/n270 ), .Z(mix_col_out[77]) );
  XOR \d/U266  ( .A(shift_row_out[69]), .B(\d/n359 ), .Z(\d/n270 ) );
  XOR \d/U265  ( .A(shift_row_out[84]), .B(shift_row_out[76]), .Z(\d/n271 ) );
  XOR \d/U264  ( .A(\d/n273 ), .B(\d/n272 ), .Z(mix_col_out[78]) );
  XOR \d/U263  ( .A(shift_row_out[70]), .B(\d/n360 ), .Z(\d/n272 ) );
  XOR \d/U262  ( .A(shift_row_out[85]), .B(shift_row_out[77]), .Z(\d/n273 ) );
  XOR \d/U261  ( .A(\d/n275 ), .B(\d/n274 ), .Z(mix_col_out[79]) );
  XOR \d/U260  ( .A(shift_row_out[71]), .B(\d/n356 ), .Z(\d/n274 ) );
  XOR \d/U259  ( .A(shift_row_out[86]), .B(shift_row_out[78]), .Z(\d/n275 ) );
  XOR \d/U258  ( .A(\d/n277 ), .B(\d/n276 ), .Z(mix_col_out[80]) );
  XOR \d/U257  ( .A(shift_row_out[64]), .B(\d/n356 ), .Z(\d/n276 ) );
  XOR \d/U256  ( .A(shift_row_out[88]), .B(shift_row_out[72]), .Z(\d/n277 ) );
  XOR \d/U255  ( .A(\d/n279 ), .B(\d/n278 ), .Z(mix_col_out[82]) );
  XOR \d/U254  ( .A(shift_row_out[66]), .B(\d/n357 ), .Z(\d/n278 ) );
  XOR \d/U253  ( .A(shift_row_out[90]), .B(shift_row_out[74]), .Z(\d/n279 ) );
  XOR \d/U252  ( .A(\d/n361 ), .B(\d/n280 ), .Z(mix_col_out[85]) );
  XOR \d/U251  ( .A(shift_row_out[93]), .B(\d/n358 ), .Z(\d/n280 ) );
  XOR \d/U250  ( .A(\d/n362 ), .B(\d/n281 ), .Z(mix_col_out[86]) );
  XOR \d/U249  ( .A(shift_row_out[94]), .B(\d/n359 ), .Z(\d/n281 ) );
  XOR \d/U248  ( .A(\d/n283 ), .B(\d/n282 ), .Z(mix_col_out[87]) );
  XOR \d/U247  ( .A(shift_row_out[71]), .B(\d/n360 ), .Z(\d/n282 ) );
  XOR \d/U246  ( .A(shift_row_out[95]), .B(shift_row_out[79]), .Z(\d/n283 ) );
  XOR \d/U245  ( .A(\d/n285 ), .B(\d/n284 ), .Z(mix_col_out[88]) );
  XOR \d/U244  ( .A(shift_row_out[64]), .B(\d/n286 ), .Z(\d/n284 ) );
  XOR \d/U243  ( .A(shift_row_out[72]), .B(shift_row_out[71]), .Z(\d/n285 ) );
  XOR \d/U242  ( .A(shift_row_out[95]), .B(shift_row_out[80]), .Z(\d/n286 ) );
  XOR \d/U241  ( .A(\d/n288 ), .B(\d/n287 ), .Z(mix_col_out[90]) );
  XOR \d/U240  ( .A(shift_row_out[65]), .B(\d/n289 ), .Z(\d/n287 ) );
  XOR \d/U239  ( .A(shift_row_out[74]), .B(shift_row_out[66]), .Z(\d/n288 ) );
  XOR \d/U238  ( .A(shift_row_out[89]), .B(shift_row_out[82]), .Z(\d/n289 ) );
  XOR \d/U237  ( .A(\d/n291 ), .B(\d/n290 ), .Z(mix_col_out[93]) );
  XOR \d/U236  ( .A(shift_row_out[68]), .B(\d/n361 ), .Z(\d/n290 ) );
  XOR \d/U235  ( .A(shift_row_out[92]), .B(shift_row_out[85]), .Z(\d/n291 ) );
  XOR \d/U234  ( .A(\d/n293 ), .B(\d/n292 ), .Z(mix_col_out[94]) );
  XOR \d/U233  ( .A(shift_row_out[69]), .B(\d/n362 ), .Z(\d/n292 ) );
  XOR \d/U232  ( .A(shift_row_out[93]), .B(shift_row_out[86]), .Z(\d/n293 ) );
  XOR \d/U231  ( .A(\d/n295 ), .B(\d/n294 ), .Z(mix_col_out[95]) );
  XOR \d/U230  ( .A(shift_row_out[70]), .B(\d/n296 ), .Z(\d/n294 ) );
  XOR \d/U229  ( .A(shift_row_out[79]), .B(shift_row_out[71]), .Z(\d/n295 ) );
  XOR \d/U228  ( .A(shift_row_out[94]), .B(shift_row_out[87]), .Z(\d/n296 ) );
  XOR \d/U227  ( .A(shift_row_out[111]), .B(\d/n297 ), .Z(\d/n364 ) );
  XOR \d/U226  ( .A(shift_row_out[120]), .B(shift_row_out[112]), .Z(\d/n297 )
         );
  XOR \d/U225  ( .A(\d/n364 ), .B(\d/n298 ), .Z(mix_col_out[96]) );
  XOR \d/U224  ( .A(shift_row_out[104]), .B(shift_row_out[103]), .Z(\d/n298 )
         );
  XOR \d/U223  ( .A(shift_row_out[105]), .B(\d/n299 ), .Z(\d/n365 ) );
  XOR \d/U222  ( .A(shift_row_out[122]), .B(shift_row_out[114]), .Z(\d/n299 )
         );
  XOR \d/U221  ( .A(\d/n365 ), .B(\d/n300 ), .Z(mix_col_out[98]) );
  XOR \d/U220  ( .A(shift_row_out[106]), .B(shift_row_out[97]), .Z(\d/n300 )
         );
  XOR \d/U219  ( .A(shift_row_out[125]), .B(shift_row_out[117]), .Z(\d/n369 )
         );
  XOR \d/U218  ( .A(\d/n363 ), .B(\d/n301 ), .Z(mix_col_out[101]) );
  XOR \d/U217  ( .A(shift_row_out[109]), .B(\d/n369 ), .Z(\d/n301 ) );
  XOR \d/U216  ( .A(shift_row_out[126]), .B(shift_row_out[118]), .Z(\d/n370 )
         );
  XOR \d/U215  ( .A(shift_row_out[109]), .B(shift_row_out[101]), .Z(\d/n371 )
         );
  XOR \d/U214  ( .A(\d/n371 ), .B(\d/n302 ), .Z(mix_col_out[102]) );
  XOR \d/U213  ( .A(shift_row_out[110]), .B(\d/n370 ), .Z(\d/n302 ) );
  XOR \d/U212  ( .A(shift_row_out[127]), .B(shift_row_out[119]), .Z(\d/n366 )
         );
  XOR \d/U211  ( .A(shift_row_out[110]), .B(shift_row_out[102]), .Z(\d/n372 )
         );
  XOR \d/U210  ( .A(\d/n372 ), .B(\d/n303 ), .Z(mix_col_out[103]) );
  XOR \d/U209  ( .A(shift_row_out[111]), .B(\d/n366 ), .Z(\d/n303 ) );
  XOR \d/U208  ( .A(\d/n364 ), .B(\d/n304 ), .Z(mix_col_out[104]) );
  XOR \d/U207  ( .A(shift_row_out[119]), .B(shift_row_out[96]), .Z(\d/n304 )
         );
  XOR \d/U206  ( .A(\d/n365 ), .B(\d/n305 ), .Z(mix_col_out[106]) );
  XOR \d/U205  ( .A(shift_row_out[113]), .B(shift_row_out[98]), .Z(\d/n305 )
         );
  XOR \d/U204  ( .A(\d/n307 ), .B(\d/n306 ), .Z(mix_col_out[109]) );
  XOR \d/U203  ( .A(shift_row_out[101]), .B(\d/n369 ), .Z(\d/n306 ) );
  XOR \d/U202  ( .A(shift_row_out[116]), .B(shift_row_out[108]), .Z(\d/n307 )
         );
  XOR \d/U201  ( .A(\d/n309 ), .B(\d/n308 ), .Z(mix_col_out[110]) );
  XOR \d/U200  ( .A(shift_row_out[102]), .B(\d/n370 ), .Z(\d/n308 ) );
  XOR \d/U199  ( .A(shift_row_out[117]), .B(shift_row_out[109]), .Z(\d/n309 )
         );
  XOR \d/U198  ( .A(\d/n311 ), .B(\d/n310 ), .Z(mix_col_out[111]) );
  XOR \d/U197  ( .A(shift_row_out[103]), .B(\d/n366 ), .Z(\d/n310 ) );
  XOR \d/U196  ( .A(shift_row_out[118]), .B(shift_row_out[110]), .Z(\d/n311 )
         );
  XOR \d/U195  ( .A(\d/n313 ), .B(\d/n312 ), .Z(mix_col_out[112]) );
  XOR \d/U194  ( .A(shift_row_out[96]), .B(\d/n366 ), .Z(\d/n312 ) );
  XOR \d/U193  ( .A(shift_row_out[120]), .B(shift_row_out[104]), .Z(\d/n313 )
         );
  XOR \d/U192  ( .A(\d/n315 ), .B(\d/n314 ), .Z(mix_col_out[114]) );
  XOR \d/U191  ( .A(shift_row_out[98]), .B(\d/n367 ), .Z(\d/n314 ) );
  XOR \d/U190  ( .A(shift_row_out[122]), .B(shift_row_out[106]), .Z(\d/n315 )
         );
  XOR \d/U189  ( .A(\d/n371 ), .B(\d/n316 ), .Z(mix_col_out[117]) );
  XOR \d/U188  ( .A(shift_row_out[125]), .B(\d/n368 ), .Z(\d/n316 ) );
  XOR \d/U187  ( .A(\d/n372 ), .B(\d/n317 ), .Z(mix_col_out[118]) );
  XOR \d/U186  ( .A(shift_row_out[126]), .B(\d/n369 ), .Z(\d/n317 ) );
  XOR \d/U185  ( .A(\d/n319 ), .B(\d/n318 ), .Z(mix_col_out[119]) );
  XOR \d/U184  ( .A(shift_row_out[103]), .B(\d/n370 ), .Z(\d/n318 ) );
  XOR \d/U183  ( .A(shift_row_out[127]), .B(shift_row_out[111]), .Z(\d/n319 )
         );
  XOR \d/U182  ( .A(\d/n321 ), .B(\d/n320 ), .Z(mix_col_out[120]) );
  XOR \d/U181  ( .A(shift_row_out[96]), .B(\d/n322 ), .Z(\d/n320 ) );
  XOR \d/U180  ( .A(shift_row_out[104]), .B(shift_row_out[103]), .Z(\d/n321 )
         );
  XOR \d/U179  ( .A(shift_row_out[127]), .B(shift_row_out[112]), .Z(\d/n322 )
         );
  XOR \d/U178  ( .A(\d/n324 ), .B(\d/n323 ), .Z(mix_col_out[122]) );
  XOR \d/U177  ( .A(shift_row_out[97]), .B(\d/n325 ), .Z(\d/n323 ) );
  XOR \d/U176  ( .A(shift_row_out[106]), .B(shift_row_out[98]), .Z(\d/n324 )
         );
  XOR \d/U175  ( .A(shift_row_out[121]), .B(shift_row_out[114]), .Z(\d/n325 )
         );
  XOR \d/U174  ( .A(\d/n327 ), .B(\d/n326 ), .Z(mix_col_out[125]) );
  XOR \d/U173  ( .A(shift_row_out[100]), .B(\d/n371 ), .Z(\d/n326 ) );
  XOR \d/U172  ( .A(shift_row_out[124]), .B(shift_row_out[117]), .Z(\d/n327 )
         );
  XOR \d/U171  ( .A(\d/n329 ), .B(\d/n328 ), .Z(mix_col_out[126]) );
  XOR \d/U170  ( .A(shift_row_out[101]), .B(\d/n372 ), .Z(\d/n328 ) );
  XOR \d/U169  ( .A(shift_row_out[125]), .B(shift_row_out[118]), .Z(\d/n329 )
         );
  XOR \d/U168  ( .A(\d/n331 ), .B(\d/n330 ), .Z(mix_col_out[127]) );
  XOR \d/U167  ( .A(shift_row_out[102]), .B(\d/n332 ), .Z(\d/n330 ) );
  XOR \d/U166  ( .A(shift_row_out[111]), .B(shift_row_out[103]), .Z(\d/n331 )
         );
  XOR \d/U165  ( .A(shift_row_out[126]), .B(shift_row_out[119]), .Z(\d/n332 )
         );
  MUX \e/a/U7005  ( .IN0(key[100]), .IN1(n2736), .SEL(key[97]), .F(n3082) );
  MUX \e/a/U7004  ( .IN0(key[100]), .IN1(n2745), .SEL(key[97]), .F(n3081) );
  MUX \e/a/U7003  ( .IN0(n2737), .IN1(n2740), .SEL(key[97]), .F(n3080) );
  MUX \e/a/U7002  ( .IN0(n2742), .IN1(n1518), .SEL(key[97]), .F(n3079) );
  MUX \e/a/U7000  ( .IN0(n2745), .IN1(n2736), .SEL(key[98]), .F(n2914) );
  MUX \e/a/U6999  ( .IN0(n2738), .IN1(n1528), .SEL(key[98]), .F(n2915) );
  MUX \e/a/U6998  ( .IN0(n1482), .IN1(n1490), .SEL(key[97]), .F(n2878) );
  MUX \e/a/U6997  ( .IN0(n2764), .IN1(n3070), .SEL(key[103]), .F(n3078) );
  MUX \e/a/U6996  ( .IN0(n2740), .IN1(n2736), .SEL(key[97]), .F(n3072) );
  MUX \e/a/U6995  ( .IN0(n1524), .IN1(n2742), .SEL(key[97]), .F(n3077) );
  MUX \e/a/U6994  ( .IN0(key[99]), .IN1(n1518), .SEL(key[97]), .F(n3076) );
  MUX \e/a/U6993  ( .IN0(n2745), .IN1(n1524), .SEL(key[97]), .F(n3075) );
  MUX \e/a/U6992  ( .IN0(key[100]), .IN1(n2742), .SEL(key[97]), .F(n3074) );
  MUX \e/a/U6991  ( .IN0(n1510), .IN1(n1494), .SEL(key[101]), .F(n2788) );
  MUX \e/a/U6990  ( .IN0(n2737), .IN1(n1490), .SEL(key[97]), .F(n3073) );
  NANDN \e/a/U6987  ( .B(n2743), .A(key[103]), .Z(n3053) );
  NAND \e/a/U6986  ( .A(key[103]), .B(n1491), .Z(n3021) );
  NAND \e/a/U6985  ( .A(key[103]), .B(n1500), .Z(n2962) );
  NAND \e/a/U6984  ( .A(key[103]), .B(n3068), .Z(n2995) );
  NAND \e/a/U6983  ( .A(key[103]), .B(n2990), .Z(n2953) );
  NAND \e/a/U6981  ( .A(n1528), .B(n1518), .Z(n3071) );
  NAND \e/a/U6980  ( .A(key[103]), .B(n3069), .Z(n3067) );
  NAND \e/a/U6979  ( .A(n600), .B(key[103]), .Z(n3047) );
  NAND \e/a/U6977  ( .A(key[98]), .B(n2745), .Z(n2907) );
  NAND \e/a/U6976  ( .A(n1518), .B(key[97]), .Z(n2862) );
  NAND \e/a/U6975  ( .A(key[103]), .B(n3072), .Z(n2861) );
  NAND \e/a/U6973  ( .A(n3071), .B(key[103]), .Z(n2877) );
  NAND \e/a/U6972  ( .A(n2895), .B(n2745), .Z(n3070) );
  NANDN \e/a/U6971  ( .B(n1482), .A(n1528), .Z(n3069) );
  NAND \e/a/U6969  ( .A(key[97]), .B(n2745), .Z(n2793) );
  NAND \e/a/U6968  ( .A(n1482), .B(n1528), .Z(n3068) );
  NAND \e/a/U6965  ( .A(key[97]), .B(n2740), .Z(n2895) );
  ANDN \e/a/U6963  ( .A(key[98]), .B(key[97]), .Z(n2923) );
  AND \e/a/U6962  ( .A(n2737), .B(n3067), .Z(n2838) );
  MUX \e/a/U6961  ( .IN0(n3066), .IN1(n3050), .SEL(key[102]), .F(\e/t[31] ) );
  MUX \e/a/U6960  ( .IN0(n3065), .IN1(n3058), .SEL(key[96]), .F(n3066) );
  MUX \e/a/U6959  ( .IN0(n3064), .IN1(n3061), .SEL(key[101]), .F(n3065) );
  MUX \e/a/U6958  ( .IN0(n3063), .IN1(n3062), .SEL(key[98]), .F(n3064) );
  MUX \e/a/U6957  ( .IN0(key[100]), .IN1(n1495), .SEL(key[103]), .F(n3063) );
  MUX \e/a/U6956  ( .IN0(n2738), .IN1(n1497), .SEL(key[103]), .F(n3062) );
  MUX \e/a/U6955  ( .IN0(n3060), .IN1(n3059), .SEL(key[98]), .F(n3061) );
  MUX \e/a/U6954  ( .IN0(n2792), .IN1(n1491), .SEL(key[103]), .F(n3060) );
  MUX \e/a/U6953  ( .IN0(n2748), .IN1(n2757), .SEL(key[103]), .F(n3059) );
  MUX \e/a/U6952  ( .IN0(n3057), .IN1(n3054), .SEL(key[101]), .F(n3058) );
  MUX \e/a/U6951  ( .IN0(n3056), .IN1(n3055), .SEL(key[98]), .F(n3057) );
  MUX \e/a/U6950  ( .IN0(n2769), .IN1(n2747), .SEL(key[103]), .F(n3056) );
  MUX \e/a/U6949  ( .IN0(n1500), .IN1(n2766), .SEL(key[103]), .F(n3055) );
  MUX \e/a/U6948  ( .IN0(n3052), .IN1(n3051), .SEL(key[98]), .F(n3054) );
  AND \e/a/U6947  ( .A(n1493), .B(n3053), .Z(n3052) );
  MUX \e/a/U6946  ( .IN0(n2752), .IN1(n599), .SEL(key[103]), .F(n3051) );
  MUX \e/a/U6945  ( .IN0(n3049), .IN1(n3041), .SEL(key[96]), .F(n3050) );
  MUX \e/a/U6944  ( .IN0(n3048), .IN1(n3044), .SEL(key[101]), .F(n3049) );
  MUX \e/a/U6943  ( .IN0(n3045), .IN1(n3046), .SEL(key[98]), .F(n3048) );
  NAND \e/a/U6942  ( .A(n2862), .B(n3047), .Z(n3046) );
  MUX \e/a/U6941  ( .IN0(n1527), .IN1(n1519), .SEL(key[103]), .F(n3045) );
  MUX \e/a/U6940  ( .IN0(n3043), .IN1(n3042), .SEL(key[98]), .F(n3044) );
  MUX \e/a/U6939  ( .IN0(n2742), .IN1(n2736), .SEL(key[103]), .F(n3043) );
  MUX \e/a/U6938  ( .IN0(n1520), .IN1(n2770), .SEL(key[103]), .F(n3042) );
  MUX \e/a/U6937  ( .IN0(n3040), .IN1(n3037), .SEL(key[101]), .F(n3041) );
  MUX \e/a/U6936  ( .IN0(n3039), .IN1(n3038), .SEL(key[98]), .F(n3040) );
  MUX \e/a/U6935  ( .IN0(n2773), .IN1(n2761), .SEL(key[103]), .F(n3039) );
  MUX \e/a/U6934  ( .IN0(n1483), .IN1(n2745), .SEL(key[103]), .F(n3038) );
  MUX \e/a/U6933  ( .IN0(n3036), .IN1(n3035), .SEL(key[98]), .F(n3037) );
  MUX \e/a/U6932  ( .IN0(n2774), .IN1(n2782), .SEL(key[103]), .F(n3036) );
  MUX \e/a/U6931  ( .IN0(n2768), .IN1(n3034), .SEL(key[103]), .F(n3035) );
  MUX \e/a/U6930  ( .IN0(n1524), .IN1(n1490), .SEL(key[97]), .F(n3034) );
  MUX \e/a/U6929  ( .IN0(n3033), .IN1(n3015), .SEL(key[102]), .F(\e/t[30] ) );
  MUX \e/a/U6928  ( .IN0(n3032), .IN1(n3023), .SEL(key[96]), .F(n3033) );
  MUX \e/a/U6927  ( .IN0(n3031), .IN1(n3026), .SEL(key[101]), .F(n3032) );
  MUX \e/a/U6926  ( .IN0(n3030), .IN1(n3028), .SEL(key[98]), .F(n3031) );
  MUX \e/a/U6925  ( .IN0(n3029), .IN1(n2749), .SEL(key[103]), .F(n3030) );
  MUX \e/a/U6924  ( .IN0(n1524), .IN1(n2736), .SEL(key[97]), .F(n3029) );
  MUX \e/a/U6923  ( .IN0(n3027), .IN1(n1512), .SEL(key[103]), .F(n3028) );
  MUX \e/a/U6922  ( .IN0(n2736), .IN1(n2737), .SEL(key[97]), .F(n3027) );
  MUX \e/a/U6921  ( .IN0(n3025), .IN1(n3024), .SEL(key[98]), .F(n3026) );
  MUX \e/a/U6920  ( .IN0(n598), .IN1(n2813), .SEL(key[103]), .F(n3025) );
  MUX \e/a/U6919  ( .IN0(n2772), .IN1(n2778), .SEL(key[103]), .F(n3024) );
  MUX \e/a/U6918  ( .IN0(n3022), .IN1(n3018), .SEL(key[101]), .F(n3023) );
  MUX \e/a/U6917  ( .IN0(n3020), .IN1(n3019), .SEL(key[98]), .F(n3022) );
  AND \e/a/U6916  ( .A(n1477), .B(n3021), .Z(n3020) );
  MUX \e/a/U6915  ( .IN0(n2848), .IN1(key[99]), .SEL(key[103]), .F(n3019) );
  MUX \e/a/U6914  ( .IN0(n3017), .IN1(n3016), .SEL(key[98]), .F(n3018) );
  MUX \e/a/U6913  ( .IN0(n1509), .IN1(n2740), .SEL(key[103]), .F(n3017) );
  MUX \e/a/U6911  ( .IN0(n3014), .IN1(n3007), .SEL(key[96]), .F(n3015) );
  MUX \e/a/U6910  ( .IN0(n3013), .IN1(n3010), .SEL(key[101]), .F(n3014) );
  MUX \e/a/U6909  ( .IN0(n3012), .IN1(n3011), .SEL(key[98]), .F(n3013) );
  MUX \e/a/U6908  ( .IN0(n1505), .IN1(n2744), .SEL(key[103]), .F(n3012) );
  MUX \e/a/U6907  ( .IN0(n2748), .IN1(n599), .SEL(key[103]), .F(n3011) );
  MUX \e/a/U6906  ( .IN0(n3009), .IN1(n3008), .SEL(key[98]), .F(n3010) );
  MUX \e/a/U6905  ( .IN0(n2762), .IN1(n1480), .SEL(key[103]), .F(n3009) );
  MUX \e/a/U6904  ( .IN0(n1495), .IN1(n1519), .SEL(key[103]), .F(n3008) );
  MUX \e/a/U6903  ( .IN0(n3006), .IN1(n3002), .SEL(key[101]), .F(n3007) );
  MUX \e/a/U6902  ( .IN0(n3005), .IN1(n3004), .SEL(key[98]), .F(n3006) );
  MUX \e/a/U6901  ( .IN0(n2753), .IN1(n1519), .SEL(key[103]), .F(n3005) );
  MUX \e/a/U6900  ( .IN0(n3003), .IN1(n2771), .SEL(key[103]), .F(n3004) );
  NANDN \e/a/U6899  ( .B(key[100]), .A(key[97]), .Z(n3003) );
  MUX \e/a/U6898  ( .IN0(n3001), .IN1(n2999), .SEL(key[98]), .F(n3002) );
  MUX \e/a/U6897  ( .IN0(n1490), .IN1(n3000), .SEL(key[103]), .F(n3001) );
  MUX \e/a/U6896  ( .IN0(n1510), .IN1(n1501), .SEL(key[97]), .F(n3000) );
  MUX \e/a/U6895  ( .IN0(n1481), .IN1(n2749), .SEL(key[103]), .F(n2999) );
  NANDN \e/a/U6894  ( .B(n1482), .A(key[97]), .Z(n2749) );
  MUX \e/a/U6893  ( .IN0(n2998), .IN1(n2977), .SEL(key[102]), .F(\e/t[29] ) );
  MUX \e/a/U6892  ( .IN0(n2997), .IN1(n2987), .SEL(key[96]), .F(n2998) );
  MUX \e/a/U6891  ( .IN0(n2996), .IN1(n2992), .SEL(key[101]), .F(n2997) );
  MUX \e/a/U6890  ( .IN0(n2993), .IN1(n2994), .SEL(key[98]), .F(n2996) );
  AND \e/a/U6889  ( .A(n2765), .B(n2995), .Z(n2994) );
  MUX \e/a/U6888  ( .IN0(n2745), .IN1(n1520), .SEL(key[103]), .F(n2993) );
  MUX \e/a/U6887  ( .IN0(n2991), .IN1(n2989), .SEL(key[98]), .F(n2992) );
  MUX \e/a/U6886  ( .IN0(n1485), .IN1(n2990), .SEL(key[103]), .F(n2991) );
  NAND \e/a/U6885  ( .A(n1501), .B(n1528), .Z(n2990) );
  MUX \e/a/U6884  ( .IN0(n2745), .IN1(n2988), .SEL(key[103]), .F(n2989) );
  NAND \e/a/U6883  ( .A(n2736), .B(n2793), .Z(n2988) );
  MUX \e/a/U6882  ( .IN0(n2986), .IN1(n2982), .SEL(key[101]), .F(n2987) );
  MUX \e/a/U6881  ( .IN0(n2985), .IN1(n2984), .SEL(key[98]), .F(n2986) );
  MUX \e/a/U6880  ( .IN0(n2756), .IN1(n1522), .SEL(key[103]), .F(n2985) );
  MUX \e/a/U6879  ( .IN0(n2778), .IN1(n2983), .SEL(key[103]), .F(n2984) );
  MUX \e/a/U6878  ( .IN0(n1518), .IN1(n1501), .SEL(key[97]), .F(n2983) );
  MUX \e/a/U6877  ( .IN0(n2981), .IN1(n2980), .SEL(key[98]), .F(n2982) );
  MUX \e/a/U6876  ( .IN0(n1516), .IN1(n597), .SEL(key[103]), .F(n2981) );
  MUX \e/a/U6875  ( .IN0(n2979), .IN1(n2978), .SEL(key[103]), .F(n2980) );
  AND \e/a/U6874  ( .A(n2742), .B(n2813), .Z(n2979) );
  MUX \e/a/U6873  ( .IN0(n1494), .IN1(n1482), .SEL(key[97]), .F(n2978) );
  MUX \e/a/U6872  ( .IN0(n2976), .IN1(n2967), .SEL(key[96]), .F(n2977) );
  MUX \e/a/U6871  ( .IN0(n2975), .IN1(n2971), .SEL(key[101]), .F(n2976) );
  MUX \e/a/U6870  ( .IN0(n2974), .IN1(n2972), .SEL(key[98]), .F(n2975) );
  MUX \e/a/U6869  ( .IN0(n2748), .IN1(n2973), .SEL(key[103]), .F(n2974) );
  NAND \e/a/U6868  ( .A(key[97]), .B(n1494), .Z(n2973) );
  MUX \e/a/U6867  ( .IN0(n1482), .IN1(n1525), .SEL(key[103]), .F(n2972) );
  MUX \e/a/U6866  ( .IN0(n2970), .IN1(n2969), .SEL(key[98]), .F(n2971) );
  MUX \e/a/U6865  ( .IN0(n2771), .IN1(n1496), .SEL(key[103]), .F(n2970) );
  MUX \e/a/U6864  ( .IN0(n2968), .IN1(n2737), .SEL(n596), .F(n2969) );
  AND \e/a/U6863  ( .A(key[103]), .B(key[99]), .Z(n2968) );
  MUX \e/a/U6862  ( .IN0(n2966), .IN1(n2963), .SEL(key[101]), .F(n2967) );
  MUX \e/a/U6861  ( .IN0(n2965), .IN1(n2964), .SEL(key[98]), .F(n2966) );
  MUX \e/a/U6860  ( .IN0(n2894), .IN1(n2737), .SEL(key[103]), .F(n2965) );
  MUX \e/a/U6859  ( .IN0(n595), .IN1(n1523), .SEL(key[103]), .F(n2964) );
  MUX \e/a/U6858  ( .IN0(n2961), .IN1(n2960), .SEL(key[98]), .F(n2963) );
  AND \e/a/U6857  ( .A(n2962), .B(n2862), .Z(n2961) );
  MUX \e/a/U6856  ( .IN0(n1484), .IN1(n1518), .SEL(key[103]), .F(n2960) );
  MUX \e/a/U6855  ( .IN0(n2959), .IN1(n2942), .SEL(key[102]), .F(\e/t[28] ) );
  MUX \e/a/U6854  ( .IN0(n2958), .IN1(n2950), .SEL(key[96]), .F(n2959) );
  MUX \e/a/U6853  ( .IN0(n2957), .IN1(n2954), .SEL(key[101]), .F(n2958) );
  MUX \e/a/U6852  ( .IN0(n2956), .IN1(n2955), .SEL(key[98]), .F(n2957) );
  MUX \e/a/U6851  ( .IN0(n1502), .IN1(n1521), .SEL(key[103]), .F(n2956) );
  MUX \e/a/U6850  ( .IN0(n2813), .IN1(n2778), .SEL(key[103]), .F(n2955) );
  NAND \e/a/U6849  ( .A(key[97]), .B(n2736), .Z(n2813) );
  MUX \e/a/U6848  ( .IN0(n2951), .IN1(n2952), .SEL(key[98]), .F(n2954) );
  AND \e/a/U6847  ( .A(n2765), .B(n2953), .Z(n2952) );
  MUX \e/a/U6846  ( .IN0(n2763), .IN1(n1504), .SEL(key[103]), .F(n2951) );
  MUX \e/a/U6845  ( .IN0(n2949), .IN1(n2946), .SEL(key[101]), .F(n2950) );
  MUX \e/a/U6844  ( .IN0(n2948), .IN1(n2947), .SEL(key[98]), .F(n2949) );
  MUX \e/a/U6843  ( .IN0(n1477), .IN1(n1511), .SEL(key[103]), .F(n2948) );
  MUX \e/a/U6842  ( .IN0(n1482), .IN1(n2745), .SEL(key[103]), .F(n2947) );
  MUX \e/a/U6841  ( .IN0(n2945), .IN1(n2943), .SEL(key[98]), .F(n2946) );
  MUX \e/a/U6840  ( .IN0(n2759), .IN1(n2944), .SEL(key[103]), .F(n2945) );
  AND \e/a/U6839  ( .A(n2745), .B(n1528), .Z(n2944) );
  MUX \e/a/U6838  ( .IN0(n1493), .IN1(n1507), .SEL(key[103]), .F(n2943) );
  MUX \e/a/U6837  ( .IN0(n2941), .IN1(n2935), .SEL(key[96]), .F(n2942) );
  MUX \e/a/U6836  ( .IN0(n2940), .IN1(n2938), .SEL(key[101]), .F(n2941) );
  MUX \e/a/U6835  ( .IN0(n2939), .IN1(n2739), .SEL(key[98]), .F(n2940) );
  MUX \e/a/U6834  ( .IN0(n2757), .IN1(n1509), .SEL(key[103]), .F(n2939) );
  MUX \e/a/U6833  ( .IN0(n2937), .IN1(n2936), .SEL(key[98]), .F(n2938) );
  MUX \e/a/U6832  ( .IN0(n594), .IN1(n1502), .SEL(key[103]), .F(n2937) );
  MUX \e/a/U6831  ( .IN0(n2767), .IN1(n2769), .SEL(key[103]), .F(n2936) );
  MUX \e/a/U6830  ( .IN0(n2934), .IN1(n2931), .SEL(key[101]), .F(n2935) );
  MUX \e/a/U6829  ( .IN0(n2933), .IN1(n2932), .SEL(key[98]), .F(n2934) );
  MUX \e/a/U6828  ( .IN0(n1483), .IN1(n2741), .SEL(key[103]), .F(n2933) );
  MUX \e/a/U6827  ( .IN0(n1518), .IN1(n2761), .SEL(key[103]), .F(n2932) );
  MUX \e/a/U6826  ( .IN0(n1474), .IN1(n2930), .SEL(key[98]), .F(n2931) );
  MUX \e/a/U6825  ( .IN0(n1489), .IN1(n2745), .SEL(key[103]), .F(n2930) );
  MUX \e/a/U6824  ( .IN0(n2929), .IN1(n2910), .SEL(key[102]), .F(\e/t[27] ) );
  MUX \e/a/U6823  ( .IN0(n2928), .IN1(n2920), .SEL(key[96]), .F(n2929) );
  MUX \e/a/U6822  ( .IN0(n2927), .IN1(n2924), .SEL(key[101]), .F(n2928) );
  MUX \e/a/U6821  ( .IN0(n2926), .IN1(n2925), .SEL(key[103]), .F(n2927) );
  MUX \e/a/U6820  ( .IN0(n2753), .IN1(n1507), .SEL(key[98]), .F(n2926) );
  MUX \e/a/U6819  ( .IN0(n597), .IN1(n1476), .SEL(key[98]), .F(n2925) );
  MUX \e/a/U6818  ( .IN0(n2922), .IN1(n2921), .SEL(key[103]), .F(n2924) );
  AND \e/a/U6817  ( .A(n2923), .B(key[100]), .Z(n2922) );
  MUX \e/a/U6816  ( .IN0(n1498), .IN1(n2764), .SEL(key[98]), .F(n2921) );
  MUX \e/a/U6815  ( .IN0(n2919), .IN1(n2916), .SEL(key[101]), .F(n2920) );
  MUX \e/a/U6814  ( .IN0(n2918), .IN1(n2917), .SEL(key[103]), .F(n2919) );
  MUX \e/a/U6813  ( .IN0(n2756), .IN1(n593), .SEL(key[98]), .F(n2918) );
  MUX \e/a/U6812  ( .IN0(n1475), .IN1(n1489), .SEL(key[98]), .F(n2917) );
  MUX \e/a/U6811  ( .IN0(n2912), .IN1(n2913), .SEL(key[103]), .F(n2916) );
  NAND \e/a/U6810  ( .A(n2914), .B(n2915), .Z(n2913) );
  MUX \e/a/U6809  ( .IN0(n1508), .IN1(n2911), .SEL(key[98]), .F(n2912) );
  MUX \e/a/U6808  ( .IN0(n1490), .IN1(n1524), .SEL(key[97]), .F(n2911) );
  MUX \e/a/U6807  ( .IN0(n2909), .IN1(n2900), .SEL(key[96]), .F(n2910) );
  MUX \e/a/U6806  ( .IN0(n2908), .IN1(n2904), .SEL(key[101]), .F(n2909) );
  MUX \e/a/U6805  ( .IN0(n2906), .IN1(n2905), .SEL(key[103]), .F(n2908) );
  NAND \e/a/U6804  ( .A(n1482), .B(n2907), .Z(n2906) );
  MUX \e/a/U6803  ( .IN0(n1523), .IN1(n1491), .SEL(key[98]), .F(n2905) );
  MUX \e/a/U6802  ( .IN0(n2903), .IN1(n2901), .SEL(key[103]), .F(n2904) );
  MUX \e/a/U6801  ( .IN0(n2748), .IN1(n2902), .SEL(key[98]), .F(n2903) );
  AND \e/a/U6800  ( .A(key[97]), .B(n1482), .Z(n2902) );
  MUX \e/a/U6799  ( .IN0(n1486), .IN1(n2765), .SEL(key[98]), .F(n2901) );
  MUX \e/a/U6798  ( .IN0(n2899), .IN1(n2893), .SEL(key[101]), .F(n2900) );
  MUX \e/a/U6797  ( .IN0(n2898), .IN1(n2896), .SEL(key[103]), .F(n2899) );
  MUX \e/a/U6796  ( .IN0(n2897), .IN1(n2737), .SEL(n2781), .F(n2898) );
  MUX \e/a/U6795  ( .IN0(key[99]), .IN1(key[100]), .SEL(key[98]), .F(n2897) );
  MUX \e/a/U6794  ( .IN0(n2765), .IN1(n2894), .SEL(key[98]), .F(n2896) );
  NAND \e/a/U6793  ( .A(n2737), .B(n2895), .Z(n2894) );
  MUX \e/a/U6792  ( .IN0(n2890), .IN1(n2891), .SEL(key[103]), .F(n2893) );
  AND \e/a/U6791  ( .A(n1506), .B(n2892), .Z(n2891) );
  MUX \e/a/U6790  ( .IN0(n1492), .IN1(n2738), .SEL(key[98]), .F(n2890) );
  MUX \e/a/U6789  ( .IN0(n2889), .IN1(n2873), .SEL(key[102]), .F(\e/t[26] ) );
  MUX \e/a/U6788  ( .IN0(n2888), .IN1(n2880), .SEL(key[96]), .F(n2889) );
  MUX \e/a/U6787  ( .IN0(n2887), .IN1(n2883), .SEL(key[101]), .F(n2888) );
  MUX \e/a/U6786  ( .IN0(n2886), .IN1(n2884), .SEL(key[98]), .F(n2887) );
  MUX \e/a/U6785  ( .IN0(n1498), .IN1(n2885), .SEL(key[103]), .F(n2886) );
  MUX \e/a/U6784  ( .IN0(n2745), .IN1(n1482), .SEL(key[97]), .F(n2885) );
  MUX \e/a/U6783  ( .IN0(n2780), .IN1(n1512), .SEL(key[103]), .F(n2884) );
  MUX \e/a/U6782  ( .IN0(n2882), .IN1(n2881), .SEL(key[98]), .F(n2883) );
  MUX \e/a/U6781  ( .IN0(n2738), .IN1(n1487), .SEL(key[103]), .F(n2882) );
  MUX \e/a/U6780  ( .IN0(n1515), .IN1(n2768), .SEL(key[103]), .F(n2881) );
  MUX \e/a/U6779  ( .IN0(n2879), .IN1(n2875), .SEL(key[101]), .F(n2880) );
  MUX \e/a/U6778  ( .IN0(n2876), .IN1(n1474), .SEL(key[98]), .F(n2879) );
  NAND \e/a/U6777  ( .A(n2877), .B(n2878), .Z(n2876) );
  MUX \e/a/U6776  ( .IN0(n595), .IN1(n2874), .SEL(n2779), .F(n2875) );
  MUX \e/a/U6775  ( .IN0(n1497), .IN1(n2750), .SEL(key[98]), .F(n2874) );
  MUX \e/a/U6774  ( .IN0(n2872), .IN1(n2864), .SEL(key[96]), .F(n2873) );
  MUX \e/a/U6773  ( .IN0(n2871), .IN1(n2868), .SEL(key[101]), .F(n2872) );
  MUX \e/a/U6772  ( .IN0(n2870), .IN1(n2869), .SEL(key[98]), .F(n2871) );
  MUX \e/a/U6771  ( .IN0(n1521), .IN1(key[97]), .SEL(key[103]), .F(n2870) );
  MUX \e/a/U6770  ( .IN0(n598), .IN1(n2751), .SEL(key[103]), .F(n2869) );
  MUX \e/a/U6769  ( .IN0(n2867), .IN1(n2866), .SEL(key[98]), .F(n2868) );
  MUX \e/a/U6768  ( .IN0(n1526), .IN1(n1520), .SEL(key[103]), .F(n2867) );
  MUX \e/a/U6767  ( .IN0(n598), .IN1(n2865), .SEL(key[103]), .F(n2866) );
  MUX \e/a/U6766  ( .IN0(n1482), .IN1(n1510), .SEL(key[97]), .F(n2865) );
  MUX \e/a/U6765  ( .IN0(n2863), .IN1(n2857), .SEL(key[101]), .F(n2864) );
  MUX \e/a/U6764  ( .IN0(n2860), .IN1(n2859), .SEL(key[98]), .F(n2863) );
  NAND \e/a/U6763  ( .A(n2861), .B(n2862), .Z(n2860) );
  MUX \e/a/U6762  ( .IN0(n2737), .IN1(n2858), .SEL(n596), .F(n2859) );
  MUX \e/a/U6761  ( .IN0(key[99]), .IN1(n1490), .SEL(key[103]), .F(n2858) );
  MUX \e/a/U6760  ( .IN0(n2856), .IN1(n2855), .SEL(key[98]), .F(n2857) );
  MUX \e/a/U6759  ( .IN0(n2778), .IN1(n1488), .SEL(key[103]), .F(n2856) );
  MUX \e/a/U6758  ( .IN0(n2774), .IN1(n2854), .SEL(key[103]), .F(n2855) );
  MUX \e/a/U6757  ( .IN0(n2740), .IN1(n2745), .SEL(key[97]), .F(n2854) );
  MUX \e/a/U6756  ( .IN0(n2853), .IN1(n2835), .SEL(key[102]), .F(\e/t[25] ) );
  MUX \e/a/U6755  ( .IN0(n2852), .IN1(n2843), .SEL(key[96]), .F(n2853) );
  MUX \e/a/U6754  ( .IN0(n2851), .IN1(n2847), .SEL(key[101]), .F(n2852) );
  MUX \e/a/U6753  ( .IN0(n2850), .IN1(n2849), .SEL(key[98]), .F(n2851) );
  MUX \e/a/U6752  ( .IN0(n1517), .IN1(n600), .SEL(key[103]), .F(n2850) );
  MUX \e/a/U6751  ( .IN0(n2848), .IN1(n594), .SEL(key[103]), .F(n2849) );
  NAND \e/a/U6750  ( .A(n1528), .B(n1494), .Z(n2848) );
  MUX \e/a/U6749  ( .IN0(n2846), .IN1(n2845), .SEL(key[98]), .F(n2847) );
  MUX \e/a/U6748  ( .IN0(n1477), .IN1(n2752), .SEL(key[103]), .F(n2846) );
  MUX \e/a/U6747  ( .IN0(n2742), .IN1(n2844), .SEL(key[103]), .F(n2845) );
  AND \e/a/U6746  ( .A(key[97]), .B(key[100]), .Z(n2844) );
  MUX \e/a/U6745  ( .IN0(n2842), .IN1(n2839), .SEL(key[101]), .F(n2843) );
  MUX \e/a/U6744  ( .IN0(n2841), .IN1(n2840), .SEL(key[98]), .F(n2842) );
  MUX \e/a/U6743  ( .IN0(n2777), .IN1(n1526), .SEL(key[103]), .F(n2841) );
  MUX \e/a/U6742  ( .IN0(n1503), .IN1(n2750), .SEL(key[103]), .F(n2840) );
  MUX \e/a/U6741  ( .IN0(n2836), .IN1(n2837), .SEL(key[98]), .F(n2839) );
  AND \e/a/U6740  ( .A(n2838), .B(n2793), .Z(n2837) );
  MUX \e/a/U6739  ( .IN0(n2755), .IN1(n2745), .SEL(key[103]), .F(n2836) );
  MUX \e/a/U6738  ( .IN0(n2834), .IN1(n2826), .SEL(key[96]), .F(n2835) );
  MUX \e/a/U6737  ( .IN0(n2833), .IN1(n2829), .SEL(key[101]), .F(n2834) );
  MUX \e/a/U6736  ( .IN0(n2832), .IN1(n2831), .SEL(key[98]), .F(n2833) );
  MUX \e/a/U6735  ( .IN0(n2744), .IN1(n1496), .SEL(key[103]), .F(n2832) );
  MUX \e/a/U6734  ( .IN0(n2830), .IN1(n1484), .SEL(key[103]), .F(n2831) );
  MUX \e/a/U6733  ( .IN0(n2742), .IN1(n1490), .SEL(key[97]), .F(n2830) );
  MUX \e/a/U6732  ( .IN0(n2828), .IN1(n2827), .SEL(key[98]), .F(n2829) );
  MUX \e/a/U6731  ( .IN0(n1521), .IN1(n1501), .SEL(key[103]), .F(n2828) );
  MUX \e/a/U6730  ( .IN0(n1517), .IN1(n1486), .SEL(key[103]), .F(n2827) );
  MUX \e/a/U6729  ( .IN0(n2825), .IN1(n2820), .SEL(key[101]), .F(n2826) );
  MUX \e/a/U6728  ( .IN0(n2824), .IN1(n2821), .SEL(key[98]), .F(n2825) );
  MUX \e/a/U6727  ( .IN0(n2822), .IN1(n2823), .SEL(key[103]), .F(n2824) );
  NAND \e/a/U6726  ( .A(n2745), .B(n2813), .Z(n2823) );
  MUX \e/a/U6725  ( .IN0(n2745), .IN1(n1490), .SEL(key[97]), .F(n2822) );
  MUX \e/a/U6724  ( .IN0(n2760), .IN1(n2758), .SEL(key[103]), .F(n2821) );
  MUX \e/a/U6723  ( .IN0(n2776), .IN1(n2819), .SEL(key[98]), .F(n2820) );
  MUX \e/a/U6722  ( .IN0(n1494), .IN1(n1520), .SEL(key[103]), .F(n2819) );
  MUX \e/a/U6721  ( .IN0(n2818), .IN1(n2801), .SEL(key[102]), .F(\e/t[24] ) );
  MUX \e/a/U6720  ( .IN0(n2817), .IN1(n2809), .SEL(key[96]), .F(n2818) );
  MUX \e/a/U6719  ( .IN0(n2816), .IN1(n2814), .SEL(key[98]), .F(n2817) );
  MUX \e/a/U6718  ( .IN0(n1475), .IN1(n2815), .SEL(key[103]), .F(n2816) );
  MUX \e/a/U6717  ( .IN0(n1515), .IN1(n1518), .SEL(key[101]), .F(n2815) );
  MUX \e/a/U6716  ( .IN0(n2811), .IN1(n2810), .SEL(key[103]), .F(n2814) );
  NAND \e/a/U6715  ( .A(n2812), .B(n2813), .Z(n2811) );
  MUX \e/a/U6714  ( .IN0(n1514), .IN1(n1528), .SEL(key[101]), .F(n2810) );
  MUX \e/a/U6713  ( .IN0(n2808), .IN1(n2804), .SEL(key[98]), .F(n2809) );
  MUX \e/a/U6712  ( .IN0(n2807), .IN1(n2805), .SEL(key[103]), .F(n2808) );
  MUX \e/a/U6711  ( .IN0(n2806), .IN1(n1478), .SEL(key[101]), .F(n2807) );
  NAND \e/a/U6710  ( .A(n1528), .B(n2737), .Z(n2806) );
  MUX \e/a/U6708  ( .IN0(n2803), .IN1(n2802), .SEL(key[103]), .F(n2804) );
  MUX \e/a/U6707  ( .IN0(n595), .IN1(n1476), .SEL(key[101]), .F(n2803) );
  MUX \e/a/U6706  ( .IN0(n1516), .IN1(n1482), .SEL(key[101]), .F(n2802) );
  MUX \e/a/U6705  ( .IN0(n2800), .IN1(n2790), .SEL(key[96]), .F(n2801) );
  MUX \e/a/U6704  ( .IN0(n2799), .IN1(n2795), .SEL(key[98]), .F(n2800) );
  MUX \e/a/U6703  ( .IN0(n2798), .IN1(n2797), .SEL(key[103]), .F(n2799) );
  MUX \e/a/U6702  ( .IN0(n593), .IN1(n1479), .SEL(key[101]), .F(n2798) );
  MUX \e/a/U6701  ( .IN0(n2796), .IN1(n1506), .SEL(key[101]), .F(n2797) );
  NAND \e/a/U6700  ( .A(n2736), .B(n2738), .Z(n2796) );
  MUX \e/a/U6699  ( .IN0(n2794), .IN1(n2791), .SEL(key[103]), .F(n2795) );
  MUX \e/a/U6698  ( .IN0(n1485), .IN1(n2792), .SEL(key[101]), .F(n2794) );
  NAND \e/a/U6697  ( .A(n2740), .B(n2793), .Z(n2792) );
  MUX \e/a/U6696  ( .IN0(n2754), .IN1(n2746), .SEL(key[101]), .F(n2791) );
  MUX \e/a/U6695  ( .IN0(n2789), .IN1(n2785), .SEL(key[98]), .F(n2790) );
  MUX \e/a/U6694  ( .IN0(n2787), .IN1(n2786), .SEL(key[103]), .F(n2789) );
  NAND \e/a/U6693  ( .A(n2788), .B(n2775), .Z(n2787) );
  MUX \e/a/U6692  ( .IN0(key[99]), .IN1(n2768), .SEL(key[101]), .F(n2786) );
  MUX \e/a/U6691  ( .IN0(n2784), .IN1(n2783), .SEL(key[103]), .F(n2785) );
  MUX \e/a/U6690  ( .IN0(n1488), .IN1(n1499), .SEL(key[101]), .F(n2784) );
  MUX \e/a/U6689  ( .IN0(n1513), .IN1(n1503), .SEL(key[101]), .F(n2783) );
  XOR \e/a/U6688  ( .A(n2737), .B(key[97]), .Z(n2782) );
  XOR \e/a/U6687  ( .A(key[97]), .B(key[98]), .Z(n2781) );
  XOR \e/a/U6686  ( .A(key[97]), .B(key[99]), .Z(n2780) );
  XOR \e/a/U6685  ( .A(key[98]), .B(key[103]), .Z(n2779) );
  XOR \e/a/U6684  ( .A(n1528), .B(n1482), .Z(n2778) );
  XOR \e/a/U6683  ( .A(key[97]), .B(n1518), .Z(n2777) );
  XOR \e/a/U6681  ( .A(key[97]), .B(key[101]), .Z(n2775) );
  NAND \e/a/U6680  ( .A(key[97]), .B(key[99]), .Z(n2774) );
  MUX \e/a/U6679  ( .IN0(n2737), .IN1(n1482), .SEL(key[97]), .F(n2773) );
  MUX \e/a/U6677  ( .IN0(key[99]), .IN1(n1510), .SEL(key[97]), .F(n2772) );
  MUX \e/a/U6676  ( .IN0(n1494), .IN1(n1510), .SEL(key[97]), .F(n2771) );
  MUX \e/a/U6675  ( .IN0(n2740), .IN1(n2742), .SEL(key[97]), .F(n2770) );
  MUX \e/a/U6674  ( .IN0(key[100]), .IN1(n1494), .SEL(key[97]), .F(n2769) );
  OR \e/a/U6673  ( .A(key[97]), .B(key[100]), .Z(n2768) );
  NAND \e/a/U6671  ( .A(n1510), .B(n1528), .Z(n2767) );
  MUX \e/a/U6670  ( .IN0(n1510), .IN1(key[100]), .SEL(key[97]), .F(n2766) );
  MUX \e/a/U6669  ( .IN0(n2736), .IN1(n2745), .SEL(key[97]), .F(n2765) );
  MUX \e/a/U6668  ( .IN0(n1524), .IN1(key[100]), .SEL(key[97]), .F(n2764) );
  MUX \e/a/U6667  ( .IN0(n1490), .IN1(n1510), .SEL(key[97]), .F(n2763) );
  MUX \e/a/U6666  ( .IN0(n2736), .IN1(key[100]), .SEL(key[97]), .F(n2762) );
  MUX \e/a/U6665  ( .IN0(n1501), .IN1(n1494), .SEL(key[97]), .F(n2761) );
  XOR \e/a/U6664  ( .A(n1490), .B(key[97]), .Z(n2760) );
  MUX \e/a/U6663  ( .IN0(n2742), .IN1(n1501), .SEL(key[97]), .F(n2759) );
  NANDN \e/a/U6662  ( .B(key[97]), .A(key[99]), .Z(n2758) );
  MUX \e/a/U6661  ( .IN0(n1482), .IN1(key[99]), .SEL(key[97]), .F(n2757) );
  NAND \e/a/U6659  ( .A(n2740), .B(n1528), .Z(n2756) );
  MUX \e/a/U6658  ( .IN0(key[100]), .IN1(n2737), .SEL(key[97]), .F(n2755) );
  MUX \e/a/U6657  ( .IN0(n1501), .IN1(key[99]), .SEL(key[97]), .F(n2754) );
  MUX \e/a/U6655  ( .IN0(key[100]), .IN1(n1518), .SEL(key[97]), .F(n2753) );
  MUX \e/a/U6654  ( .IN0(n1482), .IN1(n1524), .SEL(key[97]), .F(n2752) );
  NAND \e/a/U6653  ( .A(n2738), .B(n1482), .Z(n2751) );
  MUX \e/a/U6652  ( .IN0(n2737), .IN1(n2745), .SEL(key[97]), .F(n2750) );
  NAND \e/a/U6651  ( .A(n2749), .B(n2736), .Z(n2748) );
  MUX \e/a/U6650  ( .IN0(n2740), .IN1(n1524), .SEL(key[97]), .F(n2747) );
  MUX \e/a/U6649  ( .IN0(n1524), .IN1(n1494), .SEL(key[97]), .F(n2746) );
  NANDN \e/a/U6648  ( .B(key[99]), .A(key[100]), .Z(n2745) );
  MUX \e/a/U6647  ( .IN0(n2740), .IN1(key[99]), .SEL(key[97]), .F(n2744) );
  OR \e/a/U6646  ( .A(key[99]), .B(key[100]), .Z(n2740) );
  MUX \e/a/U6645  ( .IN0(n1482), .IN1(n1494), .SEL(key[97]), .F(n2743) );
  XOR \e/a/U6644  ( .A(n1490), .B(key[99]), .Z(n2742) );
  NANDN \e/a/U6643  ( .B(key[99]), .A(key[97]), .Z(n2741) );
  NAND \e/a/U6642  ( .A(n2740), .B(n2738), .Z(n2739) );
  NAND \e/a/U6641  ( .A(key[97]), .B(n2737), .Z(n2738) );
  NANDN \e/a/U6640  ( .B(key[100]), .A(key[99]), .Z(n2737) );
  NAND \e/a/U6639  ( .A(key[99]), .B(key[100]), .Z(n2736) );
  MUX \e/a/U6638  ( .IN0(key[124]), .IN1(n2389), .SEL(key[121]), .F(n2735) );
  MUX \e/a/U6637  ( .IN0(key[124]), .IN1(n2398), .SEL(key[121]), .F(n2734) );
  MUX \e/a/U6636  ( .IN0(n2390), .IN1(n2393), .SEL(key[121]), .F(n2733) );
  MUX \e/a/U6635  ( .IN0(n2395), .IN1(n1574), .SEL(key[121]), .F(n2732) );
  MUX \e/a/U6633  ( .IN0(n2398), .IN1(n2389), .SEL(key[122]), .F(n2567) );
  MUX \e/a/U6632  ( .IN0(n2391), .IN1(n1584), .SEL(key[122]), .F(n2568) );
  MUX \e/a/U6631  ( .IN0(n1538), .IN1(n1546), .SEL(key[121]), .F(n2531) );
  MUX \e/a/U6630  ( .IN0(n2417), .IN1(n2723), .SEL(key[127]), .F(n2731) );
  MUX \e/a/U6629  ( .IN0(n2393), .IN1(n2389), .SEL(key[121]), .F(n2725) );
  MUX \e/a/U6628  ( .IN0(n1580), .IN1(n2395), .SEL(key[121]), .F(n2730) );
  MUX \e/a/U6627  ( .IN0(key[123]), .IN1(n1574), .SEL(key[121]), .F(n2729) );
  MUX \e/a/U6626  ( .IN0(n2398), .IN1(n1580), .SEL(key[121]), .F(n2728) );
  MUX \e/a/U6625  ( .IN0(key[124]), .IN1(n2395), .SEL(key[121]), .F(n2727) );
  MUX \e/a/U6624  ( .IN0(n1566), .IN1(n1550), .SEL(key[125]), .F(n2441) );
  MUX \e/a/U6623  ( .IN0(n2390), .IN1(n1546), .SEL(key[121]), .F(n2726) );
  NANDN \e/a/U6620  ( .B(n2396), .A(key[127]), .Z(n2706) );
  NAND \e/a/U6619  ( .A(key[127]), .B(n1547), .Z(n2674) );
  NAND \e/a/U6618  ( .A(key[127]), .B(n1556), .Z(n2615) );
  NAND \e/a/U6617  ( .A(key[127]), .B(n2721), .Z(n2648) );
  NAND \e/a/U6616  ( .A(key[127]), .B(n2643), .Z(n2606) );
  NAND \e/a/U6614  ( .A(n1584), .B(n1574), .Z(n2724) );
  NAND \e/a/U6613  ( .A(key[127]), .B(n2722), .Z(n2720) );
  NAND \e/a/U6612  ( .A(n592), .B(key[127]), .Z(n2700) );
  NAND \e/a/U6610  ( .A(key[122]), .B(n2398), .Z(n2560) );
  NAND \e/a/U6609  ( .A(n1574), .B(key[121]), .Z(n2515) );
  NAND \e/a/U6608  ( .A(key[127]), .B(n2725), .Z(n2514) );
  NAND \e/a/U6606  ( .A(n2724), .B(key[127]), .Z(n2530) );
  NAND \e/a/U6605  ( .A(n2548), .B(n2398), .Z(n2723) );
  NANDN \e/a/U6604  ( .B(n1538), .A(n1584), .Z(n2722) );
  NAND \e/a/U6602  ( .A(key[121]), .B(n2398), .Z(n2446) );
  NAND \e/a/U6601  ( .A(n1538), .B(n1584), .Z(n2721) );
  NAND \e/a/U6598  ( .A(key[121]), .B(n2393), .Z(n2548) );
  ANDN \e/a/U6596  ( .A(key[122]), .B(key[121]), .Z(n2576) );
  AND \e/a/U6595  ( .A(n2390), .B(n2720), .Z(n2491) );
  MUX \e/a/U6594  ( .IN0(n2719), .IN1(n2703), .SEL(key[126]), .F(\e/t[23] ) );
  MUX \e/a/U6593  ( .IN0(n2718), .IN1(n2711), .SEL(key[120]), .F(n2719) );
  MUX \e/a/U6592  ( .IN0(n2717), .IN1(n2714), .SEL(key[125]), .F(n2718) );
  MUX \e/a/U6591  ( .IN0(n2716), .IN1(n2715), .SEL(key[122]), .F(n2717) );
  MUX \e/a/U6590  ( .IN0(key[124]), .IN1(n1551), .SEL(key[127]), .F(n2716) );
  MUX \e/a/U6589  ( .IN0(n2391), .IN1(n1553), .SEL(key[127]), .F(n2715) );
  MUX \e/a/U6588  ( .IN0(n2713), .IN1(n2712), .SEL(key[122]), .F(n2714) );
  MUX \e/a/U6587  ( .IN0(n2445), .IN1(n1547), .SEL(key[127]), .F(n2713) );
  MUX \e/a/U6586  ( .IN0(n2401), .IN1(n2410), .SEL(key[127]), .F(n2712) );
  MUX \e/a/U6585  ( .IN0(n2710), .IN1(n2707), .SEL(key[125]), .F(n2711) );
  MUX \e/a/U6584  ( .IN0(n2709), .IN1(n2708), .SEL(key[122]), .F(n2710) );
  MUX \e/a/U6583  ( .IN0(n2422), .IN1(n2400), .SEL(key[127]), .F(n2709) );
  MUX \e/a/U6582  ( .IN0(n1556), .IN1(n2419), .SEL(key[127]), .F(n2708) );
  MUX \e/a/U6581  ( .IN0(n2705), .IN1(n2704), .SEL(key[122]), .F(n2707) );
  AND \e/a/U6580  ( .A(n1549), .B(n2706), .Z(n2705) );
  MUX \e/a/U6579  ( .IN0(n2405), .IN1(n591), .SEL(key[127]), .F(n2704) );
  MUX \e/a/U6578  ( .IN0(n2702), .IN1(n2694), .SEL(key[120]), .F(n2703) );
  MUX \e/a/U6577  ( .IN0(n2701), .IN1(n2697), .SEL(key[125]), .F(n2702) );
  MUX \e/a/U6576  ( .IN0(n2698), .IN1(n2699), .SEL(key[122]), .F(n2701) );
  NAND \e/a/U6575  ( .A(n2515), .B(n2700), .Z(n2699) );
  MUX \e/a/U6574  ( .IN0(n1583), .IN1(n1575), .SEL(key[127]), .F(n2698) );
  MUX \e/a/U6573  ( .IN0(n2696), .IN1(n2695), .SEL(key[122]), .F(n2697) );
  MUX \e/a/U6572  ( .IN0(n2395), .IN1(n2389), .SEL(key[127]), .F(n2696) );
  MUX \e/a/U6571  ( .IN0(n1576), .IN1(n2423), .SEL(key[127]), .F(n2695) );
  MUX \e/a/U6570  ( .IN0(n2693), .IN1(n2690), .SEL(key[125]), .F(n2694) );
  MUX \e/a/U6569  ( .IN0(n2692), .IN1(n2691), .SEL(key[122]), .F(n2693) );
  MUX \e/a/U6568  ( .IN0(n2426), .IN1(n2414), .SEL(key[127]), .F(n2692) );
  MUX \e/a/U6567  ( .IN0(n1539), .IN1(n2398), .SEL(key[127]), .F(n2691) );
  MUX \e/a/U6566  ( .IN0(n2689), .IN1(n2688), .SEL(key[122]), .F(n2690) );
  MUX \e/a/U6565  ( .IN0(n2427), .IN1(n2435), .SEL(key[127]), .F(n2689) );
  MUX \e/a/U6564  ( .IN0(n2421), .IN1(n2687), .SEL(key[127]), .F(n2688) );
  MUX \e/a/U6563  ( .IN0(n1580), .IN1(n1546), .SEL(key[121]), .F(n2687) );
  MUX \e/a/U6562  ( .IN0(n2686), .IN1(n2668), .SEL(key[126]), .F(\e/t[22] ) );
  MUX \e/a/U6561  ( .IN0(n2685), .IN1(n2676), .SEL(key[120]), .F(n2686) );
  MUX \e/a/U6560  ( .IN0(n2684), .IN1(n2679), .SEL(key[125]), .F(n2685) );
  MUX \e/a/U6559  ( .IN0(n2683), .IN1(n2681), .SEL(key[122]), .F(n2684) );
  MUX \e/a/U6558  ( .IN0(n2682), .IN1(n2402), .SEL(key[127]), .F(n2683) );
  MUX \e/a/U6557  ( .IN0(n1580), .IN1(n2389), .SEL(key[121]), .F(n2682) );
  MUX \e/a/U6556  ( .IN0(n2680), .IN1(n1568), .SEL(key[127]), .F(n2681) );
  MUX \e/a/U6555  ( .IN0(n2389), .IN1(n2390), .SEL(key[121]), .F(n2680) );
  MUX \e/a/U6554  ( .IN0(n2678), .IN1(n2677), .SEL(key[122]), .F(n2679) );
  MUX \e/a/U6553  ( .IN0(n590), .IN1(n2466), .SEL(key[127]), .F(n2678) );
  MUX \e/a/U6552  ( .IN0(n2425), .IN1(n2431), .SEL(key[127]), .F(n2677) );
  MUX \e/a/U6551  ( .IN0(n2675), .IN1(n2671), .SEL(key[125]), .F(n2676) );
  MUX \e/a/U6550  ( .IN0(n2673), .IN1(n2672), .SEL(key[122]), .F(n2675) );
  AND \e/a/U6549  ( .A(n1533), .B(n2674), .Z(n2673) );
  MUX \e/a/U6548  ( .IN0(n2501), .IN1(key[123]), .SEL(key[127]), .F(n2672) );
  MUX \e/a/U6547  ( .IN0(n2670), .IN1(n2669), .SEL(key[122]), .F(n2671) );
  MUX \e/a/U6546  ( .IN0(n1565), .IN1(n2393), .SEL(key[127]), .F(n2670) );
  MUX \e/a/U6544  ( .IN0(n2667), .IN1(n2660), .SEL(key[120]), .F(n2668) );
  MUX \e/a/U6543  ( .IN0(n2666), .IN1(n2663), .SEL(key[125]), .F(n2667) );
  MUX \e/a/U6542  ( .IN0(n2665), .IN1(n2664), .SEL(key[122]), .F(n2666) );
  MUX \e/a/U6541  ( .IN0(n1561), .IN1(n2397), .SEL(key[127]), .F(n2665) );
  MUX \e/a/U6540  ( .IN0(n2401), .IN1(n591), .SEL(key[127]), .F(n2664) );
  MUX \e/a/U6539  ( .IN0(n2662), .IN1(n2661), .SEL(key[122]), .F(n2663) );
  MUX \e/a/U6538  ( .IN0(n2415), .IN1(n1536), .SEL(key[127]), .F(n2662) );
  MUX \e/a/U6537  ( .IN0(n1551), .IN1(n1575), .SEL(key[127]), .F(n2661) );
  MUX \e/a/U6536  ( .IN0(n2659), .IN1(n2655), .SEL(key[125]), .F(n2660) );
  MUX \e/a/U6535  ( .IN0(n2658), .IN1(n2657), .SEL(key[122]), .F(n2659) );
  MUX \e/a/U6534  ( .IN0(n2406), .IN1(n1575), .SEL(key[127]), .F(n2658) );
  MUX \e/a/U6533  ( .IN0(n2656), .IN1(n2424), .SEL(key[127]), .F(n2657) );
  NANDN \e/a/U6532  ( .B(key[124]), .A(key[121]), .Z(n2656) );
  MUX \e/a/U6531  ( .IN0(n2654), .IN1(n2652), .SEL(key[122]), .F(n2655) );
  MUX \e/a/U6530  ( .IN0(n1546), .IN1(n2653), .SEL(key[127]), .F(n2654) );
  MUX \e/a/U6529  ( .IN0(n1566), .IN1(n1557), .SEL(key[121]), .F(n2653) );
  MUX \e/a/U6528  ( .IN0(n1537), .IN1(n2402), .SEL(key[127]), .F(n2652) );
  NANDN \e/a/U6527  ( .B(n1538), .A(key[121]), .Z(n2402) );
  MUX \e/a/U6526  ( .IN0(n2651), .IN1(n2630), .SEL(key[126]), .F(\e/t[21] ) );
  MUX \e/a/U6525  ( .IN0(n2650), .IN1(n2640), .SEL(key[120]), .F(n2651) );
  MUX \e/a/U6524  ( .IN0(n2649), .IN1(n2645), .SEL(key[125]), .F(n2650) );
  MUX \e/a/U6523  ( .IN0(n2646), .IN1(n2647), .SEL(key[122]), .F(n2649) );
  AND \e/a/U6522  ( .A(n2418), .B(n2648), .Z(n2647) );
  MUX \e/a/U6521  ( .IN0(n2398), .IN1(n1576), .SEL(key[127]), .F(n2646) );
  MUX \e/a/U6520  ( .IN0(n2644), .IN1(n2642), .SEL(key[122]), .F(n2645) );
  MUX \e/a/U6519  ( .IN0(n1541), .IN1(n2643), .SEL(key[127]), .F(n2644) );
  NAND \e/a/U6518  ( .A(n1557), .B(n1584), .Z(n2643) );
  MUX \e/a/U6517  ( .IN0(n2398), .IN1(n2641), .SEL(key[127]), .F(n2642) );
  NAND \e/a/U6516  ( .A(n2389), .B(n2446), .Z(n2641) );
  MUX \e/a/U6515  ( .IN0(n2639), .IN1(n2635), .SEL(key[125]), .F(n2640) );
  MUX \e/a/U6514  ( .IN0(n2638), .IN1(n2637), .SEL(key[122]), .F(n2639) );
  MUX \e/a/U6513  ( .IN0(n2409), .IN1(n1578), .SEL(key[127]), .F(n2638) );
  MUX \e/a/U6512  ( .IN0(n2431), .IN1(n2636), .SEL(key[127]), .F(n2637) );
  MUX \e/a/U6511  ( .IN0(n1574), .IN1(n1557), .SEL(key[121]), .F(n2636) );
  MUX \e/a/U6510  ( .IN0(n2634), .IN1(n2633), .SEL(key[122]), .F(n2635) );
  MUX \e/a/U6509  ( .IN0(n1572), .IN1(n589), .SEL(key[127]), .F(n2634) );
  MUX \e/a/U6508  ( .IN0(n2632), .IN1(n2631), .SEL(key[127]), .F(n2633) );
  AND \e/a/U6507  ( .A(n2395), .B(n2466), .Z(n2632) );
  MUX \e/a/U6506  ( .IN0(n1550), .IN1(n1538), .SEL(key[121]), .F(n2631) );
  MUX \e/a/U6505  ( .IN0(n2629), .IN1(n2620), .SEL(key[120]), .F(n2630) );
  MUX \e/a/U6504  ( .IN0(n2628), .IN1(n2624), .SEL(key[125]), .F(n2629) );
  MUX \e/a/U6503  ( .IN0(n2627), .IN1(n2625), .SEL(key[122]), .F(n2628) );
  MUX \e/a/U6502  ( .IN0(n2401), .IN1(n2626), .SEL(key[127]), .F(n2627) );
  NAND \e/a/U6501  ( .A(key[121]), .B(n1550), .Z(n2626) );
  MUX \e/a/U6500  ( .IN0(n1538), .IN1(n1581), .SEL(key[127]), .F(n2625) );
  MUX \e/a/U6499  ( .IN0(n2623), .IN1(n2622), .SEL(key[122]), .F(n2624) );
  MUX \e/a/U6498  ( .IN0(n2424), .IN1(n1552), .SEL(key[127]), .F(n2623) );
  MUX \e/a/U6497  ( .IN0(n2621), .IN1(n2390), .SEL(n588), .F(n2622) );
  AND \e/a/U6496  ( .A(key[127]), .B(key[123]), .Z(n2621) );
  MUX \e/a/U6495  ( .IN0(n2619), .IN1(n2616), .SEL(key[125]), .F(n2620) );
  MUX \e/a/U6494  ( .IN0(n2618), .IN1(n2617), .SEL(key[122]), .F(n2619) );
  MUX \e/a/U6493  ( .IN0(n2547), .IN1(n2390), .SEL(key[127]), .F(n2618) );
  MUX \e/a/U6492  ( .IN0(n587), .IN1(n1579), .SEL(key[127]), .F(n2617) );
  MUX \e/a/U6491  ( .IN0(n2614), .IN1(n2613), .SEL(key[122]), .F(n2616) );
  AND \e/a/U6490  ( .A(n2615), .B(n2515), .Z(n2614) );
  MUX \e/a/U6489  ( .IN0(n1540), .IN1(n1574), .SEL(key[127]), .F(n2613) );
  MUX \e/a/U6488  ( .IN0(n2612), .IN1(n2595), .SEL(key[126]), .F(\e/t[20] ) );
  MUX \e/a/U6487  ( .IN0(n2611), .IN1(n2603), .SEL(key[120]), .F(n2612) );
  MUX \e/a/U6486  ( .IN0(n2610), .IN1(n2607), .SEL(key[125]), .F(n2611) );
  MUX \e/a/U6485  ( .IN0(n2609), .IN1(n2608), .SEL(key[122]), .F(n2610) );
  MUX \e/a/U6484  ( .IN0(n1558), .IN1(n1577), .SEL(key[127]), .F(n2609) );
  MUX \e/a/U6483  ( .IN0(n2466), .IN1(n2431), .SEL(key[127]), .F(n2608) );
  NAND \e/a/U6482  ( .A(key[121]), .B(n2389), .Z(n2466) );
  MUX \e/a/U6481  ( .IN0(n2604), .IN1(n2605), .SEL(key[122]), .F(n2607) );
  AND \e/a/U6480  ( .A(n2418), .B(n2606), .Z(n2605) );
  MUX \e/a/U6479  ( .IN0(n2416), .IN1(n1560), .SEL(key[127]), .F(n2604) );
  MUX \e/a/U6478  ( .IN0(n2602), .IN1(n2599), .SEL(key[125]), .F(n2603) );
  MUX \e/a/U6477  ( .IN0(n2601), .IN1(n2600), .SEL(key[122]), .F(n2602) );
  MUX \e/a/U6476  ( .IN0(n1533), .IN1(n1567), .SEL(key[127]), .F(n2601) );
  MUX \e/a/U6475  ( .IN0(n1538), .IN1(n2398), .SEL(key[127]), .F(n2600) );
  MUX \e/a/U6474  ( .IN0(n2598), .IN1(n2596), .SEL(key[122]), .F(n2599) );
  MUX \e/a/U6473  ( .IN0(n2412), .IN1(n2597), .SEL(key[127]), .F(n2598) );
  AND \e/a/U6472  ( .A(n2398), .B(n1584), .Z(n2597) );
  MUX \e/a/U6471  ( .IN0(n1549), .IN1(n1563), .SEL(key[127]), .F(n2596) );
  MUX \e/a/U6470  ( .IN0(n2594), .IN1(n2588), .SEL(key[120]), .F(n2595) );
  MUX \e/a/U6469  ( .IN0(n2593), .IN1(n2591), .SEL(key[125]), .F(n2594) );
  MUX \e/a/U6468  ( .IN0(n2592), .IN1(n2392), .SEL(key[122]), .F(n2593) );
  MUX \e/a/U6467  ( .IN0(n2410), .IN1(n1565), .SEL(key[127]), .F(n2592) );
  MUX \e/a/U6466  ( .IN0(n2590), .IN1(n2589), .SEL(key[122]), .F(n2591) );
  MUX \e/a/U6465  ( .IN0(n586), .IN1(n1558), .SEL(key[127]), .F(n2590) );
  MUX \e/a/U6464  ( .IN0(n2420), .IN1(n2422), .SEL(key[127]), .F(n2589) );
  MUX \e/a/U6463  ( .IN0(n2587), .IN1(n2584), .SEL(key[125]), .F(n2588) );
  MUX \e/a/U6462  ( .IN0(n2586), .IN1(n2585), .SEL(key[122]), .F(n2587) );
  MUX \e/a/U6461  ( .IN0(n1539), .IN1(n2394), .SEL(key[127]), .F(n2586) );
  MUX \e/a/U6460  ( .IN0(n1574), .IN1(n2414), .SEL(key[127]), .F(n2585) );
  MUX \e/a/U6459  ( .IN0(n1530), .IN1(n2583), .SEL(key[122]), .F(n2584) );
  MUX \e/a/U6458  ( .IN0(n1545), .IN1(n2398), .SEL(key[127]), .F(n2583) );
  MUX \e/a/U6457  ( .IN0(n2582), .IN1(n2563), .SEL(key[126]), .F(\e/t[19] ) );
  MUX \e/a/U6456  ( .IN0(n2581), .IN1(n2573), .SEL(key[120]), .F(n2582) );
  MUX \e/a/U6455  ( .IN0(n2580), .IN1(n2577), .SEL(key[125]), .F(n2581) );
  MUX \e/a/U6454  ( .IN0(n2579), .IN1(n2578), .SEL(key[127]), .F(n2580) );
  MUX \e/a/U6453  ( .IN0(n2406), .IN1(n1563), .SEL(key[122]), .F(n2579) );
  MUX \e/a/U6452  ( .IN0(n589), .IN1(n1532), .SEL(key[122]), .F(n2578) );
  MUX \e/a/U6451  ( .IN0(n2575), .IN1(n2574), .SEL(key[127]), .F(n2577) );
  AND \e/a/U6450  ( .A(n2576), .B(key[124]), .Z(n2575) );
  MUX \e/a/U6449  ( .IN0(n1554), .IN1(n2417), .SEL(key[122]), .F(n2574) );
  MUX \e/a/U6448  ( .IN0(n2572), .IN1(n2569), .SEL(key[125]), .F(n2573) );
  MUX \e/a/U6447  ( .IN0(n2571), .IN1(n2570), .SEL(key[127]), .F(n2572) );
  MUX \e/a/U6446  ( .IN0(n2409), .IN1(n585), .SEL(key[122]), .F(n2571) );
  MUX \e/a/U6445  ( .IN0(n1531), .IN1(n1545), .SEL(key[122]), .F(n2570) );
  MUX \e/a/U6444  ( .IN0(n2565), .IN1(n2566), .SEL(key[127]), .F(n2569) );
  NAND \e/a/U6443  ( .A(n2567), .B(n2568), .Z(n2566) );
  MUX \e/a/U6442  ( .IN0(n1564), .IN1(n2564), .SEL(key[122]), .F(n2565) );
  MUX \e/a/U6441  ( .IN0(n1546), .IN1(n1580), .SEL(key[121]), .F(n2564) );
  MUX \e/a/U6440  ( .IN0(n2562), .IN1(n2553), .SEL(key[120]), .F(n2563) );
  MUX \e/a/U6439  ( .IN0(n2561), .IN1(n2557), .SEL(key[125]), .F(n2562) );
  MUX \e/a/U6438  ( .IN0(n2559), .IN1(n2558), .SEL(key[127]), .F(n2561) );
  NAND \e/a/U6437  ( .A(n1538), .B(n2560), .Z(n2559) );
  MUX \e/a/U6436  ( .IN0(n1579), .IN1(n1547), .SEL(key[122]), .F(n2558) );
  MUX \e/a/U6435  ( .IN0(n2556), .IN1(n2554), .SEL(key[127]), .F(n2557) );
  MUX \e/a/U6434  ( .IN0(n2401), .IN1(n2555), .SEL(key[122]), .F(n2556) );
  AND \e/a/U6433  ( .A(key[121]), .B(n1538), .Z(n2555) );
  MUX \e/a/U6432  ( .IN0(n1542), .IN1(n2418), .SEL(key[122]), .F(n2554) );
  MUX \e/a/U6431  ( .IN0(n2552), .IN1(n2546), .SEL(key[125]), .F(n2553) );
  MUX \e/a/U6430  ( .IN0(n2551), .IN1(n2549), .SEL(key[127]), .F(n2552) );
  MUX \e/a/U6429  ( .IN0(n2550), .IN1(n2390), .SEL(n2434), .F(n2551) );
  MUX \e/a/U6428  ( .IN0(key[123]), .IN1(key[124]), .SEL(key[122]), .F(n2550)
         );
  MUX \e/a/U6427  ( .IN0(n2418), .IN1(n2547), .SEL(key[122]), .F(n2549) );
  NAND \e/a/U6426  ( .A(n2390), .B(n2548), .Z(n2547) );
  MUX \e/a/U6425  ( .IN0(n2543), .IN1(n2544), .SEL(key[127]), .F(n2546) );
  AND \e/a/U6424  ( .A(n1562), .B(n2545), .Z(n2544) );
  MUX \e/a/U6423  ( .IN0(n1548), .IN1(n2391), .SEL(key[122]), .F(n2543) );
  MUX \e/a/U6422  ( .IN0(n2542), .IN1(n2526), .SEL(key[126]), .F(\e/t[18] ) );
  MUX \e/a/U6421  ( .IN0(n2541), .IN1(n2533), .SEL(key[120]), .F(n2542) );
  MUX \e/a/U6420  ( .IN0(n2540), .IN1(n2536), .SEL(key[125]), .F(n2541) );
  MUX \e/a/U6419  ( .IN0(n2539), .IN1(n2537), .SEL(key[122]), .F(n2540) );
  MUX \e/a/U6418  ( .IN0(n1554), .IN1(n2538), .SEL(key[127]), .F(n2539) );
  MUX \e/a/U6417  ( .IN0(n2398), .IN1(n1538), .SEL(key[121]), .F(n2538) );
  MUX \e/a/U6416  ( .IN0(n2433), .IN1(n1568), .SEL(key[127]), .F(n2537) );
  MUX \e/a/U6415  ( .IN0(n2535), .IN1(n2534), .SEL(key[122]), .F(n2536) );
  MUX \e/a/U6414  ( .IN0(n2391), .IN1(n1543), .SEL(key[127]), .F(n2535) );
  MUX \e/a/U6413  ( .IN0(n1571), .IN1(n2421), .SEL(key[127]), .F(n2534) );
  MUX \e/a/U6412  ( .IN0(n2532), .IN1(n2528), .SEL(key[125]), .F(n2533) );
  MUX \e/a/U6411  ( .IN0(n2529), .IN1(n1530), .SEL(key[122]), .F(n2532) );
  NAND \e/a/U6410  ( .A(n2530), .B(n2531), .Z(n2529) );
  MUX \e/a/U6409  ( .IN0(n587), .IN1(n2527), .SEL(n2432), .F(n2528) );
  MUX \e/a/U6408  ( .IN0(n1553), .IN1(n2403), .SEL(key[122]), .F(n2527) );
  MUX \e/a/U6407  ( .IN0(n2525), .IN1(n2517), .SEL(key[120]), .F(n2526) );
  MUX \e/a/U6406  ( .IN0(n2524), .IN1(n2521), .SEL(key[125]), .F(n2525) );
  MUX \e/a/U6405  ( .IN0(n2523), .IN1(n2522), .SEL(key[122]), .F(n2524) );
  MUX \e/a/U6404  ( .IN0(n1577), .IN1(key[121]), .SEL(key[127]), .F(n2523) );
  MUX \e/a/U6403  ( .IN0(n590), .IN1(n2404), .SEL(key[127]), .F(n2522) );
  MUX \e/a/U6402  ( .IN0(n2520), .IN1(n2519), .SEL(key[122]), .F(n2521) );
  MUX \e/a/U6401  ( .IN0(n1582), .IN1(n1576), .SEL(key[127]), .F(n2520) );
  MUX \e/a/U6400  ( .IN0(n590), .IN1(n2518), .SEL(key[127]), .F(n2519) );
  MUX \e/a/U6399  ( .IN0(n1538), .IN1(n1566), .SEL(key[121]), .F(n2518) );
  MUX \e/a/U6398  ( .IN0(n2516), .IN1(n2510), .SEL(key[125]), .F(n2517) );
  MUX \e/a/U6397  ( .IN0(n2513), .IN1(n2512), .SEL(key[122]), .F(n2516) );
  NAND \e/a/U6396  ( .A(n2514), .B(n2515), .Z(n2513) );
  MUX \e/a/U6395  ( .IN0(n2390), .IN1(n2511), .SEL(n588), .F(n2512) );
  MUX \e/a/U6394  ( .IN0(key[123]), .IN1(n1546), .SEL(key[127]), .F(n2511) );
  MUX \e/a/U6393  ( .IN0(n2509), .IN1(n2508), .SEL(key[122]), .F(n2510) );
  MUX \e/a/U6392  ( .IN0(n2431), .IN1(n1544), .SEL(key[127]), .F(n2509) );
  MUX \e/a/U6391  ( .IN0(n2427), .IN1(n2507), .SEL(key[127]), .F(n2508) );
  MUX \e/a/U6390  ( .IN0(n2393), .IN1(n2398), .SEL(key[121]), .F(n2507) );
  MUX \e/a/U6389  ( .IN0(n2506), .IN1(n2488), .SEL(key[126]), .F(\e/t[17] ) );
  MUX \e/a/U6388  ( .IN0(n2505), .IN1(n2496), .SEL(key[120]), .F(n2506) );
  MUX \e/a/U6387  ( .IN0(n2504), .IN1(n2500), .SEL(key[125]), .F(n2505) );
  MUX \e/a/U6386  ( .IN0(n2503), .IN1(n2502), .SEL(key[122]), .F(n2504) );
  MUX \e/a/U6385  ( .IN0(n1573), .IN1(n592), .SEL(key[127]), .F(n2503) );
  MUX \e/a/U6384  ( .IN0(n2501), .IN1(n586), .SEL(key[127]), .F(n2502) );
  NAND \e/a/U6383  ( .A(n1584), .B(n1550), .Z(n2501) );
  MUX \e/a/U6382  ( .IN0(n2499), .IN1(n2498), .SEL(key[122]), .F(n2500) );
  MUX \e/a/U6381  ( .IN0(n1533), .IN1(n2405), .SEL(key[127]), .F(n2499) );
  MUX \e/a/U6380  ( .IN0(n2395), .IN1(n2497), .SEL(key[127]), .F(n2498) );
  AND \e/a/U6379  ( .A(key[121]), .B(key[124]), .Z(n2497) );
  MUX \e/a/U6378  ( .IN0(n2495), .IN1(n2492), .SEL(key[125]), .F(n2496) );
  MUX \e/a/U6377  ( .IN0(n2494), .IN1(n2493), .SEL(key[122]), .F(n2495) );
  MUX \e/a/U6376  ( .IN0(n2430), .IN1(n1582), .SEL(key[127]), .F(n2494) );
  MUX \e/a/U6375  ( .IN0(n1559), .IN1(n2403), .SEL(key[127]), .F(n2493) );
  MUX \e/a/U6374  ( .IN0(n2489), .IN1(n2490), .SEL(key[122]), .F(n2492) );
  AND \e/a/U6373  ( .A(n2491), .B(n2446), .Z(n2490) );
  MUX \e/a/U6372  ( .IN0(n2408), .IN1(n2398), .SEL(key[127]), .F(n2489) );
  MUX \e/a/U6371  ( .IN0(n2487), .IN1(n2479), .SEL(key[120]), .F(n2488) );
  MUX \e/a/U6370  ( .IN0(n2486), .IN1(n2482), .SEL(key[125]), .F(n2487) );
  MUX \e/a/U6369  ( .IN0(n2485), .IN1(n2484), .SEL(key[122]), .F(n2486) );
  MUX \e/a/U6368  ( .IN0(n2397), .IN1(n1552), .SEL(key[127]), .F(n2485) );
  MUX \e/a/U6367  ( .IN0(n2483), .IN1(n1540), .SEL(key[127]), .F(n2484) );
  MUX \e/a/U6366  ( .IN0(n2395), .IN1(n1546), .SEL(key[121]), .F(n2483) );
  MUX \e/a/U6365  ( .IN0(n2481), .IN1(n2480), .SEL(key[122]), .F(n2482) );
  MUX \e/a/U6364  ( .IN0(n1577), .IN1(n1557), .SEL(key[127]), .F(n2481) );
  MUX \e/a/U6363  ( .IN0(n1573), .IN1(n1542), .SEL(key[127]), .F(n2480) );
  MUX \e/a/U6362  ( .IN0(n2478), .IN1(n2473), .SEL(key[125]), .F(n2479) );
  MUX \e/a/U6361  ( .IN0(n2477), .IN1(n2474), .SEL(key[122]), .F(n2478) );
  MUX \e/a/U6360  ( .IN0(n2475), .IN1(n2476), .SEL(key[127]), .F(n2477) );
  NAND \e/a/U6359  ( .A(n2398), .B(n2466), .Z(n2476) );
  MUX \e/a/U6358  ( .IN0(n2398), .IN1(n1546), .SEL(key[121]), .F(n2475) );
  MUX \e/a/U6357  ( .IN0(n2413), .IN1(n2411), .SEL(key[127]), .F(n2474) );
  MUX \e/a/U6356  ( .IN0(n2429), .IN1(n2472), .SEL(key[122]), .F(n2473) );
  MUX \e/a/U6355  ( .IN0(n1550), .IN1(n1576), .SEL(key[127]), .F(n2472) );
  MUX \e/a/U6354  ( .IN0(n2471), .IN1(n2454), .SEL(key[126]), .F(\e/t[16] ) );
  MUX \e/a/U6353  ( .IN0(n2470), .IN1(n2462), .SEL(key[120]), .F(n2471) );
  MUX \e/a/U6352  ( .IN0(n2469), .IN1(n2467), .SEL(key[122]), .F(n2470) );
  MUX \e/a/U6351  ( .IN0(n1531), .IN1(n2468), .SEL(key[127]), .F(n2469) );
  MUX \e/a/U6350  ( .IN0(n1571), .IN1(n1574), .SEL(key[125]), .F(n2468) );
  MUX \e/a/U6349  ( .IN0(n2464), .IN1(n2463), .SEL(key[127]), .F(n2467) );
  NAND \e/a/U6348  ( .A(n2465), .B(n2466), .Z(n2464) );
  MUX \e/a/U6347  ( .IN0(n1570), .IN1(n1584), .SEL(key[125]), .F(n2463) );
  MUX \e/a/U6346  ( .IN0(n2461), .IN1(n2457), .SEL(key[122]), .F(n2462) );
  MUX \e/a/U6345  ( .IN0(n2460), .IN1(n2458), .SEL(key[127]), .F(n2461) );
  MUX \e/a/U6344  ( .IN0(n2459), .IN1(n1534), .SEL(key[125]), .F(n2460) );
  NAND \e/a/U6343  ( .A(n1584), .B(n2390), .Z(n2459) );
  MUX \e/a/U6341  ( .IN0(n2456), .IN1(n2455), .SEL(key[127]), .F(n2457) );
  MUX \e/a/U6340  ( .IN0(n587), .IN1(n1532), .SEL(key[125]), .F(n2456) );
  MUX \e/a/U6339  ( .IN0(n1572), .IN1(n1538), .SEL(key[125]), .F(n2455) );
  MUX \e/a/U6338  ( .IN0(n2453), .IN1(n2443), .SEL(key[120]), .F(n2454) );
  MUX \e/a/U6337  ( .IN0(n2452), .IN1(n2448), .SEL(key[122]), .F(n2453) );
  MUX \e/a/U6336  ( .IN0(n2451), .IN1(n2450), .SEL(key[127]), .F(n2452) );
  MUX \e/a/U6335  ( .IN0(n585), .IN1(n1535), .SEL(key[125]), .F(n2451) );
  MUX \e/a/U6334  ( .IN0(n2449), .IN1(n1562), .SEL(key[125]), .F(n2450) );
  NAND \e/a/U6333  ( .A(n2389), .B(n2391), .Z(n2449) );
  MUX \e/a/U6332  ( .IN0(n2447), .IN1(n2444), .SEL(key[127]), .F(n2448) );
  MUX \e/a/U6331  ( .IN0(n1541), .IN1(n2445), .SEL(key[125]), .F(n2447) );
  NAND \e/a/U6330  ( .A(n2393), .B(n2446), .Z(n2445) );
  MUX \e/a/U6329  ( .IN0(n2407), .IN1(n2399), .SEL(key[125]), .F(n2444) );
  MUX \e/a/U6328  ( .IN0(n2442), .IN1(n2438), .SEL(key[122]), .F(n2443) );
  MUX \e/a/U6327  ( .IN0(n2440), .IN1(n2439), .SEL(key[127]), .F(n2442) );
  NAND \e/a/U6326  ( .A(n2441), .B(n2428), .Z(n2440) );
  MUX \e/a/U6325  ( .IN0(key[123]), .IN1(n2421), .SEL(key[125]), .F(n2439) );
  MUX \e/a/U6324  ( .IN0(n2437), .IN1(n2436), .SEL(key[127]), .F(n2438) );
  MUX \e/a/U6323  ( .IN0(n1544), .IN1(n1555), .SEL(key[125]), .F(n2437) );
  MUX \e/a/U6322  ( .IN0(n1569), .IN1(n1559), .SEL(key[125]), .F(n2436) );
  XOR \e/a/U6321  ( .A(n2390), .B(key[121]), .Z(n2435) );
  XOR \e/a/U6320  ( .A(key[121]), .B(key[122]), .Z(n2434) );
  XOR \e/a/U6319  ( .A(key[121]), .B(key[123]), .Z(n2433) );
  XOR \e/a/U6318  ( .A(key[122]), .B(key[127]), .Z(n2432) );
  XOR \e/a/U6317  ( .A(n1584), .B(n1538), .Z(n2431) );
  XOR \e/a/U6316  ( .A(key[121]), .B(n1574), .Z(n2430) );
  XOR \e/a/U6314  ( .A(key[121]), .B(key[125]), .Z(n2428) );
  NAND \e/a/U6313  ( .A(key[121]), .B(key[123]), .Z(n2427) );
  MUX \e/a/U6312  ( .IN0(n2390), .IN1(n1538), .SEL(key[121]), .F(n2426) );
  MUX \e/a/U6310  ( .IN0(key[123]), .IN1(n1566), .SEL(key[121]), .F(n2425) );
  MUX \e/a/U6309  ( .IN0(n1550), .IN1(n1566), .SEL(key[121]), .F(n2424) );
  MUX \e/a/U6308  ( .IN0(n2393), .IN1(n2395), .SEL(key[121]), .F(n2423) );
  MUX \e/a/U6307  ( .IN0(key[124]), .IN1(n1550), .SEL(key[121]), .F(n2422) );
  OR \e/a/U6306  ( .A(key[121]), .B(key[124]), .Z(n2421) );
  NAND \e/a/U6304  ( .A(n1566), .B(n1584), .Z(n2420) );
  MUX \e/a/U6303  ( .IN0(n1566), .IN1(key[124]), .SEL(key[121]), .F(n2419) );
  MUX \e/a/U6302  ( .IN0(n2389), .IN1(n2398), .SEL(key[121]), .F(n2418) );
  MUX \e/a/U6301  ( .IN0(n1580), .IN1(key[124]), .SEL(key[121]), .F(n2417) );
  MUX \e/a/U6300  ( .IN0(n1546), .IN1(n1566), .SEL(key[121]), .F(n2416) );
  MUX \e/a/U6299  ( .IN0(n2389), .IN1(key[124]), .SEL(key[121]), .F(n2415) );
  MUX \e/a/U6298  ( .IN0(n1557), .IN1(n1550), .SEL(key[121]), .F(n2414) );
  XOR \e/a/U6297  ( .A(n1546), .B(key[121]), .Z(n2413) );
  MUX \e/a/U6296  ( .IN0(n2395), .IN1(n1557), .SEL(key[121]), .F(n2412) );
  NANDN \e/a/U6295  ( .B(key[121]), .A(key[123]), .Z(n2411) );
  MUX \e/a/U6294  ( .IN0(n1538), .IN1(key[123]), .SEL(key[121]), .F(n2410) );
  NAND \e/a/U6292  ( .A(n2393), .B(n1584), .Z(n2409) );
  MUX \e/a/U6291  ( .IN0(key[124]), .IN1(n2390), .SEL(key[121]), .F(n2408) );
  MUX \e/a/U6290  ( .IN0(n1557), .IN1(key[123]), .SEL(key[121]), .F(n2407) );
  MUX \e/a/U6288  ( .IN0(key[124]), .IN1(n1574), .SEL(key[121]), .F(n2406) );
  MUX \e/a/U6287  ( .IN0(n1538), .IN1(n1580), .SEL(key[121]), .F(n2405) );
  NAND \e/a/U6286  ( .A(n2391), .B(n1538), .Z(n2404) );
  MUX \e/a/U6285  ( .IN0(n2390), .IN1(n2398), .SEL(key[121]), .F(n2403) );
  NAND \e/a/U6284  ( .A(n2402), .B(n2389), .Z(n2401) );
  MUX \e/a/U6283  ( .IN0(n2393), .IN1(n1580), .SEL(key[121]), .F(n2400) );
  MUX \e/a/U6282  ( .IN0(n1580), .IN1(n1550), .SEL(key[121]), .F(n2399) );
  NANDN \e/a/U6281  ( .B(key[123]), .A(key[124]), .Z(n2398) );
  MUX \e/a/U6280  ( .IN0(n2393), .IN1(key[123]), .SEL(key[121]), .F(n2397) );
  OR \e/a/U6279  ( .A(key[123]), .B(key[124]), .Z(n2393) );
  MUX \e/a/U6278  ( .IN0(n1538), .IN1(n1550), .SEL(key[121]), .F(n2396) );
  XOR \e/a/U6277  ( .A(n1546), .B(key[123]), .Z(n2395) );
  NANDN \e/a/U6276  ( .B(key[123]), .A(key[121]), .Z(n2394) );
  NAND \e/a/U6275  ( .A(n2393), .B(n2391), .Z(n2392) );
  NAND \e/a/U6274  ( .A(key[121]), .B(n2390), .Z(n2391) );
  NANDN \e/a/U6273  ( .B(key[124]), .A(key[123]), .Z(n2390) );
  NAND \e/a/U6272  ( .A(key[123]), .B(key[124]), .Z(n2389) );
  MUX \e/a/U6271  ( .IN0(key[116]), .IN1(n2042), .SEL(key[113]), .F(n2388) );
  MUX \e/a/U6270  ( .IN0(key[116]), .IN1(n2051), .SEL(key[113]), .F(n2387) );
  MUX \e/a/U6269  ( .IN0(n2043), .IN1(n2046), .SEL(key[113]), .F(n2386) );
  MUX \e/a/U6268  ( .IN0(n2048), .IN1(n1630), .SEL(key[113]), .F(n2385) );
  MUX \e/a/U6266  ( .IN0(n2051), .IN1(n2042), .SEL(key[114]), .F(n2220) );
  MUX \e/a/U6265  ( .IN0(n2044), .IN1(n1640), .SEL(key[114]), .F(n2221) );
  MUX \e/a/U6264  ( .IN0(n1594), .IN1(n1602), .SEL(key[113]), .F(n2184) );
  MUX \e/a/U6263  ( .IN0(n2070), .IN1(n2376), .SEL(key[119]), .F(n2384) );
  MUX \e/a/U6262  ( .IN0(n2046), .IN1(n2042), .SEL(key[113]), .F(n2378) );
  MUX \e/a/U6261  ( .IN0(n1636), .IN1(n2048), .SEL(key[113]), .F(n2383) );
  MUX \e/a/U6260  ( .IN0(key[115]), .IN1(n1630), .SEL(key[113]), .F(n2382) );
  MUX \e/a/U6259  ( .IN0(n2051), .IN1(n1636), .SEL(key[113]), .F(n2381) );
  MUX \e/a/U6258  ( .IN0(key[116]), .IN1(n2048), .SEL(key[113]), .F(n2380) );
  MUX \e/a/U6257  ( .IN0(n1622), .IN1(n1606), .SEL(key[117]), .F(n2094) );
  MUX \e/a/U6256  ( .IN0(n2043), .IN1(n1602), .SEL(key[113]), .F(n2379) );
  NANDN \e/a/U6253  ( .B(n2049), .A(key[119]), .Z(n2359) );
  NAND \e/a/U6252  ( .A(key[119]), .B(n1603), .Z(n2327) );
  NAND \e/a/U6251  ( .A(key[119]), .B(n1612), .Z(n2268) );
  NAND \e/a/U6250  ( .A(key[119]), .B(n2374), .Z(n2301) );
  NAND \e/a/U6249  ( .A(key[119]), .B(n2296), .Z(n2259) );
  NAND \e/a/U6247  ( .A(n1640), .B(n1630), .Z(n2377) );
  NAND \e/a/U6246  ( .A(key[119]), .B(n2375), .Z(n2373) );
  NAND \e/a/U6245  ( .A(n584), .B(key[119]), .Z(n2353) );
  NAND \e/a/U6243  ( .A(key[114]), .B(n2051), .Z(n2213) );
  NAND \e/a/U6242  ( .A(n1630), .B(key[113]), .Z(n2168) );
  NAND \e/a/U6241  ( .A(key[119]), .B(n2378), .Z(n2167) );
  NAND \e/a/U6239  ( .A(n2377), .B(key[119]), .Z(n2183) );
  NAND \e/a/U6238  ( .A(n2201), .B(n2051), .Z(n2376) );
  NANDN \e/a/U6237  ( .B(n1594), .A(n1640), .Z(n2375) );
  NAND \e/a/U6235  ( .A(key[113]), .B(n2051), .Z(n2099) );
  NAND \e/a/U6234  ( .A(n1594), .B(n1640), .Z(n2374) );
  NAND \e/a/U6231  ( .A(key[113]), .B(n2046), .Z(n2201) );
  ANDN \e/a/U6229  ( .A(key[114]), .B(key[113]), .Z(n2229) );
  AND \e/a/U6228  ( .A(n2043), .B(n2373), .Z(n2144) );
  MUX \e/a/U6227  ( .IN0(n2372), .IN1(n2356), .SEL(key[118]), .F(\e/t[15] ) );
  MUX \e/a/U6226  ( .IN0(n2371), .IN1(n2364), .SEL(key[112]), .F(n2372) );
  MUX \e/a/U6225  ( .IN0(n2370), .IN1(n2367), .SEL(key[117]), .F(n2371) );
  MUX \e/a/U6224  ( .IN0(n2369), .IN1(n2368), .SEL(key[114]), .F(n2370) );
  MUX \e/a/U6223  ( .IN0(key[116]), .IN1(n1607), .SEL(key[119]), .F(n2369) );
  MUX \e/a/U6222  ( .IN0(n2044), .IN1(n1609), .SEL(key[119]), .F(n2368) );
  MUX \e/a/U6221  ( .IN0(n2366), .IN1(n2365), .SEL(key[114]), .F(n2367) );
  MUX \e/a/U6220  ( .IN0(n2098), .IN1(n1603), .SEL(key[119]), .F(n2366) );
  MUX \e/a/U6219  ( .IN0(n2054), .IN1(n2063), .SEL(key[119]), .F(n2365) );
  MUX \e/a/U6218  ( .IN0(n2363), .IN1(n2360), .SEL(key[117]), .F(n2364) );
  MUX \e/a/U6217  ( .IN0(n2362), .IN1(n2361), .SEL(key[114]), .F(n2363) );
  MUX \e/a/U6216  ( .IN0(n2075), .IN1(n2053), .SEL(key[119]), .F(n2362) );
  MUX \e/a/U6215  ( .IN0(n1612), .IN1(n2072), .SEL(key[119]), .F(n2361) );
  MUX \e/a/U6214  ( .IN0(n2358), .IN1(n2357), .SEL(key[114]), .F(n2360) );
  AND \e/a/U6213  ( .A(n1605), .B(n2359), .Z(n2358) );
  MUX \e/a/U6212  ( .IN0(n2058), .IN1(n583), .SEL(key[119]), .F(n2357) );
  MUX \e/a/U6211  ( .IN0(n2355), .IN1(n2347), .SEL(key[112]), .F(n2356) );
  MUX \e/a/U6210  ( .IN0(n2354), .IN1(n2350), .SEL(key[117]), .F(n2355) );
  MUX \e/a/U6209  ( .IN0(n2351), .IN1(n2352), .SEL(key[114]), .F(n2354) );
  NAND \e/a/U6208  ( .A(n2168), .B(n2353), .Z(n2352) );
  MUX \e/a/U6207  ( .IN0(n1639), .IN1(n1631), .SEL(key[119]), .F(n2351) );
  MUX \e/a/U6206  ( .IN0(n2349), .IN1(n2348), .SEL(key[114]), .F(n2350) );
  MUX \e/a/U6205  ( .IN0(n2048), .IN1(n2042), .SEL(key[119]), .F(n2349) );
  MUX \e/a/U6204  ( .IN0(n1632), .IN1(n2076), .SEL(key[119]), .F(n2348) );
  MUX \e/a/U6203  ( .IN0(n2346), .IN1(n2343), .SEL(key[117]), .F(n2347) );
  MUX \e/a/U6202  ( .IN0(n2345), .IN1(n2344), .SEL(key[114]), .F(n2346) );
  MUX \e/a/U6201  ( .IN0(n2079), .IN1(n2067), .SEL(key[119]), .F(n2345) );
  MUX \e/a/U6200  ( .IN0(n1595), .IN1(n2051), .SEL(key[119]), .F(n2344) );
  MUX \e/a/U6199  ( .IN0(n2342), .IN1(n2341), .SEL(key[114]), .F(n2343) );
  MUX \e/a/U6198  ( .IN0(n2080), .IN1(n2088), .SEL(key[119]), .F(n2342) );
  MUX \e/a/U6197  ( .IN0(n2074), .IN1(n2340), .SEL(key[119]), .F(n2341) );
  MUX \e/a/U6196  ( .IN0(n1636), .IN1(n1602), .SEL(key[113]), .F(n2340) );
  MUX \e/a/U6195  ( .IN0(n2339), .IN1(n2321), .SEL(key[118]), .F(\e/t[14] ) );
  MUX \e/a/U6194  ( .IN0(n2338), .IN1(n2329), .SEL(key[112]), .F(n2339) );
  MUX \e/a/U6193  ( .IN0(n2337), .IN1(n2332), .SEL(key[117]), .F(n2338) );
  MUX \e/a/U6192  ( .IN0(n2336), .IN1(n2334), .SEL(key[114]), .F(n2337) );
  MUX \e/a/U6191  ( .IN0(n2335), .IN1(n2055), .SEL(key[119]), .F(n2336) );
  MUX \e/a/U6190  ( .IN0(n1636), .IN1(n2042), .SEL(key[113]), .F(n2335) );
  MUX \e/a/U6189  ( .IN0(n2333), .IN1(n1624), .SEL(key[119]), .F(n2334) );
  MUX \e/a/U6188  ( .IN0(n2042), .IN1(n2043), .SEL(key[113]), .F(n2333) );
  MUX \e/a/U6187  ( .IN0(n2331), .IN1(n2330), .SEL(key[114]), .F(n2332) );
  MUX \e/a/U6186  ( .IN0(n582), .IN1(n2119), .SEL(key[119]), .F(n2331) );
  MUX \e/a/U6185  ( .IN0(n2078), .IN1(n2084), .SEL(key[119]), .F(n2330) );
  MUX \e/a/U6184  ( .IN0(n2328), .IN1(n2324), .SEL(key[117]), .F(n2329) );
  MUX \e/a/U6183  ( .IN0(n2326), .IN1(n2325), .SEL(key[114]), .F(n2328) );
  AND \e/a/U6182  ( .A(n1589), .B(n2327), .Z(n2326) );
  MUX \e/a/U6181  ( .IN0(n2154), .IN1(key[115]), .SEL(key[119]), .F(n2325) );
  MUX \e/a/U6180  ( .IN0(n2323), .IN1(n2322), .SEL(key[114]), .F(n2324) );
  MUX \e/a/U6179  ( .IN0(n1621), .IN1(n2046), .SEL(key[119]), .F(n2323) );
  MUX \e/a/U6177  ( .IN0(n2320), .IN1(n2313), .SEL(key[112]), .F(n2321) );
  MUX \e/a/U6176  ( .IN0(n2319), .IN1(n2316), .SEL(key[117]), .F(n2320) );
  MUX \e/a/U6175  ( .IN0(n2318), .IN1(n2317), .SEL(key[114]), .F(n2319) );
  MUX \e/a/U6174  ( .IN0(n1617), .IN1(n2050), .SEL(key[119]), .F(n2318) );
  MUX \e/a/U6173  ( .IN0(n2054), .IN1(n583), .SEL(key[119]), .F(n2317) );
  MUX \e/a/U6172  ( .IN0(n2315), .IN1(n2314), .SEL(key[114]), .F(n2316) );
  MUX \e/a/U6171  ( .IN0(n2068), .IN1(n1592), .SEL(key[119]), .F(n2315) );
  MUX \e/a/U6170  ( .IN0(n1607), .IN1(n1631), .SEL(key[119]), .F(n2314) );
  MUX \e/a/U6169  ( .IN0(n2312), .IN1(n2308), .SEL(key[117]), .F(n2313) );
  MUX \e/a/U6168  ( .IN0(n2311), .IN1(n2310), .SEL(key[114]), .F(n2312) );
  MUX \e/a/U6167  ( .IN0(n2059), .IN1(n1631), .SEL(key[119]), .F(n2311) );
  MUX \e/a/U6166  ( .IN0(n2309), .IN1(n2077), .SEL(key[119]), .F(n2310) );
  NANDN \e/a/U6165  ( .B(key[116]), .A(key[113]), .Z(n2309) );
  MUX \e/a/U6164  ( .IN0(n2307), .IN1(n2305), .SEL(key[114]), .F(n2308) );
  MUX \e/a/U6163  ( .IN0(n1602), .IN1(n2306), .SEL(key[119]), .F(n2307) );
  MUX \e/a/U6162  ( .IN0(n1622), .IN1(n1613), .SEL(key[113]), .F(n2306) );
  MUX \e/a/U6161  ( .IN0(n1593), .IN1(n2055), .SEL(key[119]), .F(n2305) );
  NANDN \e/a/U6160  ( .B(n1594), .A(key[113]), .Z(n2055) );
  MUX \e/a/U6159  ( .IN0(n2304), .IN1(n2283), .SEL(key[118]), .F(\e/t[13] ) );
  MUX \e/a/U6158  ( .IN0(n2303), .IN1(n2293), .SEL(key[112]), .F(n2304) );
  MUX \e/a/U6157  ( .IN0(n2302), .IN1(n2298), .SEL(key[117]), .F(n2303) );
  MUX \e/a/U6156  ( .IN0(n2299), .IN1(n2300), .SEL(key[114]), .F(n2302) );
  AND \e/a/U6155  ( .A(n2071), .B(n2301), .Z(n2300) );
  MUX \e/a/U6154  ( .IN0(n2051), .IN1(n1632), .SEL(key[119]), .F(n2299) );
  MUX \e/a/U6153  ( .IN0(n2297), .IN1(n2295), .SEL(key[114]), .F(n2298) );
  MUX \e/a/U6152  ( .IN0(n1597), .IN1(n2296), .SEL(key[119]), .F(n2297) );
  NAND \e/a/U6151  ( .A(n1613), .B(n1640), .Z(n2296) );
  MUX \e/a/U6150  ( .IN0(n2051), .IN1(n2294), .SEL(key[119]), .F(n2295) );
  NAND \e/a/U6149  ( .A(n2042), .B(n2099), .Z(n2294) );
  MUX \e/a/U6148  ( .IN0(n2292), .IN1(n2288), .SEL(key[117]), .F(n2293) );
  MUX \e/a/U6147  ( .IN0(n2291), .IN1(n2290), .SEL(key[114]), .F(n2292) );
  MUX \e/a/U6146  ( .IN0(n2062), .IN1(n1634), .SEL(key[119]), .F(n2291) );
  MUX \e/a/U6145  ( .IN0(n2084), .IN1(n2289), .SEL(key[119]), .F(n2290) );
  MUX \e/a/U6144  ( .IN0(n1630), .IN1(n1613), .SEL(key[113]), .F(n2289) );
  MUX \e/a/U6143  ( .IN0(n2287), .IN1(n2286), .SEL(key[114]), .F(n2288) );
  MUX \e/a/U6142  ( .IN0(n1628), .IN1(n581), .SEL(key[119]), .F(n2287) );
  MUX \e/a/U6141  ( .IN0(n2285), .IN1(n2284), .SEL(key[119]), .F(n2286) );
  AND \e/a/U6140  ( .A(n2048), .B(n2119), .Z(n2285) );
  MUX \e/a/U6139  ( .IN0(n1606), .IN1(n1594), .SEL(key[113]), .F(n2284) );
  MUX \e/a/U6138  ( .IN0(n2282), .IN1(n2273), .SEL(key[112]), .F(n2283) );
  MUX \e/a/U6137  ( .IN0(n2281), .IN1(n2277), .SEL(key[117]), .F(n2282) );
  MUX \e/a/U6136  ( .IN0(n2280), .IN1(n2278), .SEL(key[114]), .F(n2281) );
  MUX \e/a/U6135  ( .IN0(n2054), .IN1(n2279), .SEL(key[119]), .F(n2280) );
  NAND \e/a/U6134  ( .A(key[113]), .B(n1606), .Z(n2279) );
  MUX \e/a/U6133  ( .IN0(n1594), .IN1(n1637), .SEL(key[119]), .F(n2278) );
  MUX \e/a/U6132  ( .IN0(n2276), .IN1(n2275), .SEL(key[114]), .F(n2277) );
  MUX \e/a/U6131  ( .IN0(n2077), .IN1(n1608), .SEL(key[119]), .F(n2276) );
  MUX \e/a/U6130  ( .IN0(n2274), .IN1(n2043), .SEL(n580), .F(n2275) );
  AND \e/a/U6129  ( .A(key[119]), .B(key[115]), .Z(n2274) );
  MUX \e/a/U6128  ( .IN0(n2272), .IN1(n2269), .SEL(key[117]), .F(n2273) );
  MUX \e/a/U6127  ( .IN0(n2271), .IN1(n2270), .SEL(key[114]), .F(n2272) );
  MUX \e/a/U6126  ( .IN0(n2200), .IN1(n2043), .SEL(key[119]), .F(n2271) );
  MUX \e/a/U6125  ( .IN0(n579), .IN1(n1635), .SEL(key[119]), .F(n2270) );
  MUX \e/a/U6124  ( .IN0(n2267), .IN1(n2266), .SEL(key[114]), .F(n2269) );
  AND \e/a/U6123  ( .A(n2268), .B(n2168), .Z(n2267) );
  MUX \e/a/U6122  ( .IN0(n1596), .IN1(n1630), .SEL(key[119]), .F(n2266) );
  MUX \e/a/U6121  ( .IN0(n2265), .IN1(n2248), .SEL(key[118]), .F(\e/t[12] ) );
  MUX \e/a/U6120  ( .IN0(n2264), .IN1(n2256), .SEL(key[112]), .F(n2265) );
  MUX \e/a/U6119  ( .IN0(n2263), .IN1(n2260), .SEL(key[117]), .F(n2264) );
  MUX \e/a/U6118  ( .IN0(n2262), .IN1(n2261), .SEL(key[114]), .F(n2263) );
  MUX \e/a/U6117  ( .IN0(n1614), .IN1(n1633), .SEL(key[119]), .F(n2262) );
  MUX \e/a/U6116  ( .IN0(n2119), .IN1(n2084), .SEL(key[119]), .F(n2261) );
  NAND \e/a/U6115  ( .A(key[113]), .B(n2042), .Z(n2119) );
  MUX \e/a/U6114  ( .IN0(n2257), .IN1(n2258), .SEL(key[114]), .F(n2260) );
  AND \e/a/U6113  ( .A(n2071), .B(n2259), .Z(n2258) );
  MUX \e/a/U6112  ( .IN0(n2069), .IN1(n1616), .SEL(key[119]), .F(n2257) );
  MUX \e/a/U6111  ( .IN0(n2255), .IN1(n2252), .SEL(key[117]), .F(n2256) );
  MUX \e/a/U6110  ( .IN0(n2254), .IN1(n2253), .SEL(key[114]), .F(n2255) );
  MUX \e/a/U6109  ( .IN0(n1589), .IN1(n1623), .SEL(key[119]), .F(n2254) );
  MUX \e/a/U6108  ( .IN0(n1594), .IN1(n2051), .SEL(key[119]), .F(n2253) );
  MUX \e/a/U6107  ( .IN0(n2251), .IN1(n2249), .SEL(key[114]), .F(n2252) );
  MUX \e/a/U6106  ( .IN0(n2065), .IN1(n2250), .SEL(key[119]), .F(n2251) );
  AND \e/a/U6105  ( .A(n2051), .B(n1640), .Z(n2250) );
  MUX \e/a/U6104  ( .IN0(n1605), .IN1(n1619), .SEL(key[119]), .F(n2249) );
  MUX \e/a/U6103  ( .IN0(n2247), .IN1(n2241), .SEL(key[112]), .F(n2248) );
  MUX \e/a/U6102  ( .IN0(n2246), .IN1(n2244), .SEL(key[117]), .F(n2247) );
  MUX \e/a/U6101  ( .IN0(n2245), .IN1(n2045), .SEL(key[114]), .F(n2246) );
  MUX \e/a/U6100  ( .IN0(n2063), .IN1(n1621), .SEL(key[119]), .F(n2245) );
  MUX \e/a/U6099  ( .IN0(n2243), .IN1(n2242), .SEL(key[114]), .F(n2244) );
  MUX \e/a/U6098  ( .IN0(n578), .IN1(n1614), .SEL(key[119]), .F(n2243) );
  MUX \e/a/U6097  ( .IN0(n2073), .IN1(n2075), .SEL(key[119]), .F(n2242) );
  MUX \e/a/U6096  ( .IN0(n2240), .IN1(n2237), .SEL(key[117]), .F(n2241) );
  MUX \e/a/U6095  ( .IN0(n2239), .IN1(n2238), .SEL(key[114]), .F(n2240) );
  MUX \e/a/U6094  ( .IN0(n1595), .IN1(n2047), .SEL(key[119]), .F(n2239) );
  MUX \e/a/U6093  ( .IN0(n1630), .IN1(n2067), .SEL(key[119]), .F(n2238) );
  MUX \e/a/U6092  ( .IN0(n1586), .IN1(n2236), .SEL(key[114]), .F(n2237) );
  MUX \e/a/U6091  ( .IN0(n1601), .IN1(n2051), .SEL(key[119]), .F(n2236) );
  MUX \e/a/U6090  ( .IN0(n2235), .IN1(n2216), .SEL(key[118]), .F(\e/t[11] ) );
  MUX \e/a/U6089  ( .IN0(n2234), .IN1(n2226), .SEL(key[112]), .F(n2235) );
  MUX \e/a/U6088  ( .IN0(n2233), .IN1(n2230), .SEL(key[117]), .F(n2234) );
  MUX \e/a/U6087  ( .IN0(n2232), .IN1(n2231), .SEL(key[119]), .F(n2233) );
  MUX \e/a/U6086  ( .IN0(n2059), .IN1(n1619), .SEL(key[114]), .F(n2232) );
  MUX \e/a/U6085  ( .IN0(n581), .IN1(n1588), .SEL(key[114]), .F(n2231) );
  MUX \e/a/U6084  ( .IN0(n2228), .IN1(n2227), .SEL(key[119]), .F(n2230) );
  AND \e/a/U6083  ( .A(n2229), .B(key[116]), .Z(n2228) );
  MUX \e/a/U6082  ( .IN0(n1610), .IN1(n2070), .SEL(key[114]), .F(n2227) );
  MUX \e/a/U6081  ( .IN0(n2225), .IN1(n2222), .SEL(key[117]), .F(n2226) );
  MUX \e/a/U6080  ( .IN0(n2224), .IN1(n2223), .SEL(key[119]), .F(n2225) );
  MUX \e/a/U6079  ( .IN0(n2062), .IN1(n577), .SEL(key[114]), .F(n2224) );
  MUX \e/a/U6078  ( .IN0(n1587), .IN1(n1601), .SEL(key[114]), .F(n2223) );
  MUX \e/a/U6077  ( .IN0(n2218), .IN1(n2219), .SEL(key[119]), .F(n2222) );
  NAND \e/a/U6076  ( .A(n2220), .B(n2221), .Z(n2219) );
  MUX \e/a/U6075  ( .IN0(n1620), .IN1(n2217), .SEL(key[114]), .F(n2218) );
  MUX \e/a/U6074  ( .IN0(n1602), .IN1(n1636), .SEL(key[113]), .F(n2217) );
  MUX \e/a/U6073  ( .IN0(n2215), .IN1(n2206), .SEL(key[112]), .F(n2216) );
  MUX \e/a/U6072  ( .IN0(n2214), .IN1(n2210), .SEL(key[117]), .F(n2215) );
  MUX \e/a/U6071  ( .IN0(n2212), .IN1(n2211), .SEL(key[119]), .F(n2214) );
  NAND \e/a/U6070  ( .A(n1594), .B(n2213), .Z(n2212) );
  MUX \e/a/U6069  ( .IN0(n1635), .IN1(n1603), .SEL(key[114]), .F(n2211) );
  MUX \e/a/U6068  ( .IN0(n2209), .IN1(n2207), .SEL(key[119]), .F(n2210) );
  MUX \e/a/U6067  ( .IN0(n2054), .IN1(n2208), .SEL(key[114]), .F(n2209) );
  AND \e/a/U6066  ( .A(key[113]), .B(n1594), .Z(n2208) );
  MUX \e/a/U6065  ( .IN0(n1598), .IN1(n2071), .SEL(key[114]), .F(n2207) );
  MUX \e/a/U6064  ( .IN0(n2205), .IN1(n2199), .SEL(key[117]), .F(n2206) );
  MUX \e/a/U6063  ( .IN0(n2204), .IN1(n2202), .SEL(key[119]), .F(n2205) );
  MUX \e/a/U6062  ( .IN0(n2203), .IN1(n2043), .SEL(n2087), .F(n2204) );
  MUX \e/a/U6061  ( .IN0(key[115]), .IN1(key[116]), .SEL(key[114]), .F(n2203)
         );
  MUX \e/a/U6060  ( .IN0(n2071), .IN1(n2200), .SEL(key[114]), .F(n2202) );
  NAND \e/a/U6059  ( .A(n2043), .B(n2201), .Z(n2200) );
  MUX \e/a/U6058  ( .IN0(n2196), .IN1(n2197), .SEL(key[119]), .F(n2199) );
  AND \e/a/U6057  ( .A(n1618), .B(n2198), .Z(n2197) );
  MUX \e/a/U6056  ( .IN0(n1604), .IN1(n2044), .SEL(key[114]), .F(n2196) );
  MUX \e/a/U6055  ( .IN0(n2195), .IN1(n2179), .SEL(key[118]), .F(\e/t[10] ) );
  MUX \e/a/U6054  ( .IN0(n2194), .IN1(n2186), .SEL(key[112]), .F(n2195) );
  MUX \e/a/U6053  ( .IN0(n2193), .IN1(n2189), .SEL(key[117]), .F(n2194) );
  MUX \e/a/U6052  ( .IN0(n2192), .IN1(n2190), .SEL(key[114]), .F(n2193) );
  MUX \e/a/U6051  ( .IN0(n1610), .IN1(n2191), .SEL(key[119]), .F(n2192) );
  MUX \e/a/U6050  ( .IN0(n2051), .IN1(n1594), .SEL(key[113]), .F(n2191) );
  MUX \e/a/U6049  ( .IN0(n2086), .IN1(n1624), .SEL(key[119]), .F(n2190) );
  MUX \e/a/U6048  ( .IN0(n2188), .IN1(n2187), .SEL(key[114]), .F(n2189) );
  MUX \e/a/U6047  ( .IN0(n2044), .IN1(n1599), .SEL(key[119]), .F(n2188) );
  MUX \e/a/U6046  ( .IN0(n1627), .IN1(n2074), .SEL(key[119]), .F(n2187) );
  MUX \e/a/U6045  ( .IN0(n2185), .IN1(n2181), .SEL(key[117]), .F(n2186) );
  MUX \e/a/U6044  ( .IN0(n2182), .IN1(n1586), .SEL(key[114]), .F(n2185) );
  NAND \e/a/U6043  ( .A(n2183), .B(n2184), .Z(n2182) );
  MUX \e/a/U6042  ( .IN0(n579), .IN1(n2180), .SEL(n2085), .F(n2181) );
  MUX \e/a/U6041  ( .IN0(n1609), .IN1(n2056), .SEL(key[114]), .F(n2180) );
  MUX \e/a/U6040  ( .IN0(n2178), .IN1(n2170), .SEL(key[112]), .F(n2179) );
  MUX \e/a/U6039  ( .IN0(n2177), .IN1(n2174), .SEL(key[117]), .F(n2178) );
  MUX \e/a/U6038  ( .IN0(n2176), .IN1(n2175), .SEL(key[114]), .F(n2177) );
  MUX \e/a/U6037  ( .IN0(n1633), .IN1(key[113]), .SEL(key[119]), .F(n2176) );
  MUX \e/a/U6036  ( .IN0(n582), .IN1(n2057), .SEL(key[119]), .F(n2175) );
  MUX \e/a/U6035  ( .IN0(n2173), .IN1(n2172), .SEL(key[114]), .F(n2174) );
  MUX \e/a/U6034  ( .IN0(n1638), .IN1(n1632), .SEL(key[119]), .F(n2173) );
  MUX \e/a/U6033  ( .IN0(n582), .IN1(n2171), .SEL(key[119]), .F(n2172) );
  MUX \e/a/U6032  ( .IN0(n1594), .IN1(n1622), .SEL(key[113]), .F(n2171) );
  MUX \e/a/U6031  ( .IN0(n2169), .IN1(n2163), .SEL(key[117]), .F(n2170) );
  MUX \e/a/U6030  ( .IN0(n2166), .IN1(n2165), .SEL(key[114]), .F(n2169) );
  NAND \e/a/U6029  ( .A(n2167), .B(n2168), .Z(n2166) );
  MUX \e/a/U6028  ( .IN0(n2043), .IN1(n2164), .SEL(n580), .F(n2165) );
  MUX \e/a/U6027  ( .IN0(key[115]), .IN1(n1602), .SEL(key[119]), .F(n2164) );
  MUX \e/a/U6026  ( .IN0(n2162), .IN1(n2161), .SEL(key[114]), .F(n2163) );
  MUX \e/a/U6025  ( .IN0(n2084), .IN1(n1600), .SEL(key[119]), .F(n2162) );
  MUX \e/a/U6024  ( .IN0(n2080), .IN1(n2160), .SEL(key[119]), .F(n2161) );
  MUX \e/a/U6023  ( .IN0(n2046), .IN1(n2051), .SEL(key[113]), .F(n2160) );
  MUX \e/a/U6022  ( .IN0(n2159), .IN1(n2141), .SEL(key[118]), .F(\e/t[9] ) );
  MUX \e/a/U6021  ( .IN0(n2158), .IN1(n2149), .SEL(key[112]), .F(n2159) );
  MUX \e/a/U6020  ( .IN0(n2157), .IN1(n2153), .SEL(key[117]), .F(n2158) );
  MUX \e/a/U6019  ( .IN0(n2156), .IN1(n2155), .SEL(key[114]), .F(n2157) );
  MUX \e/a/U6018  ( .IN0(n1629), .IN1(n584), .SEL(key[119]), .F(n2156) );
  MUX \e/a/U6017  ( .IN0(n2154), .IN1(n578), .SEL(key[119]), .F(n2155) );
  NAND \e/a/U6016  ( .A(n1640), .B(n1606), .Z(n2154) );
  MUX \e/a/U6015  ( .IN0(n2152), .IN1(n2151), .SEL(key[114]), .F(n2153) );
  MUX \e/a/U6014  ( .IN0(n1589), .IN1(n2058), .SEL(key[119]), .F(n2152) );
  MUX \e/a/U6013  ( .IN0(n2048), .IN1(n2150), .SEL(key[119]), .F(n2151) );
  AND \e/a/U6012  ( .A(key[113]), .B(key[116]), .Z(n2150) );
  MUX \e/a/U6011  ( .IN0(n2148), .IN1(n2145), .SEL(key[117]), .F(n2149) );
  MUX \e/a/U6010  ( .IN0(n2147), .IN1(n2146), .SEL(key[114]), .F(n2148) );
  MUX \e/a/U6009  ( .IN0(n2083), .IN1(n1638), .SEL(key[119]), .F(n2147) );
  MUX \e/a/U6008  ( .IN0(n1615), .IN1(n2056), .SEL(key[119]), .F(n2146) );
  MUX \e/a/U6007  ( .IN0(n2142), .IN1(n2143), .SEL(key[114]), .F(n2145) );
  AND \e/a/U6006  ( .A(n2144), .B(n2099), .Z(n2143) );
  MUX \e/a/U6005  ( .IN0(n2061), .IN1(n2051), .SEL(key[119]), .F(n2142) );
  MUX \e/a/U6004  ( .IN0(n2140), .IN1(n2132), .SEL(key[112]), .F(n2141) );
  MUX \e/a/U6003  ( .IN0(n2139), .IN1(n2135), .SEL(key[117]), .F(n2140) );
  MUX \e/a/U6002  ( .IN0(n2138), .IN1(n2137), .SEL(key[114]), .F(n2139) );
  MUX \e/a/U6001  ( .IN0(n2050), .IN1(n1608), .SEL(key[119]), .F(n2138) );
  MUX \e/a/U6000  ( .IN0(n2136), .IN1(n1596), .SEL(key[119]), .F(n2137) );
  MUX \e/a/U5999  ( .IN0(n2048), .IN1(n1602), .SEL(key[113]), .F(n2136) );
  MUX \e/a/U5998  ( .IN0(n2134), .IN1(n2133), .SEL(key[114]), .F(n2135) );
  MUX \e/a/U5997  ( .IN0(n1633), .IN1(n1613), .SEL(key[119]), .F(n2134) );
  MUX \e/a/U5996  ( .IN0(n1629), .IN1(n1598), .SEL(key[119]), .F(n2133) );
  MUX \e/a/U5995  ( .IN0(n2131), .IN1(n2126), .SEL(key[117]), .F(n2132) );
  MUX \e/a/U5994  ( .IN0(n2130), .IN1(n2127), .SEL(key[114]), .F(n2131) );
  MUX \e/a/U5993  ( .IN0(n2128), .IN1(n2129), .SEL(key[119]), .F(n2130) );
  NAND \e/a/U5992  ( .A(n2051), .B(n2119), .Z(n2129) );
  MUX \e/a/U5991  ( .IN0(n2051), .IN1(n1602), .SEL(key[113]), .F(n2128) );
  MUX \e/a/U5990  ( .IN0(n2066), .IN1(n2064), .SEL(key[119]), .F(n2127) );
  MUX \e/a/U5989  ( .IN0(n2082), .IN1(n2125), .SEL(key[114]), .F(n2126) );
  MUX \e/a/U5988  ( .IN0(n1606), .IN1(n1632), .SEL(key[119]), .F(n2125) );
  MUX \e/a/U5987  ( .IN0(n2124), .IN1(n2107), .SEL(key[118]), .F(\e/t[8] ) );
  MUX \e/a/U5986  ( .IN0(n2123), .IN1(n2115), .SEL(key[112]), .F(n2124) );
  MUX \e/a/U5985  ( .IN0(n2122), .IN1(n2120), .SEL(key[114]), .F(n2123) );
  MUX \e/a/U5984  ( .IN0(n1587), .IN1(n2121), .SEL(key[119]), .F(n2122) );
  MUX \e/a/U5983  ( .IN0(n1627), .IN1(n1630), .SEL(key[117]), .F(n2121) );
  MUX \e/a/U5982  ( .IN0(n2117), .IN1(n2116), .SEL(key[119]), .F(n2120) );
  NAND \e/a/U5981  ( .A(n2118), .B(n2119), .Z(n2117) );
  MUX \e/a/U5980  ( .IN0(n1626), .IN1(n1640), .SEL(key[117]), .F(n2116) );
  MUX \e/a/U5979  ( .IN0(n2114), .IN1(n2110), .SEL(key[114]), .F(n2115) );
  MUX \e/a/U5978  ( .IN0(n2113), .IN1(n2111), .SEL(key[119]), .F(n2114) );
  MUX \e/a/U5977  ( .IN0(n2112), .IN1(n1590), .SEL(key[117]), .F(n2113) );
  NAND \e/a/U5976  ( .A(n1640), .B(n2043), .Z(n2112) );
  MUX \e/a/U5974  ( .IN0(n2109), .IN1(n2108), .SEL(key[119]), .F(n2110) );
  MUX \e/a/U5973  ( .IN0(n579), .IN1(n1588), .SEL(key[117]), .F(n2109) );
  MUX \e/a/U5972  ( .IN0(n1628), .IN1(n1594), .SEL(key[117]), .F(n2108) );
  MUX \e/a/U5971  ( .IN0(n2106), .IN1(n2096), .SEL(key[112]), .F(n2107) );
  MUX \e/a/U5970  ( .IN0(n2105), .IN1(n2101), .SEL(key[114]), .F(n2106) );
  MUX \e/a/U5969  ( .IN0(n2104), .IN1(n2103), .SEL(key[119]), .F(n2105) );
  MUX \e/a/U5968  ( .IN0(n577), .IN1(n1591), .SEL(key[117]), .F(n2104) );
  MUX \e/a/U5967  ( .IN0(n2102), .IN1(n1618), .SEL(key[117]), .F(n2103) );
  NAND \e/a/U5966  ( .A(n2042), .B(n2044), .Z(n2102) );
  MUX \e/a/U5965  ( .IN0(n2100), .IN1(n2097), .SEL(key[119]), .F(n2101) );
  MUX \e/a/U5964  ( .IN0(n1597), .IN1(n2098), .SEL(key[117]), .F(n2100) );
  NAND \e/a/U5963  ( .A(n2046), .B(n2099), .Z(n2098) );
  MUX \e/a/U5962  ( .IN0(n2060), .IN1(n2052), .SEL(key[117]), .F(n2097) );
  MUX \e/a/U5961  ( .IN0(n2095), .IN1(n2091), .SEL(key[114]), .F(n2096) );
  MUX \e/a/U5960  ( .IN0(n2093), .IN1(n2092), .SEL(key[119]), .F(n2095) );
  NAND \e/a/U5959  ( .A(n2094), .B(n2081), .Z(n2093) );
  MUX \e/a/U5958  ( .IN0(key[115]), .IN1(n2074), .SEL(key[117]), .F(n2092) );
  MUX \e/a/U5957  ( .IN0(n2090), .IN1(n2089), .SEL(key[119]), .F(n2091) );
  MUX \e/a/U5956  ( .IN0(n1600), .IN1(n1611), .SEL(key[117]), .F(n2090) );
  MUX \e/a/U5955  ( .IN0(n1625), .IN1(n1615), .SEL(key[117]), .F(n2089) );
  XOR \e/a/U5954  ( .A(n2043), .B(key[113]), .Z(n2088) );
  XOR \e/a/U5953  ( .A(key[113]), .B(key[114]), .Z(n2087) );
  XOR \e/a/U5952  ( .A(key[113]), .B(key[115]), .Z(n2086) );
  XOR \e/a/U5951  ( .A(key[114]), .B(key[119]), .Z(n2085) );
  XOR \e/a/U5950  ( .A(n1640), .B(n1594), .Z(n2084) );
  XOR \e/a/U5949  ( .A(key[113]), .B(n1630), .Z(n2083) );
  XOR \e/a/U5947  ( .A(key[113]), .B(key[117]), .Z(n2081) );
  NAND \e/a/U5946  ( .A(key[113]), .B(key[115]), .Z(n2080) );
  MUX \e/a/U5945  ( .IN0(n2043), .IN1(n1594), .SEL(key[113]), .F(n2079) );
  MUX \e/a/U5943  ( .IN0(key[115]), .IN1(n1622), .SEL(key[113]), .F(n2078) );
  MUX \e/a/U5942  ( .IN0(n1606), .IN1(n1622), .SEL(key[113]), .F(n2077) );
  MUX \e/a/U5941  ( .IN0(n2046), .IN1(n2048), .SEL(key[113]), .F(n2076) );
  MUX \e/a/U5940  ( .IN0(key[116]), .IN1(n1606), .SEL(key[113]), .F(n2075) );
  OR \e/a/U5939  ( .A(key[113]), .B(key[116]), .Z(n2074) );
  NAND \e/a/U5937  ( .A(n1622), .B(n1640), .Z(n2073) );
  MUX \e/a/U5936  ( .IN0(n1622), .IN1(key[116]), .SEL(key[113]), .F(n2072) );
  MUX \e/a/U5935  ( .IN0(n2042), .IN1(n2051), .SEL(key[113]), .F(n2071) );
  MUX \e/a/U5934  ( .IN0(n1636), .IN1(key[116]), .SEL(key[113]), .F(n2070) );
  MUX \e/a/U5933  ( .IN0(n1602), .IN1(n1622), .SEL(key[113]), .F(n2069) );
  MUX \e/a/U5932  ( .IN0(n2042), .IN1(key[116]), .SEL(key[113]), .F(n2068) );
  MUX \e/a/U5931  ( .IN0(n1613), .IN1(n1606), .SEL(key[113]), .F(n2067) );
  XOR \e/a/U5930  ( .A(n1602), .B(key[113]), .Z(n2066) );
  MUX \e/a/U5929  ( .IN0(n2048), .IN1(n1613), .SEL(key[113]), .F(n2065) );
  NANDN \e/a/U5928  ( .B(key[113]), .A(key[115]), .Z(n2064) );
  MUX \e/a/U5927  ( .IN0(n1594), .IN1(key[115]), .SEL(key[113]), .F(n2063) );
  NAND \e/a/U5925  ( .A(n2046), .B(n1640), .Z(n2062) );
  MUX \e/a/U5924  ( .IN0(key[116]), .IN1(n2043), .SEL(key[113]), .F(n2061) );
  MUX \e/a/U5923  ( .IN0(n1613), .IN1(key[115]), .SEL(key[113]), .F(n2060) );
  MUX \e/a/U5921  ( .IN0(key[116]), .IN1(n1630), .SEL(key[113]), .F(n2059) );
  MUX \e/a/U5920  ( .IN0(n1594), .IN1(n1636), .SEL(key[113]), .F(n2058) );
  NAND \e/a/U5919  ( .A(n2044), .B(n1594), .Z(n2057) );
  MUX \e/a/U5918  ( .IN0(n2043), .IN1(n2051), .SEL(key[113]), .F(n2056) );
  NAND \e/a/U5917  ( .A(n2055), .B(n2042), .Z(n2054) );
  MUX \e/a/U5916  ( .IN0(n2046), .IN1(n1636), .SEL(key[113]), .F(n2053) );
  MUX \e/a/U5915  ( .IN0(n1636), .IN1(n1606), .SEL(key[113]), .F(n2052) );
  NANDN \e/a/U5914  ( .B(key[115]), .A(key[116]), .Z(n2051) );
  MUX \e/a/U5913  ( .IN0(n2046), .IN1(key[115]), .SEL(key[113]), .F(n2050) );
  OR \e/a/U5912  ( .A(key[115]), .B(key[116]), .Z(n2046) );
  MUX \e/a/U5911  ( .IN0(n1594), .IN1(n1606), .SEL(key[113]), .F(n2049) );
  XOR \e/a/U5910  ( .A(n1602), .B(key[115]), .Z(n2048) );
  NANDN \e/a/U5909  ( .B(key[115]), .A(key[113]), .Z(n2047) );
  NAND \e/a/U5908  ( .A(n2046), .B(n2044), .Z(n2045) );
  NAND \e/a/U5907  ( .A(key[113]), .B(n2043), .Z(n2044) );
  NANDN \e/a/U5906  ( .B(key[116]), .A(key[115]), .Z(n2043) );
  NAND \e/a/U5905  ( .A(key[115]), .B(key[116]), .Z(n2042) );
  MUX \e/a/U5904  ( .IN0(key[108]), .IN1(n1696), .SEL(key[105]), .F(n2041) );
  MUX \e/a/U5903  ( .IN0(key[108]), .IN1(n1697), .SEL(key[105]), .F(n2040) );
  MUX \e/a/U5902  ( .IN0(n1699), .IN1(n1702), .SEL(key[105]), .F(n2039) );
  MUX \e/a/U5901  ( .IN0(n1719), .IN1(n1661), .SEL(key[105]), .F(n2038) );
  MUX \e/a/U5899  ( .IN0(n1697), .IN1(n1696), .SEL(key[106]), .F(n1863) );
  MUX \e/a/U5898  ( .IN0(n1698), .IN1(n1695), .SEL(key[106]), .F(n1864) );
  MUX \e/a/U5897  ( .IN0(n1688), .IN1(n1646), .SEL(key[105]), .F(n1829) );
  MUX \e/a/U5896  ( .IN0(n1726), .IN1(n2029), .SEL(key[111]), .F(n2037) );
  MUX \e/a/U5895  ( .IN0(n1702), .IN1(n1696), .SEL(key[105]), .F(n2031) );
  MUX \e/a/U5894  ( .IN0(n1691), .IN1(n1719), .SEL(key[105]), .F(n2036) );
  MUX \e/a/U5893  ( .IN0(key[107]), .IN1(n1661), .SEL(key[105]), .F(n2035) );
  MUX \e/a/U5892  ( .IN0(n1697), .IN1(n1691), .SEL(key[105]), .F(n2034) );
  MUX \e/a/U5891  ( .IN0(key[108]), .IN1(n1719), .SEL(key[105]), .F(n2033) );
  MUX \e/a/U5890  ( .IN0(n1669), .IN1(n1651), .SEL(key[109]), .F(n1747) );
  MUX \e/a/U5889  ( .IN0(n1699), .IN1(n1646), .SEL(key[105]), .F(n2032) );
  NANDN \e/a/U5886  ( .B(n1704), .A(key[111]), .Z(n2006) );
  NAND \e/a/U5885  ( .A(key[111]), .B(n1648), .Z(n1972) );
  NAND \e/a/U5884  ( .A(key[111]), .B(n1677), .Z(n1924) );
  NAND \e/a/U5883  ( .A(key[111]), .B(n2027), .Z(n1950) );
  NAND \e/a/U5882  ( .A(key[111]), .B(n1952), .Z(n1912) );
  NAND \e/a/U5880  ( .A(n1695), .B(n1661), .Z(n2030) );
  NAND \e/a/U5879  ( .A(key[111]), .B(n2028), .Z(n2026) );
  NAND \e/a/U5878  ( .A(n576), .B(key[111]), .Z(n2012) );
  NAND \e/a/U5876  ( .A(key[106]), .B(n1697), .Z(n1877) );
  NAND \e/a/U5875  ( .A(key[105]), .B(n1661), .Z(n1821) );
  NAND \e/a/U5874  ( .A(key[111]), .B(n2031), .Z(n1820) );
  NAND \e/a/U5873  ( .A(n2030), .B(key[111]), .Z(n1828) );
  NAND \e/a/U5871  ( .A(n1697), .B(n1854), .Z(n2029) );
  NANDN \e/a/U5870  ( .B(n1688), .A(n1695), .Z(n2028) );
  NAND \e/a/U5867  ( .A(key[105]), .B(n1702), .Z(n1854) );
  NAND \e/a/U5866  ( .A(n1697), .B(key[105]), .Z(n1761) );
  NAND \e/a/U5865  ( .A(n1688), .B(n1695), .Z(n2027) );
  ANDN \e/a/U5862  ( .A(key[106]), .B(key[105]), .Z(n1882) );
  AND \e/a/U5861  ( .A(n2026), .B(n1699), .Z(n1788) );
  MUX \e/a/U5860  ( .IN0(n2025), .IN1(n2009), .SEL(key[104]), .F(\e/Q[7] ) );
  MUX \e/a/U5859  ( .IN0(n2024), .IN1(n2017), .SEL(key[110]), .F(n2025) );
  MUX \e/a/U5858  ( .IN0(n2023), .IN1(n2020), .SEL(key[106]), .F(n2024) );
  MUX \e/a/U5857  ( .IN0(n2022), .IN1(n2021), .SEL(key[109]), .F(n2023) );
  MUX \e/a/U5856  ( .IN0(key[108]), .IN1(n1652), .SEL(key[111]), .F(n2022) );
  MUX \e/a/U5855  ( .IN0(n1760), .IN1(n1648), .SEL(key[111]), .F(n2021) );
  MUX \e/a/U5854  ( .IN0(n2019), .IN1(n2018), .SEL(key[109]), .F(n2020) );
  MUX \e/a/U5853  ( .IN0(n1698), .IN1(n1654), .SEL(key[111]), .F(n2019) );
  MUX \e/a/U5852  ( .IN0(n1709), .IN1(n1717), .SEL(key[111]), .F(n2018) );
  MUX \e/a/U5851  ( .IN0(n2016), .IN1(n2013), .SEL(key[106]), .F(n2017) );
  MUX \e/a/U5850  ( .IN0(n2015), .IN1(n2014), .SEL(key[109]), .F(n2016) );
  MUX \e/a/U5849  ( .IN0(n1692), .IN1(n1662), .SEL(key[111]), .F(n2015) );
  MUX \e/a/U5848  ( .IN0(n1719), .IN1(n1696), .SEL(key[111]), .F(n2014) );
  MUX \e/a/U5847  ( .IN0(n2011), .IN1(n2010), .SEL(key[109]), .F(n2013) );
  NAND \e/a/U5846  ( .A(n1821), .B(n2012), .Z(n2011) );
  MUX \e/a/U5845  ( .IN0(n1663), .IN1(n1731), .SEL(key[111]), .F(n2010) );
  MUX \e/a/U5844  ( .IN0(n2008), .IN1(n2000), .SEL(key[110]), .F(n2009) );
  MUX \e/a/U5843  ( .IN0(n2007), .IN1(n2003), .SEL(key[106]), .F(n2008) );
  MUX \e/a/U5842  ( .IN0(n2004), .IN1(n2005), .SEL(key[109]), .F(n2007) );
  AND \e/a/U5841  ( .A(n1650), .B(n2006), .Z(n2005) );
  MUX \e/a/U5840  ( .IN0(n1730), .IN1(n1707), .SEL(key[111]), .F(n2004) );
  MUX \e/a/U5839  ( .IN0(n2002), .IN1(n2001), .SEL(key[109]), .F(n2003) );
  MUX \e/a/U5838  ( .IN0(n1677), .IN1(n1727), .SEL(key[111]), .F(n2002) );
  MUX \e/a/U5837  ( .IN0(n1713), .IN1(n575), .SEL(key[111]), .F(n2001) );
  MUX \e/a/U5836  ( .IN0(n1999), .IN1(n1996), .SEL(key[106]), .F(n2000) );
  MUX \e/a/U5835  ( .IN0(n1998), .IN1(n1997), .SEL(key[109]), .F(n1999) );
  MUX \e/a/U5834  ( .IN0(n1734), .IN1(n1721), .SEL(key[111]), .F(n1998) );
  MUX \e/a/U5833  ( .IN0(n1700), .IN1(n1741), .SEL(key[111]), .F(n1997) );
  MUX \e/a/U5832  ( .IN0(n1995), .IN1(n1994), .SEL(key[109]), .F(n1996) );
  MUX \e/a/U5831  ( .IN0(n1660), .IN1(n1697), .SEL(key[111]), .F(n1995) );
  MUX \e/a/U5830  ( .IN0(n1728), .IN1(n1993), .SEL(key[111]), .F(n1994) );
  MUX \e/a/U5829  ( .IN0(n1691), .IN1(n1646), .SEL(key[105]), .F(n1993) );
  MUX \e/a/U5828  ( .IN0(n1992), .IN1(n1975), .SEL(key[104]), .F(\e/Q[6] ) );
  MUX \e/a/U5827  ( .IN0(n1991), .IN1(n1982), .SEL(key[110]), .F(n1992) );
  MUX \e/a/U5826  ( .IN0(n1990), .IN1(n1986), .SEL(key[106]), .F(n1991) );
  MUX \e/a/U5825  ( .IN0(n1989), .IN1(n1987), .SEL(key[109]), .F(n1990) );
  MUX \e/a/U5824  ( .IN0(n1988), .IN1(n1710), .SEL(key[111]), .F(n1989) );
  MUX \e/a/U5823  ( .IN0(n1691), .IN1(n1696), .SEL(key[105]), .F(n1988) );
  MUX \e/a/U5822  ( .IN0(n574), .IN1(n1772), .SEL(key[111]), .F(n1987) );
  MUX \e/a/U5821  ( .IN0(n1985), .IN1(n1983), .SEL(key[109]), .F(n1986) );
  MUX \e/a/U5820  ( .IN0(n1984), .IN1(n1664), .SEL(key[111]), .F(n1985) );
  MUX \e/a/U5819  ( .IN0(n1696), .IN1(n1699), .SEL(key[105]), .F(n1984) );
  MUX \e/a/U5818  ( .IN0(n1732), .IN1(n1738), .SEL(key[111]), .F(n1983) );
  MUX \e/a/U5817  ( .IN0(n1981), .IN1(n1978), .SEL(key[106]), .F(n1982) );
  MUX \e/a/U5816  ( .IN0(n1980), .IN1(n1979), .SEL(key[109]), .F(n1981) );
  MUX \e/a/U5815  ( .IN0(n1675), .IN1(n1705), .SEL(key[111]), .F(n1980) );
  MUX \e/a/U5814  ( .IN0(n1723), .IN1(n1687), .SEL(key[111]), .F(n1979) );
  MUX \e/a/U5813  ( .IN0(n1977), .IN1(n1976), .SEL(key[109]), .F(n1978) );
  MUX \e/a/U5812  ( .IN0(n1709), .IN1(n575), .SEL(key[111]), .F(n1977) );
  MUX \e/a/U5811  ( .IN0(n1652), .IN1(n1662), .SEL(key[111]), .F(n1976) );
  MUX \e/a/U5810  ( .IN0(n1974), .IN1(n1966), .SEL(key[110]), .F(n1975) );
  MUX \e/a/U5809  ( .IN0(n1973), .IN1(n1969), .SEL(key[106]), .F(n1974) );
  MUX \e/a/U5808  ( .IN0(n1971), .IN1(n1970), .SEL(key[109]), .F(n1973) );
  AND \e/a/U5807  ( .A(n1685), .B(n1972), .Z(n1971) );
  MUX \e/a/U5806  ( .IN0(n1668), .IN1(n1702), .SEL(key[111]), .F(n1970) );
  MUX \e/a/U5805  ( .IN0(n1968), .IN1(n1967), .SEL(key[109]), .F(n1969) );
  MUX \e/a/U5804  ( .IN0(n1805), .IN1(key[107]), .SEL(key[111]), .F(n1968) );
  MUX \e/a/U5802  ( .IN0(n1965), .IN1(n1961), .SEL(key[106]), .F(n1966) );
  MUX \e/a/U5801  ( .IN0(n1964), .IN1(n1963), .SEL(key[109]), .F(n1965) );
  MUX \e/a/U5800  ( .IN0(n1714), .IN1(n1662), .SEL(key[111]), .F(n1964) );
  MUX \e/a/U5799  ( .IN0(n1646), .IN1(n1962), .SEL(key[111]), .F(n1963) );
  MUX \e/a/U5798  ( .IN0(n1669), .IN1(n1678), .SEL(key[105]), .F(n1962) );
  MUX \e/a/U5797  ( .IN0(n1960), .IN1(n1958), .SEL(key[109]), .F(n1961) );
  MUX \e/a/U5796  ( .IN0(n1959), .IN1(n1733), .SEL(key[111]), .F(n1960) );
  NANDN \e/a/U5795  ( .B(key[108]), .A(key[105]), .Z(n1959) );
  MUX \e/a/U5794  ( .IN0(n1644), .IN1(n1710), .SEL(key[111]), .F(n1958) );
  NANDN \e/a/U5793  ( .B(n1688), .A(key[105]), .Z(n1710) );
  MUX \e/a/U5792  ( .IN0(n1957), .IN1(n1937), .SEL(key[104]), .F(\e/Q[5] ) );
  MUX \e/a/U5791  ( .IN0(n1956), .IN1(n1946), .SEL(key[110]), .F(n1957) );
  MUX \e/a/U5790  ( .IN0(n1955), .IN1(n1951), .SEL(key[106]), .F(n1956) );
  MUX \e/a/U5789  ( .IN0(n1954), .IN1(n1953), .SEL(key[109]), .F(n1955) );
  MUX \e/a/U5788  ( .IN0(n1697), .IN1(n1663), .SEL(key[111]), .F(n1954) );
  MUX \e/a/U5787  ( .IN0(n1690), .IN1(n1952), .SEL(key[111]), .F(n1953) );
  NAND \e/a/U5786  ( .A(n1678), .B(n1695), .Z(n1952) );
  MUX \e/a/U5785  ( .IN0(n1949), .IN1(n1948), .SEL(key[109]), .F(n1951) );
  AND \e/a/U5784  ( .A(n1725), .B(n1950), .Z(n1949) );
  MUX \e/a/U5783  ( .IN0(n1697), .IN1(n1947), .SEL(key[111]), .F(n1948) );
  NAND \e/a/U5782  ( .A(n1696), .B(n1761), .Z(n1947) );
  MUX \e/a/U5781  ( .IN0(n1945), .IN1(n1941), .SEL(key[106]), .F(n1946) );
  MUX \e/a/U5780  ( .IN0(n1944), .IN1(n1942), .SEL(key[109]), .F(n1945) );
  MUX \e/a/U5779  ( .IN0(n1709), .IN1(n1943), .SEL(key[111]), .F(n1944) );
  NAND \e/a/U5778  ( .A(key[105]), .B(n1651), .Z(n1943) );
  MUX \e/a/U5777  ( .IN0(n1733), .IN1(n1653), .SEL(key[111]), .F(n1942) );
  MUX \e/a/U5776  ( .IN0(n1940), .IN1(n1939), .SEL(key[109]), .F(n1941) );
  MUX \e/a/U5775  ( .IN0(n1688), .IN1(n1693), .SEL(key[111]), .F(n1940) );
  MUX \e/a/U5774  ( .IN0(n1938), .IN1(n1699), .SEL(n573), .F(n1939) );
  AND \e/a/U5773  ( .A(key[111]), .B(key[107]), .Z(n1938) );
  MUX \e/a/U5772  ( .IN0(n1936), .IN1(n1926), .SEL(key[110]), .F(n1937) );
  MUX \e/a/U5771  ( .IN0(n1935), .IN1(n1932), .SEL(key[106]), .F(n1936) );
  MUX \e/a/U5770  ( .IN0(n1934), .IN1(n1933), .SEL(key[109]), .F(n1935) );
  MUX \e/a/U5769  ( .IN0(n1716), .IN1(n1682), .SEL(key[111]), .F(n1934) );
  MUX \e/a/U5768  ( .IN0(n1658), .IN1(n572), .SEL(key[111]), .F(n1933) );
  MUX \e/a/U5767  ( .IN0(n1931), .IN1(n1929), .SEL(key[109]), .F(n1932) );
  MUX \e/a/U5766  ( .IN0(n1738), .IN1(n1930), .SEL(key[111]), .F(n1931) );
  MUX \e/a/U5765  ( .IN0(n1661), .IN1(n1678), .SEL(key[105]), .F(n1930) );
  MUX \e/a/U5764  ( .IN0(n1928), .IN1(n1927), .SEL(key[111]), .F(n1929) );
  AND \e/a/U5763  ( .A(n1719), .B(n1772), .Z(n1928) );
  MUX \e/a/U5762  ( .IN0(n1651), .IN1(n1688), .SEL(key[105]), .F(n1927) );
  MUX \e/a/U5761  ( .IN0(n1925), .IN1(n1921), .SEL(key[106]), .F(n1926) );
  MUX \e/a/U5760  ( .IN0(n1922), .IN1(n1923), .SEL(key[109]), .F(n1925) );
  AND \e/a/U5759  ( .A(n1924), .B(n1821), .Z(n1923) );
  MUX \e/a/U5758  ( .IN0(n1853), .IN1(n1699), .SEL(key[111]), .F(n1922) );
  MUX \e/a/U5757  ( .IN0(n1920), .IN1(n1919), .SEL(key[109]), .F(n1921) );
  MUX \e/a/U5756  ( .IN0(n571), .IN1(n1683), .SEL(key[111]), .F(n1920) );
  MUX \e/a/U5755  ( .IN0(n1689), .IN1(n1661), .SEL(key[111]), .F(n1919) );
  MUX \e/a/U5754  ( .IN0(n1918), .IN1(n1903), .SEL(key[104]), .F(\e/Q[4] ) );
  MUX \e/a/U5753  ( .IN0(n1917), .IN1(n1909), .SEL(key[110]), .F(n1918) );
  MUX \e/a/U5752  ( .IN0(n1916), .IN1(n1913), .SEL(key[106]), .F(n1917) );
  MUX \e/a/U5751  ( .IN0(n1915), .IN1(n1914), .SEL(key[109]), .F(n1916) );
  MUX \e/a/U5750  ( .IN0(n1670), .IN1(n1665), .SEL(key[111]), .F(n1915) );
  MUX \e/a/U5749  ( .IN0(n1724), .IN1(n1681), .SEL(key[111]), .F(n1914) );
  MUX \e/a/U5748  ( .IN0(n1910), .IN1(n1911), .SEL(key[109]), .F(n1913) );
  AND \e/a/U5747  ( .A(n1725), .B(n1912), .Z(n1911) );
  MUX \e/a/U5746  ( .IN0(n1772), .IN1(n1738), .SEL(key[111]), .F(n1910) );
  NAND \e/a/U5745  ( .A(key[105]), .B(n1696), .Z(n1772) );
  MUX \e/a/U5744  ( .IN0(n1908), .IN1(n1905), .SEL(key[106]), .F(n1909) );
  MUX \e/a/U5743  ( .IN0(n1907), .IN1(n1906), .SEL(key[109]), .F(n1908) );
  MUX \e/a/U5742  ( .IN0(n1717), .IN1(n1668), .SEL(key[111]), .F(n1907) );
  MUX \e/a/U5741  ( .IN0(n570), .IN1(n1670), .SEL(key[111]), .F(n1906) );
  MUX \e/a/U5740  ( .IN0(n1701), .IN1(n1904), .SEL(key[109]), .F(n1905) );
  MUX \e/a/U5739  ( .IN0(n1729), .IN1(n1730), .SEL(key[111]), .F(n1904) );
  MUX \e/a/U5738  ( .IN0(n1902), .IN1(n1894), .SEL(key[110]), .F(n1903) );
  MUX \e/a/U5737  ( .IN0(n1901), .IN1(n1897), .SEL(key[106]), .F(n1902) );
  MUX \e/a/U5736  ( .IN0(n1900), .IN1(n1899), .SEL(key[109]), .F(n1901) );
  MUX \e/a/U5735  ( .IN0(n1685), .IN1(n1671), .SEL(key[111]), .F(n1900) );
  MUX \e/a/U5734  ( .IN0(n1718), .IN1(n1898), .SEL(key[111]), .F(n1899) );
  AND \e/a/U5733  ( .A(n1697), .B(n1695), .Z(n1898) );
  MUX \e/a/U5732  ( .IN0(n1896), .IN1(n1895), .SEL(key[109]), .F(n1897) );
  MUX \e/a/U5731  ( .IN0(n1688), .IN1(n1697), .SEL(key[111]), .F(n1896) );
  MUX \e/a/U5730  ( .IN0(n1650), .IN1(n1666), .SEL(key[111]), .F(n1895) );
  MUX \e/a/U5729  ( .IN0(n1893), .IN1(n1891), .SEL(key[106]), .F(n1894) );
  MUX \e/a/U5728  ( .IN0(n1892), .IN1(n1641), .SEL(key[109]), .F(n1893) );
  MUX \e/a/U5727  ( .IN0(n1660), .IN1(n1703), .SEL(key[111]), .F(n1892) );
  MUX \e/a/U5726  ( .IN0(n1890), .IN1(n1889), .SEL(key[109]), .F(n1891) );
  MUX \e/a/U5725  ( .IN0(n1661), .IN1(n1721), .SEL(key[111]), .F(n1890) );
  MUX \e/a/U5724  ( .IN0(n1645), .IN1(n1697), .SEL(key[111]), .F(n1889) );
  MUX \e/a/U5723  ( .IN0(n1888), .IN1(n1870), .SEL(key[104]), .F(\e/Q[3] ) );
  MUX \e/a/U5722  ( .IN0(n1887), .IN1(n1879), .SEL(key[110]), .F(n1888) );
  MUX \e/a/U5721  ( .IN0(n1886), .IN1(n1883), .SEL(key[109]), .F(n1887) );
  MUX \e/a/U5720  ( .IN0(n1885), .IN1(n1884), .SEL(key[111]), .F(n1886) );
  MUX \e/a/U5719  ( .IN0(n1714), .IN1(n1666), .SEL(key[106]), .F(n1885) );
  MUX \e/a/U5718  ( .IN0(n572), .IN1(n1684), .SEL(key[106]), .F(n1884) );
  MUX \e/a/U5717  ( .IN0(n1881), .IN1(n1880), .SEL(key[111]), .F(n1883) );
  AND \e/a/U5716  ( .A(n1882), .B(key[108]), .Z(n1881) );
  MUX \e/a/U5715  ( .IN0(n1655), .IN1(n1726), .SEL(key[106]), .F(n1880) );
  MUX \e/a/U5714  ( .IN0(n1878), .IN1(n1874), .SEL(key[109]), .F(n1879) );
  MUX \e/a/U5713  ( .IN0(n1876), .IN1(n1875), .SEL(key[111]), .F(n1878) );
  NAND \e/a/U5712  ( .A(n1688), .B(n1877), .Z(n1876) );
  MUX \e/a/U5711  ( .IN0(n1683), .IN1(n1648), .SEL(key[106]), .F(n1875) );
  MUX \e/a/U5710  ( .IN0(n1873), .IN1(n1871), .SEL(key[111]), .F(n1874) );
  MUX \e/a/U5709  ( .IN0(n1709), .IN1(n1872), .SEL(key[106]), .F(n1873) );
  AND \e/a/U5708  ( .A(key[105]), .B(n1688), .Z(n1872) );
  MUX \e/a/U5707  ( .IN0(n1676), .IN1(n1725), .SEL(key[106]), .F(n1871) );
  MUX \e/a/U5706  ( .IN0(n1869), .IN1(n1859), .SEL(key[110]), .F(n1870) );
  MUX \e/a/U5705  ( .IN0(n1868), .IN1(n1865), .SEL(key[109]), .F(n1869) );
  MUX \e/a/U5704  ( .IN0(n1867), .IN1(n1866), .SEL(key[111]), .F(n1868) );
  MUX \e/a/U5703  ( .IN0(n1716), .IN1(n569), .SEL(key[106]), .F(n1867) );
  MUX \e/a/U5702  ( .IN0(n1647), .IN1(n1645), .SEL(key[106]), .F(n1866) );
  MUX \e/a/U5701  ( .IN0(n1861), .IN1(n1862), .SEL(key[111]), .F(n1865) );
  NAND \e/a/U5700  ( .A(n1863), .B(n1864), .Z(n1862) );
  MUX \e/a/U5699  ( .IN0(n1667), .IN1(n1860), .SEL(key[106]), .F(n1861) );
  MUX \e/a/U5698  ( .IN0(n1646), .IN1(n1691), .SEL(key[105]), .F(n1860) );
  MUX \e/a/U5697  ( .IN0(n1858), .IN1(n1852), .SEL(key[109]), .F(n1859) );
  MUX \e/a/U5696  ( .IN0(n1857), .IN1(n1855), .SEL(key[111]), .F(n1858) );
  MUX \e/a/U5695  ( .IN0(n1856), .IN1(n1699), .SEL(n1740), .F(n1857) );
  MUX \e/a/U5694  ( .IN0(key[107]), .IN1(key[108]), .SEL(key[106]), .F(n1856)
         );
  MUX \e/a/U5693  ( .IN0(n1725), .IN1(n1853), .SEL(key[106]), .F(n1855) );
  NAND \e/a/U5692  ( .A(n1699), .B(n1854), .Z(n1853) );
  MUX \e/a/U5691  ( .IN0(n1849), .IN1(n1850), .SEL(key[111]), .F(n1852) );
  AND \e/a/U5690  ( .A(n1657), .B(n1851), .Z(n1850) );
  MUX \e/a/U5689  ( .IN0(n1649), .IN1(n1698), .SEL(key[106]), .F(n1849) );
  MUX \e/a/U5688  ( .IN0(n1848), .IN1(n1832), .SEL(key[104]), .F(\e/Q[2] ) );
  MUX \e/a/U5687  ( .IN0(n1847), .IN1(n1839), .SEL(key[110]), .F(n1848) );
  MUX \e/a/U5686  ( .IN0(n1846), .IN1(n1842), .SEL(key[106]), .F(n1847) );
  MUX \e/a/U5685  ( .IN0(n1845), .IN1(n1843), .SEL(key[109]), .F(n1846) );
  MUX \e/a/U5684  ( .IN0(n1655), .IN1(n1844), .SEL(key[111]), .F(n1845) );
  MUX \e/a/U5683  ( .IN0(n1697), .IN1(n1688), .SEL(key[105]), .F(n1844) );
  MUX \e/a/U5682  ( .IN0(n1698), .IN1(n1642), .SEL(key[111]), .F(n1843) );
  MUX \e/a/U5681  ( .IN0(n1841), .IN1(n1840), .SEL(key[109]), .F(n1842) );
  MUX \e/a/U5680  ( .IN0(n1739), .IN1(n1664), .SEL(key[111]), .F(n1841) );
  MUX \e/a/U5679  ( .IN0(n1674), .IN1(n1728), .SEL(key[111]), .F(n1840) );
  MUX \e/a/U5678  ( .IN0(n1838), .IN1(n1835), .SEL(key[106]), .F(n1839) );
  MUX \e/a/U5677  ( .IN0(n1837), .IN1(n1836), .SEL(key[109]), .F(n1838) );
  MUX \e/a/U5676  ( .IN0(n1665), .IN1(key[105]), .SEL(key[111]), .F(n1837) );
  MUX \e/a/U5675  ( .IN0(n1694), .IN1(n1663), .SEL(key[111]), .F(n1836) );
  MUX \e/a/U5674  ( .IN0(n574), .IN1(n1834), .SEL(key[111]), .F(n1835) );
  MUX \e/a/U5673  ( .IN0(n1712), .IN1(n1833), .SEL(key[109]), .F(n1834) );
  MUX \e/a/U5672  ( .IN0(n1688), .IN1(n1669), .SEL(key[105]), .F(n1833) );
  MUX \e/a/U5671  ( .IN0(n1831), .IN1(n1823), .SEL(key[110]), .F(n1832) );
  MUX \e/a/U5670  ( .IN0(n1830), .IN1(n1825), .SEL(key[106]), .F(n1831) );
  MUX \e/a/U5669  ( .IN0(n1827), .IN1(n1826), .SEL(key[109]), .F(n1830) );
  NAND \e/a/U5668  ( .A(n1828), .B(n1829), .Z(n1827) );
  MUX \e/a/U5667  ( .IN0(n571), .IN1(n1654), .SEL(key[111]), .F(n1826) );
  MUX \e/a/U5666  ( .IN0(n1641), .IN1(n1824), .SEL(key[109]), .F(n1825) );
  MUX \e/a/U5665  ( .IN0(n1711), .IN1(n571), .SEL(key[111]), .F(n1824) );
  MUX \e/a/U5664  ( .IN0(n1822), .IN1(n1817), .SEL(key[106]), .F(n1823) );
  MUX \e/a/U5663  ( .IN0(n1819), .IN1(n1818), .SEL(key[109]), .F(n1822) );
  NAND \e/a/U5662  ( .A(n1820), .B(n1821), .Z(n1819) );
  MUX \e/a/U5661  ( .IN0(n1738), .IN1(n1643), .SEL(key[111]), .F(n1818) );
  MUX \e/a/U5660  ( .IN0(n1816), .IN1(n1814), .SEL(key[109]), .F(n1817) );
  MUX \e/a/U5659  ( .IN0(n1699), .IN1(n1815), .SEL(n573), .F(n1816) );
  MUX \e/a/U5658  ( .IN0(key[107]), .IN1(n1646), .SEL(key[111]), .F(n1815) );
  MUX \e/a/U5657  ( .IN0(n1700), .IN1(n1813), .SEL(key[111]), .F(n1814) );
  MUX \e/a/U5656  ( .IN0(n1702), .IN1(n1697), .SEL(key[105]), .F(n1813) );
  MUX \e/a/U5655  ( .IN0(n1812), .IN1(n1794), .SEL(key[104]), .F(\e/Q[1] ) );
  MUX \e/a/U5654  ( .IN0(n1811), .IN1(n1802), .SEL(key[110]), .F(n1812) );
  MUX \e/a/U5653  ( .IN0(n1810), .IN1(n1807), .SEL(key[106]), .F(n1811) );
  MUX \e/a/U5652  ( .IN0(n1809), .IN1(n1808), .SEL(key[109]), .F(n1810) );
  MUX \e/a/U5651  ( .IN0(n1659), .IN1(n576), .SEL(key[111]), .F(n1809) );
  MUX \e/a/U5650  ( .IN0(n1685), .IN1(n1713), .SEL(key[111]), .F(n1808) );
  MUX \e/a/U5649  ( .IN0(n1806), .IN1(n1804), .SEL(key[109]), .F(n1807) );
  MUX \e/a/U5648  ( .IN0(n1805), .IN1(n570), .SEL(key[111]), .F(n1806) );
  NAND \e/a/U5647  ( .A(n1695), .B(n1651), .Z(n1805) );
  MUX \e/a/U5646  ( .IN0(n1719), .IN1(n1803), .SEL(key[111]), .F(n1804) );
  AND \e/a/U5645  ( .A(key[105]), .B(key[108]), .Z(n1803) );
  MUX \e/a/U5644  ( .IN0(n1801), .IN1(n1798), .SEL(key[106]), .F(n1802) );
  MUX \e/a/U5643  ( .IN0(n1800), .IN1(n1799), .SEL(key[109]), .F(n1801) );
  MUX \e/a/U5642  ( .IN0(n1705), .IN1(n1653), .SEL(key[111]), .F(n1800) );
  MUX \e/a/U5641  ( .IN0(n1665), .IN1(n1678), .SEL(key[111]), .F(n1799) );
  MUX \e/a/U5640  ( .IN0(n1797), .IN1(n1795), .SEL(key[109]), .F(n1798) );
  MUX \e/a/U5639  ( .IN0(n1796), .IN1(n1689), .SEL(key[111]), .F(n1797) );
  MUX \e/a/U5638  ( .IN0(n1719), .IN1(n1646), .SEL(key[105]), .F(n1796) );
  MUX \e/a/U5637  ( .IN0(n1659), .IN1(n1676), .SEL(key[111]), .F(n1795) );
  MUX \e/a/U5636  ( .IN0(n1793), .IN1(n1785), .SEL(key[110]), .F(n1794) );
  MUX \e/a/U5635  ( .IN0(n1792), .IN1(n1789), .SEL(key[106]), .F(n1793) );
  MUX \e/a/U5634  ( .IN0(n1791), .IN1(n1790), .SEL(key[109]), .F(n1792) );
  MUX \e/a/U5633  ( .IN0(n1737), .IN1(n1694), .SEL(key[111]), .F(n1791) );
  MUX \e/a/U5632  ( .IN0(n1715), .IN1(n1697), .SEL(key[111]), .F(n1790) );
  MUX \e/a/U5631  ( .IN0(n1786), .IN1(n1787), .SEL(key[109]), .F(n1789) );
  AND \e/a/U5630  ( .A(n1788), .B(n1761), .Z(n1787) );
  MUX \e/a/U5629  ( .IN0(n1679), .IN1(n1711), .SEL(key[111]), .F(n1786) );
  MUX \e/a/U5628  ( .IN0(n1784), .IN1(n1780), .SEL(key[106]), .F(n1785) );
  MUX \e/a/U5627  ( .IN0(n1783), .IN1(n1736), .SEL(key[109]), .F(n1784) );
  MUX \e/a/U5626  ( .IN0(n1781), .IN1(n1782), .SEL(key[111]), .F(n1783) );
  NAND \e/a/U5625  ( .A(n1697), .B(n1772), .Z(n1782) );
  MUX \e/a/U5624  ( .IN0(n1697), .IN1(n1646), .SEL(key[105]), .F(n1781) );
  MUX \e/a/U5623  ( .IN0(n1779), .IN1(n1778), .SEL(key[109]), .F(n1780) );
  MUX \e/a/U5622  ( .IN0(n1722), .IN1(n1720), .SEL(key[111]), .F(n1779) );
  MUX \e/a/U5621  ( .IN0(n1651), .IN1(n1663), .SEL(key[111]), .F(n1778) );
  MUX \e/a/U5620  ( .IN0(n1777), .IN1(n1758), .SEL(key[104]), .F(\e/Q[0] ) );
  MUX \e/a/U5619  ( .IN0(n1776), .IN1(n1768), .SEL(key[110]), .F(n1777) );
  MUX \e/a/U5618  ( .IN0(n1775), .IN1(n1773), .SEL(key[106]), .F(n1776) );
  MUX \e/a/U5617  ( .IN0(n1647), .IN1(n1774), .SEL(key[111]), .F(n1775) );
  MUX \e/a/U5616  ( .IN0(n1674), .IN1(n1661), .SEL(key[109]), .F(n1774) );
  MUX \e/a/U5615  ( .IN0(n1770), .IN1(n1769), .SEL(key[111]), .F(n1773) );
  NAND \e/a/U5614  ( .A(n1771), .B(n1772), .Z(n1770) );
  MUX \e/a/U5613  ( .IN0(n1673), .IN1(n1695), .SEL(key[109]), .F(n1769) );
  MUX \e/a/U5612  ( .IN0(n1767), .IN1(n1763), .SEL(key[106]), .F(n1768) );
  MUX \e/a/U5611  ( .IN0(n1766), .IN1(n1765), .SEL(key[111]), .F(n1767) );
  MUX \e/a/U5610  ( .IN0(n569), .IN1(n1686), .SEL(key[109]), .F(n1766) );
  MUX \e/a/U5609  ( .IN0(n1764), .IN1(n1657), .SEL(key[109]), .F(n1765) );
  NAND \e/a/U5608  ( .A(n1696), .B(n1698), .Z(n1764) );
  MUX \e/a/U5607  ( .IN0(n1762), .IN1(n1759), .SEL(key[111]), .F(n1763) );
  MUX \e/a/U5606  ( .IN0(n1690), .IN1(n1760), .SEL(key[109]), .F(n1762) );
  NAND \e/a/U5605  ( .A(n1702), .B(n1761), .Z(n1760) );
  MUX \e/a/U5604  ( .IN0(n1680), .IN1(n1706), .SEL(key[109]), .F(n1759) );
  MUX \e/a/U5603  ( .IN0(n1757), .IN1(n1749), .SEL(key[110]), .F(n1758) );
  MUX \e/a/U5602  ( .IN0(n1756), .IN1(n1752), .SEL(key[106]), .F(n1757) );
  MUX \e/a/U5601  ( .IN0(n1755), .IN1(n1753), .SEL(key[111]), .F(n1756) );
  MUX \e/a/U5600  ( .IN0(n1754), .IN1(n1656), .SEL(key[109]), .F(n1755) );
  NAND \e/a/U5599  ( .A(n1695), .B(n1699), .Z(n1754) );
  MUX \e/a/U5597  ( .IN0(n1751), .IN1(n1750), .SEL(key[111]), .F(n1752) );
  MUX \e/a/U5596  ( .IN0(n571), .IN1(n1684), .SEL(key[109]), .F(n1751) );
  MUX \e/a/U5595  ( .IN0(n1658), .IN1(n1688), .SEL(key[109]), .F(n1750) );
  MUX \e/a/U5594  ( .IN0(n1748), .IN1(n1744), .SEL(key[106]), .F(n1749) );
  MUX \e/a/U5593  ( .IN0(n1746), .IN1(n1745), .SEL(key[111]), .F(n1748) );
  NAND \e/a/U5592  ( .A(n1747), .B(n1735), .Z(n1746) );
  MUX \e/a/U5591  ( .IN0(key[107]), .IN1(n1728), .SEL(key[109]), .F(n1745) );
  MUX \e/a/U5590  ( .IN0(n1743), .IN1(n1742), .SEL(key[111]), .F(n1744) );
  MUX \e/a/U5589  ( .IN0(n1643), .IN1(n1708), .SEL(key[109]), .F(n1743) );
  MUX \e/a/U5588  ( .IN0(n1672), .IN1(n1679), .SEL(key[109]), .F(n1742) );
  XOR \e/a/U5587  ( .A(n1699), .B(key[105]), .Z(n1741) );
  XOR \e/a/U5586  ( .A(key[105]), .B(key[106]), .Z(n1740) );
  XOR \e/a/U5585  ( .A(key[105]), .B(key[107]), .Z(n1739) );
  XOR \e/a/U5584  ( .A(n1695), .B(n1688), .Z(n1738) );
  XOR \e/a/U5583  ( .A(key[105]), .B(n1661), .Z(n1737) );
  XOR \e/a/U5581  ( .A(n1691), .B(key[108]), .Z(n1719) );
  XOR \e/a/U5580  ( .A(key[109]), .B(key[105]), .Z(n1735) );
  MUX \e/a/U5579  ( .IN0(n1699), .IN1(n1688), .SEL(key[105]), .F(n1734) );
  MUX \e/a/U5577  ( .IN0(n1651), .IN1(n1669), .SEL(key[105]), .F(n1733) );
  MUX \e/a/U5576  ( .IN0(key[107]), .IN1(n1669), .SEL(key[105]), .F(n1732) );
  MUX \e/a/U5575  ( .IN0(n1702), .IN1(n1719), .SEL(key[105]), .F(n1731) );
  MUX \e/a/U5574  ( .IN0(key[108]), .IN1(n1651), .SEL(key[105]), .F(n1730) );
  NAND \e/a/U5573  ( .A(n1669), .B(n1695), .Z(n1729) );
  OR \e/a/U5572  ( .A(key[108]), .B(key[105]), .Z(n1728) );
  MUX \e/a/U5570  ( .IN0(n1669), .IN1(key[108]), .SEL(key[105]), .F(n1727) );
  MUX \e/a/U5569  ( .IN0(n1691), .IN1(key[108]), .SEL(key[105]), .F(n1726) );
  MUX \e/a/U5568  ( .IN0(n1696), .IN1(n1697), .SEL(key[105]), .F(n1725) );
  MUX \e/a/U5567  ( .IN0(n1646), .IN1(n1669), .SEL(key[105]), .F(n1724) );
  MUX \e/a/U5566  ( .IN0(n1696), .IN1(key[108]), .SEL(key[105]), .F(n1723) );
  XOR \e/a/U5565  ( .A(n1695), .B(key[108]), .Z(n1722) );
  MUX \e/a/U5564  ( .IN0(n1678), .IN1(n1651), .SEL(key[105]), .F(n1721) );
  NANDN \e/a/U5563  ( .B(key[105]), .A(key[107]), .Z(n1720) );
  MUX \e/a/U5562  ( .IN0(n1719), .IN1(n1678), .SEL(key[105]), .F(n1718) );
  MUX \e/a/U5561  ( .IN0(n1688), .IN1(key[107]), .SEL(key[105]), .F(n1717) );
  NAND \e/a/U5559  ( .A(n1702), .B(n1695), .Z(n1716) );
  MUX \e/a/U5558  ( .IN0(key[108]), .IN1(n1699), .SEL(key[105]), .F(n1715) );
  MUX \e/a/U5557  ( .IN0(key[108]), .IN1(n1661), .SEL(key[105]), .F(n1714) );
  MUX \e/a/U5556  ( .IN0(n1688), .IN1(n1691), .SEL(key[105]), .F(n1713) );
  NAND \e/a/U5555  ( .A(n1698), .B(n1688), .Z(n1712) );
  MUX \e/a/U5554  ( .IN0(n1699), .IN1(n1697), .SEL(key[105]), .F(n1711) );
  NAND \e/a/U5553  ( .A(n1710), .B(n1696), .Z(n1709) );
  MUX \e/a/U5552  ( .IN0(n1699), .IN1(n1691), .SEL(key[105]), .F(n1708) );
  NANDN \e/a/U5550  ( .B(key[108]), .A(key[107]), .Z(n1699) );
  MUX \e/a/U5549  ( .IN0(n1702), .IN1(n1691), .SEL(key[105]), .F(n1707) );
  MUX \e/a/U5548  ( .IN0(n1691), .IN1(n1651), .SEL(key[105]), .F(n1706) );
  MUX \e/a/U5547  ( .IN0(n1702), .IN1(key[107]), .SEL(key[105]), .F(n1705) );
  OR \e/a/U5546  ( .A(key[108]), .B(key[107]), .Z(n1702) );
  MUX \e/a/U5545  ( .IN0(n1688), .IN1(n1651), .SEL(key[105]), .F(n1704) );
  NANDN \e/a/U5544  ( .B(key[107]), .A(key[105]), .Z(n1703) );
  NAND \e/a/U5543  ( .A(n1702), .B(n1698), .Z(n1701) );
  NAND \e/a/U5542  ( .A(key[105]), .B(key[107]), .Z(n1700) );
  NAND \e/a/U5541  ( .A(key[105]), .B(n1699), .Z(n1698) );
  NANDN \e/a/U5540  ( .B(key[107]), .A(key[108]), .Z(n1697) );
  NAND \e/a/U5539  ( .A(key[108]), .B(key[107]), .Z(n1696) );
  MUX U659 ( .IN0(msg[99]), .IN1(\b/n5446 ), .SEL(msg[97]), .F(\b/n260 ) );
  MUX U660 ( .IN0(msg[107]), .IN1(\b/n5802 ), .SEL(msg[105]), .F(\b/n181 ) );
  MUX U661 ( .IN0(msg[75]), .IN1(\b/n4367 ), .SEL(msg[73]), .F(\b/n464 ) );
  MUX U662 ( .IN0(msg[43]), .IN1(\b/n2931 ), .SEL(msg[41]), .F(\b/n748 ) );
  MUX U663 ( .IN0(key[107]), .IN1(n1699), .SEL(key[105]), .F(n1677) );
  MUX U664 ( .IN0(n1702), .IN1(key[108]), .SEL(key[105]), .F(n1645) );
  MUX U665 ( .IN0(msg[91]), .IN1(\b/n5085 ), .SEL(msg[89]), .F(\b/n322 ) );
  MUX U666 ( .IN0(msg[51]), .IN1(\b/n3290 ), .SEL(msg[49]), .F(\b/n677 ) );
  MUX U667 ( .IN0(\b/n1501 ), .IN1(msg[12]), .SEL(msg[9]), .F(\b/n1014 ) );
  MUX U668 ( .IN0(\b/n3298 ), .IN1(\b/n3293 ), .SEL(msg[49]), .F(\b/n685 ) );
  MUX U669 ( .IN0(\b/n5088 ), .IN1(msg[92]), .SEL(msg[89]), .F(\b/n306 ) );
  MUX U670 ( .IN0(\b/n5449 ), .IN1(msg[100]), .SEL(msg[97]), .F(\b/n219 ) );
  MUX U671 ( .IN0(msg[59]), .IN1(\b/n3649 ), .SEL(msg[57]), .F(\b/n606 ) );
  MUX U672 ( .IN0(msg[19]), .IN1(\b/n1854 ), .SEL(msg[17]), .F(\b/n961 ) );
  MUX U673 ( .IN0(\b/n5805 ), .IN1(msg[108]), .SEL(msg[105]), .F(\b/n165 ) );
  MUX U674 ( .IN0(\b/n1862 ), .IN1(\b/n1857 ), .SEL(msg[17]), .F(\b/n969 ) );
  MUX U675 ( .IN0(\b/n3652 ), .IN1(msg[60]), .SEL(msg[57]), .F(\b/n590 ) );
  MUX U676 ( .IN0(\b/n4011 ), .IN1(msg[68]), .SEL(msg[65]), .F(\b/n519 ) );
  MUX U677 ( .IN0(msg[67]), .IN1(\b/n4008 ), .SEL(msg[65]), .F(\b/n535 ) );
  MUX U678 ( .IN0(msg[27]), .IN1(\b/n2213 ), .SEL(msg[25]), .F(\b/n890 ) );
  MUX U679 ( .IN0(msg[115]), .IN1(\b/n6161 ), .SEL(msg[113]), .F(\b/n110 ) );
  MUX U680 ( .IN0(\b/n4370 ), .IN1(msg[76]), .SEL(msg[73]), .F(\b/n448 ) );
  MUX U681 ( .IN0(\b/n6169 ), .IN1(\b/n6164 ), .SEL(msg[113]), .F(\b/n118 ) );
  MUX U682 ( .IN0(\b/n2216 ), .IN1(msg[28]), .SEL(msg[25]), .F(\b/n874 ) );
  MUX U683 ( .IN0(\b/n2575 ), .IN1(msg[36]), .SEL(msg[33]), .F(\b/n803 ) );
  MUX U684 ( .IN0(msg[35]), .IN1(\b/n2572 ), .SEL(msg[33]), .F(\b/n819 ) );
  MUX U685 ( .IN0(msg[123]), .IN1(\b/n6520 ), .SEL(msg[121]), .F(\b/n39 ) );
  MUX U686 ( .IN0(msg[83]), .IN1(\b/n4726 ), .SEL(msg[81]), .F(\b/n393 ) );
  MUX U687 ( .IN0(\b/n2934 ), .IN1(msg[44]), .SEL(msg[41]), .F(\b/n732 ) );
  MUX U688 ( .IN0(\b/n4734 ), .IN1(\b/n4729 ), .SEL(msg[81]), .F(\b/n401 ) );
  MUX U689 ( .IN0(\b/n6523 ), .IN1(msg[124]), .SEL(msg[121]), .F(\b/n23 ) );
  MUX U690 ( .IN0(\b/n1139 ), .IN1(msg[4]), .SEL(msg[1]), .F(\b/n1086 ) );
  MUX U691 ( .IN0(msg[3]), .IN1(\b/n1136 ), .SEL(msg[1]), .F(\b/n1102 ) );
  MUX U692 ( .IN0(\b/n1494 ), .IN1(msg[11]), .SEL(msg[9]), .F(\b/n1018 ) );
  MUX U693 ( .IN0(\b/n1535 ), .IN1(\b/n1538 ), .SEL(msg[15]), .F(n528) );
  IV U694 ( .A(n528), .Z(\b/n1770 ) );
  MUX U695 ( .IN0(\b/n5485 ), .IN1(\b/n5471 ), .SEL(msg[103]), .F(n529) );
  IV U696 ( .A(n529), .Z(\b/n5718 ) );
  MUX U697 ( .IN0(\b/n5801 ), .IN1(msg[107]), .SEL(msg[105]), .F(\b/n169 ) );
  MUX U698 ( .IN0(\b/n4366 ), .IN1(msg[75]), .SEL(msg[73]), .F(\b/n452 ) );
  MUX U699 ( .IN0(\b/n2930 ), .IN1(msg[43]), .SEL(msg[41]), .F(\b/n736 ) );
  MUX U700 ( .IN0(key[99]), .IN1(n2737), .SEL(key[97]), .F(n1500) );
  MUX U701 ( .IN0(n2740), .IN1(key[100]), .SEL(key[97]), .F(n1489) );
  MUX U702 ( .IN0(key[123]), .IN1(n2390), .SEL(key[121]), .F(n1556) );
  MUX U703 ( .IN0(n2393), .IN1(key[124]), .SEL(key[121]), .F(n1545) );
  MUX U704 ( .IN0(key[115]), .IN1(n2043), .SEL(key[113]), .F(n1612) );
  MUX U705 ( .IN0(n2046), .IN1(key[116]), .SEL(key[113]), .F(n1601) );
  MUX U706 ( .IN0(n1696), .IN1(key[107]), .SEL(key[105]), .F(n1648) );
  MUX U707 ( .IN0(n1697), .IN1(n1702), .SEL(key[105]), .F(n1657) );
  MUX U708 ( .IN0(msg[11]), .IN1(\b/n1497 ), .SEL(msg[9]), .F(\b/n1050 ) );
  MUX U709 ( .IN0(\b/n3293 ), .IN1(msg[52]), .SEL(msg[49]), .F(\b/n661 ) );
  MUX U710 ( .IN0(\b/n5093 ), .IN1(\b/n5088 ), .SEL(msg[89]), .F(\b/n330 ) );
  MUX U711 ( .IN0(\b/n1495 ), .IN1(\b/n1501 ), .SEL(msg[9]), .F(\b/n1029 ) );
  MUX U712 ( .IN0(\b/n5444 ), .IN1(\b/n5449 ), .SEL(msg[97]), .F(\b/n236 ) );
  MUX U713 ( .IN0(\b/n1857 ), .IN1(msg[20]), .SEL(msg[17]), .F(\b/n945 ) );
  MUX U714 ( .IN0(\b/n3657 ), .IN1(\b/n3652 ), .SEL(msg[57]), .F(\b/n614 ) );
  MUX U715 ( .IN0(\b/n5810 ), .IN1(\b/n5805 ), .SEL(msg[105]), .F(\b/n189 ) );
  MUX U716 ( .IN0(\b/n4016 ), .IN1(\b/n4011 ), .SEL(msg[65]), .F(\b/n543 ) );
  MUX U717 ( .IN0(\b/n6164 ), .IN1(msg[116]), .SEL(msg[113]), .F(\b/n94 ) );
  MUX U718 ( .IN0(\b/n2221 ), .IN1(\b/n2216 ), .SEL(msg[25]), .F(\b/n898 ) );
  MUX U719 ( .IN0(\b/n4375 ), .IN1(\b/n4370 ), .SEL(msg[73]), .F(\b/n472 ) );
  MUX U720 ( .IN0(\b/n2580 ), .IN1(\b/n2575 ), .SEL(msg[33]), .F(\b/n827 ) );
  MUX U721 ( .IN0(\b/n4729 ), .IN1(msg[84]), .SEL(msg[81]), .F(\b/n377 ) );
  MUX U722 ( .IN0(\b/n6528 ), .IN1(\b/n6523 ), .SEL(msg[121]), .F(\b/n47 ) );
  MUX U723 ( .IN0(\b/n2939 ), .IN1(\b/n2934 ), .SEL(msg[41]), .F(\b/n756 ) );
  MUX U724 ( .IN0(\b/n1144 ), .IN1(\b/n1139 ), .SEL(msg[1]), .F(\b/n1110 ) );
  MUX U725 ( .IN0(\b/n5084 ), .IN1(msg[91]), .SEL(msg[89]), .F(\b/n310 ) );
  MUX U726 ( .IN0(\b/n5125 ), .IN1(\b/n5110 ), .SEL(msg[95]), .F(n530) );
  IV U727 ( .A(n530), .Z(\b/n5368 ) );
  MUX U728 ( .IN0(\b/n3304 ), .IN1(\b/n3303 ), .SEL(msg[53]), .F(n531) );
  IV U729 ( .A(n531), .Z(\b/n3362 ) );
  MUX U730 ( .IN0(\b/n3289 ), .IN1(msg[51]), .SEL(msg[49]), .F(\b/n665 ) );
  XNOR U731 ( .A(msg[103]), .B(\b/n5470 ), .Z(\b/n5487 ) );
  MUX U732 ( .IN0(\b/n3648 ), .IN1(msg[59]), .SEL(msg[57]), .F(\b/n594 ) );
  MUX U733 ( .IN0(\b/n3689 ), .IN1(\b/n3674 ), .SEL(msg[63]), .F(n532) );
  IV U734 ( .A(n532), .Z(\b/n3932 ) );
  MUX U735 ( .IN0(\b/n1868 ), .IN1(\b/n1867 ), .SEL(msg[21]), .F(n533) );
  IV U736 ( .A(n533), .Z(\b/n1926 ) );
  MUX U737 ( .IN0(\b/n1853 ), .IN1(msg[19]), .SEL(msg[17]), .F(\b/n949 ) );
  MUX U738 ( .IN0(\b/n5842 ), .IN1(\b/n5827 ), .SEL(msg[111]), .F(n534) );
  IV U739 ( .A(n534), .Z(\b/n6085 ) );
  MUX U740 ( .IN0(\b/n4048 ), .IN1(\b/n4033 ), .SEL(msg[71]), .F(n535) );
  IV U741 ( .A(n535), .Z(\b/n4291 ) );
  XNOR U742 ( .A(msg[71]), .B(\b/n4034 ), .Z(\b/n4051 ) );
  MUX U743 ( .IN0(\b/n2212 ), .IN1(msg[27]), .SEL(msg[25]), .F(\b/n878 ) );
  MUX U744 ( .IN0(\b/n2253 ), .IN1(\b/n2238 ), .SEL(msg[31]), .F(n536) );
  IV U745 ( .A(n536), .Z(\b/n2496 ) );
  MUX U746 ( .IN0(\b/n6175 ), .IN1(\b/n6174 ), .SEL(msg[117]), .F(n537) );
  IV U747 ( .A(n537), .Z(\b/n6233 ) );
  MUX U748 ( .IN0(\b/n6160 ), .IN1(msg[115]), .SEL(msg[113]), .F(\b/n98 ) );
  MUX U749 ( .IN0(\b/n4407 ), .IN1(\b/n4392 ), .SEL(msg[79]), .F(n538) );
  IV U750 ( .A(n538), .Z(\b/n4650 ) );
  MUX U751 ( .IN0(\b/n2612 ), .IN1(\b/n2597 ), .SEL(msg[39]), .F(n539) );
  IV U752 ( .A(n539), .Z(\b/n2855 ) );
  XNOR U753 ( .A(msg[39]), .B(\b/n2598 ), .Z(\b/n2615 ) );
  MUX U754 ( .IN0(\b/n6519 ), .IN1(msg[123]), .SEL(msg[121]), .F(\b/n27 ) );
  MUX U755 ( .IN0(\b/n6560 ), .IN1(\b/n6545 ), .SEL(msg[127]), .F(n540) );
  IV U756 ( .A(n540), .Z(\b/n6803 ) );
  MUX U757 ( .IN0(\b/n4740 ), .IN1(\b/n4739 ), .SEL(msg[85]), .F(n541) );
  IV U758 ( .A(n541), .Z(\b/n4798 ) );
  XNOR U759 ( .A(msg[87]), .B(\b/n4752 ), .Z(\b/n4769 ) );
  MUX U760 ( .IN0(\b/n2971 ), .IN1(\b/n2956 ), .SEL(msg[47]), .F(n542) );
  IV U761 ( .A(n542), .Z(\b/n3214 ) );
  MUX U762 ( .IN0(\b/n1176 ), .IN1(\b/n1161 ), .SEL(msg[7]), .F(n543) );
  IV U763 ( .A(n543), .Z(\b/n1419 ) );
  MUX U764 ( .IN0(\b/n1135 ), .IN1(msg[3]), .SEL(msg[1]), .F(\b/n1090 ) );
  MUX U765 ( .IN0(n2745), .IN1(n2740), .SEL(key[97]), .F(n1506) );
  MUX U766 ( .IN0(n2398), .IN1(n2393), .SEL(key[121]), .F(n1562) );
  MUX U767 ( .IN0(n2051), .IN1(n2046), .SEL(key[113]), .F(n1618) );
  MUX U768 ( .IN0(n1734), .IN1(n1722), .SEL(key[111]), .F(n544) );
  IV U769 ( .A(n544), .Z(n1967) );
  NANDN U770 ( .B(\b/n1504 ), .A(msg[13]), .Z(\b/n1574 ) );
  NANDN U771 ( .B(\b/n5453 ), .A(msg[101]), .Z(\b/n5522 ) );
  NANDN U772 ( .B(\b/n5811 ), .A(msg[109]), .Z(\b/n5881 ) );
  NANDN U773 ( .B(\b/n4017 ), .A(msg[69]), .Z(\b/n4087 ) );
  NANDN U774 ( .B(\b/n4376 ), .A(msg[77]), .Z(\b/n4446 ) );
  NANDN U775 ( .B(\b/n2581 ), .A(msg[37]), .Z(\b/n2651 ) );
  NANDN U776 ( .B(\b/n4735 ), .A(msg[85]), .Z(\b/n4805 ) );
  NANDN U777 ( .B(\b/n2940 ), .A(msg[45]), .Z(\b/n3010 ) );
  MUX U778 ( .IN0(n2736), .IN1(key[99]), .SEL(key[97]), .F(n1491) );
  MUX U779 ( .IN0(n2773), .IN1(n2760), .SEL(key[103]), .F(n545) );
  IV U780 ( .A(n545), .Z(n3016) );
  MUX U781 ( .IN0(n2389), .IN1(key[123]), .SEL(key[121]), .F(n1547) );
  MUX U782 ( .IN0(n2426), .IN1(n2413), .SEL(key[127]), .F(n546) );
  IV U783 ( .A(n546), .Z(n2669) );
  MUX U784 ( .IN0(n2042), .IN1(key[115]), .SEL(key[113]), .F(n1603) );
  MUX U785 ( .IN0(n2079), .IN1(n2066), .SEL(key[119]), .F(n547) );
  IV U786 ( .A(n547), .Z(n2322) );
  XNOR U787 ( .A(key[111]), .B(n1721), .Z(n1736) );
  MUX U788 ( .IN0(counter[0]), .IN1(n548), .SEL(counter[3]), .F(n1400) );
  IV U789 ( .A(counter[1]), .Z(n548) );
  XNOR U790 ( .A(msg[95]), .B(\b/n5111 ), .Z(\b/n5128 ) );
  MUX U791 ( .IN0(\b/n5099 ), .IN1(\b/n5098 ), .SEL(msg[93]), .F(n549) );
  IV U792 ( .A(n549), .Z(\b/n5157 ) );
  MUX U793 ( .IN0(\b/n3330 ), .IN1(\b/n3315 ), .SEL(msg[55]), .F(n550) );
  IV U794 ( .A(n550), .Z(\b/n3573 ) );
  XNOR U795 ( .A(msg[55]), .B(\b/n3316 ), .Z(\b/n3333 ) );
  NAND U796 ( .A(\b/n1530 ), .B(msg[10]), .Z(\b/n1654 ) );
  NAND U797 ( .A(\b/n3326 ), .B(msg[50]), .Z(\b/n3449 ) );
  NAND U798 ( .A(\b/n5121 ), .B(msg[90]), .Z(\b/n5244 ) );
  NAND U799 ( .A(\b/n5481 ), .B(msg[98]), .Z(\b/n5602 ) );
  XNOR U800 ( .A(msg[15]), .B(\b/n1521 ), .Z(\b/n1537 ) );
  MUX U801 ( .IN0(\b/n5443 ), .IN1(msg[99]), .SEL(msg[97]), .F(\b/n224 ) );
  MUX U802 ( .IN0(\b/n1511 ), .IN1(\b/n1510 ), .SEL(msg[13]), .F(n551) );
  IV U803 ( .A(n551), .Z(\b/n1556 ) );
  MUX U804 ( .IN0(\b/n5460 ), .IN1(\b/n5459 ), .SEL(msg[101]), .F(n552) );
  IV U805 ( .A(n552), .Z(\b/n5504 ) );
  XNOR U806 ( .A(msg[63]), .B(\b/n3675 ), .Z(\b/n3692 ) );
  MUX U807 ( .IN0(\b/n3663 ), .IN1(\b/n3662 ), .SEL(msg[61]), .F(n553) );
  IV U808 ( .A(n553), .Z(\b/n3721 ) );
  MUX U809 ( .IN0(\b/n1894 ), .IN1(\b/n1879 ), .SEL(msg[23]), .F(n554) );
  IV U810 ( .A(n554), .Z(\b/n2137 ) );
  XNOR U811 ( .A(msg[23]), .B(\b/n1880 ), .Z(\b/n1897 ) );
  NAND U812 ( .A(\b/n5838 ), .B(msg[106]), .Z(\b/n5961 ) );
  NAND U813 ( .A(\b/n1890 ), .B(msg[18]), .Z(\b/n2013 ) );
  NAND U814 ( .A(\b/n3685 ), .B(msg[58]), .Z(\b/n3808 ) );
  NAND U815 ( .A(\b/n4044 ), .B(msg[66]), .Z(\b/n4167 ) );
  XNOR U816 ( .A(msg[111]), .B(\b/n5828 ), .Z(\b/n5845 ) );
  MUX U817 ( .IN0(\b/n4007 ), .IN1(msg[67]), .SEL(msg[65]), .F(\b/n523 ) );
  MUX U818 ( .IN0(\b/n5816 ), .IN1(\b/n5815 ), .SEL(msg[109]), .F(n555) );
  IV U819 ( .A(n555), .Z(\b/n5874 ) );
  MUX U820 ( .IN0(\b/n4022 ), .IN1(\b/n4021 ), .SEL(msg[69]), .F(n556) );
  IV U821 ( .A(n556), .Z(\b/n4080 ) );
  XNOR U822 ( .A(msg[31]), .B(\b/n2239 ), .Z(\b/n2256 ) );
  MUX U823 ( .IN0(\b/n2227 ), .IN1(\b/n2226 ), .SEL(msg[29]), .F(n557) );
  IV U824 ( .A(n557), .Z(\b/n2285 ) );
  MUX U825 ( .IN0(\b/n6201 ), .IN1(\b/n6186 ), .SEL(msg[119]), .F(n558) );
  IV U826 ( .A(n558), .Z(\b/n6444 ) );
  XNOR U827 ( .A(msg[119]), .B(\b/n6187 ), .Z(\b/n6204 ) );
  NAND U828 ( .A(\b/n4403 ), .B(msg[74]), .Z(\b/n4526 ) );
  NAND U829 ( .A(\b/n6197 ), .B(msg[114]), .Z(\b/n6320 ) );
  NAND U830 ( .A(\b/n2249 ), .B(msg[26]), .Z(\b/n2372 ) );
  NAND U831 ( .A(\b/n2608 ), .B(msg[34]), .Z(\b/n2731 ) );
  XNOR U832 ( .A(msg[79]), .B(\b/n4393 ), .Z(\b/n4410 ) );
  MUX U833 ( .IN0(\b/n2571 ), .IN1(msg[35]), .SEL(msg[33]), .F(\b/n807 ) );
  MUX U834 ( .IN0(\b/n4381 ), .IN1(\b/n4380 ), .SEL(msg[77]), .F(n559) );
  IV U835 ( .A(n559), .Z(\b/n4439 ) );
  MUX U836 ( .IN0(\b/n2586 ), .IN1(\b/n2585 ), .SEL(msg[37]), .F(n560) );
  IV U837 ( .A(n560), .Z(\b/n2644 ) );
  XNOR U838 ( .A(msg[127]), .B(\b/n6546 ), .Z(\b/n6563 ) );
  MUX U839 ( .IN0(\b/n6534 ), .IN1(\b/n6533 ), .SEL(msg[125]), .F(n561) );
  IV U840 ( .A(n561), .Z(\b/n6592 ) );
  MUX U841 ( .IN0(\b/n4766 ), .IN1(\b/n4751 ), .SEL(msg[87]), .F(n562) );
  IV U842 ( .A(n562), .Z(\b/n5009 ) );
  MUX U843 ( .IN0(\b/n4725 ), .IN1(msg[83]), .SEL(msg[81]), .F(\b/n381 ) );
  NAND U844 ( .A(\b/n2967 ), .B(msg[42]), .Z(\b/n3090 ) );
  NAND U845 ( .A(\b/n4762 ), .B(msg[82]), .Z(\b/n4885 ) );
  NAND U846 ( .A(\b/n6556 ), .B(msg[122]), .Z(\b/n6679 ) );
  NAND U847 ( .A(\b/n1172 ), .B(msg[2]), .Z(\b/n1295 ) );
  XNOR U848 ( .A(msg[47]), .B(\b/n2957 ), .Z(\b/n2974 ) );
  XNOR U849 ( .A(msg[7]), .B(\b/n1162 ), .Z(\b/n1179 ) );
  MUX U850 ( .IN0(\b/n2945 ), .IN1(\b/n2944 ), .SEL(msg[45]), .F(n563) );
  IV U851 ( .A(n563), .Z(\b/n3003 ) );
  MUX U852 ( .IN0(\b/n1150 ), .IN1(\b/n1149 ), .SEL(msg[5]), .F(n564) );
  IV U853 ( .A(n564), .Z(\b/n1208 ) );
  NAND U854 ( .A(n1731), .B(key[106]), .Z(n1851) );
  NANDN U855 ( .B(\b/n5094 ), .A(msg[93]), .Z(\b/n5164 ) );
  NANDN U856 ( .B(\b/n3299 ), .A(msg[53]), .Z(\b/n3369 ) );
  NANDN U857 ( .B(\b/n3658 ), .A(msg[61]), .Z(\b/n3728 ) );
  NANDN U858 ( .B(\b/n1863 ), .A(msg[21]), .Z(\b/n1933 ) );
  NANDN U859 ( .B(\b/n2222 ), .A(msg[29]), .Z(\b/n2292 ) );
  NANDN U860 ( .B(\b/n6170 ), .A(msg[117]), .Z(\b/n6240 ) );
  NANDN U861 ( .B(\b/n6529 ), .A(msg[125]), .Z(\b/n6599 ) );
  NANDN U862 ( .B(\b/n1145 ), .A(msg[5]), .Z(\b/n1215 ) );
  NAND U863 ( .A(n2770), .B(key[98]), .Z(n2892) );
  XNOR U864 ( .A(key[103]), .B(n2761), .Z(n2776) );
  MUX U865 ( .IN0(n2751), .IN1(n2750), .SEL(key[101]), .F(n565) );
  IV U866 ( .A(n565), .Z(n2805) );
  NAND U867 ( .A(n2423), .B(key[122]), .Z(n2545) );
  XNOR U868 ( .A(key[127]), .B(n2414), .Z(n2429) );
  MUX U869 ( .IN0(n2404), .IN1(n2403), .SEL(key[125]), .F(n566) );
  IV U870 ( .A(n566), .Z(n2458) );
  NAND U871 ( .A(n2076), .B(key[114]), .Z(n2198) );
  XNOR U872 ( .A(key[119]), .B(n2067), .Z(n2082) );
  MUX U873 ( .IN0(n2057), .IN1(n2056), .SEL(key[117]), .F(n567) );
  IV U874 ( .A(n567), .Z(n2111) );
  NANDN U875 ( .B(n1706), .A(key[109]), .Z(n1771) );
  MUX U876 ( .IN0(n1712), .IN1(n1711), .SEL(key[109]), .F(n568) );
  IV U877 ( .A(n568), .Z(n1753) );
  NANDN U878 ( .B(n2746), .A(key[101]), .Z(n2812) );
  NANDN U879 ( .B(n2399), .A(key[125]), .Z(n2465) );
  NANDN U880 ( .B(n2052), .A(key[117]), .Z(n2118) );
  XOR U881 ( .A(n1455), .B(n1456), .Z(\d/n384 ) );
  XOR U882 ( .A(n1439), .B(n1440), .Z(\d/n396 ) );
  XOR U883 ( .A(n1423), .B(n1424), .Z(\d/n408 ) );
  XOR U884 ( .A(n1411), .B(n1412), .Z(\d/n417 ) );
  MUX U885 ( .IN0(n1391), .IN1(counter[3]), .SEL(counter[0]), .F(n1405) );
  NOR U886 ( .A(key[105]), .B(key[107]), .Z(n569) );
  AND U887 ( .A(n1699), .B(n1772), .Z(n570) );
  AND U888 ( .A(n1696), .B(n1854), .Z(n571) );
  XNOR U889 ( .A(n1702), .B(key[105]), .Z(n572) );
  XNOR U890 ( .A(n1695), .B(key[111]), .Z(n573) );
  AND U891 ( .A(n1678), .B(key[105]), .Z(n574) );
  AND U892 ( .A(n1761), .B(n1688), .Z(n575) );
  XNOR U893 ( .A(n1696), .B(key[105]), .Z(n576) );
  NOR U894 ( .A(key[113]), .B(key[115]), .Z(n577) );
  AND U895 ( .A(n2043), .B(n2119), .Z(n578) );
  AND U896 ( .A(n2042), .B(n2201), .Z(n579) );
  XNOR U897 ( .A(n1585), .B(key[113]), .Z(n580) );
  XNOR U898 ( .A(n2046), .B(key[113]), .Z(n581) );
  AND U899 ( .A(key[113]), .B(n1613), .Z(n582) );
  AND U900 ( .A(n1594), .B(n2099), .Z(n583) );
  XNOR U901 ( .A(n2042), .B(key[113]), .Z(n584) );
  NOR U902 ( .A(key[121]), .B(key[123]), .Z(n585) );
  AND U903 ( .A(n2390), .B(n2466), .Z(n586) );
  AND U904 ( .A(n2389), .B(n2548), .Z(n587) );
  XNOR U905 ( .A(n1529), .B(key[121]), .Z(n588) );
  XNOR U906 ( .A(n2393), .B(key[121]), .Z(n589) );
  AND U907 ( .A(key[121]), .B(n1557), .Z(n590) );
  AND U908 ( .A(n1538), .B(n2446), .Z(n591) );
  XNOR U909 ( .A(n2389), .B(key[121]), .Z(n592) );
  NOR U910 ( .A(key[97]), .B(key[99]), .Z(n593) );
  AND U911 ( .A(n2737), .B(n2813), .Z(n594) );
  AND U912 ( .A(n2736), .B(n2895), .Z(n595) );
  XNOR U913 ( .A(n1473), .B(key[97]), .Z(n596) );
  XNOR U914 ( .A(n2740), .B(key[97]), .Z(n597) );
  AND U915 ( .A(key[97]), .B(n1501), .Z(n598) );
  AND U916 ( .A(n1482), .B(n2793), .Z(n599) );
  XNOR U917 ( .A(n2736), .B(key[97]), .Z(n600) );
  NOR U918 ( .A(msg[1]), .B(msg[3]), .Z(n601) );
  AND U919 ( .A(\b/n1136 ), .B(\b/n1216 ), .Z(n602) );
  AND U920 ( .A(\b/n1135 ), .B(\b/n1298 ), .Z(n603) );
  XNOR U921 ( .A(\b/n1065 ), .B(msg[1]), .Z(n604) );
  XNOR U922 ( .A(\b/n1139 ), .B(msg[1]), .Z(n605) );
  AND U923 ( .A(msg[1]), .B(\b/n1104 ), .Z(n606) );
  AND U924 ( .A(\b/n1077 ), .B(\b/n1196 ), .Z(n607) );
  XNOR U925 ( .A(\b/n1135 ), .B(msg[1]), .Z(n608) );
  NOR U926 ( .A(msg[11]), .B(msg[9]), .Z(n609) );
  AND U927 ( .A(\b/n1497 ), .B(\b/n1575 ), .Z(n610) );
  AND U928 ( .A(\b/n1494 ), .B(\b/n1657 ), .Z(n611) );
  XNOR U929 ( .A(\b/n1501 ), .B(msg[9]), .Z(n612) );
  XNOR U930 ( .A(\b/n1063 ), .B(msg[15]), .Z(n613) );
  AND U931 ( .A(\b/n1052 ), .B(msg[9]), .Z(n614) );
  AND U932 ( .A(\b/n1564 ), .B(\b/n1007 ), .Z(n615) );
  XNOR U933 ( .A(\b/n1494 ), .B(msg[9]), .Z(n616) );
  NOR U934 ( .A(msg[17]), .B(msg[19]), .Z(n617) );
  AND U935 ( .A(\b/n1854 ), .B(\b/n1934 ), .Z(n618) );
  AND U936 ( .A(\b/n1853 ), .B(\b/n2016 ), .Z(n619) );
  XNOR U937 ( .A(\b/n924 ), .B(msg[17]), .Z(n620) );
  XNOR U938 ( .A(\b/n1857 ), .B(msg[17]), .Z(n621) );
  AND U939 ( .A(msg[17]), .B(\b/n963 ), .Z(n622) );
  AND U940 ( .A(\b/n936 ), .B(\b/n1914 ), .Z(n623) );
  XNOR U941 ( .A(\b/n1853 ), .B(msg[17]), .Z(n624) );
  NOR U942 ( .A(msg[25]), .B(msg[27]), .Z(n625) );
  AND U943 ( .A(\b/n2213 ), .B(\b/n2293 ), .Z(n626) );
  AND U944 ( .A(\b/n2212 ), .B(\b/n2375 ), .Z(n627) );
  XNOR U945 ( .A(\b/n853 ), .B(msg[25]), .Z(n628) );
  XNOR U946 ( .A(\b/n2216 ), .B(msg[25]), .Z(n629) );
  AND U947 ( .A(msg[25]), .B(\b/n892 ), .Z(n630) );
  AND U948 ( .A(\b/n865 ), .B(\b/n2273 ), .Z(n631) );
  XNOR U949 ( .A(\b/n2212 ), .B(msg[25]), .Z(n632) );
  NOR U950 ( .A(msg[33]), .B(msg[35]), .Z(n633) );
  AND U951 ( .A(\b/n2572 ), .B(\b/n2652 ), .Z(n634) );
  AND U952 ( .A(\b/n2571 ), .B(\b/n2734 ), .Z(n635) );
  XNOR U953 ( .A(\b/n782 ), .B(msg[33]), .Z(n636) );
  XNOR U954 ( .A(\b/n2575 ), .B(msg[33]), .Z(n637) );
  AND U955 ( .A(msg[33]), .B(\b/n821 ), .Z(n638) );
  AND U956 ( .A(\b/n794 ), .B(\b/n2632 ), .Z(n639) );
  XNOR U957 ( .A(\b/n2571 ), .B(msg[33]), .Z(n640) );
  NOR U958 ( .A(msg[41]), .B(msg[43]), .Z(n641) );
  AND U959 ( .A(\b/n2931 ), .B(\b/n3011 ), .Z(n642) );
  AND U960 ( .A(\b/n2930 ), .B(\b/n3093 ), .Z(n643) );
  XNOR U961 ( .A(\b/n711 ), .B(msg[41]), .Z(n644) );
  XNOR U962 ( .A(\b/n2934 ), .B(msg[41]), .Z(n645) );
  AND U963 ( .A(msg[41]), .B(\b/n750 ), .Z(n646) );
  AND U964 ( .A(\b/n723 ), .B(\b/n2991 ), .Z(n647) );
  XNOR U965 ( .A(\b/n2930 ), .B(msg[41]), .Z(n648) );
  NOR U966 ( .A(msg[49]), .B(msg[51]), .Z(n649) );
  AND U967 ( .A(\b/n3290 ), .B(\b/n3370 ), .Z(n650) );
  AND U968 ( .A(\b/n3289 ), .B(\b/n3452 ), .Z(n651) );
  XNOR U969 ( .A(\b/n640 ), .B(msg[49]), .Z(n652) );
  XNOR U970 ( .A(\b/n3293 ), .B(msg[49]), .Z(n653) );
  AND U971 ( .A(msg[49]), .B(\b/n679 ), .Z(n654) );
  AND U972 ( .A(\b/n652 ), .B(\b/n3350 ), .Z(n655) );
  XNOR U973 ( .A(\b/n3289 ), .B(msg[49]), .Z(n656) );
  NOR U974 ( .A(msg[57]), .B(msg[59]), .Z(n657) );
  AND U975 ( .A(\b/n3649 ), .B(\b/n3729 ), .Z(n658) );
  AND U976 ( .A(\b/n3648 ), .B(\b/n3811 ), .Z(n659) );
  XNOR U977 ( .A(\b/n569 ), .B(msg[57]), .Z(n660) );
  XNOR U978 ( .A(\b/n3652 ), .B(msg[57]), .Z(n661) );
  AND U979 ( .A(msg[57]), .B(\b/n608 ), .Z(n662) );
  AND U980 ( .A(\b/n581 ), .B(\b/n3709 ), .Z(n663) );
  XNOR U981 ( .A(\b/n3648 ), .B(msg[57]), .Z(n664) );
  NOR U982 ( .A(msg[65]), .B(msg[67]), .Z(n665) );
  AND U983 ( .A(\b/n4008 ), .B(\b/n4088 ), .Z(n666) );
  AND U984 ( .A(\b/n4007 ), .B(\b/n4170 ), .Z(n667) );
  XNOR U985 ( .A(\b/n498 ), .B(msg[65]), .Z(n668) );
  XNOR U986 ( .A(\b/n4011 ), .B(msg[65]), .Z(n669) );
  AND U987 ( .A(msg[65]), .B(\b/n537 ), .Z(n670) );
  AND U988 ( .A(\b/n510 ), .B(\b/n4068 ), .Z(n671) );
  XNOR U989 ( .A(\b/n4007 ), .B(msg[65]), .Z(n672) );
  NOR U990 ( .A(msg[73]), .B(msg[75]), .Z(n673) );
  AND U991 ( .A(\b/n4367 ), .B(\b/n4447 ), .Z(n674) );
  AND U992 ( .A(\b/n4366 ), .B(\b/n4529 ), .Z(n675) );
  XNOR U993 ( .A(\b/n427 ), .B(msg[73]), .Z(n676) );
  XNOR U994 ( .A(\b/n4370 ), .B(msg[73]), .Z(n677) );
  AND U995 ( .A(msg[73]), .B(\b/n466 ), .Z(n678) );
  AND U996 ( .A(\b/n439 ), .B(\b/n4427 ), .Z(n679) );
  XNOR U997 ( .A(\b/n4366 ), .B(msg[73]), .Z(n680) );
  NOR U998 ( .A(msg[81]), .B(msg[83]), .Z(n681) );
  AND U999 ( .A(\b/n4726 ), .B(\b/n4806 ), .Z(n682) );
  AND U1000 ( .A(\b/n4725 ), .B(\b/n4888 ), .Z(n683) );
  XNOR U1001 ( .A(\b/n356 ), .B(msg[81]), .Z(n684) );
  XNOR U1002 ( .A(\b/n4729 ), .B(msg[81]), .Z(n685) );
  AND U1003 ( .A(msg[81]), .B(\b/n395 ), .Z(n686) );
  AND U1004 ( .A(\b/n368 ), .B(\b/n4786 ), .Z(n687) );
  XNOR U1005 ( .A(\b/n4725 ), .B(msg[81]), .Z(n688) );
  NOR U1006 ( .A(msg[89]), .B(msg[91]), .Z(n689) );
  AND U1007 ( .A(\b/n5085 ), .B(\b/n5165 ), .Z(n690) );
  AND U1008 ( .A(\b/n5084 ), .B(\b/n5247 ), .Z(n691) );
  XNOR U1009 ( .A(\b/n285 ), .B(msg[89]), .Z(n692) );
  XNOR U1010 ( .A(\b/n5088 ), .B(msg[89]), .Z(n693) );
  AND U1011 ( .A(msg[89]), .B(\b/n324 ), .Z(n694) );
  AND U1012 ( .A(\b/n297 ), .B(\b/n5145 ), .Z(n695) );
  XNOR U1013 ( .A(\b/n5084 ), .B(msg[89]), .Z(n696) );
  NOR U1014 ( .A(msg[97]), .B(msg[99]), .Z(n697) );
  AND U1015 ( .A(\b/n5446 ), .B(\b/n5523 ), .Z(n698) );
  AND U1016 ( .A(\b/n5443 ), .B(\b/n5605 ), .Z(n699) );
  XNOR U1017 ( .A(\b/n5449 ), .B(msg[97]), .Z(n700) );
  XNOR U1018 ( .A(\b/n283 ), .B(msg[103]), .Z(n701) );
  AND U1019 ( .A(\b/n262 ), .B(msg[97]), .Z(n702) );
  AND U1020 ( .A(\b/n5512 ), .B(\b/n275 ), .Z(n703) );
  XNOR U1021 ( .A(\b/n5443 ), .B(msg[97]), .Z(n704) );
  NOR U1022 ( .A(msg[105]), .B(msg[107]), .Z(n705) );
  AND U1023 ( .A(\b/n5802 ), .B(\b/n5882 ), .Z(n706) );
  AND U1024 ( .A(\b/n5801 ), .B(\b/n5964 ), .Z(n707) );
  XNOR U1025 ( .A(\b/n144 ), .B(msg[105]), .Z(n708) );
  XNOR U1026 ( .A(\b/n5805 ), .B(msg[105]), .Z(n709) );
  AND U1027 ( .A(msg[105]), .B(\b/n183 ), .Z(n710) );
  AND U1028 ( .A(\b/n156 ), .B(\b/n5862 ), .Z(n711) );
  XNOR U1029 ( .A(\b/n5801 ), .B(msg[105]), .Z(n712) );
  NOR U1030 ( .A(msg[113]), .B(msg[115]), .Z(n713) );
  AND U1031 ( .A(\b/n6161 ), .B(\b/n6241 ), .Z(n714) );
  AND U1032 ( .A(\b/n6160 ), .B(\b/n6323 ), .Z(n715) );
  XNOR U1033 ( .A(\b/n73 ), .B(msg[113]), .Z(n716) );
  XNOR U1034 ( .A(\b/n6164 ), .B(msg[113]), .Z(n717) );
  AND U1035 ( .A(msg[113]), .B(\b/n112 ), .Z(n718) );
  AND U1036 ( .A(\b/n85 ), .B(\b/n6221 ), .Z(n719) );
  XNOR U1037 ( .A(\b/n6160 ), .B(msg[113]), .Z(n720) );
  NOR U1038 ( .A(msg[121]), .B(msg[123]), .Z(n721) );
  AND U1039 ( .A(\b/n6520 ), .B(\b/n6600 ), .Z(n722) );
  AND U1040 ( .A(\b/n6519 ), .B(\b/n6682 ), .Z(n723) );
  XNOR U1041 ( .A(\b/n2 ), .B(msg[121]), .Z(n724) );
  XNOR U1042 ( .A(\b/n6523 ), .B(msg[121]), .Z(n725) );
  AND U1043 ( .A(msg[121]), .B(\b/n41 ), .Z(n726) );
  AND U1044 ( .A(\b/n14 ), .B(\b/n6580 ), .Z(n727) );
  XNOR U1045 ( .A(\b/n6519 ), .B(msg[121]), .Z(n728) );
  XNOR U1046 ( .A(key[103]), .B(\e/n118 ), .Z(n729) );
  XNOR U1047 ( .A(key[102]), .B(\e/n117 ), .Z(n730) );
  XNOR U1048 ( .A(key[101]), .B(\e/n116 ), .Z(n731) );
  XNOR U1049 ( .A(key[100]), .B(\e/n115 ), .Z(n732) );
  XNOR U1050 ( .A(key[99]), .B(\e/n114 ), .Z(n733) );
  XNOR U1051 ( .A(key[98]), .B(\e/n113 ), .Z(n734) );
  XNOR U1052 ( .A(key[97]), .B(\e/n112 ), .Z(n735) );
  XNOR U1053 ( .A(key[96]), .B(\e/n111 ), .Z(n736) );
  XOR U1054 ( .A(n737), .B(key[9]), .Z(o[9]) );
  NAND U1055 ( .A(n738), .B(n739), .Z(n737) );
  NANDN U1056 ( .B(\b/n1063 ), .A(n740), .Z(n739) );
  AND U1057 ( .A(n741), .B(n742), .Z(n738) );
  NANDN U1058 ( .B(\d/n424 ), .A(n743), .Z(n742) );
  NAND U1059 ( .A(n744), .B(shift_row_out[9]), .Z(n741) );
  XNOR U1060 ( .A(n745), .B(n1524), .Z(o[99]) );
  NAND U1061 ( .A(n746), .B(n747), .Z(n745) );
  NANDN U1062 ( .B(\b/n278 ), .A(n740), .Z(n747) );
  AND U1063 ( .A(n748), .B(n749), .Z(n746) );
  NANDN U1064 ( .B(\d/n458 ), .A(n743), .Z(n749) );
  NAND U1065 ( .A(n744), .B(shift_row_out[99]), .Z(n748) );
  XOR U1066 ( .A(n750), .B(key[98]), .Z(o[98]) );
  NAND U1067 ( .A(n751), .B(n752), .Z(n750) );
  NAND U1068 ( .A(n740), .B(msg[98]), .Z(n752) );
  AND U1069 ( .A(n753), .B(n754), .Z(n751) );
  NAND U1070 ( .A(n743), .B(mix_col_out[98]), .Z(n754) );
  NAND U1071 ( .A(n744), .B(shift_row_out[98]), .Z(n753) );
  XNOR U1072 ( .A(n755), .B(n1528), .Z(o[97]) );
  NAND U1073 ( .A(n756), .B(n757), .Z(n755) );
  NANDN U1074 ( .B(\b/n283 ), .A(n740), .Z(n757) );
  AND U1075 ( .A(n758), .B(n759), .Z(n756) );
  NANDN U1076 ( .B(\d/n457 ), .A(n743), .Z(n759) );
  NAND U1077 ( .A(n744), .B(shift_row_out[97]), .Z(n758) );
  XOR U1078 ( .A(n760), .B(key[96]), .Z(o[96]) );
  NAND U1079 ( .A(n761), .B(n762), .Z(n760) );
  NAND U1080 ( .A(n740), .B(msg[96]), .Z(n762) );
  AND U1081 ( .A(n763), .B(n764), .Z(n761) );
  NAND U1082 ( .A(n743), .B(mix_col_out[96]), .Z(n764) );
  NAND U1083 ( .A(n744), .B(shift_row_out[96]), .Z(n763) );
  XOR U1084 ( .A(n765), .B(key[95]), .Z(o[95]) );
  NAND U1085 ( .A(n766), .B(n767), .Z(n765) );
  NANDN U1086 ( .B(\b/n285 ), .A(n740), .Z(n767) );
  AND U1087 ( .A(n768), .B(n769), .Z(n766) );
  NAND U1088 ( .A(n743), .B(mix_col_out[95]), .Z(n769) );
  NAND U1089 ( .A(n744), .B(shift_row_out[95]), .Z(n768) );
  XOR U1090 ( .A(n770), .B(key[94]), .Z(o[94]) );
  NAND U1091 ( .A(n771), .B(n772), .Z(n770) );
  NAND U1092 ( .A(n740), .B(msg[94]), .Z(n772) );
  AND U1093 ( .A(n773), .B(n774), .Z(n771) );
  NAND U1094 ( .A(n743), .B(mix_col_out[94]), .Z(n774) );
  NAND U1095 ( .A(n744), .B(shift_row_out[94]), .Z(n773) );
  XOR U1096 ( .A(n775), .B(key[93]), .Z(o[93]) );
  NAND U1097 ( .A(n776), .B(n777), .Z(n775) );
  NAND U1098 ( .A(n740), .B(msg[93]), .Z(n777) );
  AND U1099 ( .A(n778), .B(n779), .Z(n776) );
  NAND U1100 ( .A(n743), .B(mix_col_out[93]), .Z(n779) );
  NAND U1101 ( .A(n744), .B(shift_row_out[93]), .Z(n778) );
  XOR U1102 ( .A(n780), .B(key[92]), .Z(o[92]) );
  NAND U1103 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U1104 ( .B(\b/n307 ), .A(n740), .Z(n782) );
  AND U1105 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U1106 ( .B(\d/n456 ), .A(n743), .Z(n784) );
  NAND U1107 ( .A(n744), .B(shift_row_out[92]), .Z(n783) );
  XOR U1108 ( .A(n785), .B(key[91]), .Z(o[91]) );
  NAND U1109 ( .A(n786), .B(n787), .Z(n785) );
  NANDN U1110 ( .B(\b/n349 ), .A(n740), .Z(n787) );
  AND U1111 ( .A(n788), .B(n789), .Z(n786) );
  NANDN U1112 ( .B(\d/n455 ), .A(n743), .Z(n789) );
  NAND U1113 ( .A(n744), .B(shift_row_out[91]), .Z(n788) );
  XOR U1114 ( .A(n790), .B(key[90]), .Z(o[90]) );
  NAND U1115 ( .A(n791), .B(n792), .Z(n790) );
  NAND U1116 ( .A(n740), .B(msg[90]), .Z(n792) );
  AND U1117 ( .A(n793), .B(n794), .Z(n791) );
  NAND U1118 ( .A(n743), .B(mix_col_out[90]), .Z(n794) );
  NAND U1119 ( .A(n744), .B(shift_row_out[90]), .Z(n793) );
  XOR U1120 ( .A(n795), .B(key[8]), .Z(o[8]) );
  NAND U1121 ( .A(n796), .B(n797), .Z(n795) );
  NAND U1122 ( .A(n740), .B(msg[8]), .Z(n797) );
  AND U1123 ( .A(n798), .B(n799), .Z(n796) );
  NAND U1124 ( .A(n743), .B(mix_col_out[8]), .Z(n799) );
  NAND U1125 ( .A(n744), .B(shift_row_out[8]), .Z(n798) );
  XOR U1126 ( .A(n800), .B(key[89]), .Z(o[89]) );
  NAND U1127 ( .A(n801), .B(n802), .Z(n800) );
  NANDN U1128 ( .B(\b/n354 ), .A(n740), .Z(n802) );
  AND U1129 ( .A(n803), .B(n804), .Z(n801) );
  NANDN U1130 ( .B(\d/n454 ), .A(n743), .Z(n804) );
  NAND U1131 ( .A(n744), .B(shift_row_out[89]), .Z(n803) );
  XOR U1132 ( .A(n805), .B(key[88]), .Z(o[88]) );
  NAND U1133 ( .A(n806), .B(n807), .Z(n805) );
  NAND U1134 ( .A(n740), .B(msg[88]), .Z(n807) );
  AND U1135 ( .A(n808), .B(n809), .Z(n806) );
  NAND U1136 ( .A(n743), .B(mix_col_out[88]), .Z(n809) );
  NAND U1137 ( .A(n744), .B(shift_row_out[88]), .Z(n808) );
  XOR U1138 ( .A(n810), .B(key[87]), .Z(o[87]) );
  NAND U1139 ( .A(n811), .B(n812), .Z(n810) );
  NANDN U1140 ( .B(\b/n356 ), .A(n740), .Z(n812) );
  AND U1141 ( .A(n813), .B(n814), .Z(n811) );
  NAND U1142 ( .A(n743), .B(mix_col_out[87]), .Z(n814) );
  NANDN U1143 ( .B(n815), .A(n744), .Z(n813) );
  XOR U1144 ( .A(n816), .B(key[86]), .Z(o[86]) );
  NAND U1145 ( .A(n817), .B(n818), .Z(n816) );
  NAND U1146 ( .A(n740), .B(msg[86]), .Z(n818) );
  AND U1147 ( .A(n819), .B(n820), .Z(n817) );
  NAND U1148 ( .A(n743), .B(mix_col_out[86]), .Z(n820) );
  NAND U1149 ( .A(n744), .B(shift_row_out[86]), .Z(n819) );
  XOR U1150 ( .A(n821), .B(key[85]), .Z(o[85]) );
  NAND U1151 ( .A(n822), .B(n823), .Z(n821) );
  NAND U1152 ( .A(n740), .B(msg[85]), .Z(n823) );
  AND U1153 ( .A(n824), .B(n825), .Z(n822) );
  NAND U1154 ( .A(n743), .B(mix_col_out[85]), .Z(n825) );
  NAND U1155 ( .A(n744), .B(shift_row_out[85]), .Z(n824) );
  XOR U1156 ( .A(n826), .B(key[84]), .Z(o[84]) );
  NAND U1157 ( .A(n827), .B(n828), .Z(n826) );
  NANDN U1158 ( .B(\b/n378 ), .A(n740), .Z(n828) );
  AND U1159 ( .A(n829), .B(n830), .Z(n827) );
  NANDN U1160 ( .B(\d/n453 ), .A(n743), .Z(n830) );
  NAND U1161 ( .A(n744), .B(shift_row_out[84]), .Z(n829) );
  XOR U1162 ( .A(n831), .B(key[83]), .Z(o[83]) );
  NAND U1163 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U1164 ( .B(\b/n420 ), .A(n740), .Z(n833) );
  AND U1165 ( .A(n834), .B(n835), .Z(n832) );
  NANDN U1166 ( .B(\d/n452 ), .A(n743), .Z(n835) );
  NAND U1167 ( .A(n744), .B(shift_row_out[83]), .Z(n834) );
  XOR U1168 ( .A(n836), .B(key[82]), .Z(o[82]) );
  NAND U1169 ( .A(n837), .B(n838), .Z(n836) );
  NAND U1170 ( .A(n740), .B(msg[82]), .Z(n838) );
  AND U1171 ( .A(n839), .B(n840), .Z(n837) );
  NAND U1172 ( .A(n743), .B(mix_col_out[82]), .Z(n840) );
  NAND U1173 ( .A(n744), .B(shift_row_out[82]), .Z(n839) );
  XOR U1174 ( .A(n841), .B(key[81]), .Z(o[81]) );
  NAND U1175 ( .A(n842), .B(n843), .Z(n841) );
  NANDN U1176 ( .B(\b/n425 ), .A(n740), .Z(n843) );
  AND U1177 ( .A(n844), .B(n845), .Z(n842) );
  NANDN U1178 ( .B(\d/n451 ), .A(n743), .Z(n845) );
  NAND U1179 ( .A(n744), .B(shift_row_out[81]), .Z(n844) );
  XOR U1180 ( .A(n846), .B(key[80]), .Z(o[80]) );
  NAND U1181 ( .A(n847), .B(n848), .Z(n846) );
  NAND U1182 ( .A(n740), .B(msg[80]), .Z(n848) );
  AND U1183 ( .A(n849), .B(n850), .Z(n847) );
  NAND U1184 ( .A(n743), .B(mix_col_out[80]), .Z(n850) );
  NAND U1185 ( .A(n744), .B(shift_row_out[80]), .Z(n849) );
  XOR U1186 ( .A(n851), .B(key[7]), .Z(o[7]) );
  NAND U1187 ( .A(n852), .B(n853), .Z(n851) );
  NANDN U1188 ( .B(\b/n1065 ), .A(n740), .Z(n853) );
  AND U1189 ( .A(n854), .B(n855), .Z(n852) );
  NAND U1190 ( .A(n743), .B(mix_col_out[7]), .Z(n855) );
  NAND U1191 ( .A(n744), .B(shift_row_out[7]), .Z(n854) );
  XOR U1192 ( .A(n856), .B(key[79]), .Z(o[79]) );
  NAND U1193 ( .A(n857), .B(n858), .Z(n856) );
  NANDN U1194 ( .B(\b/n427 ), .A(n740), .Z(n858) );
  AND U1195 ( .A(n859), .B(n860), .Z(n857) );
  NAND U1196 ( .A(n743), .B(mix_col_out[79]), .Z(n860) );
  NANDN U1197 ( .B(n861), .A(n744), .Z(n859) );
  XOR U1198 ( .A(n862), .B(key[78]), .Z(o[78]) );
  NAND U1199 ( .A(n863), .B(n864), .Z(n862) );
  NAND U1200 ( .A(n740), .B(msg[78]), .Z(n864) );
  AND U1201 ( .A(n865), .B(n866), .Z(n863) );
  NAND U1202 ( .A(n743), .B(mix_col_out[78]), .Z(n866) );
  NAND U1203 ( .A(n744), .B(shift_row_out[78]), .Z(n865) );
  XOR U1204 ( .A(n867), .B(key[77]), .Z(o[77]) );
  NAND U1205 ( .A(n868), .B(n869), .Z(n867) );
  NAND U1206 ( .A(n740), .B(msg[77]), .Z(n869) );
  AND U1207 ( .A(n870), .B(n871), .Z(n868) );
  NAND U1208 ( .A(n743), .B(mix_col_out[77]), .Z(n871) );
  NAND U1209 ( .A(n744), .B(shift_row_out[77]), .Z(n870) );
  XOR U1210 ( .A(n872), .B(key[76]), .Z(o[76]) );
  NAND U1211 ( .A(n873), .B(n874), .Z(n872) );
  NANDN U1212 ( .B(\b/n449 ), .A(n740), .Z(n874) );
  AND U1213 ( .A(n875), .B(n876), .Z(n873) );
  NANDN U1214 ( .B(\d/n450 ), .A(n743), .Z(n876) );
  NAND U1215 ( .A(n744), .B(shift_row_out[76]), .Z(n875) );
  XOR U1216 ( .A(n877), .B(key[75]), .Z(o[75]) );
  NAND U1217 ( .A(n878), .B(n879), .Z(n877) );
  NANDN U1218 ( .B(\b/n491 ), .A(n740), .Z(n879) );
  AND U1219 ( .A(n880), .B(n881), .Z(n878) );
  NANDN U1220 ( .B(\d/n449 ), .A(n743), .Z(n881) );
  NAND U1221 ( .A(n744), .B(shift_row_out[75]), .Z(n880) );
  XOR U1222 ( .A(n882), .B(key[74]), .Z(o[74]) );
  NAND U1223 ( .A(n883), .B(n884), .Z(n882) );
  NAND U1224 ( .A(n740), .B(msg[74]), .Z(n884) );
  AND U1225 ( .A(n885), .B(n886), .Z(n883) );
  NAND U1226 ( .A(n743), .B(mix_col_out[74]), .Z(n886) );
  NAND U1227 ( .A(n744), .B(shift_row_out[74]), .Z(n885) );
  XOR U1228 ( .A(n887), .B(key[73]), .Z(o[73]) );
  NAND U1229 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U1230 ( .B(\b/n496 ), .A(n740), .Z(n889) );
  AND U1231 ( .A(n890), .B(n891), .Z(n888) );
  NANDN U1232 ( .B(\d/n448 ), .A(n743), .Z(n891) );
  NAND U1233 ( .A(n744), .B(shift_row_out[73]), .Z(n890) );
  XOR U1234 ( .A(n892), .B(key[72]), .Z(o[72]) );
  NAND U1235 ( .A(n893), .B(n894), .Z(n892) );
  NAND U1236 ( .A(n740), .B(msg[72]), .Z(n894) );
  AND U1237 ( .A(n895), .B(n896), .Z(n893) );
  NAND U1238 ( .A(n743), .B(mix_col_out[72]), .Z(n896) );
  NAND U1239 ( .A(n744), .B(shift_row_out[72]), .Z(n895) );
  XOR U1240 ( .A(n897), .B(key[71]), .Z(o[71]) );
  NAND U1241 ( .A(n898), .B(n899), .Z(n897) );
  NANDN U1242 ( .B(\b/n498 ), .A(n740), .Z(n899) );
  AND U1243 ( .A(n900), .B(n901), .Z(n898) );
  NAND U1244 ( .A(n743), .B(mix_col_out[71]), .Z(n901) );
  NAND U1245 ( .A(n744), .B(shift_row_out[71]), .Z(n900) );
  XOR U1246 ( .A(n902), .B(key[70]), .Z(o[70]) );
  NAND U1247 ( .A(n903), .B(n904), .Z(n902) );
  NAND U1248 ( .A(n740), .B(msg[70]), .Z(n904) );
  AND U1249 ( .A(n905), .B(n906), .Z(n903) );
  NAND U1250 ( .A(n743), .B(mix_col_out[70]), .Z(n906) );
  NAND U1251 ( .A(n744), .B(shift_row_out[70]), .Z(n905) );
  XOR U1252 ( .A(n907), .B(key[6]), .Z(o[6]) );
  NAND U1253 ( .A(n908), .B(n909), .Z(n907) );
  NAND U1254 ( .A(n740), .B(msg[6]), .Z(n909) );
  AND U1255 ( .A(n910), .B(n911), .Z(n908) );
  NAND U1256 ( .A(n743), .B(mix_col_out[6]), .Z(n911) );
  NAND U1257 ( .A(n744), .B(shift_row_out[6]), .Z(n910) );
  XOR U1258 ( .A(n912), .B(key[69]), .Z(o[69]) );
  NAND U1259 ( .A(n913), .B(n914), .Z(n912) );
  NAND U1260 ( .A(n740), .B(msg[69]), .Z(n914) );
  AND U1261 ( .A(n915), .B(n916), .Z(n913) );
  NAND U1262 ( .A(n743), .B(mix_col_out[69]), .Z(n916) );
  NAND U1263 ( .A(n744), .B(shift_row_out[69]), .Z(n915) );
  XOR U1264 ( .A(n917), .B(key[68]), .Z(o[68]) );
  NAND U1265 ( .A(n918), .B(n919), .Z(n917) );
  NANDN U1266 ( .B(\b/n520 ), .A(n740), .Z(n919) );
  AND U1267 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1268 ( .B(\d/n447 ), .A(n743), .Z(n921) );
  NAND U1269 ( .A(n744), .B(shift_row_out[68]), .Z(n920) );
  XOR U1270 ( .A(n922), .B(key[67]), .Z(o[67]) );
  NAND U1271 ( .A(n923), .B(n924), .Z(n922) );
  NANDN U1272 ( .B(\b/n562 ), .A(n740), .Z(n924) );
  AND U1273 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1274 ( .B(\d/n446 ), .A(n743), .Z(n926) );
  NAND U1275 ( .A(shift_row_out[67]), .B(n744), .Z(n925) );
  XOR U1276 ( .A(n927), .B(key[66]), .Z(o[66]) );
  NAND U1277 ( .A(n928), .B(n929), .Z(n927) );
  NAND U1278 ( .A(n740), .B(msg[66]), .Z(n929) );
  AND U1279 ( .A(n930), .B(n931), .Z(n928) );
  NAND U1280 ( .A(n743), .B(mix_col_out[66]), .Z(n931) );
  NAND U1281 ( .A(shift_row_out[66]), .B(n744), .Z(n930) );
  XOR U1282 ( .A(n932), .B(key[65]), .Z(o[65]) );
  NAND U1283 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U1284 ( .B(\b/n567 ), .A(n740), .Z(n934) );
  AND U1285 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U1286 ( .B(\d/n445 ), .A(n743), .Z(n936) );
  NAND U1287 ( .A(n744), .B(shift_row_out[65]), .Z(n935) );
  XOR U1288 ( .A(n937), .B(key[64]), .Z(o[64]) );
  NAND U1289 ( .A(n938), .B(n939), .Z(n937) );
  NAND U1290 ( .A(n740), .B(msg[64]), .Z(n939) );
  AND U1291 ( .A(n940), .B(n941), .Z(n938) );
  NAND U1292 ( .A(n743), .B(mix_col_out[64]), .Z(n941) );
  NAND U1293 ( .A(shift_row_out[64]), .B(n744), .Z(n940) );
  XOR U1294 ( .A(n942), .B(key[63]), .Z(o[63]) );
  NAND U1295 ( .A(n943), .B(n944), .Z(n942) );
  NANDN U1296 ( .B(\b/n569 ), .A(n740), .Z(n944) );
  AND U1297 ( .A(n945), .B(n946), .Z(n943) );
  NAND U1298 ( .A(n743), .B(mix_col_out[63]), .Z(n946) );
  NAND U1299 ( .A(n744), .B(shift_row_out[63]), .Z(n945) );
  XOR U1300 ( .A(n947), .B(key[62]), .Z(o[62]) );
  NAND U1301 ( .A(n948), .B(n949), .Z(n947) );
  NAND U1302 ( .A(n740), .B(msg[62]), .Z(n949) );
  AND U1303 ( .A(n950), .B(n951), .Z(n948) );
  NAND U1304 ( .A(n743), .B(mix_col_out[62]), .Z(n951) );
  NAND U1305 ( .A(n744), .B(shift_row_out[62]), .Z(n950) );
  XOR U1306 ( .A(n952), .B(key[61]), .Z(o[61]) );
  NAND U1307 ( .A(n953), .B(n954), .Z(n952) );
  NAND U1308 ( .A(n740), .B(msg[61]), .Z(n954) );
  AND U1309 ( .A(n955), .B(n956), .Z(n953) );
  NAND U1310 ( .A(n743), .B(mix_col_out[61]), .Z(n956) );
  NAND U1311 ( .A(n744), .B(shift_row_out[61]), .Z(n955) );
  XOR U1312 ( .A(n957), .B(key[60]), .Z(o[60]) );
  NAND U1313 ( .A(n958), .B(n959), .Z(n957) );
  NANDN U1314 ( .B(\b/n591 ), .A(n740), .Z(n959) );
  AND U1315 ( .A(n960), .B(n961), .Z(n958) );
  NANDN U1316 ( .B(\d/n444 ), .A(n743), .Z(n961) );
  NAND U1317 ( .A(n744), .B(shift_row_out[60]), .Z(n960) );
  XOR U1318 ( .A(n962), .B(key[5]), .Z(o[5]) );
  NAND U1319 ( .A(n963), .B(n964), .Z(n962) );
  NAND U1320 ( .A(n740), .B(msg[5]), .Z(n964) );
  AND U1321 ( .A(n965), .B(n966), .Z(n963) );
  NAND U1322 ( .A(n743), .B(mix_col_out[5]), .Z(n966) );
  NAND U1323 ( .A(n744), .B(shift_row_out[5]), .Z(n965) );
  XOR U1324 ( .A(n967), .B(key[59]), .Z(o[59]) );
  NAND U1325 ( .A(n968), .B(n969), .Z(n967) );
  NANDN U1326 ( .B(\b/n633 ), .A(n740), .Z(n969) );
  AND U1327 ( .A(n970), .B(n971), .Z(n968) );
  NANDN U1328 ( .B(\d/n443 ), .A(n743), .Z(n971) );
  NAND U1329 ( .A(n744), .B(shift_row_out[59]), .Z(n970) );
  XOR U1330 ( .A(n972), .B(key[58]), .Z(o[58]) );
  NAND U1331 ( .A(n973), .B(n974), .Z(n972) );
  NAND U1332 ( .A(n740), .B(msg[58]), .Z(n974) );
  AND U1333 ( .A(n975), .B(n976), .Z(n973) );
  NAND U1334 ( .A(n743), .B(mix_col_out[58]), .Z(n976) );
  NAND U1335 ( .A(n744), .B(shift_row_out[58]), .Z(n975) );
  XOR U1336 ( .A(n977), .B(key[57]), .Z(o[57]) );
  NAND U1337 ( .A(n978), .B(n979), .Z(n977) );
  NANDN U1338 ( .B(\b/n638 ), .A(n740), .Z(n979) );
  AND U1339 ( .A(n980), .B(n981), .Z(n978) );
  NANDN U1340 ( .B(\d/n442 ), .A(n743), .Z(n981) );
  NAND U1341 ( .A(n744), .B(shift_row_out[57]), .Z(n980) );
  XOR U1342 ( .A(n982), .B(key[56]), .Z(o[56]) );
  NAND U1343 ( .A(n983), .B(n984), .Z(n982) );
  NAND U1344 ( .A(n740), .B(msg[56]), .Z(n984) );
  AND U1345 ( .A(n985), .B(n986), .Z(n983) );
  NAND U1346 ( .A(n743), .B(mix_col_out[56]), .Z(n986) );
  NAND U1347 ( .A(n744), .B(shift_row_out[56]), .Z(n985) );
  XOR U1348 ( .A(n987), .B(key[55]), .Z(o[55]) );
  NAND U1349 ( .A(n988), .B(n989), .Z(n987) );
  NANDN U1350 ( .B(\b/n640 ), .A(n740), .Z(n989) );
  AND U1351 ( .A(n990), .B(n991), .Z(n988) );
  NAND U1352 ( .A(n743), .B(mix_col_out[55]), .Z(n991) );
  NANDN U1353 ( .B(n992), .A(n744), .Z(n990) );
  XOR U1354 ( .A(n993), .B(key[54]), .Z(o[54]) );
  NAND U1355 ( .A(n994), .B(n995), .Z(n993) );
  NAND U1356 ( .A(n740), .B(msg[54]), .Z(n995) );
  AND U1357 ( .A(n996), .B(n997), .Z(n994) );
  NAND U1358 ( .A(n743), .B(mix_col_out[54]), .Z(n997) );
  NAND U1359 ( .A(n744), .B(shift_row_out[54]), .Z(n996) );
  XOR U1360 ( .A(n998), .B(key[53]), .Z(o[53]) );
  NAND U1361 ( .A(n999), .B(n1000), .Z(n998) );
  NAND U1362 ( .A(n740), .B(msg[53]), .Z(n1000) );
  AND U1363 ( .A(n1001), .B(n1002), .Z(n999) );
  NAND U1364 ( .A(n743), .B(mix_col_out[53]), .Z(n1002) );
  NAND U1365 ( .A(n744), .B(shift_row_out[53]), .Z(n1001) );
  XOR U1366 ( .A(n1003), .B(key[52]), .Z(o[52]) );
  NAND U1367 ( .A(n1004), .B(n1005), .Z(n1003) );
  NANDN U1368 ( .B(\b/n662 ), .A(n740), .Z(n1005) );
  AND U1369 ( .A(n1006), .B(n1007), .Z(n1004) );
  NANDN U1370 ( .B(\d/n441 ), .A(n743), .Z(n1007) );
  NAND U1371 ( .A(n744), .B(shift_row_out[52]), .Z(n1006) );
  XOR U1372 ( .A(n1008), .B(key[51]), .Z(o[51]) );
  NAND U1373 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U1374 ( .B(\b/n704 ), .A(n740), .Z(n1010) );
  AND U1375 ( .A(n1011), .B(n1012), .Z(n1009) );
  NANDN U1376 ( .B(\d/n440 ), .A(n743), .Z(n1012) );
  NAND U1377 ( .A(n744), .B(shift_row_out[51]), .Z(n1011) );
  XOR U1378 ( .A(n1013), .B(key[50]), .Z(o[50]) );
  NAND U1379 ( .A(n1014), .B(n1015), .Z(n1013) );
  NAND U1380 ( .A(n740), .B(msg[50]), .Z(n1015) );
  AND U1381 ( .A(n1016), .B(n1017), .Z(n1014) );
  NAND U1382 ( .A(n743), .B(mix_col_out[50]), .Z(n1017) );
  NAND U1383 ( .A(n744), .B(shift_row_out[50]), .Z(n1016) );
  XOR U1384 ( .A(n1018), .B(key[4]), .Z(o[4]) );
  NAND U1385 ( .A(n1019), .B(n1020), .Z(n1018) );
  NANDN U1386 ( .B(\b/n1087 ), .A(n740), .Z(n1020) );
  AND U1387 ( .A(n1021), .B(n1022), .Z(n1019) );
  NANDN U1388 ( .B(\d/n423 ), .A(n743), .Z(n1022) );
  NAND U1389 ( .A(n744), .B(shift_row_out[4]), .Z(n1021) );
  XOR U1390 ( .A(n1023), .B(key[49]), .Z(o[49]) );
  NAND U1391 ( .A(n1024), .B(n1025), .Z(n1023) );
  NANDN U1392 ( .B(\b/n709 ), .A(n740), .Z(n1025) );
  AND U1393 ( .A(n1026), .B(n1027), .Z(n1024) );
  NANDN U1394 ( .B(\d/n439 ), .A(n743), .Z(n1027) );
  NAND U1395 ( .A(n744), .B(shift_row_out[49]), .Z(n1026) );
  XOR U1396 ( .A(n1028), .B(key[48]), .Z(o[48]) );
  NAND U1397 ( .A(n1029), .B(n1030), .Z(n1028) );
  NAND U1398 ( .A(n740), .B(msg[48]), .Z(n1030) );
  AND U1399 ( .A(n1031), .B(n1032), .Z(n1029) );
  NAND U1400 ( .A(n743), .B(mix_col_out[48]), .Z(n1032) );
  NAND U1401 ( .A(n744), .B(shift_row_out[48]), .Z(n1031) );
  XOR U1402 ( .A(n1033), .B(key[47]), .Z(o[47]) );
  NAND U1403 ( .A(n1034), .B(n1035), .Z(n1033) );
  NANDN U1404 ( .B(\b/n711 ), .A(n740), .Z(n1035) );
  AND U1405 ( .A(n1036), .B(n1037), .Z(n1034) );
  NAND U1406 ( .A(n743), .B(mix_col_out[47]), .Z(n1037) );
  NANDN U1407 ( .B(n1038), .A(n744), .Z(n1036) );
  XOR U1408 ( .A(n1039), .B(key[46]), .Z(o[46]) );
  NAND U1409 ( .A(n1040), .B(n1041), .Z(n1039) );
  NAND U1410 ( .A(n740), .B(msg[46]), .Z(n1041) );
  AND U1411 ( .A(n1042), .B(n1043), .Z(n1040) );
  NAND U1412 ( .A(n743), .B(mix_col_out[46]), .Z(n1043) );
  NAND U1413 ( .A(n744), .B(shift_row_out[46]), .Z(n1042) );
  XOR U1414 ( .A(n1044), .B(key[45]), .Z(o[45]) );
  NAND U1415 ( .A(n1045), .B(n1046), .Z(n1044) );
  NAND U1416 ( .A(n740), .B(msg[45]), .Z(n1046) );
  AND U1417 ( .A(n1047), .B(n1048), .Z(n1045) );
  NAND U1418 ( .A(n743), .B(mix_col_out[45]), .Z(n1048) );
  NAND U1419 ( .A(n744), .B(shift_row_out[45]), .Z(n1047) );
  XOR U1420 ( .A(n1049), .B(key[44]), .Z(o[44]) );
  NAND U1421 ( .A(n1050), .B(n1051), .Z(n1049) );
  NANDN U1422 ( .B(\b/n733 ), .A(n740), .Z(n1051) );
  AND U1423 ( .A(n1052), .B(n1053), .Z(n1050) );
  NANDN U1424 ( .B(\d/n438 ), .A(n743), .Z(n1053) );
  NAND U1425 ( .A(n744), .B(shift_row_out[44]), .Z(n1052) );
  XOR U1426 ( .A(n1054), .B(key[43]), .Z(o[43]) );
  NAND U1427 ( .A(n1055), .B(n1056), .Z(n1054) );
  NANDN U1428 ( .B(\b/n775 ), .A(n740), .Z(n1056) );
  AND U1429 ( .A(n1057), .B(n1058), .Z(n1055) );
  NANDN U1430 ( .B(\d/n437 ), .A(n743), .Z(n1058) );
  NAND U1431 ( .A(n744), .B(shift_row_out[43]), .Z(n1057) );
  XOR U1432 ( .A(n1059), .B(key[42]), .Z(o[42]) );
  NAND U1433 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U1434 ( .A(n740), .B(msg[42]), .Z(n1061) );
  AND U1435 ( .A(n1062), .B(n1063), .Z(n1060) );
  NAND U1436 ( .A(n743), .B(mix_col_out[42]), .Z(n1063) );
  NAND U1437 ( .A(n744), .B(shift_row_out[42]), .Z(n1062) );
  XOR U1438 ( .A(n1064), .B(key[41]), .Z(o[41]) );
  NAND U1439 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U1440 ( .B(\b/n780 ), .A(n740), .Z(n1066) );
  AND U1441 ( .A(n1067), .B(n1068), .Z(n1065) );
  NANDN U1442 ( .B(\d/n436 ), .A(n743), .Z(n1068) );
  NAND U1443 ( .A(n744), .B(shift_row_out[41]), .Z(n1067) );
  XOR U1444 ( .A(n1069), .B(key[40]), .Z(o[40]) );
  NAND U1445 ( .A(n1070), .B(n1071), .Z(n1069) );
  NAND U1446 ( .A(n740), .B(msg[40]), .Z(n1071) );
  AND U1447 ( .A(n1072), .B(n1073), .Z(n1070) );
  NAND U1448 ( .A(n743), .B(mix_col_out[40]), .Z(n1073) );
  NAND U1449 ( .A(n744), .B(shift_row_out[40]), .Z(n1072) );
  XOR U1450 ( .A(n1074), .B(key[3]), .Z(o[3]) );
  NAND U1451 ( .A(n1075), .B(n1076), .Z(n1074) );
  NANDN U1452 ( .B(\b/n1129 ), .A(n740), .Z(n1076) );
  AND U1453 ( .A(n1077), .B(n1078), .Z(n1075) );
  NANDN U1454 ( .B(\d/n422 ), .A(n743), .Z(n1078) );
  NAND U1455 ( .A(n744), .B(shift_row_out[3]), .Z(n1077) );
  XOR U1456 ( .A(n1079), .B(key[39]), .Z(o[39]) );
  NAND U1457 ( .A(n1080), .B(n1081), .Z(n1079) );
  NANDN U1458 ( .B(\b/n782 ), .A(n740), .Z(n1081) );
  AND U1459 ( .A(n1082), .B(n1083), .Z(n1080) );
  NAND U1460 ( .A(n743), .B(mix_col_out[39]), .Z(n1083) );
  NAND U1461 ( .A(n744), .B(shift_row_out[39]), .Z(n1082) );
  XOR U1462 ( .A(n1084), .B(key[38]), .Z(o[38]) );
  NAND U1463 ( .A(n1085), .B(n1086), .Z(n1084) );
  NAND U1464 ( .A(n740), .B(msg[38]), .Z(n1086) );
  AND U1465 ( .A(n1087), .B(n1088), .Z(n1085) );
  NAND U1466 ( .A(n743), .B(mix_col_out[38]), .Z(n1088) );
  NAND U1467 ( .A(n744), .B(shift_row_out[38]), .Z(n1087) );
  XOR U1468 ( .A(n1089), .B(key[37]), .Z(o[37]) );
  NAND U1469 ( .A(n1090), .B(n1091), .Z(n1089) );
  NAND U1470 ( .A(n740), .B(msg[37]), .Z(n1091) );
  AND U1471 ( .A(n1092), .B(n1093), .Z(n1090) );
  NAND U1472 ( .A(n743), .B(mix_col_out[37]), .Z(n1093) );
  NAND U1473 ( .A(n744), .B(shift_row_out[37]), .Z(n1092) );
  XOR U1474 ( .A(n1094), .B(key[36]), .Z(o[36]) );
  NAND U1475 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1476 ( .B(\b/n804 ), .A(n740), .Z(n1096) );
  AND U1477 ( .A(n1097), .B(n1098), .Z(n1095) );
  NANDN U1478 ( .B(\d/n435 ), .A(n743), .Z(n1098) );
  NAND U1479 ( .A(n744), .B(shift_row_out[36]), .Z(n1097) );
  XOR U1480 ( .A(n1099), .B(key[35]), .Z(o[35]) );
  NAND U1481 ( .A(n1100), .B(n1101), .Z(n1099) );
  NANDN U1482 ( .B(\b/n846 ), .A(n740), .Z(n1101) );
  AND U1483 ( .A(n1102), .B(n1103), .Z(n1100) );
  NANDN U1484 ( .B(\d/n434 ), .A(n743), .Z(n1103) );
  NAND U1485 ( .A(shift_row_out[35]), .B(n744), .Z(n1102) );
  XOR U1486 ( .A(n1104), .B(key[34]), .Z(o[34]) );
  NAND U1487 ( .A(n1105), .B(n1106), .Z(n1104) );
  NAND U1488 ( .A(n740), .B(msg[34]), .Z(n1106) );
  AND U1489 ( .A(n1107), .B(n1108), .Z(n1105) );
  NAND U1490 ( .A(n743), .B(mix_col_out[34]), .Z(n1108) );
  NAND U1491 ( .A(shift_row_out[34]), .B(n744), .Z(n1107) );
  XOR U1492 ( .A(n1109), .B(key[33]), .Z(o[33]) );
  NAND U1493 ( .A(n1110), .B(n1111), .Z(n1109) );
  NANDN U1494 ( .B(\b/n851 ), .A(n740), .Z(n1111) );
  AND U1495 ( .A(n1112), .B(n1113), .Z(n1110) );
  NANDN U1496 ( .B(\d/n433 ), .A(n743), .Z(n1113) );
  NAND U1497 ( .A(n744), .B(shift_row_out[33]), .Z(n1112) );
  XOR U1498 ( .A(n1114), .B(key[32]), .Z(o[32]) );
  NAND U1499 ( .A(n1115), .B(n1116), .Z(n1114) );
  NAND U1500 ( .A(n740), .B(msg[32]), .Z(n1116) );
  AND U1501 ( .A(n1117), .B(n1118), .Z(n1115) );
  NAND U1502 ( .A(n743), .B(mix_col_out[32]), .Z(n1118) );
  NAND U1503 ( .A(shift_row_out[32]), .B(n744), .Z(n1117) );
  XOR U1504 ( .A(n1119), .B(key[31]), .Z(o[31]) );
  NAND U1505 ( .A(n1120), .B(n1121), .Z(n1119) );
  NANDN U1506 ( .B(\b/n853 ), .A(n740), .Z(n1121) );
  AND U1507 ( .A(n1122), .B(n1123), .Z(n1120) );
  NAND U1508 ( .A(n743), .B(mix_col_out[31]), .Z(n1123) );
  NANDN U1509 ( .B(n1124), .A(n744), .Z(n1122) );
  XOR U1510 ( .A(n1125), .B(key[30]), .Z(o[30]) );
  NAND U1511 ( .A(n1126), .B(n1127), .Z(n1125) );
  NAND U1512 ( .A(n740), .B(msg[30]), .Z(n1127) );
  AND U1513 ( .A(n1128), .B(n1129), .Z(n1126) );
  NAND U1514 ( .A(n743), .B(mix_col_out[30]), .Z(n1129) );
  NAND U1515 ( .A(n744), .B(shift_row_out[30]), .Z(n1128) );
  XOR U1516 ( .A(n1130), .B(key[2]), .Z(o[2]) );
  NAND U1517 ( .A(n1131), .B(n1132), .Z(n1130) );
  NAND U1518 ( .A(n740), .B(msg[2]), .Z(n1132) );
  AND U1519 ( .A(n1133), .B(n1134), .Z(n1131) );
  NAND U1520 ( .A(n743), .B(mix_col_out[2]), .Z(n1134) );
  NAND U1521 ( .A(n744), .B(shift_row_out[2]), .Z(n1133) );
  XOR U1522 ( .A(n1135), .B(key[29]), .Z(o[29]) );
  NAND U1523 ( .A(n1136), .B(n1137), .Z(n1135) );
  NAND U1524 ( .A(n740), .B(msg[29]), .Z(n1137) );
  AND U1525 ( .A(n1138), .B(n1139), .Z(n1136) );
  NAND U1526 ( .A(n743), .B(mix_col_out[29]), .Z(n1139) );
  NAND U1527 ( .A(n744), .B(shift_row_out[29]), .Z(n1138) );
  XOR U1528 ( .A(n1140), .B(key[28]), .Z(o[28]) );
  NAND U1529 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1530 ( .B(\b/n875 ), .A(n740), .Z(n1142) );
  AND U1531 ( .A(n1143), .B(n1144), .Z(n1141) );
  NANDN U1532 ( .B(\d/n432 ), .A(n743), .Z(n1144) );
  NAND U1533 ( .A(n744), .B(shift_row_out[28]), .Z(n1143) );
  XOR U1534 ( .A(n1145), .B(key[27]), .Z(o[27]) );
  NAND U1535 ( .A(n1146), .B(n1147), .Z(n1145) );
  NANDN U1536 ( .B(\b/n917 ), .A(n740), .Z(n1147) );
  AND U1537 ( .A(n1148), .B(n1149), .Z(n1146) );
  NANDN U1538 ( .B(\d/n431 ), .A(n743), .Z(n1149) );
  NAND U1539 ( .A(n744), .B(shift_row_out[27]), .Z(n1148) );
  XOR U1540 ( .A(n1150), .B(key[26]), .Z(o[26]) );
  NAND U1541 ( .A(n1151), .B(n1152), .Z(n1150) );
  NAND U1542 ( .A(n740), .B(msg[26]), .Z(n1152) );
  AND U1543 ( .A(n1153), .B(n1154), .Z(n1151) );
  NAND U1544 ( .A(n743), .B(mix_col_out[26]), .Z(n1154) );
  NAND U1545 ( .A(n744), .B(shift_row_out[26]), .Z(n1153) );
  XOR U1546 ( .A(n1155), .B(key[25]), .Z(o[25]) );
  NAND U1547 ( .A(n1156), .B(n1157), .Z(n1155) );
  NANDN U1548 ( .B(\b/n922 ), .A(n740), .Z(n1157) );
  AND U1549 ( .A(n1158), .B(n1159), .Z(n1156) );
  NANDN U1550 ( .B(\d/n430 ), .A(n743), .Z(n1159) );
  NAND U1551 ( .A(n744), .B(shift_row_out[25]), .Z(n1158) );
  XOR U1552 ( .A(n1160), .B(key[24]), .Z(o[24]) );
  NAND U1553 ( .A(n1161), .B(n1162), .Z(n1160) );
  NAND U1554 ( .A(n740), .B(msg[24]), .Z(n1162) );
  AND U1555 ( .A(n1163), .B(n1164), .Z(n1161) );
  NAND U1556 ( .A(n743), .B(mix_col_out[24]), .Z(n1164) );
  NAND U1557 ( .A(n744), .B(shift_row_out[24]), .Z(n1163) );
  XOR U1558 ( .A(n1165), .B(key[23]), .Z(o[23]) );
  NAND U1559 ( .A(n1166), .B(n1167), .Z(n1165) );
  NANDN U1560 ( .B(\b/n924 ), .A(n740), .Z(n1167) );
  AND U1561 ( .A(n1168), .B(n1169), .Z(n1166) );
  NAND U1562 ( .A(n743), .B(mix_col_out[23]), .Z(n1169) );
  NANDN U1563 ( .B(n1170), .A(n744), .Z(n1168) );
  XOR U1564 ( .A(n1171), .B(key[22]), .Z(o[22]) );
  NAND U1565 ( .A(n1172), .B(n1173), .Z(n1171) );
  NAND U1566 ( .A(n740), .B(msg[22]), .Z(n1173) );
  AND U1567 ( .A(n1174), .B(n1175), .Z(n1172) );
  NAND U1568 ( .A(n743), .B(mix_col_out[22]), .Z(n1175) );
  NAND U1569 ( .A(n744), .B(shift_row_out[22]), .Z(n1174) );
  XOR U1570 ( .A(n1176), .B(key[21]), .Z(o[21]) );
  NAND U1571 ( .A(n1177), .B(n1178), .Z(n1176) );
  NAND U1572 ( .A(n740), .B(msg[21]), .Z(n1178) );
  AND U1573 ( .A(n1179), .B(n1180), .Z(n1177) );
  NAND U1574 ( .A(n743), .B(mix_col_out[21]), .Z(n1180) );
  NAND U1575 ( .A(n744), .B(shift_row_out[21]), .Z(n1179) );
  XOR U1576 ( .A(n1181), .B(key[20]), .Z(o[20]) );
  NAND U1577 ( .A(n1182), .B(n1183), .Z(n1181) );
  NANDN U1578 ( .B(\b/n946 ), .A(n740), .Z(n1183) );
  AND U1579 ( .A(n1184), .B(n1185), .Z(n1182) );
  NANDN U1580 ( .B(\d/n429 ), .A(n743), .Z(n1185) );
  NAND U1581 ( .A(n744), .B(shift_row_out[20]), .Z(n1184) );
  XOR U1582 ( .A(n1186), .B(key[1]), .Z(o[1]) );
  NAND U1583 ( .A(n1187), .B(n1188), .Z(n1186) );
  NANDN U1584 ( .B(\b/n1134 ), .A(n740), .Z(n1188) );
  AND U1585 ( .A(n1189), .B(n1190), .Z(n1187) );
  NANDN U1586 ( .B(\d/n421 ), .A(n743), .Z(n1190) );
  NAND U1587 ( .A(n744), .B(shift_row_out[1]), .Z(n1189) );
  XOR U1588 ( .A(n1191), .B(key[19]), .Z(o[19]) );
  NAND U1589 ( .A(n1192), .B(n1193), .Z(n1191) );
  NANDN U1590 ( .B(\b/n988 ), .A(n740), .Z(n1193) );
  AND U1591 ( .A(n1194), .B(n1195), .Z(n1192) );
  NANDN U1592 ( .B(\d/n428 ), .A(n743), .Z(n1195) );
  NAND U1593 ( .A(n744), .B(shift_row_out[19]), .Z(n1194) );
  XOR U1594 ( .A(n1196), .B(key[18]), .Z(o[18]) );
  NAND U1595 ( .A(n1197), .B(n1198), .Z(n1196) );
  NAND U1596 ( .A(n740), .B(msg[18]), .Z(n1198) );
  AND U1597 ( .A(n1199), .B(n1200), .Z(n1197) );
  NAND U1598 ( .A(n743), .B(mix_col_out[18]), .Z(n1200) );
  NAND U1599 ( .A(n744), .B(shift_row_out[18]), .Z(n1199) );
  XOR U1600 ( .A(n1201), .B(key[17]), .Z(o[17]) );
  NAND U1601 ( .A(n1202), .B(n1203), .Z(n1201) );
  NANDN U1602 ( .B(\b/n993 ), .A(n740), .Z(n1203) );
  AND U1603 ( .A(n1204), .B(n1205), .Z(n1202) );
  NANDN U1604 ( .B(\d/n427 ), .A(n743), .Z(n1205) );
  NAND U1605 ( .A(n744), .B(shift_row_out[17]), .Z(n1204) );
  XOR U1606 ( .A(n1206), .B(key[16]), .Z(o[16]) );
  NAND U1607 ( .A(n1207), .B(n1208), .Z(n1206) );
  NAND U1608 ( .A(n740), .B(msg[16]), .Z(n1208) );
  AND U1609 ( .A(n1209), .B(n1210), .Z(n1207) );
  NAND U1610 ( .A(n743), .B(mix_col_out[16]), .Z(n1210) );
  NAND U1611 ( .A(shift_row_out[16]), .B(n744), .Z(n1209) );
  XOR U1612 ( .A(n1211), .B(key[15]), .Z(o[15]) );
  NAND U1613 ( .A(n1212), .B(n1213), .Z(n1211) );
  NAND U1614 ( .A(n740), .B(msg[15]), .Z(n1213) );
  AND U1615 ( .A(n1214), .B(n1215), .Z(n1212) );
  NAND U1616 ( .A(n743), .B(mix_col_out[15]), .Z(n1215) );
  NAND U1617 ( .A(n744), .B(shift_row_out[15]), .Z(n1214) );
  XOR U1618 ( .A(n1216), .B(key[14]), .Z(o[14]) );
  NAND U1619 ( .A(n1217), .B(n1218), .Z(n1216) );
  NAND U1620 ( .A(n740), .B(msg[14]), .Z(n1218) );
  AND U1621 ( .A(n1219), .B(n1220), .Z(n1217) );
  NAND U1622 ( .A(n743), .B(mix_col_out[14]), .Z(n1220) );
  NAND U1623 ( .A(n744), .B(shift_row_out[14]), .Z(n1219) );
  XOR U1624 ( .A(n1221), .B(key[13]), .Z(o[13]) );
  NAND U1625 ( .A(n1222), .B(n1223), .Z(n1221) );
  NAND U1626 ( .A(n740), .B(msg[13]), .Z(n1223) );
  AND U1627 ( .A(n1224), .B(n1225), .Z(n1222) );
  NAND U1628 ( .A(n743), .B(mix_col_out[13]), .Z(n1225) );
  NAND U1629 ( .A(n744), .B(shift_row_out[13]), .Z(n1224) );
  XOR U1630 ( .A(n1226), .B(key[12]), .Z(o[12]) );
  NAND U1631 ( .A(n1227), .B(n1228), .Z(n1226) );
  NANDN U1632 ( .B(\b/n1015 ), .A(n740), .Z(n1228) );
  AND U1633 ( .A(n1229), .B(n1230), .Z(n1227) );
  NANDN U1634 ( .B(\d/n426 ), .A(n743), .Z(n1230) );
  NAND U1635 ( .A(n744), .B(shift_row_out[12]), .Z(n1229) );
  XNOR U1636 ( .A(n1231), .B(n1529), .Z(o[127]) );
  NAND U1637 ( .A(n1232), .B(n1233), .Z(n1231) );
  NANDN U1638 ( .B(\b/n2 ), .A(n740), .Z(n1233) );
  AND U1639 ( .A(n1234), .B(n1235), .Z(n1232) );
  NAND U1640 ( .A(n743), .B(mix_col_out[127]), .Z(n1235) );
  NAND U1641 ( .A(n744), .B(shift_row_out[127]), .Z(n1234) );
  XOR U1642 ( .A(n1236), .B(key[126]), .Z(o[126]) );
  NAND U1643 ( .A(n1237), .B(n1238), .Z(n1236) );
  NAND U1644 ( .A(n740), .B(msg[126]), .Z(n1238) );
  AND U1645 ( .A(n1239), .B(n1240), .Z(n1237) );
  NAND U1646 ( .A(n743), .B(mix_col_out[126]), .Z(n1240) );
  NAND U1647 ( .A(n744), .B(shift_row_out[126]), .Z(n1239) );
  XOR U1648 ( .A(n1241), .B(key[125]), .Z(o[125]) );
  NAND U1649 ( .A(n1242), .B(n1243), .Z(n1241) );
  NAND U1650 ( .A(n740), .B(msg[125]), .Z(n1243) );
  AND U1651 ( .A(n1244), .B(n1245), .Z(n1242) );
  NAND U1652 ( .A(n743), .B(mix_col_out[125]), .Z(n1245) );
  NAND U1653 ( .A(n744), .B(shift_row_out[125]), .Z(n1244) );
  XNOR U1654 ( .A(n1246), .B(n1546), .Z(o[124]) );
  NAND U1655 ( .A(n1247), .B(n1248), .Z(n1246) );
  NANDN U1656 ( .B(\b/n24 ), .A(n740), .Z(n1248) );
  AND U1657 ( .A(n1249), .B(n1250), .Z(n1247) );
  NANDN U1658 ( .B(\d/n468 ), .A(n743), .Z(n1250) );
  NAND U1659 ( .A(n744), .B(shift_row_out[124]), .Z(n1249) );
  XNOR U1660 ( .A(n1251), .B(n1580), .Z(o[123]) );
  NAND U1661 ( .A(n1252), .B(n1253), .Z(n1251) );
  NANDN U1662 ( .B(\b/n66 ), .A(n740), .Z(n1253) );
  AND U1663 ( .A(n1254), .B(n1255), .Z(n1252) );
  NANDN U1664 ( .B(\d/n467 ), .A(n743), .Z(n1255) );
  NAND U1665 ( .A(n744), .B(shift_row_out[123]), .Z(n1254) );
  XOR U1666 ( .A(n1256), .B(key[122]), .Z(o[122]) );
  NAND U1667 ( .A(n1257), .B(n1258), .Z(n1256) );
  NAND U1668 ( .A(n740), .B(msg[122]), .Z(n1258) );
  AND U1669 ( .A(n1259), .B(n1260), .Z(n1257) );
  NAND U1670 ( .A(n743), .B(mix_col_out[122]), .Z(n1260) );
  NAND U1671 ( .A(n744), .B(shift_row_out[122]), .Z(n1259) );
  XNOR U1672 ( .A(n1261), .B(n1584), .Z(o[121]) );
  NAND U1673 ( .A(n1262), .B(n1263), .Z(n1261) );
  NANDN U1674 ( .B(\b/n71 ), .A(n740), .Z(n1263) );
  AND U1675 ( .A(n1264), .B(n1265), .Z(n1262) );
  NANDN U1676 ( .B(\d/n466 ), .A(n743), .Z(n1265) );
  NAND U1677 ( .A(n744), .B(shift_row_out[121]), .Z(n1264) );
  XOR U1678 ( .A(n1266), .B(key[120]), .Z(o[120]) );
  NAND U1679 ( .A(n1267), .B(n1268), .Z(n1266) );
  NAND U1680 ( .A(n740), .B(msg[120]), .Z(n1268) );
  AND U1681 ( .A(n1269), .B(n1270), .Z(n1267) );
  NAND U1682 ( .A(n743), .B(mix_col_out[120]), .Z(n1270) );
  NAND U1683 ( .A(n744), .B(shift_row_out[120]), .Z(n1269) );
  XOR U1684 ( .A(n1271), .B(key[11]), .Z(o[11]) );
  NAND U1685 ( .A(n1272), .B(n1273), .Z(n1271) );
  NANDN U1686 ( .B(\b/n1058 ), .A(n740), .Z(n1273) );
  AND U1687 ( .A(n1274), .B(n1275), .Z(n1272) );
  NANDN U1688 ( .B(\d/n425 ), .A(n743), .Z(n1275) );
  NAND U1689 ( .A(shift_row_out[11]), .B(n744), .Z(n1274) );
  XNOR U1690 ( .A(n1276), .B(n1585), .Z(o[119]) );
  NAND U1691 ( .A(n1277), .B(n1278), .Z(n1276) );
  NANDN U1692 ( .B(\b/n73 ), .A(n740), .Z(n1278) );
  AND U1693 ( .A(n1279), .B(n1280), .Z(n1277) );
  NAND U1694 ( .A(n743), .B(mix_col_out[119]), .Z(n1280) );
  NANDN U1695 ( .B(n1281), .A(n744), .Z(n1279) );
  XOR U1696 ( .A(n1282), .B(key[118]), .Z(o[118]) );
  NAND U1697 ( .A(n1283), .B(n1284), .Z(n1282) );
  NAND U1698 ( .A(n740), .B(msg[118]), .Z(n1284) );
  AND U1699 ( .A(n1285), .B(n1286), .Z(n1283) );
  NAND U1700 ( .A(n743), .B(mix_col_out[118]), .Z(n1286) );
  NAND U1701 ( .A(n744), .B(shift_row_out[118]), .Z(n1285) );
  XOR U1702 ( .A(n1287), .B(key[117]), .Z(o[117]) );
  NAND U1703 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1704 ( .A(n740), .B(msg[117]), .Z(n1289) );
  AND U1705 ( .A(n1290), .B(n1291), .Z(n1288) );
  NAND U1706 ( .A(n743), .B(mix_col_out[117]), .Z(n1291) );
  NAND U1707 ( .A(n744), .B(shift_row_out[117]), .Z(n1290) );
  XNOR U1708 ( .A(n1292), .B(n1602), .Z(o[116]) );
  NAND U1709 ( .A(n1293), .B(n1294), .Z(n1292) );
  NANDN U1710 ( .B(\b/n95 ), .A(n740), .Z(n1294) );
  AND U1711 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1712 ( .B(\d/n465 ), .A(n743), .Z(n1296) );
  NAND U1713 ( .A(n744), .B(shift_row_out[116]), .Z(n1295) );
  XNOR U1714 ( .A(n1297), .B(n1636), .Z(o[115]) );
  NAND U1715 ( .A(n1298), .B(n1299), .Z(n1297) );
  NANDN U1716 ( .B(\b/n137 ), .A(n740), .Z(n1299) );
  AND U1717 ( .A(n1300), .B(n1301), .Z(n1298) );
  NANDN U1718 ( .B(\d/n464 ), .A(n743), .Z(n1301) );
  NAND U1719 ( .A(n744), .B(shift_row_out[115]), .Z(n1300) );
  XOR U1720 ( .A(n1302), .B(key[114]), .Z(o[114]) );
  NAND U1721 ( .A(n1303), .B(n1304), .Z(n1302) );
  NAND U1722 ( .A(n740), .B(msg[114]), .Z(n1304) );
  AND U1723 ( .A(n1305), .B(n1306), .Z(n1303) );
  NAND U1724 ( .A(n743), .B(mix_col_out[114]), .Z(n1306) );
  NAND U1725 ( .A(n744), .B(shift_row_out[114]), .Z(n1305) );
  XNOR U1726 ( .A(n1307), .B(n1640), .Z(o[113]) );
  NAND U1727 ( .A(n1308), .B(n1309), .Z(n1307) );
  NANDN U1728 ( .B(\b/n142 ), .A(n740), .Z(n1309) );
  AND U1729 ( .A(n1310), .B(n1311), .Z(n1308) );
  NANDN U1730 ( .B(\d/n463 ), .A(n743), .Z(n1311) );
  NAND U1731 ( .A(n744), .B(shift_row_out[113]), .Z(n1310) );
  XOR U1732 ( .A(n1312), .B(key[112]), .Z(o[112]) );
  NAND U1733 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1734 ( .A(n740), .B(msg[112]), .Z(n1314) );
  AND U1735 ( .A(n1315), .B(n1316), .Z(n1313) );
  NAND U1736 ( .A(n743), .B(mix_col_out[112]), .Z(n1316) );
  NAND U1737 ( .A(n744), .B(shift_row_out[112]), .Z(n1315) );
  XOR U1738 ( .A(n1317), .B(key[111]), .Z(o[111]) );
  NAND U1739 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1740 ( .B(\b/n144 ), .A(n740), .Z(n1319) );
  AND U1741 ( .A(n1320), .B(n1321), .Z(n1318) );
  NAND U1742 ( .A(n743), .B(mix_col_out[111]), .Z(n1321) );
  NANDN U1743 ( .B(n1322), .A(n744), .Z(n1320) );
  XOR U1744 ( .A(n1323), .B(key[110]), .Z(o[110]) );
  NAND U1745 ( .A(n1324), .B(n1325), .Z(n1323) );
  NAND U1746 ( .A(n740), .B(msg[110]), .Z(n1325) );
  AND U1747 ( .A(n1326), .B(n1327), .Z(n1324) );
  NAND U1748 ( .A(n743), .B(mix_col_out[110]), .Z(n1327) );
  NAND U1749 ( .A(n744), .B(shift_row_out[110]), .Z(n1326) );
  XOR U1750 ( .A(n1328), .B(key[10]), .Z(o[10]) );
  NAND U1751 ( .A(n1329), .B(n1330), .Z(n1328) );
  NAND U1752 ( .A(n740), .B(msg[10]), .Z(n1330) );
  AND U1753 ( .A(n1331), .B(n1332), .Z(n1329) );
  NAND U1754 ( .A(n743), .B(mix_col_out[10]), .Z(n1332) );
  NAND U1755 ( .A(shift_row_out[10]), .B(n744), .Z(n1331) );
  XOR U1756 ( .A(n1333), .B(key[109]), .Z(o[109]) );
  NAND U1757 ( .A(n1334), .B(n1335), .Z(n1333) );
  NAND U1758 ( .A(n740), .B(msg[109]), .Z(n1335) );
  AND U1759 ( .A(n1336), .B(n1337), .Z(n1334) );
  NAND U1760 ( .A(n743), .B(mix_col_out[109]), .Z(n1337) );
  NAND U1761 ( .A(n744), .B(shift_row_out[109]), .Z(n1336) );
  XNOR U1762 ( .A(n1338), .B(n1646), .Z(o[108]) );
  NAND U1763 ( .A(n1339), .B(n1340), .Z(n1338) );
  NANDN U1764 ( .B(\b/n166 ), .A(n740), .Z(n1340) );
  AND U1765 ( .A(n1341), .B(n1342), .Z(n1339) );
  NANDN U1766 ( .B(\d/n462 ), .A(n743), .Z(n1342) );
  NAND U1767 ( .A(n744), .B(shift_row_out[108]), .Z(n1341) );
  XNOR U1768 ( .A(n1343), .B(n1691), .Z(o[107]) );
  NAND U1769 ( .A(n1344), .B(n1345), .Z(n1343) );
  NANDN U1770 ( .B(\b/n208 ), .A(n740), .Z(n1345) );
  AND U1771 ( .A(n1346), .B(n1347), .Z(n1344) );
  NANDN U1772 ( .B(\d/n461 ), .A(n743), .Z(n1347) );
  NAND U1773 ( .A(shift_row_out[107]), .B(n744), .Z(n1346) );
  XOR U1774 ( .A(n1348), .B(key[106]), .Z(o[106]) );
  NAND U1775 ( .A(n1349), .B(n1350), .Z(n1348) );
  NAND U1776 ( .A(n740), .B(msg[106]), .Z(n1350) );
  AND U1777 ( .A(n1351), .B(n1352), .Z(n1349) );
  NAND U1778 ( .A(n743), .B(mix_col_out[106]), .Z(n1352) );
  NAND U1779 ( .A(shift_row_out[106]), .B(n744), .Z(n1351) );
  XNOR U1780 ( .A(n1353), .B(n1695), .Z(o[105]) );
  NAND U1781 ( .A(n1354), .B(n1355), .Z(n1353) );
  NANDN U1782 ( .B(\b/n213 ), .A(n740), .Z(n1355) );
  AND U1783 ( .A(n1356), .B(n1357), .Z(n1354) );
  NANDN U1784 ( .B(\d/n460 ), .A(n743), .Z(n1357) );
  NAND U1785 ( .A(n744), .B(shift_row_out[105]), .Z(n1356) );
  XOR U1786 ( .A(n1358), .B(key[104]), .Z(o[104]) );
  NAND U1787 ( .A(n1359), .B(n1360), .Z(n1358) );
  NAND U1788 ( .A(n740), .B(msg[104]), .Z(n1360) );
  AND U1789 ( .A(n1361), .B(n1362), .Z(n1359) );
  NAND U1790 ( .A(n743), .B(mix_col_out[104]), .Z(n1362) );
  NAND U1791 ( .A(shift_row_out[104]), .B(n744), .Z(n1361) );
  XNOR U1792 ( .A(n1363), .B(n1473), .Z(o[103]) );
  NAND U1793 ( .A(n1364), .B(n1365), .Z(n1363) );
  NAND U1794 ( .A(n740), .B(msg[103]), .Z(n1365) );
  AND U1795 ( .A(n1366), .B(n1367), .Z(n1364) );
  NAND U1796 ( .A(n743), .B(mix_col_out[103]), .Z(n1367) );
  NAND U1797 ( .A(n744), .B(shift_row_out[103]), .Z(n1366) );
  XOR U1798 ( .A(n1368), .B(key[102]), .Z(o[102]) );
  NAND U1799 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1800 ( .A(n740), .B(msg[102]), .Z(n1370) );
  AND U1801 ( .A(n1371), .B(n1372), .Z(n1369) );
  NAND U1802 ( .A(n743), .B(mix_col_out[102]), .Z(n1372) );
  NAND U1803 ( .A(n744), .B(shift_row_out[102]), .Z(n1371) );
  XOR U1804 ( .A(n1373), .B(key[101]), .Z(o[101]) );
  NAND U1805 ( .A(n1374), .B(n1375), .Z(n1373) );
  NAND U1806 ( .A(n740), .B(msg[101]), .Z(n1375) );
  AND U1807 ( .A(n1376), .B(n1377), .Z(n1374) );
  NAND U1808 ( .A(n743), .B(mix_col_out[101]), .Z(n1377) );
  NAND U1809 ( .A(n744), .B(shift_row_out[101]), .Z(n1376) );
  XNOR U1810 ( .A(n1378), .B(n1490), .Z(o[100]) );
  NAND U1811 ( .A(n1379), .B(n1380), .Z(n1378) );
  NANDN U1812 ( .B(\b/n220 ), .A(n740), .Z(n1380) );
  AND U1813 ( .A(n1381), .B(n1382), .Z(n1379) );
  NANDN U1814 ( .B(\d/n459 ), .A(n743), .Z(n1382) );
  NAND U1815 ( .A(n744), .B(shift_row_out[100]), .Z(n1381) );
  XOR U1816 ( .A(n1383), .B(key[0]), .Z(o[0]) );
  NAND U1817 ( .A(n1384), .B(n1385), .Z(n1383) );
  NAND U1818 ( .A(n740), .B(msg[0]), .Z(n1385) );
  AND U1819 ( .A(n1386), .B(n1387), .Z(n1384) );
  NAND U1820 ( .A(n743), .B(mix_col_out[0]), .Z(n1387) );
  NOR U1821 ( .A(n740), .B(n744), .Z(n743) );
  AND U1822 ( .A(n1388), .B(n1389), .Z(n740) );
  ANDN U1823 ( .A(n1390), .B(counter[3]), .Z(n1389) );
  NAND U1824 ( .A(shift_row_out[0]), .B(n744), .Z(n1386) );
  AND U1825 ( .A(n1391), .B(counter[3]), .Z(n744) );
  XOR U1826 ( .A(key[9]), .B(\e/t[9] ), .Z(nextKey[9]) );
  XOR U1827 ( .A(key[8]), .B(\e/t[8] ), .Z(nextKey[8]) );
  IV U1828 ( .A(\e/n102 ), .Z(nextKey[7]) );
  IV U1829 ( .A(\e/n118 ), .Z(nextKey[71]) );
  IV U1830 ( .A(\e/n117 ), .Z(nextKey[70]) );
  IV U1831 ( .A(\e/n101 ), .Z(nextKey[6]) );
  IV U1832 ( .A(\e/n116 ), .Z(nextKey[69]) );
  IV U1833 ( .A(\e/n115 ), .Z(nextKey[68]) );
  IV U1834 ( .A(\e/n114 ), .Z(nextKey[67]) );
  IV U1835 ( .A(\e/n113 ), .Z(nextKey[66]) );
  IV U1836 ( .A(\e/n112 ), .Z(nextKey[65]) );
  IV U1837 ( .A(\e/n111 ), .Z(nextKey[64]) );
  IV U1838 ( .A(\e/n100 ), .Z(nextKey[5]) );
  IV U1839 ( .A(\e/n99 ), .Z(nextKey[4]) );
  IV U1840 ( .A(\e/n98 ), .Z(nextKey[3]) );
  IV U1841 ( .A(\e/n110 ), .Z(nextKey[39]) );
  IV U1842 ( .A(\e/n109 ), .Z(nextKey[38]) );
  IV U1843 ( .A(\e/n108 ), .Z(nextKey[37]) );
  IV U1844 ( .A(\e/n107 ), .Z(nextKey[36]) );
  IV U1845 ( .A(\e/n106 ), .Z(nextKey[35]) );
  IV U1846 ( .A(\e/n105 ), .Z(nextKey[34]) );
  IV U1847 ( .A(\e/n104 ), .Z(nextKey[33]) );
  IV U1848 ( .A(\e/n103 ), .Z(nextKey[32]) );
  XOR U1849 ( .A(key[31]), .B(\e/t[31] ), .Z(nextKey[31]) );
  XOR U1850 ( .A(key[30]), .B(\e/t[30] ), .Z(nextKey[30]) );
  IV U1851 ( .A(\e/n97 ), .Z(nextKey[2]) );
  XOR U1852 ( .A(key[29]), .B(\e/t[29] ), .Z(nextKey[29]) );
  XOR U1853 ( .A(key[28]), .B(\e/t[28] ), .Z(nextKey[28]) );
  XOR U1854 ( .A(key[27]), .B(\e/t[27] ), .Z(nextKey[27]) );
  XOR U1855 ( .A(key[26]), .B(\e/t[26] ), .Z(nextKey[26]) );
  XOR U1856 ( .A(key[25]), .B(\e/t[25] ), .Z(nextKey[25]) );
  XOR U1857 ( .A(key[24]), .B(\e/t[24] ), .Z(nextKey[24]) );
  XOR U1858 ( .A(key[23]), .B(\e/t[23] ), .Z(nextKey[23]) );
  XOR U1859 ( .A(key[22]), .B(\e/t[22] ), .Z(nextKey[22]) );
  XOR U1860 ( .A(key[21]), .B(\e/t[21] ), .Z(nextKey[21]) );
  XOR U1861 ( .A(key[20]), .B(\e/t[20] ), .Z(nextKey[20]) );
  IV U1862 ( .A(\e/n96 ), .Z(nextKey[1]) );
  XOR U1863 ( .A(key[19]), .B(\e/t[19] ), .Z(nextKey[19]) );
  XOR U1864 ( .A(key[18]), .B(\e/t[18] ), .Z(nextKey[18]) );
  XOR U1865 ( .A(key[17]), .B(\e/t[17] ), .Z(nextKey[17]) );
  XOR U1866 ( .A(key[16]), .B(\e/t[16] ), .Z(nextKey[16]) );
  XOR U1867 ( .A(key[15]), .B(\e/t[15] ), .Z(nextKey[15]) );
  XOR U1868 ( .A(key[14]), .B(\e/t[14] ), .Z(nextKey[14]) );
  XOR U1869 ( .A(key[13]), .B(\e/t[13] ), .Z(nextKey[13]) );
  XOR U1870 ( .A(key[12]), .B(\e/t[12] ), .Z(nextKey[12]) );
  XOR U1871 ( .A(key[11]), .B(\e/t[11] ), .Z(nextKey[11]) );
  XOR U1872 ( .A(key[10]), .B(\e/t[10] ), .Z(nextKey[10]) );
  IV U1873 ( .A(\e/n95 ), .Z(nextKey[0]) );
  NANDN U1874 ( .B(n1390), .A(n1392), .Z(\e/n94 ) );
  ANDN U1875 ( .A(counter[0]), .B(n1393), .Z(n1392) );
  NANDN U1876 ( .B(n1390), .A(n1394), .Z(\e/n93 ) );
  ANDN U1877 ( .A(n7), .B(n1393), .Z(n1394) );
  AND U1878 ( .A(n1395), .B(n1396), .Z(\e/n92 ) );
  NANDN U1879 ( .B(n7), .A(counter[3]), .Z(n1396) );
  NANDN U1880 ( .B(n1390), .A(n1397), .Z(n1395) );
  ANDN U1881 ( .A(n1393), .B(n7), .Z(n1397) );
  ANDN U1882 ( .A(n1398), .B(n1399), .Z(\e/n91 ) );
  NANDN U1883 ( .B(n1390), .A(n1388), .Z(n1398) );
  ANDN U1884 ( .A(n7), .B(counter[1]), .Z(n1388) );
  NAND U1885 ( .A(n1400), .B(n1401), .Z(\e/n90 ) );
  NOR U1886 ( .A(counter[2]), .B(n1402), .Z(n1401) );
  NAND U1887 ( .A(n1405), .B(n1406), .Z(\e/n89 ) );
  NOR U1888 ( .A(counter[2]), .B(n1403), .Z(n1406) );
  AND U1889 ( .A(counter[3]), .B(counter[1]), .Z(n1403) );
  IV U1890 ( .A(counter[0]), .Z(n7) );
  NOR U1891 ( .A(n1402), .B(n1399), .Z(\e/n88 ) );
  AND U1892 ( .A(counter[3]), .B(n1393), .Z(n1399) );
  ANDN U1893 ( .A(counter[0]), .B(n1391), .Z(n1402) );
  OR U1894 ( .A(n1391), .B(counter[0]), .Z(\e/n87 ) );
  NANDN U1895 ( .B(counter[1]), .A(n1390), .Z(n1391) );
  IV U1896 ( .A(n2422), .Z(n1548) );
  IV U1897 ( .A(key[124]), .Z(n1546) );
  IV U1898 ( .A(n2726), .Z(n1544) );
  IV U1899 ( .A(n2416), .Z(n1543) );
  IV U1900 ( .A(n2412), .Z(n1542) );
  IV U1901 ( .A(n2748), .Z(n1478) );
  IV U1902 ( .A(n2727), .Z(n1541) );
  IV U1903 ( .A(n2730), .Z(n1540) );
  IV U1904 ( .A(n2732), .Z(n1539) );
  IV U1905 ( .A(n2395), .Z(n1538) );
  IV U1906 ( .A(n2531), .Z(n1537) );
  IV U1907 ( .A(n2722), .Z(n1536) );
  IV U1908 ( .A(n2721), .Z(n1535) );
  IV U1909 ( .A(n2401), .Z(n1534) );
  IV U1910 ( .A(n2410), .Z(n1533) );
  IV U1911 ( .A(n2405), .Z(n1532) );
  IV U1912 ( .A(n2396), .Z(n1531) );
  IV U1913 ( .A(n2731), .Z(n1530) );
  IV U1914 ( .A(key[127]), .Z(n1529) );
  IV U1915 ( .A(key[97]), .Z(n1528) );
  IV U1916 ( .A(n2757), .Z(n1477) );
  IV U1917 ( .A(n2774), .Z(n1527) );
  IV U1918 ( .A(n2758), .Z(n1526) );
  IV U1919 ( .A(n2741), .Z(n1525) );
  IV U1920 ( .A(key[99]), .Z(n1524) );
  IV U1921 ( .A(n2768), .Z(n1523) );
  IV U1922 ( .A(n2764), .Z(n1522) );
  IV U1923 ( .A(n2793), .Z(n1521) );
  IV U1924 ( .A(n3075), .Z(n1520) );
  IV U1925 ( .A(n3081), .Z(n1519) );
  IV U1926 ( .A(n2745), .Z(n1518) );
  IV U1927 ( .A(n2752), .Z(n1476) );
  IV U1928 ( .A(n3076), .Z(n1517) );
  IV U1929 ( .A(n2753), .Z(n1516) );
  IV U1930 ( .A(n2744), .Z(n1515) );
  IV U1931 ( .A(n2747), .Z(n1514) );
  IV U1932 ( .A(n2756), .Z(n1513) );
  IV U1933 ( .A(n3070), .Z(n1512) );
  IV U1934 ( .A(n2895), .Z(n1511) );
  IV U1935 ( .A(n2740), .Z(n1510) );
  IV U1936 ( .A(n2772), .Z(n1509) );
  IV U1937 ( .A(n2767), .Z(n1508) );
  IV U1938 ( .A(n2766), .Z(n1507) );
  IV U1939 ( .A(n2739), .Z(n1505) );
  IV U1940 ( .A(n2738), .Z(n1504) );
  IV U1941 ( .A(n2755), .Z(n1503) );
  IV U1942 ( .A(n3080), .Z(n1502) );
  IV U1943 ( .A(n2737), .Z(n1501) );
  IV U1944 ( .A(n2743), .Z(n1475) );
  IV U1945 ( .A(n2754), .Z(n1499) );
  IV U1946 ( .A(n2762), .Z(n1498) );
  IV U1947 ( .A(n2765), .Z(n1497) );
  IV U1948 ( .A(n3072), .Z(n1496) );
  IV U1949 ( .A(n3082), .Z(n1495) );
  IV U1950 ( .A(n2736), .Z(n1494) );
  IV U1951 ( .A(n3078), .Z(n1474) );
  IV U1952 ( .A(n2771), .Z(n1493) );
  IV U1953 ( .A(key[105]), .Z(n1695) );
  IV U1954 ( .A(n1720), .Z(n1694) );
  IV U1955 ( .A(n1703), .Z(n1693) );
  IV U1956 ( .A(n2769), .Z(n1492) );
  IV U1957 ( .A(n1700), .Z(n1692) );
  IV U1958 ( .A(key[107]), .Z(n1691) );
  IV U1959 ( .A(n2033), .Z(n1690) );
  IV U1960 ( .A(n2036), .Z(n1689) );
  IV U1961 ( .A(n1719), .Z(n1688) );
  IV U1962 ( .A(n2028), .Z(n1687) );
  IV U1963 ( .A(n2027), .Z(n1686) );
  IV U1964 ( .A(n1717), .Z(n1685) );
  IV U1965 ( .A(n1713), .Z(n1684) );
  IV U1966 ( .A(n1728), .Z(n1683) );
  IV U1967 ( .A(n1726), .Z(n1682) );
  IV U1968 ( .A(n1698), .Z(n1681) );
  IV U1969 ( .A(n1708), .Z(n1680) );
  IV U1970 ( .A(n1715), .Z(n1679) );
  IV U1971 ( .A(n1699), .Z(n1678) );
  IV U1972 ( .A(n1718), .Z(n1676) );
  IV U1973 ( .A(n1701), .Z(n1675) );
  IV U1974 ( .A(n1705), .Z(n1674) );
  IV U1975 ( .A(n1707), .Z(n1673) );
  IV U1976 ( .A(n1716), .Z(n1672) );
  IV U1977 ( .A(n1854), .Z(n1671) );
  IV U1978 ( .A(n2039), .Z(n1670) );
  IV U1979 ( .A(n1702), .Z(n1669) );
  IV U1980 ( .A(n1732), .Z(n1668) );
  IV U1981 ( .A(n1729), .Z(n1667) );
  IV U1982 ( .A(n1727), .Z(n1666) );
  IV U1983 ( .A(n1761), .Z(n1665) );
  IV U1984 ( .A(n2029), .Z(n1664) );
  IV U1985 ( .A(n2034), .Z(n1663) );
  IV U1986 ( .A(n2040), .Z(n1662) );
  IV U1987 ( .A(n1697), .Z(n1661) );
  IV U1988 ( .A(key[100]), .Z(n1490) );
  IV U1989 ( .A(n2038), .Z(n1660) );
  IV U1990 ( .A(n2035), .Z(n1659) );
  IV U1991 ( .A(n1714), .Z(n1658) );
  IV U1992 ( .A(n1709), .Z(n1656) );
  IV U1993 ( .A(n1723), .Z(n1655) );
  IV U1994 ( .A(n1725), .Z(n1654) );
  IV U1995 ( .A(n2031), .Z(n1653) );
  IV U1996 ( .A(n2041), .Z(n1652) );
  IV U1997 ( .A(n1696), .Z(n1651) );
  IV U1998 ( .A(n1733), .Z(n1650) );
  IV U1999 ( .A(n1730), .Z(n1649) );
  IV U2000 ( .A(n1704), .Z(n1647) );
  IV U2001 ( .A(key[108]), .Z(n1646) );
  IV U2002 ( .A(n3073), .Z(n1488) );
  IV U2003 ( .A(n1829), .Z(n1644) );
  IV U2004 ( .A(n2032), .Z(n1643) );
  IV U2005 ( .A(n1724), .Z(n1642) );
  IV U2006 ( .A(n2037), .Z(n1641) );
  IV U2007 ( .A(key[113]), .Z(n1640) );
  IV U2008 ( .A(n2080), .Z(n1639) );
  IV U2009 ( .A(n2064), .Z(n1638) );
  IV U2010 ( .A(n2763), .Z(n1487) );
  IV U2011 ( .A(n2047), .Z(n1637) );
  IV U2012 ( .A(key[115]), .Z(n1636) );
  IV U2013 ( .A(n2074), .Z(n1635) );
  IV U2014 ( .A(n2070), .Z(n1634) );
  IV U2015 ( .A(n2099), .Z(n1633) );
  IV U2016 ( .A(n2381), .Z(n1632) );
  IV U2017 ( .A(n2387), .Z(n1631) );
  IV U2018 ( .A(n2051), .Z(n1630) );
  IV U2019 ( .A(n2382), .Z(n1629) );
  IV U2020 ( .A(n2059), .Z(n1628) );
  IV U2021 ( .A(key[103]), .Z(n1473) );
  IV U2022 ( .A(n2050), .Z(n1627) );
  IV U2023 ( .A(n2053), .Z(n1626) );
  IV U2024 ( .A(n2062), .Z(n1625) );
  IV U2025 ( .A(n2376), .Z(n1624) );
  IV U2026 ( .A(n2201), .Z(n1623) );
  IV U2027 ( .A(n2046), .Z(n1622) );
  IV U2028 ( .A(n2078), .Z(n1621) );
  IV U2029 ( .A(n2073), .Z(n1620) );
  IV U2030 ( .A(n2072), .Z(n1619) );
  IV U2031 ( .A(n2759), .Z(n1486) );
  IV U2032 ( .A(n2045), .Z(n1617) );
  IV U2033 ( .A(n2044), .Z(n1616) );
  IV U2034 ( .A(n2061), .Z(n1615) );
  IV U2035 ( .A(n2386), .Z(n1614) );
  IV U2036 ( .A(n2043), .Z(n1613) );
  IV U2037 ( .A(n2060), .Z(n1611) );
  IV U2038 ( .A(n2068), .Z(n1610) );
  IV U2039 ( .A(n2071), .Z(n1609) );
  IV U2040 ( .A(n2378), .Z(n1608) );
  IV U2041 ( .A(n2388), .Z(n1607) );
  IV U2042 ( .A(n2042), .Z(n1606) );
  IV U2043 ( .A(n2077), .Z(n1605) );
  IV U2044 ( .A(n2075), .Z(n1604) );
  IV U2045 ( .A(n3074), .Z(n1485) );
  IV U2046 ( .A(key[116]), .Z(n1602) );
  IV U2047 ( .A(n2379), .Z(n1600) );
  IV U2048 ( .A(n2069), .Z(n1599) );
  IV U2049 ( .A(n2065), .Z(n1598) );
  IV U2050 ( .A(n3077), .Z(n1484) );
  IV U2051 ( .A(n2380), .Z(n1597) );
  IV U2052 ( .A(n2383), .Z(n1596) );
  IV U2053 ( .A(n2385), .Z(n1595) );
  IV U2054 ( .A(n2048), .Z(n1594) );
  IV U2055 ( .A(n2184), .Z(n1593) );
  IV U2056 ( .A(n2375), .Z(n1592) );
  IV U2057 ( .A(n2374), .Z(n1591) );
  IV U2058 ( .A(n2054), .Z(n1590) );
  IV U2059 ( .A(n3079), .Z(n1483) );
  IV U2060 ( .A(n2063), .Z(n1589) );
  IV U2061 ( .A(n2058), .Z(n1588) );
  IV U2062 ( .A(n2049), .Z(n1587) );
  IV U2063 ( .A(n2384), .Z(n1586) );
  IV U2064 ( .A(key[119]), .Z(n1585) );
  IV U2065 ( .A(key[121]), .Z(n1584) );
  IV U2066 ( .A(n2427), .Z(n1583) );
  IV U2067 ( .A(n2742), .Z(n1482) );
  IV U2068 ( .A(n2411), .Z(n1582) );
  IV U2069 ( .A(n2394), .Z(n1581) );
  IV U2070 ( .A(key[123]), .Z(n1580) );
  IV U2071 ( .A(n2421), .Z(n1579) );
  IV U2072 ( .A(n2417), .Z(n1578) );
  IV U2073 ( .A(n2446), .Z(n1577) );
  IV U2074 ( .A(n2728), .Z(n1576) );
  IV U2075 ( .A(n2734), .Z(n1575) );
  IV U2076 ( .A(n2398), .Z(n1574) );
  IV U2077 ( .A(n2729), .Z(n1573) );
  IV U2078 ( .A(n2878), .Z(n1481) );
  IV U2079 ( .A(n2406), .Z(n1572) );
  IV U2080 ( .A(n2397), .Z(n1571) );
  IV U2081 ( .A(n2400), .Z(n1570) );
  IV U2082 ( .A(n2409), .Z(n1569) );
  IV U2083 ( .A(n2723), .Z(n1568) );
  IV U2084 ( .A(n2548), .Z(n1567) );
  IV U2085 ( .A(n2393), .Z(n1566) );
  IV U2086 ( .A(n2425), .Z(n1565) );
  IV U2087 ( .A(n2420), .Z(n1564) );
  IV U2088 ( .A(n2419), .Z(n1563) );
  IV U2089 ( .A(n2392), .Z(n1561) );
  IV U2090 ( .A(n2391), .Z(n1560) );
  IV U2091 ( .A(n2408), .Z(n1559) );
  IV U2092 ( .A(n2733), .Z(n1558) );
  IV U2093 ( .A(n2390), .Z(n1557) );
  IV U2094 ( .A(n3069), .Z(n1480) );
  IV U2095 ( .A(n2407), .Z(n1555) );
  IV U2096 ( .A(n2415), .Z(n1554) );
  IV U2097 ( .A(n2418), .Z(n1553) );
  IV U2098 ( .A(n2725), .Z(n1552) );
  IV U2099 ( .A(n2735), .Z(n1551) );
  IV U2100 ( .A(n2389), .Z(n1550) );
  IV U2101 ( .A(n2424), .Z(n1549) );
  IV U2102 ( .A(n3068), .Z(n1479) );
  XNOR U2103 ( .A(n1407), .B(n1408), .Z(\d/n420 ) );
  XNOR U2104 ( .A(shift_row_out[0]), .B(shift_row_out[8]), .Z(n1407) );
  XNOR U2105 ( .A(n1409), .B(n1408), .Z(\d/n419 ) );
  XNOR U2106 ( .A(shift_row_out[10]), .B(shift_row_out[2]), .Z(n1409) );
  XNOR U2107 ( .A(n1410), .B(n1408), .Z(\d/n418 ) );
  XNOR U2108 ( .A(shift_row_out[15]), .B(shift_row_out[7]), .Z(n1408) );
  XNOR U2109 ( .A(shift_row_out[11]), .B(shift_row_out[3]), .Z(n1410) );
  XNOR U2110 ( .A(shift_row_out[16]), .B(shift_row_out[8]), .Z(n1411) );
  XOR U2111 ( .A(n1413), .B(n1412), .Z(\d/n416 ) );
  XNOR U2112 ( .A(shift_row_out[10]), .B(shift_row_out[18]), .Z(n1413) );
  XOR U2113 ( .A(n1414), .B(n1412), .Z(\d/n415 ) );
  XOR U2114 ( .A(shift_row_out[15]), .B(shift_row_out[23]), .Z(n1412) );
  XNOR U2115 ( .A(shift_row_out[11]), .B(shift_row_out[19]), .Z(n1414) );
  XOR U2116 ( .A(n1415), .B(n1416), .Z(\d/n414 ) );
  XNOR U2117 ( .A(shift_row_out[16]), .B(shift_row_out[24]), .Z(n1415) );
  XOR U2118 ( .A(n1417), .B(n1416), .Z(\d/n413 ) );
  XNOR U2119 ( .A(shift_row_out[18]), .B(shift_row_out[26]), .Z(n1417) );
  XOR U2120 ( .A(n1418), .B(n1416), .Z(\d/n412 ) );
  XOR U2121 ( .A(n1170), .B(n1124), .Z(n1416) );
  IV U2122 ( .A(shift_row_out[23]), .Z(n1170) );
  XNOR U2123 ( .A(shift_row_out[19]), .B(shift_row_out[27]), .Z(n1418) );
  XNOR U2124 ( .A(n1419), .B(n1420), .Z(\d/n411 ) );
  XNOR U2125 ( .A(shift_row_out[0]), .B(shift_row_out[24]), .Z(n1419) );
  XNOR U2126 ( .A(n1421), .B(n1420), .Z(\d/n410 ) );
  XNOR U2127 ( .A(shift_row_out[26]), .B(shift_row_out[2]), .Z(n1421) );
  XNOR U2128 ( .A(n1422), .B(n1420), .Z(\d/n409 ) );
  XOR U2129 ( .A(n1124), .B(shift_row_out[7]), .Z(n1420) );
  IV U2130 ( .A(shift_row_out[31]), .Z(n1124) );
  XNOR U2131 ( .A(shift_row_out[27]), .B(shift_row_out[3]), .Z(n1422) );
  XNOR U2132 ( .A(shift_row_out[32]), .B(shift_row_out[40]), .Z(n1423) );
  XOR U2133 ( .A(n1425), .B(n1424), .Z(\d/n407 ) );
  XNOR U2134 ( .A(shift_row_out[34]), .B(shift_row_out[42]), .Z(n1425) );
  XOR U2135 ( .A(n1426), .B(n1424), .Z(\d/n406 ) );
  XOR U2136 ( .A(shift_row_out[39]), .B(shift_row_out[47]), .Z(n1424) );
  XNOR U2137 ( .A(shift_row_out[35]), .B(shift_row_out[43]), .Z(n1426) );
  XOR U2138 ( .A(n1427), .B(n1428), .Z(\d/n405 ) );
  XNOR U2139 ( .A(shift_row_out[40]), .B(shift_row_out[48]), .Z(n1427) );
  XOR U2140 ( .A(n1429), .B(n1428), .Z(\d/n404 ) );
  XNOR U2141 ( .A(shift_row_out[42]), .B(shift_row_out[50]), .Z(n1429) );
  XOR U2142 ( .A(n1430), .B(n1428), .Z(\d/n403 ) );
  XOR U2143 ( .A(n1038), .B(n992), .Z(n1428) );
  IV U2144 ( .A(shift_row_out[47]), .Z(n1038) );
  XNOR U2145 ( .A(shift_row_out[43]), .B(shift_row_out[51]), .Z(n1430) );
  XNOR U2146 ( .A(n1431), .B(n1432), .Z(\d/n402 ) );
  XNOR U2147 ( .A(shift_row_out[48]), .B(shift_row_out[56]), .Z(n1431) );
  XNOR U2148 ( .A(n1433), .B(n1432), .Z(\d/n401 ) );
  XNOR U2149 ( .A(shift_row_out[50]), .B(shift_row_out[58]), .Z(n1433) );
  XNOR U2150 ( .A(n1434), .B(n1432), .Z(\d/n400 ) );
  XOR U2151 ( .A(n992), .B(shift_row_out[63]), .Z(n1432) );
  IV U2152 ( .A(shift_row_out[55]), .Z(n992) );
  XNOR U2153 ( .A(shift_row_out[51]), .B(shift_row_out[59]), .Z(n1434) );
  XNOR U2154 ( .A(n1435), .B(n1436), .Z(\d/n399 ) );
  XNOR U2155 ( .A(shift_row_out[32]), .B(shift_row_out[56]), .Z(n1435) );
  XNOR U2156 ( .A(n1437), .B(n1436), .Z(\d/n398 ) );
  XNOR U2157 ( .A(shift_row_out[34]), .B(shift_row_out[58]), .Z(n1437) );
  XNOR U2158 ( .A(n1438), .B(n1436), .Z(\d/n397 ) );
  XNOR U2159 ( .A(shift_row_out[39]), .B(shift_row_out[63]), .Z(n1436) );
  XNOR U2160 ( .A(shift_row_out[35]), .B(shift_row_out[59]), .Z(n1438) );
  XNOR U2161 ( .A(shift_row_out[64]), .B(shift_row_out[72]), .Z(n1439) );
  XOR U2162 ( .A(n1441), .B(n1440), .Z(\d/n395 ) );
  XNOR U2163 ( .A(shift_row_out[66]), .B(shift_row_out[74]), .Z(n1441) );
  XOR U2164 ( .A(n1442), .B(n1440), .Z(\d/n394 ) );
  XOR U2165 ( .A(shift_row_out[71]), .B(shift_row_out[79]), .Z(n1440) );
  XNOR U2166 ( .A(shift_row_out[67]), .B(shift_row_out[75]), .Z(n1442) );
  XOR U2167 ( .A(n1443), .B(n1444), .Z(\d/n393 ) );
  XNOR U2168 ( .A(shift_row_out[72]), .B(shift_row_out[80]), .Z(n1443) );
  XOR U2169 ( .A(n1445), .B(n1444), .Z(\d/n392 ) );
  XNOR U2170 ( .A(shift_row_out[74]), .B(shift_row_out[82]), .Z(n1445) );
  XOR U2171 ( .A(n1446), .B(n1444), .Z(\d/n391 ) );
  XOR U2172 ( .A(n861), .B(n815), .Z(n1444) );
  IV U2173 ( .A(shift_row_out[79]), .Z(n861) );
  XNOR U2174 ( .A(shift_row_out[75]), .B(shift_row_out[83]), .Z(n1446) );
  XNOR U2175 ( .A(n1447), .B(n1448), .Z(\d/n390 ) );
  XNOR U2176 ( .A(shift_row_out[80]), .B(shift_row_out[88]), .Z(n1447) );
  XNOR U2177 ( .A(n1449), .B(n1448), .Z(\d/n389 ) );
  XNOR U2178 ( .A(shift_row_out[82]), .B(shift_row_out[90]), .Z(n1449) );
  XNOR U2179 ( .A(n1450), .B(n1448), .Z(\d/n388 ) );
  XOR U2180 ( .A(n815), .B(shift_row_out[95]), .Z(n1448) );
  IV U2181 ( .A(shift_row_out[87]), .Z(n815) );
  XNOR U2182 ( .A(shift_row_out[83]), .B(shift_row_out[91]), .Z(n1450) );
  XNOR U2183 ( .A(n1451), .B(n1452), .Z(\d/n387 ) );
  XNOR U2184 ( .A(shift_row_out[64]), .B(shift_row_out[88]), .Z(n1451) );
  XNOR U2185 ( .A(n1453), .B(n1452), .Z(\d/n386 ) );
  XNOR U2186 ( .A(shift_row_out[66]), .B(shift_row_out[90]), .Z(n1453) );
  XNOR U2187 ( .A(n1454), .B(n1452), .Z(\d/n385 ) );
  XNOR U2188 ( .A(shift_row_out[71]), .B(shift_row_out[95]), .Z(n1452) );
  XNOR U2189 ( .A(shift_row_out[67]), .B(shift_row_out[91]), .Z(n1454) );
  XNOR U2190 ( .A(shift_row_out[104]), .B(shift_row_out[96]), .Z(n1455) );
  XOR U2191 ( .A(n1457), .B(n1456), .Z(\d/n383 ) );
  XNOR U2192 ( .A(shift_row_out[106]), .B(shift_row_out[98]), .Z(n1457) );
  XOR U2193 ( .A(n1458), .B(n1456), .Z(\d/n382 ) );
  XOR U2194 ( .A(shift_row_out[103]), .B(shift_row_out[111]), .Z(n1456) );
  XNOR U2195 ( .A(shift_row_out[107]), .B(shift_row_out[99]), .Z(n1458) );
  XOR U2196 ( .A(n1459), .B(n1460), .Z(\d/n381 ) );
  XNOR U2197 ( .A(shift_row_out[104]), .B(shift_row_out[112]), .Z(n1459) );
  XOR U2198 ( .A(n1461), .B(n1460), .Z(\d/n380 ) );
  XNOR U2199 ( .A(shift_row_out[106]), .B(shift_row_out[114]), .Z(n1461) );
  XOR U2200 ( .A(n1462), .B(n1460), .Z(\d/n379 ) );
  XOR U2201 ( .A(n1322), .B(n1281), .Z(n1460) );
  IV U2202 ( .A(shift_row_out[111]), .Z(n1322) );
  XNOR U2203 ( .A(shift_row_out[107]), .B(shift_row_out[115]), .Z(n1462) );
  XNOR U2204 ( .A(n1463), .B(n1464), .Z(\d/n378 ) );
  XNOR U2205 ( .A(shift_row_out[112]), .B(shift_row_out[120]), .Z(n1463) );
  XNOR U2206 ( .A(n1465), .B(n1464), .Z(\d/n377 ) );
  XNOR U2207 ( .A(shift_row_out[114]), .B(shift_row_out[122]), .Z(n1465) );
  XNOR U2208 ( .A(n1466), .B(n1464), .Z(\d/n376 ) );
  XOR U2209 ( .A(n1281), .B(shift_row_out[127]), .Z(n1464) );
  IV U2210 ( .A(shift_row_out[119]), .Z(n1281) );
  XNOR U2211 ( .A(shift_row_out[115]), .B(shift_row_out[123]), .Z(n1466) );
  XNOR U2212 ( .A(n1467), .B(n1468), .Z(\d/n375 ) );
  XNOR U2213 ( .A(shift_row_out[120]), .B(shift_row_out[96]), .Z(n1467) );
  XNOR U2214 ( .A(n1469), .B(n1468), .Z(\d/n374 ) );
  XNOR U2215 ( .A(shift_row_out[122]), .B(shift_row_out[98]), .Z(n1469) );
  XNOR U2216 ( .A(n1470), .B(n1468), .Z(\d/n373 ) );
  XNOR U2217 ( .A(shift_row_out[103]), .B(shift_row_out[127]), .Z(n1468) );
  XNOR U2218 ( .A(shift_row_out[123]), .B(shift_row_out[99]), .Z(n1470) );
  IV U2219 ( .A(\b/n1512 ), .Z(\b/n999 ) );
  IV U2220 ( .A(\b/n1502 ), .Z(\b/n997 ) );
  IV U2221 ( .A(\b/n1523 ), .Z(\b/n996 ) );
  IV U2222 ( .A(\b/n1847 ), .Z(\b/n995 ) );
  IV U2223 ( .A(msg[17]), .Z(\b/n993 ) );
  IV U2224 ( .A(\b/n1895 ), .Z(\b/n991 ) );
  IV U2225 ( .A(\b/n1877 ), .Z(\b/n990 ) );
  IV U2226 ( .A(\b/n6196 ), .Z(\b/n99 ) );
  IV U2227 ( .A(\b/n1858 ), .Z(\b/n989 ) );
  IV U2228 ( .A(msg[19]), .Z(\b/n988 ) );
  IV U2229 ( .A(\b/n1888 ), .Z(\b/n987 ) );
  IV U2230 ( .A(\b/n1883 ), .Z(\b/n986 ) );
  IV U2231 ( .A(\b/n1914 ), .Z(\b/n985 ) );
  IV U2232 ( .A(\b/n2203 ), .Z(\b/n984 ) );
  IV U2233 ( .A(\b/n2210 ), .Z(\b/n983 ) );
  IV U2234 ( .A(\b/n1862 ), .Z(\b/n982 ) );
  IV U2235 ( .A(\b/n2204 ), .Z(\b/n981 ) );
  IV U2236 ( .A(\b/n1870 ), .Z(\b/n980 ) );
  IV U2237 ( .A(\b/n1861 ), .Z(\b/n979 ) );
  IV U2238 ( .A(\b/n1864 ), .Z(\b/n978 ) );
  IV U2239 ( .A(\b/n1874 ), .Z(\b/n977 ) );
  IV U2240 ( .A(\b/n2194 ), .Z(\b/n976 ) );
  IV U2241 ( .A(\b/n2016 ), .Z(\b/n975 ) );
  IV U2242 ( .A(\b/n1857 ), .Z(\b/n973 ) );
  IV U2243 ( .A(\b/n1892 ), .Z(\b/n972 ) );
  IV U2244 ( .A(\b/n1886 ), .Z(\b/n971 ) );
  IV U2245 ( .A(\b/n1885 ), .Z(\b/n970 ) );
  IV U2246 ( .A(\b/n1856 ), .Z(\b/n968 ) );
  IV U2247 ( .A(\b/n1855 ), .Z(\b/n967 ) );
  IV U2248 ( .A(\b/n1873 ), .Z(\b/n965 ) );
  IV U2249 ( .A(\b/n2209 ), .Z(\b/n964 ) );
  IV U2250 ( .A(\b/n1854 ), .Z(\b/n963 ) );
  IV U2251 ( .A(\b/n1872 ), .Z(\b/n960 ) );
  IV U2252 ( .A(\b/n1881 ), .Z(\b/n958 ) );
  IV U2253 ( .A(\b/n1884 ), .Z(\b/n957 ) );
  IV U2254 ( .A(\b/n2197 ), .Z(\b/n954 ) );
  IV U2255 ( .A(\b/n2211 ), .Z(\b/n953 ) );
  IV U2256 ( .A(\b/n1853 ), .Z(\b/n952 ) );
  IV U2257 ( .A(\b/n1891 ), .Z(\b/n951 ) );
  IV U2258 ( .A(\b/n1889 ), .Z(\b/n950 ) );
  IV U2259 ( .A(msg[116]), .Z(\b/n95 ) );
  IV U2260 ( .A(msg[20]), .Z(\b/n946 ) );
  IV U2261 ( .A(\b/n2201 ), .Z(\b/n944 ) );
  IV U2262 ( .A(\b/n1882 ), .Z(\b/n943 ) );
  IV U2263 ( .A(\b/n1878 ), .Z(\b/n941 ) );
  IV U2264 ( .A(\b/n2202 ), .Z(\b/n939 ) );
  IV U2265 ( .A(\b/n2205 ), .Z(\b/n938 ) );
  IV U2266 ( .A(\b/n2208 ), .Z(\b/n937 ) );
  IV U2267 ( .A(\b/n1859 ), .Z(\b/n936 ) );
  IV U2268 ( .A(\b/n1999 ), .Z(\b/n935 ) );
  IV U2269 ( .A(\b/n2193 ), .Z(\b/n933 ) );
  IV U2270 ( .A(\b/n2191 ), .Z(\b/n932 ) );
  IV U2271 ( .A(\b/n1865 ), .Z(\b/n931 ) );
  IV U2272 ( .A(\b/n6508 ), .Z(\b/n93 ) );
  IV U2273 ( .A(\b/n1876 ), .Z(\b/n929 ) );
  IV U2274 ( .A(\b/n1869 ), .Z(\b/n928 ) );
  IV U2275 ( .A(\b/n1860 ), .Z(\b/n926 ) );
  IV U2276 ( .A(\b/n2206 ), .Z(\b/n925 ) );
  IV U2277 ( .A(msg[23]), .Z(\b/n924 ) );
  IV U2278 ( .A(msg[25]), .Z(\b/n922 ) );
  IV U2279 ( .A(\b/n2254 ), .Z(\b/n920 ) );
  IV U2280 ( .A(\b/n6189 ), .Z(\b/n92 ) );
  IV U2281 ( .A(\b/n2236 ), .Z(\b/n919 ) );
  IV U2282 ( .A(\b/n2217 ), .Z(\b/n918 ) );
  IV U2283 ( .A(msg[27]), .Z(\b/n917 ) );
  IV U2284 ( .A(\b/n2247 ), .Z(\b/n916 ) );
  IV U2285 ( .A(\b/n2242 ), .Z(\b/n915 ) );
  IV U2286 ( .A(\b/n2273 ), .Z(\b/n914 ) );
  IV U2287 ( .A(\b/n2562 ), .Z(\b/n913 ) );
  IV U2288 ( .A(\b/n2569 ), .Z(\b/n912 ) );
  IV U2289 ( .A(\b/n2221 ), .Z(\b/n911 ) );
  IV U2290 ( .A(\b/n2563 ), .Z(\b/n910 ) );
  IV U2291 ( .A(\b/n2229 ), .Z(\b/n909 ) );
  IV U2292 ( .A(\b/n2220 ), .Z(\b/n908 ) );
  IV U2293 ( .A(\b/n2223 ), .Z(\b/n907 ) );
  IV U2294 ( .A(\b/n2233 ), .Z(\b/n906 ) );
  IV U2295 ( .A(\b/n2553 ), .Z(\b/n905 ) );
  IV U2296 ( .A(\b/n2375 ), .Z(\b/n904 ) );
  IV U2297 ( .A(\b/n2216 ), .Z(\b/n902 ) );
  IV U2298 ( .A(\b/n2251 ), .Z(\b/n901 ) );
  IV U2299 ( .A(\b/n2245 ), .Z(\b/n900 ) );
  IV U2300 ( .A(\b/n6185 ), .Z(\b/n90 ) );
  IV U2301 ( .A(\b/n6531 ), .Z(\b/n9 ) );
  IV U2302 ( .A(\b/n2244 ), .Z(\b/n899 ) );
  IV U2303 ( .A(\b/n2215 ), .Z(\b/n897 ) );
  IV U2304 ( .A(\b/n2214 ), .Z(\b/n896 ) );
  IV U2305 ( .A(\b/n2232 ), .Z(\b/n894 ) );
  IV U2306 ( .A(\b/n2568 ), .Z(\b/n893 ) );
  IV U2307 ( .A(\b/n2213 ), .Z(\b/n892 ) );
  IV U2308 ( .A(\b/n2231 ), .Z(\b/n889 ) );
  IV U2309 ( .A(\b/n2240 ), .Z(\b/n887 ) );
  IV U2310 ( .A(\b/n2243 ), .Z(\b/n886 ) );
  IV U2311 ( .A(\b/n2556 ), .Z(\b/n883 ) );
  IV U2312 ( .A(\b/n2570 ), .Z(\b/n882 ) );
  IV U2313 ( .A(\b/n2212 ), .Z(\b/n881 ) );
  IV U2314 ( .A(\b/n2250 ), .Z(\b/n880 ) );
  IV U2315 ( .A(\b/n6509 ), .Z(\b/n88 ) );
  IV U2316 ( .A(\b/n2248 ), .Z(\b/n879 ) );
  IV U2317 ( .A(msg[28]), .Z(\b/n875 ) );
  IV U2318 ( .A(\b/n2560 ), .Z(\b/n873 ) );
  IV U2319 ( .A(\b/n2241 ), .Z(\b/n872 ) );
  IV U2320 ( .A(\b/n2237 ), .Z(\b/n870 ) );
  IV U2321 ( .A(\b/n6512 ), .Z(\b/n87 ) );
  IV U2322 ( .A(\b/n2561 ), .Z(\b/n868 ) );
  IV U2323 ( .A(\b/n2564 ), .Z(\b/n867 ) );
  IV U2324 ( .A(\b/n2567 ), .Z(\b/n866 ) );
  IV U2325 ( .A(\b/n2218 ), .Z(\b/n865 ) );
  IV U2326 ( .A(\b/n2358 ), .Z(\b/n864 ) );
  IV U2327 ( .A(\b/n2552 ), .Z(\b/n862 ) );
  IV U2328 ( .A(\b/n2550 ), .Z(\b/n861 ) );
  IV U2329 ( .A(\b/n2224 ), .Z(\b/n860 ) );
  IV U2330 ( .A(\b/n6515 ), .Z(\b/n86 ) );
  IV U2331 ( .A(\b/n2235 ), .Z(\b/n858 ) );
  IV U2332 ( .A(\b/n2228 ), .Z(\b/n857 ) );
  IV U2333 ( .A(\b/n2219 ), .Z(\b/n855 ) );
  IV U2334 ( .A(\b/n2565 ), .Z(\b/n854 ) );
  IV U2335 ( .A(msg[31]), .Z(\b/n853 ) );
  IV U2336 ( .A(msg[33]), .Z(\b/n851 ) );
  IV U2337 ( .A(\b/n6166 ), .Z(\b/n85 ) );
  IV U2338 ( .A(\b/n2613 ), .Z(\b/n849 ) );
  IV U2339 ( .A(\b/n2595 ), .Z(\b/n848 ) );
  IV U2340 ( .A(\b/n2576 ), .Z(\b/n847 ) );
  IV U2341 ( .A(msg[35]), .Z(\b/n846 ) );
  IV U2342 ( .A(\b/n2606 ), .Z(\b/n845 ) );
  IV U2343 ( .A(\b/n2601 ), .Z(\b/n844 ) );
  IV U2344 ( .A(\b/n2632 ), .Z(\b/n843 ) );
  IV U2345 ( .A(\b/n2921 ), .Z(\b/n842 ) );
  IV U2346 ( .A(\b/n2928 ), .Z(\b/n841 ) );
  IV U2347 ( .A(\b/n2580 ), .Z(\b/n840 ) );
  IV U2348 ( .A(\b/n6306 ), .Z(\b/n84 ) );
  IV U2349 ( .A(\b/n2922 ), .Z(\b/n839 ) );
  IV U2350 ( .A(\b/n2588 ), .Z(\b/n838 ) );
  IV U2351 ( .A(\b/n2579 ), .Z(\b/n837 ) );
  IV U2352 ( .A(\b/n2582 ), .Z(\b/n836 ) );
  IV U2353 ( .A(\b/n2592 ), .Z(\b/n835 ) );
  IV U2354 ( .A(\b/n2912 ), .Z(\b/n834 ) );
  IV U2355 ( .A(\b/n2734 ), .Z(\b/n833 ) );
  IV U2356 ( .A(\b/n2575 ), .Z(\b/n831 ) );
  IV U2357 ( .A(\b/n2610 ), .Z(\b/n830 ) );
  IV U2358 ( .A(\b/n2604 ), .Z(\b/n829 ) );
  IV U2359 ( .A(\b/n2603 ), .Z(\b/n828 ) );
  IV U2360 ( .A(\b/n2574 ), .Z(\b/n826 ) );
  IV U2361 ( .A(\b/n2573 ), .Z(\b/n825 ) );
  IV U2362 ( .A(\b/n2591 ), .Z(\b/n823 ) );
  IV U2363 ( .A(\b/n2927 ), .Z(\b/n822 ) );
  IV U2364 ( .A(\b/n2572 ), .Z(\b/n821 ) );
  IV U2365 ( .A(\b/n6500 ), .Z(\b/n82 ) );
  IV U2366 ( .A(\b/n2590 ), .Z(\b/n818 ) );
  IV U2367 ( .A(\b/n2599 ), .Z(\b/n816 ) );
  IV U2368 ( .A(\b/n2602 ), .Z(\b/n815 ) );
  IV U2369 ( .A(\b/n2915 ), .Z(\b/n812 ) );
  IV U2370 ( .A(\b/n2929 ), .Z(\b/n811 ) );
  IV U2371 ( .A(\b/n2571 ), .Z(\b/n810 ) );
  IV U2372 ( .A(\b/n6498 ), .Z(\b/n81 ) );
  IV U2373 ( .A(\b/n2609 ), .Z(\b/n809 ) );
  IV U2374 ( .A(\b/n2607 ), .Z(\b/n808 ) );
  IV U2375 ( .A(msg[36]), .Z(\b/n804 ) );
  IV U2376 ( .A(\b/n2919 ), .Z(\b/n802 ) );
  IV U2377 ( .A(\b/n2600 ), .Z(\b/n801 ) );
  IV U2378 ( .A(\b/n6172 ), .Z(\b/n80 ) );
  IV U2379 ( .A(\b/n2596 ), .Z(\b/n799 ) );
  IV U2380 ( .A(\b/n2920 ), .Z(\b/n797 ) );
  IV U2381 ( .A(\b/n2923 ), .Z(\b/n796 ) );
  IV U2382 ( .A(\b/n2926 ), .Z(\b/n795 ) );
  IV U2383 ( .A(\b/n2577 ), .Z(\b/n794 ) );
  IV U2384 ( .A(\b/n2717 ), .Z(\b/n793 ) );
  IV U2385 ( .A(\b/n2911 ), .Z(\b/n791 ) );
  IV U2386 ( .A(\b/n2909 ), .Z(\b/n790 ) );
  IV U2387 ( .A(\b/n2583 ), .Z(\b/n789 ) );
  IV U2388 ( .A(\b/n2594 ), .Z(\b/n787 ) );
  IV U2389 ( .A(\b/n2587 ), .Z(\b/n786 ) );
  IV U2390 ( .A(\b/n2578 ), .Z(\b/n784 ) );
  IV U2391 ( .A(\b/n2924 ), .Z(\b/n783 ) );
  IV U2392 ( .A(msg[39]), .Z(\b/n782 ) );
  IV U2393 ( .A(msg[41]), .Z(\b/n780 ) );
  IV U2394 ( .A(\b/n6183 ), .Z(\b/n78 ) );
  IV U2395 ( .A(\b/n2972 ), .Z(\b/n778 ) );
  IV U2396 ( .A(\b/n2954 ), .Z(\b/n777 ) );
  IV U2397 ( .A(\b/n2935 ), .Z(\b/n776 ) );
  IV U2398 ( .A(msg[43]), .Z(\b/n775 ) );
  IV U2399 ( .A(\b/n2965 ), .Z(\b/n774 ) );
  IV U2400 ( .A(\b/n2960 ), .Z(\b/n773 ) );
  IV U2401 ( .A(\b/n2991 ), .Z(\b/n772 ) );
  IV U2402 ( .A(\b/n3280 ), .Z(\b/n771 ) );
  IV U2403 ( .A(\b/n3287 ), .Z(\b/n770 ) );
  IV U2404 ( .A(\b/n6176 ), .Z(\b/n77 ) );
  IV U2405 ( .A(\b/n2939 ), .Z(\b/n769 ) );
  IV U2406 ( .A(\b/n3281 ), .Z(\b/n768 ) );
  IV U2407 ( .A(\b/n2947 ), .Z(\b/n767 ) );
  IV U2408 ( .A(\b/n2938 ), .Z(\b/n766 ) );
  IV U2409 ( .A(\b/n2941 ), .Z(\b/n765 ) );
  IV U2410 ( .A(\b/n2951 ), .Z(\b/n764 ) );
  IV U2411 ( .A(\b/n3271 ), .Z(\b/n763 ) );
  IV U2412 ( .A(\b/n3093 ), .Z(\b/n762 ) );
  IV U2413 ( .A(\b/n2934 ), .Z(\b/n760 ) );
  IV U2414 ( .A(\b/n2969 ), .Z(\b/n759 ) );
  IV U2415 ( .A(\b/n2963 ), .Z(\b/n758 ) );
  IV U2416 ( .A(\b/n2962 ), .Z(\b/n757 ) );
  IV U2417 ( .A(\b/n2933 ), .Z(\b/n755 ) );
  IV U2418 ( .A(\b/n2932 ), .Z(\b/n754 ) );
  IV U2419 ( .A(\b/n2950 ), .Z(\b/n752 ) );
  IV U2420 ( .A(\b/n3286 ), .Z(\b/n751 ) );
  IV U2421 ( .A(\b/n2931 ), .Z(\b/n750 ) );
  IV U2422 ( .A(\b/n6167 ), .Z(\b/n75 ) );
  IV U2423 ( .A(\b/n2949 ), .Z(\b/n747 ) );
  IV U2424 ( .A(\b/n2958 ), .Z(\b/n745 ) );
  IV U2425 ( .A(\b/n2961 ), .Z(\b/n744 ) );
  IV U2426 ( .A(\b/n3274 ), .Z(\b/n741 ) );
  IV U2427 ( .A(\b/n3288 ), .Z(\b/n740 ) );
  IV U2428 ( .A(\b/n6513 ), .Z(\b/n74 ) );
  IV U2429 ( .A(\b/n2930 ), .Z(\b/n739 ) );
  IV U2430 ( .A(\b/n2968 ), .Z(\b/n738 ) );
  IV U2431 ( .A(\b/n2966 ), .Z(\b/n737 ) );
  IV U2432 ( .A(msg[44]), .Z(\b/n733 ) );
  IV U2433 ( .A(\b/n3278 ), .Z(\b/n731 ) );
  IV U2434 ( .A(\b/n2959 ), .Z(\b/n730 ) );
  IV U2435 ( .A(msg[119]), .Z(\b/n73 ) );
  IV U2436 ( .A(\b/n2955 ), .Z(\b/n728 ) );
  IV U2437 ( .A(\b/n3279 ), .Z(\b/n726 ) );
  IV U2438 ( .A(\b/n3282 ), .Z(\b/n725 ) );
  IV U2439 ( .A(\b/n3285 ), .Z(\b/n724 ) );
  IV U2440 ( .A(\b/n2936 ), .Z(\b/n723 ) );
  IV U2441 ( .A(\b/n3076 ), .Z(\b/n722 ) );
  IV U2442 ( .A(\b/n3270 ), .Z(\b/n720 ) );
  IV U2443 ( .A(\b/n3268 ), .Z(\b/n719 ) );
  IV U2444 ( .A(\b/n2942 ), .Z(\b/n718 ) );
  IV U2445 ( .A(\b/n2953 ), .Z(\b/n716 ) );
  IV U2446 ( .A(\b/n2946 ), .Z(\b/n715 ) );
  IV U2447 ( .A(\b/n2937 ), .Z(\b/n713 ) );
  IV U2448 ( .A(\b/n3283 ), .Z(\b/n712 ) );
  IV U2449 ( .A(msg[47]), .Z(\b/n711 ) );
  IV U2450 ( .A(msg[121]), .Z(\b/n71 ) );
  IV U2451 ( .A(msg[49]), .Z(\b/n709 ) );
  IV U2452 ( .A(\b/n3331 ), .Z(\b/n707 ) );
  IV U2453 ( .A(\b/n3313 ), .Z(\b/n706 ) );
  IV U2454 ( .A(\b/n3294 ), .Z(\b/n705 ) );
  IV U2455 ( .A(msg[51]), .Z(\b/n704 ) );
  IV U2456 ( .A(\b/n3324 ), .Z(\b/n703 ) );
  IV U2457 ( .A(\b/n3319 ), .Z(\b/n702 ) );
  IV U2458 ( .A(\b/n3350 ), .Z(\b/n701 ) );
  IV U2459 ( .A(\b/n3639 ), .Z(\b/n700 ) );
  IV U2460 ( .A(\b/n6542 ), .Z(\b/n7 ) );
  IV U2461 ( .A(\b/n3646 ), .Z(\b/n699 ) );
  IV U2462 ( .A(\b/n3298 ), .Z(\b/n698 ) );
  IV U2463 ( .A(\b/n3640 ), .Z(\b/n697 ) );
  IV U2464 ( .A(\b/n3306 ), .Z(\b/n696 ) );
  IV U2465 ( .A(\b/n3297 ), .Z(\b/n695 ) );
  IV U2466 ( .A(\b/n3300 ), .Z(\b/n694 ) );
  IV U2467 ( .A(\b/n3310 ), .Z(\b/n693 ) );
  IV U2468 ( .A(\b/n3630 ), .Z(\b/n692 ) );
  IV U2469 ( .A(\b/n3452 ), .Z(\b/n691 ) );
  IV U2470 ( .A(\b/n6561 ), .Z(\b/n69 ) );
  IV U2471 ( .A(\b/n3293 ), .Z(\b/n689 ) );
  IV U2472 ( .A(\b/n3328 ), .Z(\b/n688 ) );
  IV U2473 ( .A(\b/n3322 ), .Z(\b/n687 ) );
  IV U2474 ( .A(\b/n3321 ), .Z(\b/n686 ) );
  IV U2475 ( .A(\b/n3292 ), .Z(\b/n684 ) );
  IV U2476 ( .A(\b/n3291 ), .Z(\b/n683 ) );
  IV U2477 ( .A(\b/n3309 ), .Z(\b/n681 ) );
  IV U2478 ( .A(\b/n3645 ), .Z(\b/n680 ) );
  IV U2479 ( .A(\b/n6543 ), .Z(\b/n68 ) );
  IV U2480 ( .A(\b/n3290 ), .Z(\b/n679 ) );
  IV U2481 ( .A(\b/n3308 ), .Z(\b/n676 ) );
  IV U2482 ( .A(\b/n3317 ), .Z(\b/n674 ) );
  IV U2483 ( .A(\b/n3320 ), .Z(\b/n673 ) );
  IV U2484 ( .A(\b/n3633 ), .Z(\b/n670 ) );
  IV U2485 ( .A(\b/n6524 ), .Z(\b/n67 ) );
  IV U2486 ( .A(\b/n3647 ), .Z(\b/n669 ) );
  IV U2487 ( .A(\b/n3289 ), .Z(\b/n668 ) );
  IV U2488 ( .A(\b/n3327 ), .Z(\b/n667 ) );
  IV U2489 ( .A(\b/n3325 ), .Z(\b/n666 ) );
  IV U2490 ( .A(msg[52]), .Z(\b/n662 ) );
  IV U2491 ( .A(\b/n3637 ), .Z(\b/n660 ) );
  IV U2492 ( .A(msg[123]), .Z(\b/n66 ) );
  IV U2493 ( .A(\b/n3318 ), .Z(\b/n659 ) );
  IV U2494 ( .A(\b/n3314 ), .Z(\b/n657 ) );
  IV U2495 ( .A(\b/n3638 ), .Z(\b/n655 ) );
  IV U2496 ( .A(\b/n3641 ), .Z(\b/n654 ) );
  IV U2497 ( .A(\b/n3644 ), .Z(\b/n653 ) );
  IV U2498 ( .A(\b/n3295 ), .Z(\b/n652 ) );
  IV U2499 ( .A(\b/n3435 ), .Z(\b/n651 ) );
  IV U2500 ( .A(\b/n6554 ), .Z(\b/n65 ) );
  IV U2501 ( .A(\b/n3629 ), .Z(\b/n649 ) );
  IV U2502 ( .A(\b/n3627 ), .Z(\b/n648 ) );
  IV U2503 ( .A(\b/n3301 ), .Z(\b/n647 ) );
  IV U2504 ( .A(\b/n3312 ), .Z(\b/n645 ) );
  IV U2505 ( .A(\b/n3305 ), .Z(\b/n644 ) );
  IV U2506 ( .A(\b/n3296 ), .Z(\b/n642 ) );
  IV U2507 ( .A(\b/n3642 ), .Z(\b/n641 ) );
  IV U2508 ( .A(msg[55]), .Z(\b/n640 ) );
  IV U2509 ( .A(\b/n6549 ), .Z(\b/n64 ) );
  IV U2510 ( .A(msg[57]), .Z(\b/n638 ) );
  IV U2511 ( .A(\b/n3690 ), .Z(\b/n636 ) );
  IV U2512 ( .A(\b/n3672 ), .Z(\b/n635 ) );
  IV U2513 ( .A(\b/n3653 ), .Z(\b/n634 ) );
  IV U2514 ( .A(msg[59]), .Z(\b/n633 ) );
  IV U2515 ( .A(\b/n3683 ), .Z(\b/n632 ) );
  IV U2516 ( .A(\b/n3678 ), .Z(\b/n631 ) );
  IV U2517 ( .A(\b/n3709 ), .Z(\b/n630 ) );
  IV U2518 ( .A(\b/n6580 ), .Z(\b/n63 ) );
  IV U2519 ( .A(\b/n3998 ), .Z(\b/n629 ) );
  IV U2520 ( .A(\b/n4005 ), .Z(\b/n628 ) );
  IV U2521 ( .A(\b/n3657 ), .Z(\b/n627 ) );
  IV U2522 ( .A(\b/n3999 ), .Z(\b/n626 ) );
  IV U2523 ( .A(\b/n3665 ), .Z(\b/n625 ) );
  IV U2524 ( .A(\b/n3656 ), .Z(\b/n624 ) );
  IV U2525 ( .A(\b/n3659 ), .Z(\b/n623 ) );
  IV U2526 ( .A(\b/n3669 ), .Z(\b/n622 ) );
  IV U2527 ( .A(\b/n3989 ), .Z(\b/n621 ) );
  IV U2528 ( .A(\b/n3811 ), .Z(\b/n620 ) );
  IV U2529 ( .A(\b/n6869 ), .Z(\b/n62 ) );
  IV U2530 ( .A(\b/n3652 ), .Z(\b/n618 ) );
  IV U2531 ( .A(\b/n3687 ), .Z(\b/n617 ) );
  IV U2532 ( .A(\b/n3681 ), .Z(\b/n616 ) );
  IV U2533 ( .A(\b/n3680 ), .Z(\b/n615 ) );
  IV U2534 ( .A(\b/n3651 ), .Z(\b/n613 ) );
  IV U2535 ( .A(\b/n3650 ), .Z(\b/n612 ) );
  IV U2536 ( .A(\b/n3668 ), .Z(\b/n610 ) );
  IV U2537 ( .A(\b/n6876 ), .Z(\b/n61 ) );
  IV U2538 ( .A(\b/n4004 ), .Z(\b/n609 ) );
  IV U2539 ( .A(\b/n3649 ), .Z(\b/n608 ) );
  IV U2540 ( .A(\b/n3667 ), .Z(\b/n605 ) );
  IV U2541 ( .A(\b/n3676 ), .Z(\b/n603 ) );
  IV U2542 ( .A(\b/n3679 ), .Z(\b/n602 ) );
  IV U2543 ( .A(\b/n6528 ), .Z(\b/n60 ) );
  IV U2544 ( .A(\b/n6535 ), .Z(\b/n6 ) );
  IV U2545 ( .A(\b/n3992 ), .Z(\b/n599 ) );
  IV U2546 ( .A(\b/n4006 ), .Z(\b/n598 ) );
  IV U2547 ( .A(\b/n3648 ), .Z(\b/n597 ) );
  IV U2548 ( .A(\b/n3686 ), .Z(\b/n596 ) );
  IV U2549 ( .A(\b/n3684 ), .Z(\b/n595 ) );
  IV U2550 ( .A(msg[60]), .Z(\b/n591 ) );
  IV U2551 ( .A(\b/n6870 ), .Z(\b/n59 ) );
  IV U2552 ( .A(\b/n3996 ), .Z(\b/n589 ) );
  IV U2553 ( .A(\b/n3677 ), .Z(\b/n588 ) );
  IV U2554 ( .A(\b/n3673 ), .Z(\b/n586 ) );
  IV U2555 ( .A(\b/n3997 ), .Z(\b/n584 ) );
  IV U2556 ( .A(\b/n4000 ), .Z(\b/n583 ) );
  IV U2557 ( .A(\b/n4003 ), .Z(\b/n582 ) );
  IV U2558 ( .A(\b/n3654 ), .Z(\b/n581 ) );
  IV U2559 ( .A(\b/n3794 ), .Z(\b/n580 ) );
  IV U2560 ( .A(\b/n6536 ), .Z(\b/n58 ) );
  IV U2561 ( .A(\b/n3988 ), .Z(\b/n578 ) );
  IV U2562 ( .A(\b/n3986 ), .Z(\b/n577 ) );
  IV U2563 ( .A(\b/n3660 ), .Z(\b/n576 ) );
  IV U2564 ( .A(\b/n3671 ), .Z(\b/n574 ) );
  IV U2565 ( .A(\b/n3664 ), .Z(\b/n573 ) );
  IV U2566 ( .A(\b/n3655 ), .Z(\b/n571 ) );
  IV U2567 ( .A(\b/n4001 ), .Z(\b/n570 ) );
  IV U2568 ( .A(\b/n6527 ), .Z(\b/n57 ) );
  IV U2569 ( .A(msg[63]), .Z(\b/n569 ) );
  IV U2570 ( .A(msg[65]), .Z(\b/n567 ) );
  IV U2571 ( .A(\b/n4049 ), .Z(\b/n565 ) );
  IV U2572 ( .A(\b/n4031 ), .Z(\b/n564 ) );
  IV U2573 ( .A(\b/n4012 ), .Z(\b/n563 ) );
  IV U2574 ( .A(msg[67]), .Z(\b/n562 ) );
  IV U2575 ( .A(\b/n4042 ), .Z(\b/n561 ) );
  IV U2576 ( .A(\b/n4037 ), .Z(\b/n560 ) );
  IV U2577 ( .A(\b/n6530 ), .Z(\b/n56 ) );
  IV U2578 ( .A(\b/n4068 ), .Z(\b/n559 ) );
  IV U2579 ( .A(\b/n4357 ), .Z(\b/n558 ) );
  IV U2580 ( .A(\b/n4364 ), .Z(\b/n557 ) );
  IV U2581 ( .A(\b/n4016 ), .Z(\b/n556 ) );
  IV U2582 ( .A(\b/n4358 ), .Z(\b/n555 ) );
  IV U2583 ( .A(\b/n4024 ), .Z(\b/n554 ) );
  IV U2584 ( .A(\b/n4015 ), .Z(\b/n553 ) );
  IV U2585 ( .A(\b/n4018 ), .Z(\b/n552 ) );
  IV U2586 ( .A(\b/n4028 ), .Z(\b/n551 ) );
  IV U2587 ( .A(\b/n4348 ), .Z(\b/n550 ) );
  IV U2588 ( .A(\b/n6540 ), .Z(\b/n55 ) );
  IV U2589 ( .A(\b/n4170 ), .Z(\b/n549 ) );
  IV U2590 ( .A(\b/n4011 ), .Z(\b/n547 ) );
  IV U2591 ( .A(\b/n4046 ), .Z(\b/n546 ) );
  IV U2592 ( .A(\b/n4040 ), .Z(\b/n545 ) );
  IV U2593 ( .A(\b/n4039 ), .Z(\b/n544 ) );
  IV U2594 ( .A(\b/n4010 ), .Z(\b/n542 ) );
  IV U2595 ( .A(\b/n4009 ), .Z(\b/n541 ) );
  IV U2596 ( .A(\b/n6860 ), .Z(\b/n54 ) );
  IV U2597 ( .A(\b/n4027 ), .Z(\b/n539 ) );
  IV U2598 ( .A(\b/n4363 ), .Z(\b/n538 ) );
  IV U2599 ( .A(\b/n4008 ), .Z(\b/n537 ) );
  IV U2600 ( .A(\b/n4026 ), .Z(\b/n534 ) );
  IV U2601 ( .A(\b/n4035 ), .Z(\b/n532 ) );
  IV U2602 ( .A(\b/n4038 ), .Z(\b/n531 ) );
  IV U2603 ( .A(\b/n6682 ), .Z(\b/n53 ) );
  IV U2604 ( .A(\b/n4351 ), .Z(\b/n528 ) );
  IV U2605 ( .A(\b/n4365 ), .Z(\b/n527 ) );
  IV U2606 ( .A(\b/n4007 ), .Z(\b/n526 ) );
  IV U2607 ( .A(\b/n4045 ), .Z(\b/n525 ) );
  IV U2608 ( .A(\b/n4043 ), .Z(\b/n524 ) );
  IV U2609 ( .A(msg[68]), .Z(\b/n520 ) );
  IV U2610 ( .A(\b/n4355 ), .Z(\b/n518 ) );
  IV U2611 ( .A(\b/n4036 ), .Z(\b/n517 ) );
  IV U2612 ( .A(\b/n4032 ), .Z(\b/n515 ) );
  IV U2613 ( .A(\b/n4356 ), .Z(\b/n513 ) );
  IV U2614 ( .A(\b/n4359 ), .Z(\b/n512 ) );
  IV U2615 ( .A(\b/n4362 ), .Z(\b/n511 ) );
  IV U2616 ( .A(\b/n4013 ), .Z(\b/n510 ) );
  IV U2617 ( .A(\b/n6523 ), .Z(\b/n51 ) );
  IV U2618 ( .A(\b/n4153 ), .Z(\b/n509 ) );
  IV U2619 ( .A(\b/n4347 ), .Z(\b/n507 ) );
  IV U2620 ( .A(\b/n4345 ), .Z(\b/n506 ) );
  IV U2621 ( .A(\b/n4019 ), .Z(\b/n505 ) );
  IV U2622 ( .A(\b/n4030 ), .Z(\b/n503 ) );
  IV U2623 ( .A(\b/n4023 ), .Z(\b/n502 ) );
  IV U2624 ( .A(\b/n4014 ), .Z(\b/n500 ) );
  IV U2625 ( .A(\b/n6558 ), .Z(\b/n50 ) );
  IV U2626 ( .A(\b/n4360 ), .Z(\b/n499 ) );
  IV U2627 ( .A(msg[71]), .Z(\b/n498 ) );
  IV U2628 ( .A(msg[73]), .Z(\b/n496 ) );
  IV U2629 ( .A(\b/n4408 ), .Z(\b/n494 ) );
  IV U2630 ( .A(\b/n4390 ), .Z(\b/n493 ) );
  IV U2631 ( .A(\b/n4371 ), .Z(\b/n492 ) );
  IV U2632 ( .A(msg[75]), .Z(\b/n491 ) );
  IV U2633 ( .A(\b/n4401 ), .Z(\b/n490 ) );
  IV U2634 ( .A(\b/n6552 ), .Z(\b/n49 ) );
  IV U2635 ( .A(\b/n4396 ), .Z(\b/n489 ) );
  IV U2636 ( .A(\b/n4427 ), .Z(\b/n488 ) );
  IV U2637 ( .A(\b/n4716 ), .Z(\b/n487 ) );
  IV U2638 ( .A(\b/n4723 ), .Z(\b/n486 ) );
  IV U2639 ( .A(\b/n4375 ), .Z(\b/n485 ) );
  IV U2640 ( .A(\b/n4717 ), .Z(\b/n484 ) );
  IV U2641 ( .A(\b/n4383 ), .Z(\b/n483 ) );
  IV U2642 ( .A(\b/n4374 ), .Z(\b/n482 ) );
  IV U2643 ( .A(\b/n4377 ), .Z(\b/n481 ) );
  IV U2644 ( .A(\b/n4387 ), .Z(\b/n480 ) );
  IV U2645 ( .A(\b/n6551 ), .Z(\b/n48 ) );
  IV U2646 ( .A(\b/n4707 ), .Z(\b/n479 ) );
  IV U2647 ( .A(\b/n4529 ), .Z(\b/n478 ) );
  IV U2648 ( .A(\b/n4370 ), .Z(\b/n476 ) );
  IV U2649 ( .A(\b/n4405 ), .Z(\b/n475 ) );
  IV U2650 ( .A(\b/n4399 ), .Z(\b/n474 ) );
  IV U2651 ( .A(\b/n4398 ), .Z(\b/n473 ) );
  IV U2652 ( .A(\b/n4369 ), .Z(\b/n471 ) );
  IV U2653 ( .A(\b/n4368 ), .Z(\b/n470 ) );
  IV U2654 ( .A(\b/n4386 ), .Z(\b/n468 ) );
  IV U2655 ( .A(\b/n4722 ), .Z(\b/n467 ) );
  IV U2656 ( .A(\b/n4367 ), .Z(\b/n466 ) );
  IV U2657 ( .A(\b/n4385 ), .Z(\b/n463 ) );
  IV U2658 ( .A(\b/n4394 ), .Z(\b/n461 ) );
  IV U2659 ( .A(\b/n4397 ), .Z(\b/n460 ) );
  IV U2660 ( .A(\b/n6522 ), .Z(\b/n46 ) );
  IV U2661 ( .A(\b/n4710 ), .Z(\b/n457 ) );
  IV U2662 ( .A(\b/n4724 ), .Z(\b/n456 ) );
  IV U2663 ( .A(\b/n4366 ), .Z(\b/n455 ) );
  IV U2664 ( .A(\b/n4404 ), .Z(\b/n454 ) );
  IV U2665 ( .A(\b/n4402 ), .Z(\b/n453 ) );
  IV U2666 ( .A(\b/n6521 ), .Z(\b/n45 ) );
  IV U2667 ( .A(msg[76]), .Z(\b/n449 ) );
  IV U2668 ( .A(\b/n4714 ), .Z(\b/n447 ) );
  IV U2669 ( .A(\b/n4395 ), .Z(\b/n446 ) );
  IV U2670 ( .A(\b/n4391 ), .Z(\b/n444 ) );
  IV U2671 ( .A(\b/n4715 ), .Z(\b/n442 ) );
  IV U2672 ( .A(\b/n4718 ), .Z(\b/n441 ) );
  IV U2673 ( .A(\b/n4721 ), .Z(\b/n440 ) );
  IV U2674 ( .A(\b/n4372 ), .Z(\b/n439 ) );
  IV U2675 ( .A(\b/n4512 ), .Z(\b/n438 ) );
  IV U2676 ( .A(\b/n4706 ), .Z(\b/n436 ) );
  IV U2677 ( .A(\b/n4704 ), .Z(\b/n435 ) );
  IV U2678 ( .A(\b/n4378 ), .Z(\b/n434 ) );
  IV U2679 ( .A(\b/n4389 ), .Z(\b/n432 ) );
  IV U2680 ( .A(\b/n4382 ), .Z(\b/n431 ) );
  IV U2681 ( .A(\b/n6539 ), .Z(\b/n43 ) );
  IV U2682 ( .A(\b/n4373 ), .Z(\b/n429 ) );
  IV U2683 ( .A(\b/n4719 ), .Z(\b/n428 ) );
  IV U2684 ( .A(msg[79]), .Z(\b/n427 ) );
  IV U2685 ( .A(msg[81]), .Z(\b/n425 ) );
  IV U2686 ( .A(\b/n4767 ), .Z(\b/n423 ) );
  IV U2687 ( .A(\b/n4749 ), .Z(\b/n422 ) );
  IV U2688 ( .A(\b/n4730 ), .Z(\b/n421 ) );
  IV U2689 ( .A(msg[83]), .Z(\b/n420 ) );
  IV U2690 ( .A(\b/n6875 ), .Z(\b/n42 ) );
  IV U2691 ( .A(\b/n4760 ), .Z(\b/n419 ) );
  IV U2692 ( .A(\b/n4755 ), .Z(\b/n418 ) );
  IV U2693 ( .A(\b/n4786 ), .Z(\b/n417 ) );
  IV U2694 ( .A(\b/n5075 ), .Z(\b/n416 ) );
  IV U2695 ( .A(\b/n5082 ), .Z(\b/n415 ) );
  IV U2696 ( .A(\b/n4734 ), .Z(\b/n414 ) );
  IV U2697 ( .A(\b/n5076 ), .Z(\b/n413 ) );
  IV U2698 ( .A(\b/n4742 ), .Z(\b/n412 ) );
  IV U2699 ( .A(\b/n4733 ), .Z(\b/n411 ) );
  IV U2700 ( .A(\b/n4736 ), .Z(\b/n410 ) );
  IV U2701 ( .A(\b/n6520 ), .Z(\b/n41 ) );
  IV U2702 ( .A(\b/n4746 ), .Z(\b/n409 ) );
  IV U2703 ( .A(\b/n5066 ), .Z(\b/n408 ) );
  IV U2704 ( .A(\b/n4888 ), .Z(\b/n407 ) );
  IV U2705 ( .A(\b/n4729 ), .Z(\b/n405 ) );
  IV U2706 ( .A(\b/n4764 ), .Z(\b/n404 ) );
  IV U2707 ( .A(\b/n4758 ), .Z(\b/n403 ) );
  IV U2708 ( .A(\b/n4757 ), .Z(\b/n402 ) );
  IV U2709 ( .A(\b/n4728 ), .Z(\b/n400 ) );
  IV U2710 ( .A(\b/n6526 ), .Z(\b/n4 ) );
  IV U2711 ( .A(\b/n4727 ), .Z(\b/n399 ) );
  IV U2712 ( .A(\b/n4745 ), .Z(\b/n397 ) );
  IV U2713 ( .A(\b/n5081 ), .Z(\b/n396 ) );
  IV U2714 ( .A(\b/n4726 ), .Z(\b/n395 ) );
  IV U2715 ( .A(\b/n4744 ), .Z(\b/n392 ) );
  IV U2716 ( .A(\b/n4753 ), .Z(\b/n390 ) );
  IV U2717 ( .A(\b/n4756 ), .Z(\b/n389 ) );
  IV U2718 ( .A(\b/n5069 ), .Z(\b/n386 ) );
  IV U2719 ( .A(\b/n5083 ), .Z(\b/n385 ) );
  IV U2720 ( .A(\b/n4725 ), .Z(\b/n384 ) );
  IV U2721 ( .A(\b/n4763 ), .Z(\b/n383 ) );
  IV U2722 ( .A(\b/n4761 ), .Z(\b/n382 ) );
  IV U2723 ( .A(\b/n6538 ), .Z(\b/n38 ) );
  IV U2724 ( .A(msg[84]), .Z(\b/n378 ) );
  IV U2725 ( .A(\b/n5073 ), .Z(\b/n376 ) );
  IV U2726 ( .A(\b/n4754 ), .Z(\b/n375 ) );
  IV U2727 ( .A(\b/n4750 ), .Z(\b/n373 ) );
  IV U2728 ( .A(\b/n5074 ), .Z(\b/n371 ) );
  IV U2729 ( .A(\b/n5077 ), .Z(\b/n370 ) );
  IV U2730 ( .A(\b/n5080 ), .Z(\b/n369 ) );
  IV U2731 ( .A(\b/n4731 ), .Z(\b/n368 ) );
  IV U2732 ( .A(\b/n4871 ), .Z(\b/n367 ) );
  IV U2733 ( .A(\b/n5065 ), .Z(\b/n365 ) );
  IV U2734 ( .A(\b/n5063 ), .Z(\b/n364 ) );
  IV U2735 ( .A(\b/n4737 ), .Z(\b/n363 ) );
  IV U2736 ( .A(\b/n4748 ), .Z(\b/n361 ) );
  IV U2737 ( .A(\b/n4741 ), .Z(\b/n360 ) );
  IV U2738 ( .A(\b/n6547 ), .Z(\b/n36 ) );
  IV U2739 ( .A(\b/n4732 ), .Z(\b/n358 ) );
  IV U2740 ( .A(\b/n5078 ), .Z(\b/n357 ) );
  IV U2741 ( .A(msg[87]), .Z(\b/n356 ) );
  IV U2742 ( .A(msg[89]), .Z(\b/n354 ) );
  IV U2743 ( .A(\b/n5126 ), .Z(\b/n352 ) );
  IV U2744 ( .A(\b/n5108 ), .Z(\b/n351 ) );
  IV U2745 ( .A(\b/n5089 ), .Z(\b/n350 ) );
  IV U2746 ( .A(\b/n6550 ), .Z(\b/n35 ) );
  IV U2747 ( .A(msg[91]), .Z(\b/n349 ) );
  IV U2748 ( .A(\b/n5119 ), .Z(\b/n348 ) );
  IV U2749 ( .A(\b/n5114 ), .Z(\b/n347 ) );
  IV U2750 ( .A(\b/n5145 ), .Z(\b/n346 ) );
  IV U2751 ( .A(\b/n5434 ), .Z(\b/n345 ) );
  IV U2752 ( .A(\b/n5441 ), .Z(\b/n344 ) );
  IV U2753 ( .A(\b/n5093 ), .Z(\b/n343 ) );
  IV U2754 ( .A(\b/n5435 ), .Z(\b/n342 ) );
  IV U2755 ( .A(\b/n5101 ), .Z(\b/n341 ) );
  IV U2756 ( .A(\b/n5092 ), .Z(\b/n340 ) );
  IV U2757 ( .A(\b/n5095 ), .Z(\b/n339 ) );
  IV U2758 ( .A(\b/n5105 ), .Z(\b/n338 ) );
  IV U2759 ( .A(\b/n5425 ), .Z(\b/n337 ) );
  IV U2760 ( .A(\b/n5247 ), .Z(\b/n336 ) );
  IV U2761 ( .A(\b/n5088 ), .Z(\b/n334 ) );
  IV U2762 ( .A(\b/n5123 ), .Z(\b/n333 ) );
  IV U2763 ( .A(\b/n5117 ), .Z(\b/n332 ) );
  IV U2764 ( .A(\b/n5116 ), .Z(\b/n331 ) );
  IV U2765 ( .A(\b/n5087 ), .Z(\b/n329 ) );
  IV U2766 ( .A(\b/n5086 ), .Z(\b/n328 ) );
  IV U2767 ( .A(\b/n5104 ), .Z(\b/n326 ) );
  IV U2768 ( .A(\b/n5440 ), .Z(\b/n325 ) );
  IV U2769 ( .A(\b/n5085 ), .Z(\b/n324 ) );
  IV U2770 ( .A(\b/n5103 ), .Z(\b/n321 ) );
  IV U2771 ( .A(\b/n6863 ), .Z(\b/n32 ) );
  IV U2772 ( .A(\b/n5112 ), .Z(\b/n319 ) );
  IV U2773 ( .A(\b/n5115 ), .Z(\b/n318 ) );
  IV U2774 ( .A(\b/n5428 ), .Z(\b/n315 ) );
  IV U2775 ( .A(\b/n5442 ), .Z(\b/n314 ) );
  IV U2776 ( .A(\b/n5084 ), .Z(\b/n313 ) );
  IV U2777 ( .A(\b/n5122 ), .Z(\b/n312 ) );
  IV U2778 ( .A(\b/n5120 ), .Z(\b/n311 ) );
  IV U2779 ( .A(\b/n6877 ), .Z(\b/n31 ) );
  IV U2780 ( .A(msg[92]), .Z(\b/n307 ) );
  IV U2781 ( .A(\b/n5432 ), .Z(\b/n305 ) );
  IV U2782 ( .A(\b/n5113 ), .Z(\b/n304 ) );
  IV U2783 ( .A(\b/n5109 ), .Z(\b/n302 ) );
  IV U2784 ( .A(\b/n5433 ), .Z(\b/n300 ) );
  IV U2785 ( .A(\b/n6519 ), .Z(\b/n30 ) );
  IV U2786 ( .A(\b/n6872 ), .Z(\b/n3 ) );
  IV U2787 ( .A(\b/n5436 ), .Z(\b/n299 ) );
  IV U2788 ( .A(\b/n5439 ), .Z(\b/n298 ) );
  IV U2789 ( .A(\b/n5090 ), .Z(\b/n297 ) );
  IV U2790 ( .A(\b/n5230 ), .Z(\b/n296 ) );
  IV U2791 ( .A(\b/n5424 ), .Z(\b/n294 ) );
  IV U2792 ( .A(\b/n5422 ), .Z(\b/n293 ) );
  IV U2793 ( .A(\b/n5096 ), .Z(\b/n292 ) );
  IV U2794 ( .A(\b/n5107 ), .Z(\b/n290 ) );
  IV U2795 ( .A(\b/n6557 ), .Z(\b/n29 ) );
  IV U2796 ( .A(\b/n5100 ), .Z(\b/n289 ) );
  IV U2797 ( .A(\b/n5091 ), .Z(\b/n287 ) );
  IV U2798 ( .A(\b/n5437 ), .Z(\b/n286 ) );
  IV U2799 ( .A(msg[95]), .Z(\b/n285 ) );
  IV U2800 ( .A(msg[97]), .Z(\b/n283 ) );
  IV U2801 ( .A(\b/n5469 ), .Z(\b/n281 ) );
  IV U2802 ( .A(\b/n5450 ), .Z(\b/n280 ) );
  IV U2803 ( .A(\b/n6555 ), .Z(\b/n28 ) );
  IV U2804 ( .A(\b/n5447 ), .Z(\b/n279 ) );
  IV U2805 ( .A(msg[99]), .Z(\b/n278 ) );
  IV U2806 ( .A(\b/n5791 ), .Z(\b/n277 ) );
  IV U2807 ( .A(\b/n5794 ), .Z(\b/n276 ) );
  IV U2808 ( .A(\b/n5468 ), .Z(\b/n275 ) );
  IV U2809 ( .A(\b/n5782 ), .Z(\b/n274 ) );
  IV U2810 ( .A(\b/n5779 ), .Z(\b/n273 ) );
  IV U2811 ( .A(\b/n5466 ), .Z(\b/n272 ) );
  IV U2812 ( .A(\b/n5461 ), .Z(\b/n271 ) );
  IV U2813 ( .A(\b/n5478 ), .Z(\b/n270 ) );
  IV U2814 ( .A(\b/n5475 ), .Z(\b/n269 ) );
  IV U2815 ( .A(\b/n5445 ), .Z(\b/n266 ) );
  IV U2816 ( .A(\b/n5456 ), .Z(\b/n265 ) );
  IV U2817 ( .A(\b/n5463 ), .Z(\b/n264 ) );
  IV U2818 ( .A(\b/n5446 ), .Z(\b/n262 ) );
  IV U2819 ( .A(\b/n5467 ), .Z(\b/n259 ) );
  IV U2820 ( .A(\b/n5448 ), .Z(\b/n258 ) );
  IV U2821 ( .A(\b/n5452 ), .Z(\b/n257 ) );
  IV U2822 ( .A(\b/n5454 ), .Z(\b/n256 ) );
  IV U2823 ( .A(\b/n5464 ), .Z(\b/n255 ) );
  IV U2824 ( .A(\b/n5605 ), .Z(\b/n253 ) );
  IV U2825 ( .A(\b/n5798 ), .Z(\b/n251 ) );
  IV U2826 ( .A(\b/n5449 ), .Z(\b/n250 ) );
  IV U2827 ( .A(\b/n5482 ), .Z(\b/n249 ) );
  IV U2828 ( .A(\b/n5479 ), .Z(\b/n248 ) );
  IV U2829 ( .A(\b/n5476 ), .Z(\b/n247 ) );
  IV U2830 ( .A(\b/n5512 ), .Z(\b/n244 ) );
  IV U2831 ( .A(\b/n5783 ), .Z(\b/n243 ) );
  IV U2832 ( .A(\b/n5792 ), .Z(\b/n242 ) );
  IV U2833 ( .A(\b/n5799 ), .Z(\b/n241 ) );
  IV U2834 ( .A(\b/n5444 ), .Z(\b/n240 ) );
  IV U2835 ( .A(msg[124]), .Z(\b/n24 ) );
  IV U2836 ( .A(\b/n5797 ), .Z(\b/n239 ) );
  IV U2837 ( .A(\b/n5793 ), .Z(\b/n238 ) );
  IV U2838 ( .A(\b/n5462 ), .Z(\b/n237 ) );
  IV U2839 ( .A(\b/n5457 ), .Z(\b/n235 ) );
  IV U2840 ( .A(\b/n5472 ), .Z(\b/n233 ) );
  IV U2841 ( .A(\b/n5474 ), .Z(\b/n232 ) );
  IV U2842 ( .A(\b/n5786 ), .Z(\b/n229 ) );
  IV U2843 ( .A(\b/n5800 ), .Z(\b/n228 ) );
  IV U2844 ( .A(\b/n5443 ), .Z(\b/n227 ) );
  IV U2845 ( .A(\b/n5483 ), .Z(\b/n226 ) );
  IV U2846 ( .A(\b/n5480 ), .Z(\b/n225 ) );
  IV U2847 ( .A(\b/n5451 ), .Z(\b/n221 ) );
  IV U2848 ( .A(msg[100]), .Z(\b/n220 ) );
  IV U2849 ( .A(\b/n6867 ), .Z(\b/n22 ) );
  IV U2850 ( .A(\b/n5580 ), .Z(\b/n218 ) );
  IV U2851 ( .A(\b/n5790 ), .Z(\b/n217 ) );
  IV U2852 ( .A(\b/n5473 ), .Z(\b/n216 ) );
  IV U2853 ( .A(\b/n5795 ), .Z(\b/n215 ) );
  IV U2854 ( .A(msg[105]), .Z(\b/n213 ) );
  IV U2855 ( .A(\b/n5843 ), .Z(\b/n211 ) );
  IV U2856 ( .A(\b/n5825 ), .Z(\b/n210 ) );
  IV U2857 ( .A(\b/n6548 ), .Z(\b/n21 ) );
  IV U2858 ( .A(\b/n5806 ), .Z(\b/n209 ) );
  IV U2859 ( .A(msg[107]), .Z(\b/n208 ) );
  IV U2860 ( .A(\b/n5836 ), .Z(\b/n207 ) );
  IV U2861 ( .A(\b/n5831 ), .Z(\b/n206 ) );
  IV U2862 ( .A(\b/n5862 ), .Z(\b/n205 ) );
  IV U2863 ( .A(\b/n6151 ), .Z(\b/n204 ) );
  IV U2864 ( .A(\b/n6158 ), .Z(\b/n203 ) );
  IV U2865 ( .A(\b/n5810 ), .Z(\b/n202 ) );
  IV U2866 ( .A(\b/n6152 ), .Z(\b/n201 ) );
  IV U2867 ( .A(\b/n5818 ), .Z(\b/n200 ) );
  IV U2868 ( .A(msg[127]), .Z(\b/n2 ) );
  IV U2869 ( .A(\b/n5809 ), .Z(\b/n199 ) );
  IV U2870 ( .A(\b/n5812 ), .Z(\b/n198 ) );
  IV U2871 ( .A(\b/n5822 ), .Z(\b/n197 ) );
  IV U2872 ( .A(\b/n6142 ), .Z(\b/n196 ) );
  IV U2873 ( .A(\b/n5964 ), .Z(\b/n195 ) );
  IV U2874 ( .A(\b/n5805 ), .Z(\b/n193 ) );
  IV U2875 ( .A(\b/n5840 ), .Z(\b/n192 ) );
  IV U2876 ( .A(\b/n5834 ), .Z(\b/n191 ) );
  IV U2877 ( .A(\b/n5833 ), .Z(\b/n190 ) );
  IV U2878 ( .A(\b/n6544 ), .Z(\b/n19 ) );
  IV U2879 ( .A(\b/n5804 ), .Z(\b/n188 ) );
  IV U2880 ( .A(\b/n5803 ), .Z(\b/n187 ) );
  IV U2881 ( .A(\b/n5821 ), .Z(\b/n185 ) );
  IV U2882 ( .A(\b/n6157 ), .Z(\b/n184 ) );
  IV U2883 ( .A(\b/n5802 ), .Z(\b/n183 ) );
  IV U2884 ( .A(\b/n5820 ), .Z(\b/n180 ) );
  IV U2885 ( .A(\b/n5829 ), .Z(\b/n178 ) );
  IV U2886 ( .A(\b/n5832 ), .Z(\b/n177 ) );
  IV U2887 ( .A(\b/n6145 ), .Z(\b/n174 ) );
  IV U2888 ( .A(\b/n6159 ), .Z(\b/n173 ) );
  IV U2889 ( .A(\b/n5801 ), .Z(\b/n172 ) );
  IV U2890 ( .A(\b/n5839 ), .Z(\b/n171 ) );
  IV U2891 ( .A(\b/n5837 ), .Z(\b/n170 ) );
  IV U2892 ( .A(\b/n6868 ), .Z(\b/n17 ) );
  IV U2893 ( .A(msg[108]), .Z(\b/n166 ) );
  IV U2894 ( .A(\b/n6149 ), .Z(\b/n164 ) );
  IV U2895 ( .A(\b/n5830 ), .Z(\b/n163 ) );
  IV U2896 ( .A(\b/n5826 ), .Z(\b/n161 ) );
  IV U2897 ( .A(\b/n6871 ), .Z(\b/n16 ) );
  IV U2898 ( .A(\b/n6150 ), .Z(\b/n159 ) );
  IV U2899 ( .A(\b/n6153 ), .Z(\b/n158 ) );
  IV U2900 ( .A(\b/n6156 ), .Z(\b/n157 ) );
  IV U2901 ( .A(\b/n5807 ), .Z(\b/n156 ) );
  IV U2902 ( .A(\b/n5947 ), .Z(\b/n155 ) );
  IV U2903 ( .A(\b/n6141 ), .Z(\b/n153 ) );
  IV U2904 ( .A(\b/n6139 ), .Z(\b/n152 ) );
  IV U2905 ( .A(\b/n5813 ), .Z(\b/n151 ) );
  IV U2906 ( .A(\b/n6874 ), .Z(\b/n15 ) );
  IV U2907 ( .A(\b/n5824 ), .Z(\b/n149 ) );
  IV U2908 ( .A(\b/n5817 ), .Z(\b/n148 ) );
  IV U2909 ( .A(\b/n5808 ), .Z(\b/n146 ) );
  IV U2910 ( .A(\b/n6154 ), .Z(\b/n145 ) );
  IV U2911 ( .A(msg[111]), .Z(\b/n144 ) );
  IV U2912 ( .A(msg[113]), .Z(\b/n142 ) );
  IV U2913 ( .A(\b/n6202 ), .Z(\b/n140 ) );
  IV U2914 ( .A(\b/n6525 ), .Z(\b/n14 ) );
  IV U2915 ( .A(\b/n6184 ), .Z(\b/n139 ) );
  IV U2916 ( .A(\b/n6165 ), .Z(\b/n138 ) );
  IV U2917 ( .A(msg[115]), .Z(\b/n137 ) );
  IV U2918 ( .A(\b/n6195 ), .Z(\b/n136 ) );
  IV U2919 ( .A(\b/n6190 ), .Z(\b/n135 ) );
  IV U2920 ( .A(\b/n6221 ), .Z(\b/n134 ) );
  IV U2921 ( .A(\b/n6510 ), .Z(\b/n133 ) );
  IV U2922 ( .A(\b/n6517 ), .Z(\b/n132 ) );
  IV U2923 ( .A(\b/n6169 ), .Z(\b/n131 ) );
  IV U2924 ( .A(\b/n6511 ), .Z(\b/n130 ) );
  IV U2925 ( .A(\b/n6665 ), .Z(\b/n13 ) );
  IV U2926 ( .A(\b/n6177 ), .Z(\b/n129 ) );
  IV U2927 ( .A(\b/n6168 ), .Z(\b/n128 ) );
  IV U2928 ( .A(\b/n6171 ), .Z(\b/n127 ) );
  IV U2929 ( .A(\b/n6181 ), .Z(\b/n126 ) );
  IV U2930 ( .A(\b/n6501 ), .Z(\b/n125 ) );
  IV U2931 ( .A(\b/n6323 ), .Z(\b/n124 ) );
  IV U2932 ( .A(\b/n6164 ), .Z(\b/n122 ) );
  IV U2933 ( .A(\b/n6199 ), .Z(\b/n121 ) );
  IV U2934 ( .A(\b/n6193 ), .Z(\b/n120 ) );
  IV U2935 ( .A(\b/n6192 ), .Z(\b/n119 ) );
  IV U2936 ( .A(\b/n6163 ), .Z(\b/n117 ) );
  IV U2937 ( .A(\b/n6162 ), .Z(\b/n116 ) );
  IV U2938 ( .A(\b/n6180 ), .Z(\b/n114 ) );
  IV U2939 ( .A(msg[1]), .Z(\b/n1134 ) );
  IV U2940 ( .A(\b/n1177 ), .Z(\b/n1132 ) );
  IV U2941 ( .A(\b/n1159 ), .Z(\b/n1131 ) );
  IV U2942 ( .A(\b/n1140 ), .Z(\b/n1130 ) );
  IV U2943 ( .A(\b/n6516 ), .Z(\b/n113 ) );
  IV U2944 ( .A(msg[3]), .Z(\b/n1129 ) );
  IV U2945 ( .A(\b/n1170 ), .Z(\b/n1128 ) );
  IV U2946 ( .A(\b/n1165 ), .Z(\b/n1127 ) );
  IV U2947 ( .A(\b/n1196 ), .Z(\b/n1126 ) );
  IV U2948 ( .A(\b/n1485 ), .Z(\b/n1125 ) );
  IV U2949 ( .A(\b/n1492 ), .Z(\b/n1124 ) );
  IV U2950 ( .A(\b/n1144 ), .Z(\b/n1123 ) );
  IV U2951 ( .A(\b/n1486 ), .Z(\b/n1122 ) );
  IV U2952 ( .A(\b/n1152 ), .Z(\b/n1121 ) );
  IV U2953 ( .A(\b/n1143 ), .Z(\b/n1120 ) );
  IV U2954 ( .A(\b/n6161 ), .Z(\b/n112 ) );
  IV U2955 ( .A(\b/n1146 ), .Z(\b/n1119 ) );
  IV U2956 ( .A(\b/n1156 ), .Z(\b/n1118 ) );
  IV U2957 ( .A(\b/n1476 ), .Z(\b/n1117 ) );
  IV U2958 ( .A(\b/n1298 ), .Z(\b/n1116 ) );
  IV U2959 ( .A(\b/n1139 ), .Z(\b/n1114 ) );
  IV U2960 ( .A(\b/n1174 ), .Z(\b/n1113 ) );
  IV U2961 ( .A(\b/n1168 ), .Z(\b/n1112 ) );
  IV U2962 ( .A(\b/n1167 ), .Z(\b/n1111 ) );
  IV U2963 ( .A(\b/n1138 ), .Z(\b/n1109 ) );
  IV U2964 ( .A(\b/n1137 ), .Z(\b/n1108 ) );
  IV U2965 ( .A(\b/n1155 ), .Z(\b/n1106 ) );
  IV U2966 ( .A(\b/n1491 ), .Z(\b/n1105 ) );
  IV U2967 ( .A(\b/n1136 ), .Z(\b/n1104 ) );
  IV U2968 ( .A(\b/n1154 ), .Z(\b/n1101 ) );
  IV U2969 ( .A(\b/n6859 ), .Z(\b/n11 ) );
  IV U2970 ( .A(\b/n1163 ), .Z(\b/n1099 ) );
  IV U2971 ( .A(\b/n1166 ), .Z(\b/n1098 ) );
  IV U2972 ( .A(\b/n1479 ), .Z(\b/n1095 ) );
  IV U2973 ( .A(\b/n1493 ), .Z(\b/n1094 ) );
  IV U2974 ( .A(\b/n1135 ), .Z(\b/n1093 ) );
  IV U2975 ( .A(\b/n1173 ), .Z(\b/n1092 ) );
  IV U2976 ( .A(\b/n1171 ), .Z(\b/n1091 ) );
  IV U2977 ( .A(\b/n6179 ), .Z(\b/n109 ) );
  IV U2978 ( .A(msg[4]), .Z(\b/n1087 ) );
  IV U2979 ( .A(\b/n1483 ), .Z(\b/n1085 ) );
  IV U2980 ( .A(\b/n1164 ), .Z(\b/n1084 ) );
  IV U2981 ( .A(\b/n1160 ), .Z(\b/n1082 ) );
  IV U2982 ( .A(\b/n1484 ), .Z(\b/n1080 ) );
  IV U2983 ( .A(\b/n1487 ), .Z(\b/n1079 ) );
  IV U2984 ( .A(\b/n1490 ), .Z(\b/n1078 ) );
  IV U2985 ( .A(\b/n1141 ), .Z(\b/n1077 ) );
  IV U2986 ( .A(\b/n1281 ), .Z(\b/n1076 ) );
  IV U2987 ( .A(\b/n1475 ), .Z(\b/n1074 ) );
  IV U2988 ( .A(\b/n1473 ), .Z(\b/n1073 ) );
  IV U2989 ( .A(\b/n1147 ), .Z(\b/n1072 ) );
  IV U2990 ( .A(\b/n1158 ), .Z(\b/n1070 ) );
  IV U2991 ( .A(\b/n6188 ), .Z(\b/n107 ) );
  IV U2992 ( .A(\b/n1151 ), .Z(\b/n1069 ) );
  IV U2993 ( .A(\b/n1142 ), .Z(\b/n1067 ) );
  IV U2994 ( .A(\b/n1488 ), .Z(\b/n1066 ) );
  IV U2995 ( .A(msg[7]), .Z(\b/n1065 ) );
  IV U2996 ( .A(msg[9]), .Z(\b/n1063 ) );
  IV U2997 ( .A(\b/n1533 ), .Z(\b/n1061 ) );
  IV U2998 ( .A(\b/n1520 ), .Z(\b/n1060 ) );
  IV U2999 ( .A(\b/n6191 ), .Z(\b/n106 ) );
  IV U3000 ( .A(\b/n1499 ), .Z(\b/n1059 ) );
  IV U3001 ( .A(msg[11]), .Z(\b/n1058 ) );
  IV U3002 ( .A(\b/n1524 ), .Z(\b/n1056 ) );
  IV U3003 ( .A(\b/n1496 ), .Z(\b/n1055 ) );
  IV U3004 ( .A(\b/n1507 ), .Z(\b/n1054 ) );
  IV U3005 ( .A(\b/n1514 ), .Z(\b/n1053 ) );
  IV U3006 ( .A(\b/n1497 ), .Z(\b/n1052 ) );
  IV U3007 ( .A(\b/n1500 ), .Z(\b/n1049 ) );
  IV U3008 ( .A(\b/n1503 ), .Z(\b/n1048 ) );
  IV U3009 ( .A(\b/n1505 ), .Z(\b/n1047 ) );
  IV U3010 ( .A(\b/n1515 ), .Z(\b/n1046 ) );
  IV U3011 ( .A(\b/n1657 ), .Z(\b/n1045 ) );
  IV U3012 ( .A(\b/n1850 ), .Z(\b/n1043 ) );
  IV U3013 ( .A(\b/n1501 ), .Z(\b/n1042 ) );
  IV U3014 ( .A(\b/n1531 ), .Z(\b/n1041 ) );
  IV U3015 ( .A(\b/n1528 ), .Z(\b/n1040 ) );
  IV U3016 ( .A(\b/n1526 ), .Z(\b/n1039 ) );
  IV U3017 ( .A(\b/n1498 ), .Z(\b/n1038 ) );
  IV U3018 ( .A(\b/n1564 ), .Z(\b/n1036 ) );
  IV U3019 ( .A(\b/n1835 ), .Z(\b/n1035 ) );
  IV U3020 ( .A(\b/n1844 ), .Z(\b/n1034 ) );
  IV U3021 ( .A(\b/n1851 ), .Z(\b/n1033 ) );
  IV U3022 ( .A(\b/n1495 ), .Z(\b/n1032 ) );
  IV U3023 ( .A(\b/n1845 ), .Z(\b/n1031 ) );
  IV U3024 ( .A(\b/n1513 ), .Z(\b/n1030 ) );
  IV U3025 ( .A(\b/n6504 ), .Z(\b/n103 ) );
  IV U3026 ( .A(\b/n1522 ), .Z(\b/n1027 ) );
  IV U3027 ( .A(\b/n1525 ), .Z(\b/n1026 ) );
  IV U3028 ( .A(\b/n1838 ), .Z(\b/n1023 ) );
  IV U3029 ( .A(\b/n1852 ), .Z(\b/n1022 ) );
  IV U3030 ( .A(\b/n1494 ), .Z(\b/n1021 ) );
  IV U3031 ( .A(\b/n1532 ), .Z(\b/n1020 ) );
  IV U3032 ( .A(\b/n6518 ), .Z(\b/n102 ) );
  IV U3033 ( .A(\b/n1529 ), .Z(\b/n1019 ) );
  IV U3034 ( .A(msg[12]), .Z(\b/n1015 ) );
  IV U3035 ( .A(\b/n1842 ), .Z(\b/n1013 ) );
  IV U3036 ( .A(\b/n1518 ), .Z(\b/n1012 ) );
  IV U3037 ( .A(\b/n1843 ), .Z(\b/n1010 ) );
  IV U3038 ( .A(\b/n6160 ), .Z(\b/n101 ) );
  IV U3039 ( .A(\b/n1846 ), .Z(\b/n1009 ) );
  IV U3040 ( .A(\b/n1849 ), .Z(\b/n1008 ) );
  IV U3041 ( .A(\b/n1519 ), .Z(\b/n1007 ) );
  IV U3042 ( .A(\b/n1631 ), .Z(\b/n1006 ) );
  IV U3043 ( .A(\b/n1834 ), .Z(\b/n1004 ) );
  IV U3044 ( .A(\b/n1831 ), .Z(\b/n1003 ) );
  IV U3045 ( .A(\b/n1508 ), .Z(\b/n1002 ) );
  IV U3046 ( .A(\b/n1517 ), .Z(\b/n1000 ) );
  IV U3047 ( .A(\b/n6198 ), .Z(\b/n100 ) );
  IV U3048 ( .A(\b/n6857 ), .Z(\b/n10 ) );
  XNOR U3049 ( .A(n1404), .B(n1471), .Z(N7) );
  NOR U3050 ( .A(n1390), .B(n1472), .Z(n1471) );
  IV U3051 ( .A(counter[2]), .Z(n1390) );
  IV U3052 ( .A(counter[3]), .Z(n1404) );
  XNOR U3053 ( .A(counter[2]), .B(n1472), .Z(N6) );
  NANDN U3054 ( .B(n1393), .A(counter[0]), .Z(n1472) );
  XNOR U3055 ( .A(n1393), .B(counter[0]), .Z(N5) );
  IV U3056 ( .A(counter[1]), .Z(n1393) );
endmodule

