
module compare_N16384_CC256 ( clk, rst, x, y, g, e );
  input [63:0] x;
  input [63:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  OR U10 ( .A(n290), .B(n291), .Z(n8) );
  ANDN U11 ( .B(n8), .A(n274), .Z(n9) );
  NOR U12 ( .A(n292), .B(n9), .Z(n10) );
  NANDN U13 ( .A(y[15]), .B(x[15]), .Z(n11) );
  AND U14 ( .A(n10), .B(n11), .Z(n12) );
  NANDN U15 ( .A(y[17]), .B(x[17]), .Z(n13) );
  NANDN U16 ( .A(n12), .B(n293), .Z(n14) );
  NAND U17 ( .A(n13), .B(n14), .Z(n15) );
  OR U18 ( .A(n294), .B(n15), .Z(n16) );
  ANDN U19 ( .B(n16), .A(n273), .Z(n17) );
  NOR U20 ( .A(n295), .B(n17), .Z(n18) );
  NANDN U21 ( .A(y[19]), .B(x[19]), .Z(n19) );
  AND U22 ( .A(n18), .B(n19), .Z(n20) );
  OR U23 ( .A(n272), .B(n20), .Z(n21) );
  NANDN U24 ( .A(y[21]), .B(x[21]), .Z(n22) );
  AND U25 ( .A(n21), .B(n22), .Z(n23) );
  NANDN U26 ( .A(n296), .B(n23), .Z(n297) );
  OR U27 ( .A(n311), .B(n312), .Z(n24) );
  NAND U28 ( .A(n313), .B(n24), .Z(n25) );
  ANDN U29 ( .B(n25), .A(n314), .Z(n26) );
  NANDN U30 ( .A(y[41]), .B(x[41]), .Z(n27) );
  NAND U31 ( .A(n26), .B(n27), .Z(n28) );
  NANDN U32 ( .A(n264), .B(n28), .Z(n29) );
  ANDN U33 ( .B(n29), .A(n315), .Z(n30) );
  NANDN U34 ( .A(y[43]), .B(x[43]), .Z(n31) );
  AND U35 ( .A(n30), .B(n31), .Z(n32) );
  OR U36 ( .A(n263), .B(n32), .Z(n33) );
  ANDN U37 ( .B(n33), .A(n316), .Z(n34) );
  NANDN U38 ( .A(y[45]), .B(x[45]), .Z(n35) );
  NAND U39 ( .A(n34), .B(n35), .Z(n36) );
  ANDN U40 ( .B(n36), .A(n262), .Z(n37) );
  NOR U41 ( .A(n317), .B(n37), .Z(n38) );
  NANDN U42 ( .A(y[47]), .B(x[47]), .Z(n39) );
  NAND U43 ( .A(n38), .B(n39), .Z(n318) );
  XOR U44 ( .A(x[1]), .B(n279), .Z(n40) );
  NANDN U45 ( .A(y[1]), .B(n40), .Z(n41) );
  ANDN U46 ( .B(n41), .A(n280), .Z(n42) );
  NAND U47 ( .A(n279), .B(x[1]), .Z(n43) );
  AND U48 ( .A(n42), .B(n43), .Z(n44) );
  NANDN U49 ( .A(n44), .B(n281), .Z(n45) );
  NANDN U50 ( .A(y[3]), .B(x[3]), .Z(n46) );
  AND U51 ( .A(n45), .B(n46), .Z(n47) );
  NANDN U52 ( .A(n282), .B(n47), .Z(n48) );
  NANDN U53 ( .A(n278), .B(n48), .Z(n283) );
  NAND U54 ( .A(n298), .B(n297), .Z(n49) );
  NANDN U55 ( .A(y[23]), .B(x[23]), .Z(n50) );
  NAND U56 ( .A(n49), .B(n50), .Z(n51) );
  OR U57 ( .A(n299), .B(n51), .Z(n52) );
  AND U58 ( .A(n300), .B(n52), .Z(n53) );
  NOR U59 ( .A(n301), .B(n53), .Z(n54) );
  NANDN U60 ( .A(y[25]), .B(x[25]), .Z(n55) );
  NAND U61 ( .A(n54), .B(n55), .Z(n56) );
  NANDN U62 ( .A(n270), .B(n56), .Z(n57) );
  NANDN U63 ( .A(y[27]), .B(x[27]), .Z(n58) );
  NAND U64 ( .A(n57), .B(n58), .Z(n59) );
  OR U65 ( .A(n302), .B(n59), .Z(n60) );
  ANDN U66 ( .B(n60), .A(n269), .Z(n61) );
  NOR U67 ( .A(n303), .B(n61), .Z(n62) );
  NANDN U68 ( .A(y[29]), .B(x[29]), .Z(n63) );
  NAND U69 ( .A(n62), .B(n63), .Z(n64) );
  NANDN U70 ( .A(n268), .B(n64), .Z(n304) );
  NAND U71 ( .A(n319), .B(n318), .Z(n65) );
  ANDN U72 ( .B(n65), .A(n320), .Z(n66) );
  NANDN U73 ( .A(y[49]), .B(x[49]), .Z(n67) );
  NAND U74 ( .A(n66), .B(n67), .Z(n68) );
  NANDN U75 ( .A(n261), .B(n68), .Z(n69) );
  ANDN U76 ( .B(n69), .A(n321), .Z(n70) );
  NANDN U77 ( .A(y[51]), .B(x[51]), .Z(n71) );
  AND U78 ( .A(n70), .B(n71), .Z(n72) );
  OR U79 ( .A(n260), .B(n72), .Z(n73) );
  ANDN U80 ( .B(n73), .A(n322), .Z(n74) );
  NANDN U81 ( .A(y[53]), .B(x[53]), .Z(n75) );
  NAND U82 ( .A(n74), .B(n75), .Z(n76) );
  ANDN U83 ( .B(n76), .A(n259), .Z(n77) );
  NOR U84 ( .A(n323), .B(n77), .Z(n78) );
  NANDN U85 ( .A(y[55]), .B(x[55]), .Z(n79) );
  NAND U86 ( .A(n78), .B(n79), .Z(n80) );
  NAND U87 ( .A(n324), .B(n80), .Z(n325) );
  NOR U88 ( .A(n285), .B(n284), .Z(n81) );
  NAND U89 ( .A(n283), .B(n81), .Z(n82) );
  NANDN U90 ( .A(n277), .B(n82), .Z(n83) );
  ANDN U91 ( .B(n83), .A(n286), .Z(n84) );
  NANDN U92 ( .A(y[7]), .B(x[7]), .Z(n85) );
  AND U93 ( .A(n84), .B(n85), .Z(n86) );
  NANDN U94 ( .A(y[9]), .B(x[9]), .Z(n87) );
  NANDN U95 ( .A(n86), .B(n287), .Z(n88) );
  NAND U96 ( .A(n87), .B(n88), .Z(n89) );
  OR U97 ( .A(n288), .B(n89), .Z(n90) );
  ANDN U98 ( .B(n90), .A(n276), .Z(n91) );
  NOR U99 ( .A(n289), .B(n91), .Z(n92) );
  NANDN U100 ( .A(y[11]), .B(x[11]), .Z(n93) );
  NAND U101 ( .A(n92), .B(n93), .Z(n94) );
  NANDN U102 ( .A(n275), .B(n94), .Z(n95) );
  NANDN U103 ( .A(y[13]), .B(x[13]), .Z(n96) );
  NAND U104 ( .A(n95), .B(n96), .Z(n291) );
  ANDN U105 ( .B(n304), .A(n305), .Z(n97) );
  NANDN U106 ( .A(y[31]), .B(x[31]), .Z(n98) );
  AND U107 ( .A(n97), .B(n98), .Z(n99) );
  NANDN U108 ( .A(n99), .B(n306), .Z(n100) );
  ANDN U109 ( .B(n100), .A(n307), .Z(n101) );
  NANDN U110 ( .A(y[33]), .B(x[33]), .Z(n102) );
  NAND U111 ( .A(n101), .B(n102), .Z(n103) );
  NANDN U112 ( .A(n267), .B(n103), .Z(n104) );
  ANDN U113 ( .B(n104), .A(n308), .Z(n105) );
  NANDN U114 ( .A(y[35]), .B(x[35]), .Z(n106) );
  AND U115 ( .A(n105), .B(n106), .Z(n107) );
  OR U116 ( .A(n266), .B(n107), .Z(n108) );
  ANDN U117 ( .B(n108), .A(n309), .Z(n109) );
  NANDN U118 ( .A(y[37]), .B(x[37]), .Z(n110) );
  NAND U119 ( .A(n109), .B(n110), .Z(n111) );
  NANDN U120 ( .A(n265), .B(n111), .Z(n112) );
  NANDN U121 ( .A(n310), .B(n112), .Z(n312) );
  AND U122 ( .A(e), .B(n330), .Z(n113) );
  NOR U123 ( .A(n327), .B(n326), .Z(n114) );
  NAND U124 ( .A(n325), .B(n114), .Z(n115) );
  ANDN U125 ( .B(n115), .A(n258), .Z(n116) );
  NOR U126 ( .A(n328), .B(n116), .Z(n117) );
  NANDN U127 ( .A(y[59]), .B(x[59]), .Z(n118) );
  NAND U128 ( .A(n117), .B(n118), .Z(n119) );
  ANDN U129 ( .B(n119), .A(n257), .Z(n120) );
  NOR U130 ( .A(n329), .B(n120), .Z(n121) );
  NANDN U131 ( .A(y[61]), .B(x[61]), .Z(n122) );
  NAND U132 ( .A(n121), .B(n122), .Z(n123) );
  NANDN U133 ( .A(n256), .B(n123), .Z(n124) );
  NANDN U134 ( .A(y[63]), .B(x[63]), .Z(n125) );
  NAND U135 ( .A(n124), .B(n125), .Z(n126) );
  NAND U136 ( .A(n126), .B(n113), .Z(n127) );
  NANDN U137 ( .A(n113), .B(g), .Z(n128) );
  NAND U138 ( .A(n127), .B(n128), .Z(n4) );
  IV U139 ( .A(ebreg), .Z(e) );
  XNOR U140 ( .A(y[21]), .B(x[21]), .Z(n130) );
  NANDN U141 ( .A(x[20]), .B(y[20]), .Z(n129) );
  NAND U142 ( .A(n130), .B(n129), .Z(n272) );
  XNOR U143 ( .A(y[17]), .B(x[17]), .Z(n132) );
  NANDN U144 ( .A(x[16]), .B(y[16]), .Z(n131) );
  AND U145 ( .A(n132), .B(n131), .Z(n293) );
  XNOR U146 ( .A(y[19]), .B(x[19]), .Z(n134) );
  NANDN U147 ( .A(x[18]), .B(y[18]), .Z(n133) );
  NAND U148 ( .A(n134), .B(n133), .Z(n273) );
  ANDN U149 ( .B(n293), .A(n273), .Z(n137) );
  XNOR U150 ( .A(y[23]), .B(x[23]), .Z(n136) );
  NANDN U151 ( .A(x[22]), .B(y[22]), .Z(n135) );
  NAND U152 ( .A(n136), .B(n135), .Z(n271) );
  ANDN U153 ( .B(n137), .A(n271), .Z(n138) );
  NANDN U154 ( .A(n272), .B(n138), .Z(n175) );
  XNOR U155 ( .A(y[7]), .B(x[7]), .Z(n140) );
  NANDN U156 ( .A(x[6]), .B(y[6]), .Z(n139) );
  NAND U157 ( .A(n140), .B(n139), .Z(n277) );
  XNOR U158 ( .A(y[3]), .B(x[3]), .Z(n142) );
  NANDN U159 ( .A(x[2]), .B(y[2]), .Z(n141) );
  AND U160 ( .A(n142), .B(n141), .Z(n281) );
  XNOR U161 ( .A(y[5]), .B(x[5]), .Z(n144) );
  NANDN U162 ( .A(x[4]), .B(y[4]), .Z(n143) );
  NAND U163 ( .A(n144), .B(n143), .Z(n278) );
  ANDN U164 ( .B(n281), .A(n278), .Z(n148) );
  XNOR U165 ( .A(y[1]), .B(x[1]), .Z(n146) );
  NANDN U166 ( .A(x[0]), .B(y[0]), .Z(n145) );
  NAND U167 ( .A(n146), .B(n145), .Z(n147) );
  ANDN U168 ( .B(n148), .A(n147), .Z(n149) );
  NANDN U169 ( .A(n277), .B(n149), .Z(n161) );
  XNOR U170 ( .A(y[13]), .B(x[13]), .Z(n151) );
  NANDN U171 ( .A(x[12]), .B(y[12]), .Z(n150) );
  NAND U172 ( .A(n151), .B(n150), .Z(n275) );
  XNOR U173 ( .A(y[9]), .B(x[9]), .Z(n153) );
  NANDN U174 ( .A(x[8]), .B(y[8]), .Z(n152) );
  AND U175 ( .A(n153), .B(n152), .Z(n287) );
  XNOR U176 ( .A(y[11]), .B(x[11]), .Z(n155) );
  NANDN U177 ( .A(x[10]), .B(y[10]), .Z(n154) );
  NAND U178 ( .A(n155), .B(n154), .Z(n276) );
  ANDN U179 ( .B(n287), .A(n276), .Z(n158) );
  XNOR U180 ( .A(y[15]), .B(x[15]), .Z(n157) );
  NANDN U181 ( .A(x[14]), .B(y[14]), .Z(n156) );
  NAND U182 ( .A(n157), .B(n156), .Z(n274) );
  ANDN U183 ( .B(n158), .A(n274), .Z(n159) );
  NANDN U184 ( .A(n275), .B(n159), .Z(n160) );
  NOR U185 ( .A(n161), .B(n160), .Z(n173) );
  XNOR U186 ( .A(y[29]), .B(x[29]), .Z(n163) );
  NANDN U187 ( .A(x[28]), .B(y[28]), .Z(n162) );
  NAND U188 ( .A(n163), .B(n162), .Z(n269) );
  XNOR U189 ( .A(y[25]), .B(x[25]), .Z(n165) );
  NANDN U190 ( .A(x[24]), .B(y[24]), .Z(n164) );
  AND U191 ( .A(n165), .B(n164), .Z(n300) );
  XNOR U192 ( .A(y[27]), .B(x[27]), .Z(n167) );
  NANDN U193 ( .A(x[26]), .B(y[26]), .Z(n166) );
  NAND U194 ( .A(n167), .B(n166), .Z(n270) );
  ANDN U195 ( .B(n300), .A(n270), .Z(n170) );
  XNOR U196 ( .A(y[31]), .B(x[31]), .Z(n169) );
  NANDN U197 ( .A(x[30]), .B(y[30]), .Z(n168) );
  NAND U198 ( .A(n169), .B(n168), .Z(n268) );
  ANDN U199 ( .B(n170), .A(n268), .Z(n171) );
  NANDN U200 ( .A(n269), .B(n171), .Z(n172) );
  ANDN U201 ( .B(n173), .A(n172), .Z(n174) );
  NANDN U202 ( .A(n175), .B(n174), .Z(n255) );
  XNOR U203 ( .A(x[45]), .B(y[45]), .Z(n177) );
  NANDN U204 ( .A(x[44]), .B(y[44]), .Z(n176) );
  NAND U205 ( .A(n177), .B(n176), .Z(n263) );
  XNOR U206 ( .A(x[41]), .B(y[41]), .Z(n179) );
  NANDN U207 ( .A(x[40]), .B(y[40]), .Z(n178) );
  AND U208 ( .A(n179), .B(n178), .Z(n313) );
  XNOR U209 ( .A(x[43]), .B(y[43]), .Z(n181) );
  NANDN U210 ( .A(x[42]), .B(y[42]), .Z(n180) );
  NAND U211 ( .A(n181), .B(n180), .Z(n264) );
  ANDN U212 ( .B(n313), .A(n264), .Z(n184) );
  XNOR U213 ( .A(x[47]), .B(y[47]), .Z(n183) );
  NANDN U214 ( .A(x[46]), .B(y[46]), .Z(n182) );
  NAND U215 ( .A(n183), .B(n182), .Z(n262) );
  ANDN U216 ( .B(n184), .A(n262), .Z(n185) );
  NANDN U217 ( .A(n263), .B(n185), .Z(n197) );
  XNOR U218 ( .A(x[37]), .B(y[37]), .Z(n187) );
  NANDN U219 ( .A(x[36]), .B(y[36]), .Z(n186) );
  NAND U220 ( .A(n187), .B(n186), .Z(n266) );
  XNOR U221 ( .A(x[33]), .B(y[33]), .Z(n189) );
  NANDN U222 ( .A(x[32]), .B(y[32]), .Z(n188) );
  AND U223 ( .A(n189), .B(n188), .Z(n306) );
  XNOR U224 ( .A(x[35]), .B(y[35]), .Z(n191) );
  NANDN U225 ( .A(x[34]), .B(y[34]), .Z(n190) );
  NAND U226 ( .A(n191), .B(n190), .Z(n267) );
  ANDN U227 ( .B(n306), .A(n267), .Z(n194) );
  XNOR U228 ( .A(x[39]), .B(y[39]), .Z(n193) );
  NANDN U229 ( .A(x[38]), .B(y[38]), .Z(n192) );
  NAND U230 ( .A(n193), .B(n192), .Z(n265) );
  ANDN U231 ( .B(n194), .A(n265), .Z(n195) );
  NANDN U232 ( .A(n266), .B(n195), .Z(n196) );
  NOR U233 ( .A(n197), .B(n196), .Z(n253) );
  ANDN U234 ( .B(x[60]), .A(y[60]), .Z(n328) );
  ANDN U235 ( .B(x[56]), .A(y[56]), .Z(n323) );
  ANDN U236 ( .B(x[58]), .A(y[58]), .Z(n326) );
  NOR U237 ( .A(n323), .B(n326), .Z(n198) );
  ANDN U238 ( .B(x[62]), .A(y[62]), .Z(n329) );
  ANDN U239 ( .B(n198), .A(n329), .Z(n199) );
  NANDN U240 ( .A(n328), .B(n199), .Z(n211) );
  ANDN U241 ( .B(x[44]), .A(y[44]), .Z(n315) );
  ANDN U242 ( .B(x[40]), .A(y[40]), .Z(n310) );
  ANDN U243 ( .B(x[42]), .A(y[42]), .Z(n314) );
  NOR U244 ( .A(n310), .B(n314), .Z(n200) );
  ANDN U245 ( .B(x[46]), .A(y[46]), .Z(n316) );
  ANDN U246 ( .B(n200), .A(n316), .Z(n201) );
  NANDN U247 ( .A(n315), .B(n201), .Z(n205) );
  ANDN U248 ( .B(x[36]), .A(y[36]), .Z(n308) );
  ANDN U249 ( .B(x[32]), .A(y[32]), .Z(n305) );
  ANDN U250 ( .B(x[34]), .A(y[34]), .Z(n307) );
  NOR U251 ( .A(n305), .B(n307), .Z(n202) );
  ANDN U252 ( .B(x[38]), .A(y[38]), .Z(n309) );
  ANDN U253 ( .B(n202), .A(n309), .Z(n203) );
  NANDN U254 ( .A(n308), .B(n203), .Z(n204) );
  NOR U255 ( .A(n205), .B(n204), .Z(n209) );
  ANDN U256 ( .B(x[52]), .A(y[52]), .Z(n321) );
  ANDN U257 ( .B(x[48]), .A(y[48]), .Z(n317) );
  ANDN U258 ( .B(x[50]), .A(y[50]), .Z(n320) );
  NOR U259 ( .A(n317), .B(n320), .Z(n206) );
  ANDN U260 ( .B(x[54]), .A(y[54]), .Z(n322) );
  ANDN U261 ( .B(n206), .A(n322), .Z(n207) );
  NANDN U262 ( .A(n321), .B(n207), .Z(n208) );
  ANDN U263 ( .B(n209), .A(n208), .Z(n210) );
  NANDN U264 ( .A(n211), .B(n210), .Z(n251) );
  XNOR U265 ( .A(x[61]), .B(y[61]), .Z(n213) );
  NANDN U266 ( .A(x[60]), .B(y[60]), .Z(n212) );
  NAND U267 ( .A(n213), .B(n212), .Z(n257) );
  XNOR U268 ( .A(x[57]), .B(y[57]), .Z(n215) );
  NANDN U269 ( .A(x[56]), .B(y[56]), .Z(n214) );
  AND U270 ( .A(n215), .B(n214), .Z(n324) );
  XNOR U271 ( .A(x[59]), .B(y[59]), .Z(n217) );
  NANDN U272 ( .A(x[58]), .B(y[58]), .Z(n216) );
  NAND U273 ( .A(n217), .B(n216), .Z(n258) );
  ANDN U274 ( .B(n324), .A(n258), .Z(n220) );
  XNOR U275 ( .A(x[63]), .B(y[63]), .Z(n219) );
  NANDN U276 ( .A(x[62]), .B(y[62]), .Z(n218) );
  NAND U277 ( .A(n219), .B(n218), .Z(n256) );
  ANDN U278 ( .B(n220), .A(n256), .Z(n221) );
  NANDN U279 ( .A(n257), .B(n221), .Z(n233) );
  XNOR U280 ( .A(x[53]), .B(y[53]), .Z(n223) );
  NANDN U281 ( .A(x[52]), .B(y[52]), .Z(n222) );
  NAND U282 ( .A(n223), .B(n222), .Z(n260) );
  XNOR U283 ( .A(x[49]), .B(y[49]), .Z(n225) );
  NANDN U284 ( .A(x[48]), .B(y[48]), .Z(n224) );
  AND U285 ( .A(n225), .B(n224), .Z(n319) );
  XNOR U286 ( .A(x[51]), .B(y[51]), .Z(n227) );
  NANDN U287 ( .A(x[50]), .B(y[50]), .Z(n226) );
  NAND U288 ( .A(n227), .B(n226), .Z(n261) );
  ANDN U289 ( .B(n319), .A(n261), .Z(n230) );
  XNOR U290 ( .A(x[55]), .B(y[55]), .Z(n229) );
  NANDN U291 ( .A(x[54]), .B(y[54]), .Z(n228) );
  NAND U292 ( .A(n229), .B(n228), .Z(n259) );
  ANDN U293 ( .B(n230), .A(n259), .Z(n231) );
  NANDN U294 ( .A(n260), .B(n231), .Z(n232) );
  NOR U295 ( .A(n233), .B(n232), .Z(n249) );
  ANDN U296 ( .B(x[28]), .A(y[28]), .Z(n302) );
  ANDN U297 ( .B(x[24]), .A(y[24]), .Z(n299) );
  ANDN U298 ( .B(x[26]), .A(y[26]), .Z(n301) );
  NOR U299 ( .A(n299), .B(n301), .Z(n234) );
  ANDN U300 ( .B(x[30]), .A(y[30]), .Z(n303) );
  ANDN U301 ( .B(n234), .A(n303), .Z(n235) );
  NANDN U302 ( .A(n302), .B(n235), .Z(n247) );
  ANDN U303 ( .B(x[12]), .A(y[12]), .Z(n289) );
  ANDN U304 ( .B(x[8]), .A(y[8]), .Z(n286) );
  ANDN U305 ( .B(x[10]), .A(y[10]), .Z(n288) );
  NOR U306 ( .A(n286), .B(n288), .Z(n236) );
  ANDN U307 ( .B(x[14]), .A(y[14]), .Z(n290) );
  ANDN U308 ( .B(n236), .A(n290), .Z(n237) );
  NANDN U309 ( .A(n289), .B(n237), .Z(n241) );
  ANDN U310 ( .B(x[2]), .A(y[2]), .Z(n280) );
  ANDN U311 ( .B(x[4]), .A(y[4]), .Z(n282) );
  ANDN U312 ( .B(x[0]), .A(y[0]), .Z(n279) );
  NOR U313 ( .A(n282), .B(n279), .Z(n238) );
  ANDN U314 ( .B(x[6]), .A(y[6]), .Z(n285) );
  ANDN U315 ( .B(n238), .A(n285), .Z(n239) );
  NANDN U316 ( .A(n280), .B(n239), .Z(n240) );
  NOR U317 ( .A(n241), .B(n240), .Z(n245) );
  ANDN U318 ( .B(x[20]), .A(y[20]), .Z(n295) );
  ANDN U319 ( .B(x[16]), .A(y[16]), .Z(n292) );
  ANDN U320 ( .B(x[18]), .A(y[18]), .Z(n294) );
  NOR U321 ( .A(n292), .B(n294), .Z(n242) );
  ANDN U322 ( .B(x[22]), .A(y[22]), .Z(n296) );
  ANDN U323 ( .B(n242), .A(n296), .Z(n243) );
  NANDN U324 ( .A(n295), .B(n243), .Z(n244) );
  ANDN U325 ( .B(n245), .A(n244), .Z(n246) );
  NANDN U326 ( .A(n247), .B(n246), .Z(n248) );
  ANDN U327 ( .B(n249), .A(n248), .Z(n250) );
  NANDN U328 ( .A(n251), .B(n250), .Z(n252) );
  ANDN U329 ( .B(n253), .A(n252), .Z(n254) );
  NANDN U330 ( .A(n255), .B(n254), .Z(n330) );
  NANDN U331 ( .A(n330), .B(e), .Z(n5) );
  IV U332 ( .A(n271), .Z(n298) );
  ANDN U333 ( .B(x[5]), .A(y[5]), .Z(n284) );
  ANDN U334 ( .B(x[39]), .A(y[39]), .Z(n311) );
  ANDN U335 ( .B(x[57]), .A(y[57]), .Z(n327) );
endmodule

