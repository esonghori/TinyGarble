
module mult_N64_CC16 ( clk, rst, a, b, c );
  input [63:0] a;
  input [3:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587;
  wire   [127:0] sreg;

  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U7 ( .A(sreg[66]), .B(n465), .Z(n1) );
  XOR U8 ( .A(n465), .B(sreg[66]), .Z(n2) );
  NANDN U9 ( .A(n466), .B(n2), .Z(n3) );
  NAND U10 ( .A(n1), .B(n3), .Z(n484) );
  NAND U11 ( .A(sreg[70]), .B(n541), .Z(n4) );
  XOR U12 ( .A(n541), .B(sreg[70]), .Z(n5) );
  NANDN U13 ( .A(n542), .B(n5), .Z(n6) );
  NAND U14 ( .A(n4), .B(n6), .Z(n560) );
  NAND U15 ( .A(sreg[74]), .B(n617), .Z(n7) );
  XOR U16 ( .A(n617), .B(sreg[74]), .Z(n8) );
  NANDN U17 ( .A(n618), .B(n8), .Z(n9) );
  NAND U18 ( .A(n7), .B(n9), .Z(n636) );
  NAND U19 ( .A(sreg[78]), .B(n693), .Z(n10) );
  XOR U20 ( .A(n693), .B(sreg[78]), .Z(n11) );
  NANDN U21 ( .A(n694), .B(n11), .Z(n12) );
  NAND U22 ( .A(n10), .B(n12), .Z(n712) );
  NAND U23 ( .A(sreg[82]), .B(n769), .Z(n13) );
  XOR U24 ( .A(n769), .B(sreg[82]), .Z(n14) );
  NANDN U25 ( .A(n770), .B(n14), .Z(n15) );
  NAND U26 ( .A(n13), .B(n15), .Z(n788) );
  NAND U27 ( .A(sreg[86]), .B(n845), .Z(n16) );
  XOR U28 ( .A(n845), .B(sreg[86]), .Z(n17) );
  NANDN U29 ( .A(n846), .B(n17), .Z(n18) );
  NAND U30 ( .A(n16), .B(n18), .Z(n864) );
  NAND U31 ( .A(sreg[90]), .B(n921), .Z(n19) );
  XOR U32 ( .A(n921), .B(sreg[90]), .Z(n20) );
  NANDN U33 ( .A(n922), .B(n20), .Z(n21) );
  NAND U34 ( .A(n19), .B(n21), .Z(n940) );
  NAND U35 ( .A(sreg[94]), .B(n997), .Z(n22) );
  XOR U36 ( .A(n997), .B(sreg[94]), .Z(n23) );
  NANDN U37 ( .A(n998), .B(n23), .Z(n24) );
  NAND U38 ( .A(n22), .B(n24), .Z(n1016) );
  NAND U39 ( .A(sreg[98]), .B(n1073), .Z(n25) );
  XOR U40 ( .A(n1073), .B(sreg[98]), .Z(n26) );
  NANDN U41 ( .A(n1074), .B(n26), .Z(n27) );
  NAND U42 ( .A(n25), .B(n27), .Z(n1092) );
  NAND U43 ( .A(sreg[102]), .B(n1149), .Z(n28) );
  XOR U44 ( .A(n1149), .B(sreg[102]), .Z(n29) );
  NANDN U45 ( .A(n1150), .B(n29), .Z(n30) );
  NAND U46 ( .A(n28), .B(n30), .Z(n1168) );
  NAND U47 ( .A(sreg[106]), .B(n1225), .Z(n31) );
  XOR U48 ( .A(n1225), .B(sreg[106]), .Z(n32) );
  NANDN U49 ( .A(n1226), .B(n32), .Z(n33) );
  NAND U50 ( .A(n31), .B(n33), .Z(n1244) );
  NAND U51 ( .A(sreg[110]), .B(n1301), .Z(n34) );
  XOR U52 ( .A(n1301), .B(sreg[110]), .Z(n35) );
  NANDN U53 ( .A(n1302), .B(n35), .Z(n36) );
  NAND U54 ( .A(n34), .B(n36), .Z(n1320) );
  NAND U55 ( .A(sreg[114]), .B(n1377), .Z(n37) );
  XOR U56 ( .A(n1377), .B(sreg[114]), .Z(n38) );
  NANDN U57 ( .A(n1378), .B(n38), .Z(n39) );
  NAND U58 ( .A(n37), .B(n39), .Z(n1396) );
  NAND U59 ( .A(sreg[118]), .B(n1453), .Z(n40) );
  XOR U60 ( .A(n1453), .B(sreg[118]), .Z(n41) );
  NANDN U61 ( .A(n1454), .B(n41), .Z(n42) );
  NAND U62 ( .A(n40), .B(n42), .Z(n1472) );
  AND U63 ( .A(b[1]), .B(a[62]), .Z(n1545) );
  XOR U64 ( .A(n443), .B(n442), .Z(n43) );
  NANDN U65 ( .A(n444), .B(n43), .Z(n44) );
  NAND U66 ( .A(n443), .B(n442), .Z(n45) );
  AND U67 ( .A(n44), .B(n45), .Z(n458) );
  XNOR U68 ( .A(n493), .B(n494), .Z(n495) );
  XNOR U69 ( .A(n512), .B(n513), .Z(n514) );
  XNOR U70 ( .A(n569), .B(n570), .Z(n571) );
  XNOR U71 ( .A(n588), .B(n589), .Z(n590) );
  XNOR U72 ( .A(n645), .B(n646), .Z(n647) );
  XNOR U73 ( .A(n664), .B(n665), .Z(n666) );
  XNOR U74 ( .A(n721), .B(n722), .Z(n723) );
  XNOR U75 ( .A(n740), .B(n741), .Z(n742) );
  XNOR U76 ( .A(n797), .B(n798), .Z(n799) );
  XNOR U77 ( .A(n816), .B(n817), .Z(n818) );
  XNOR U78 ( .A(n873), .B(n874), .Z(n875) );
  XNOR U79 ( .A(n892), .B(n893), .Z(n894) );
  XNOR U80 ( .A(n949), .B(n950), .Z(n951) );
  XNOR U81 ( .A(n968), .B(n969), .Z(n970) );
  XNOR U82 ( .A(n1025), .B(n1026), .Z(n1027) );
  XNOR U83 ( .A(n1044), .B(n1045), .Z(n1046) );
  XNOR U84 ( .A(n1101), .B(n1102), .Z(n1103) );
  XNOR U85 ( .A(n1120), .B(n1121), .Z(n1122) );
  XNOR U86 ( .A(n1177), .B(n1178), .Z(n1179) );
  XNOR U87 ( .A(n1196), .B(n1197), .Z(n1198) );
  XNOR U88 ( .A(n1253), .B(n1254), .Z(n1255) );
  XNOR U89 ( .A(n1272), .B(n1273), .Z(n1274) );
  XNOR U90 ( .A(n1329), .B(n1330), .Z(n1331) );
  XNOR U91 ( .A(n1348), .B(n1349), .Z(n1350) );
  XNOR U92 ( .A(n1405), .B(n1406), .Z(n1407) );
  XNOR U93 ( .A(n1424), .B(n1425), .Z(n1426) );
  XNOR U94 ( .A(n1481), .B(n1482), .Z(n1483) );
  XNOR U95 ( .A(n1500), .B(n1501), .Z(n1502) );
  NAND U96 ( .A(sreg[62]), .B(n377), .Z(n46) );
  XOR U97 ( .A(n377), .B(sreg[62]), .Z(n47) );
  NANDN U98 ( .A(n378), .B(n47), .Z(n48) );
  NAND U99 ( .A(n46), .B(n48), .Z(n400) );
  NAND U100 ( .A(sreg[122]), .B(n1513), .Z(n49) );
  XOR U101 ( .A(n1513), .B(sreg[122]), .Z(n50) );
  NANDN U102 ( .A(n1514), .B(n50), .Z(n51) );
  NAND U103 ( .A(n49), .B(n51), .Z(n1548) );
  NAND U104 ( .A(sreg[67]), .B(n484), .Z(n52) );
  XOR U105 ( .A(n484), .B(sreg[67]), .Z(n53) );
  NANDN U106 ( .A(n485), .B(n53), .Z(n54) );
  NAND U107 ( .A(n52), .B(n54), .Z(n503) );
  NAND U108 ( .A(sreg[71]), .B(n560), .Z(n55) );
  XOR U109 ( .A(n560), .B(sreg[71]), .Z(n56) );
  NANDN U110 ( .A(n561), .B(n56), .Z(n57) );
  NAND U111 ( .A(n55), .B(n57), .Z(n579) );
  NAND U112 ( .A(sreg[75]), .B(n636), .Z(n58) );
  XOR U113 ( .A(n636), .B(sreg[75]), .Z(n59) );
  NANDN U114 ( .A(n637), .B(n59), .Z(n60) );
  NAND U115 ( .A(n58), .B(n60), .Z(n655) );
  NAND U116 ( .A(sreg[79]), .B(n712), .Z(n61) );
  XOR U117 ( .A(n712), .B(sreg[79]), .Z(n62) );
  NANDN U118 ( .A(n713), .B(n62), .Z(n63) );
  NAND U119 ( .A(n61), .B(n63), .Z(n731) );
  NAND U120 ( .A(sreg[83]), .B(n788), .Z(n64) );
  XOR U121 ( .A(n788), .B(sreg[83]), .Z(n65) );
  NANDN U122 ( .A(n789), .B(n65), .Z(n66) );
  NAND U123 ( .A(n64), .B(n66), .Z(n807) );
  NAND U124 ( .A(sreg[87]), .B(n864), .Z(n67) );
  XOR U125 ( .A(n864), .B(sreg[87]), .Z(n68) );
  NANDN U126 ( .A(n865), .B(n68), .Z(n69) );
  NAND U127 ( .A(n67), .B(n69), .Z(n883) );
  NAND U128 ( .A(sreg[91]), .B(n940), .Z(n70) );
  XOR U129 ( .A(n940), .B(sreg[91]), .Z(n71) );
  NANDN U130 ( .A(n941), .B(n71), .Z(n72) );
  NAND U131 ( .A(n70), .B(n72), .Z(n959) );
  NAND U132 ( .A(sreg[95]), .B(n1016), .Z(n73) );
  XOR U133 ( .A(n1016), .B(sreg[95]), .Z(n74) );
  NANDN U134 ( .A(n1017), .B(n74), .Z(n75) );
  NAND U135 ( .A(n73), .B(n75), .Z(n1035) );
  NAND U136 ( .A(sreg[99]), .B(n1092), .Z(n76) );
  XOR U137 ( .A(n1092), .B(sreg[99]), .Z(n77) );
  NANDN U138 ( .A(n1093), .B(n77), .Z(n78) );
  NAND U139 ( .A(n76), .B(n78), .Z(n1111) );
  NAND U140 ( .A(sreg[103]), .B(n1168), .Z(n79) );
  XOR U141 ( .A(n1168), .B(sreg[103]), .Z(n80) );
  NANDN U142 ( .A(n1169), .B(n80), .Z(n81) );
  NAND U143 ( .A(n79), .B(n81), .Z(n1187) );
  NAND U144 ( .A(sreg[107]), .B(n1244), .Z(n82) );
  XOR U145 ( .A(n1244), .B(sreg[107]), .Z(n83) );
  NANDN U146 ( .A(n1245), .B(n83), .Z(n84) );
  NAND U147 ( .A(n82), .B(n84), .Z(n1263) );
  NAND U148 ( .A(sreg[111]), .B(n1320), .Z(n85) );
  XOR U149 ( .A(n1320), .B(sreg[111]), .Z(n86) );
  NANDN U150 ( .A(n1321), .B(n86), .Z(n87) );
  NAND U151 ( .A(n85), .B(n87), .Z(n1339) );
  NAND U152 ( .A(sreg[115]), .B(n1396), .Z(n88) );
  XOR U153 ( .A(n1396), .B(sreg[115]), .Z(n89) );
  NANDN U154 ( .A(n1397), .B(n89), .Z(n90) );
  NAND U155 ( .A(n88), .B(n90), .Z(n1415) );
  NAND U156 ( .A(sreg[119]), .B(n1472), .Z(n91) );
  XOR U157 ( .A(n1472), .B(sreg[119]), .Z(n92) );
  NANDN U158 ( .A(n1473), .B(n92), .Z(n93) );
  NAND U159 ( .A(n91), .B(n93), .Z(n1491) );
  XNOR U160 ( .A(n436), .B(n437), .Z(n438) );
  XNOR U161 ( .A(n455), .B(n456), .Z(n457) );
  XNOR U162 ( .A(n474), .B(n475), .Z(n476) );
  NAND U163 ( .A(n501), .B(n499), .Z(n94) );
  XOR U164 ( .A(n499), .B(n501), .Z(n95) );
  NANDN U165 ( .A(n500), .B(n95), .Z(n96) );
  NAND U166 ( .A(n94), .B(n96), .Z(n515) );
  XNOR U167 ( .A(n531), .B(n532), .Z(n533) );
  XNOR U168 ( .A(n550), .B(n551), .Z(n552) );
  NAND U169 ( .A(n577), .B(n575), .Z(n97) );
  XOR U170 ( .A(n575), .B(n577), .Z(n98) );
  NANDN U171 ( .A(n576), .B(n98), .Z(n99) );
  NAND U172 ( .A(n97), .B(n99), .Z(n591) );
  XNOR U173 ( .A(n607), .B(n608), .Z(n609) );
  XNOR U174 ( .A(n626), .B(n627), .Z(n628) );
  NAND U175 ( .A(n653), .B(n651), .Z(n100) );
  XOR U176 ( .A(n651), .B(n653), .Z(n101) );
  NANDN U177 ( .A(n652), .B(n101), .Z(n102) );
  NAND U178 ( .A(n100), .B(n102), .Z(n667) );
  XNOR U179 ( .A(n683), .B(n684), .Z(n685) );
  XNOR U180 ( .A(n702), .B(n703), .Z(n704) );
  NAND U181 ( .A(n729), .B(n727), .Z(n103) );
  XOR U182 ( .A(n727), .B(n729), .Z(n104) );
  NANDN U183 ( .A(n728), .B(n104), .Z(n105) );
  NAND U184 ( .A(n103), .B(n105), .Z(n743) );
  XNOR U185 ( .A(n759), .B(n760), .Z(n761) );
  XNOR U186 ( .A(n778), .B(n779), .Z(n780) );
  NAND U187 ( .A(n805), .B(n803), .Z(n106) );
  XOR U188 ( .A(n803), .B(n805), .Z(n107) );
  NANDN U189 ( .A(n804), .B(n107), .Z(n108) );
  NAND U190 ( .A(n106), .B(n108), .Z(n819) );
  XNOR U191 ( .A(n835), .B(n836), .Z(n837) );
  XNOR U192 ( .A(n854), .B(n855), .Z(n856) );
  NAND U193 ( .A(n881), .B(n879), .Z(n109) );
  XOR U194 ( .A(n879), .B(n881), .Z(n110) );
  NANDN U195 ( .A(n880), .B(n110), .Z(n111) );
  NAND U196 ( .A(n109), .B(n111), .Z(n895) );
  XNOR U197 ( .A(n911), .B(n912), .Z(n913) );
  XNOR U198 ( .A(n930), .B(n931), .Z(n932) );
  NAND U199 ( .A(n957), .B(n955), .Z(n112) );
  XOR U200 ( .A(n955), .B(n957), .Z(n113) );
  NANDN U201 ( .A(n956), .B(n113), .Z(n114) );
  NAND U202 ( .A(n112), .B(n114), .Z(n971) );
  XNOR U203 ( .A(n987), .B(n988), .Z(n989) );
  XNOR U204 ( .A(n1006), .B(n1007), .Z(n1008) );
  NAND U205 ( .A(n1033), .B(n1031), .Z(n115) );
  XOR U206 ( .A(n1031), .B(n1033), .Z(n116) );
  NANDN U207 ( .A(n1032), .B(n116), .Z(n117) );
  NAND U208 ( .A(n115), .B(n117), .Z(n1047) );
  XNOR U209 ( .A(n1063), .B(n1064), .Z(n1065) );
  XNOR U210 ( .A(n1082), .B(n1083), .Z(n1084) );
  NAND U211 ( .A(n1109), .B(n1107), .Z(n118) );
  XOR U212 ( .A(n1107), .B(n1109), .Z(n119) );
  NANDN U213 ( .A(n1108), .B(n119), .Z(n120) );
  NAND U214 ( .A(n118), .B(n120), .Z(n1123) );
  XNOR U215 ( .A(n1139), .B(n1140), .Z(n1141) );
  XNOR U216 ( .A(n1158), .B(n1159), .Z(n1160) );
  NAND U217 ( .A(n1185), .B(n1183), .Z(n121) );
  XOR U218 ( .A(n1183), .B(n1185), .Z(n122) );
  NANDN U219 ( .A(n1184), .B(n122), .Z(n123) );
  NAND U220 ( .A(n121), .B(n123), .Z(n1199) );
  XNOR U221 ( .A(n1215), .B(n1216), .Z(n1217) );
  XNOR U222 ( .A(n1234), .B(n1235), .Z(n1236) );
  NAND U223 ( .A(n1261), .B(n1259), .Z(n124) );
  XOR U224 ( .A(n1259), .B(n1261), .Z(n125) );
  NANDN U225 ( .A(n1260), .B(n125), .Z(n126) );
  NAND U226 ( .A(n124), .B(n126), .Z(n1275) );
  XNOR U227 ( .A(n1291), .B(n1292), .Z(n1293) );
  XNOR U228 ( .A(n1310), .B(n1311), .Z(n1312) );
  NAND U229 ( .A(n1337), .B(n1335), .Z(n127) );
  XOR U230 ( .A(n1335), .B(n1337), .Z(n128) );
  NANDN U231 ( .A(n1336), .B(n128), .Z(n129) );
  NAND U232 ( .A(n127), .B(n129), .Z(n1351) );
  XNOR U233 ( .A(n1367), .B(n1368), .Z(n1369) );
  XNOR U234 ( .A(n1386), .B(n1387), .Z(n1388) );
  NAND U235 ( .A(n1413), .B(n1411), .Z(n130) );
  XOR U236 ( .A(n1411), .B(n1413), .Z(n131) );
  NANDN U237 ( .A(n1412), .B(n131), .Z(n132) );
  NAND U238 ( .A(n130), .B(n132), .Z(n1427) );
  XNOR U239 ( .A(n1443), .B(n1444), .Z(n1445) );
  XNOR U240 ( .A(n1462), .B(n1463), .Z(n1464) );
  NAND U241 ( .A(n1489), .B(n1487), .Z(n133) );
  XOR U242 ( .A(n1487), .B(n1489), .Z(n134) );
  NANDN U243 ( .A(n1488), .B(n134), .Z(n135) );
  NAND U244 ( .A(n133), .B(n135), .Z(n1503) );
  XNOR U245 ( .A(n1521), .B(n1522), .Z(n1523) );
  NAND U246 ( .A(n1547), .B(n1546), .Z(n136) );
  XOR U247 ( .A(n1546), .B(n1547), .Z(n137) );
  NAND U248 ( .A(n137), .B(n1545), .Z(n138) );
  NAND U249 ( .A(n136), .B(n138), .Z(n1567) );
  XOR U250 ( .A(n428), .B(n427), .Z(n139) );
  NANDN U251 ( .A(sreg[64]), .B(n139), .Z(n140) );
  NAND U252 ( .A(n428), .B(n427), .Z(n141) );
  AND U253 ( .A(n140), .B(n141), .Z(n446) );
  NAND U254 ( .A(sreg[68]), .B(n503), .Z(n142) );
  XOR U255 ( .A(n503), .B(sreg[68]), .Z(n143) );
  NANDN U256 ( .A(n504), .B(n143), .Z(n144) );
  NAND U257 ( .A(n142), .B(n144), .Z(n522) );
  NAND U258 ( .A(sreg[72]), .B(n579), .Z(n145) );
  XOR U259 ( .A(n579), .B(sreg[72]), .Z(n146) );
  NANDN U260 ( .A(n580), .B(n146), .Z(n147) );
  NAND U261 ( .A(n145), .B(n147), .Z(n598) );
  NAND U262 ( .A(sreg[76]), .B(n655), .Z(n148) );
  XOR U263 ( .A(n655), .B(sreg[76]), .Z(n149) );
  NANDN U264 ( .A(n656), .B(n149), .Z(n150) );
  NAND U265 ( .A(n148), .B(n150), .Z(n674) );
  NAND U266 ( .A(sreg[80]), .B(n731), .Z(n151) );
  XOR U267 ( .A(n731), .B(sreg[80]), .Z(n152) );
  NANDN U268 ( .A(n732), .B(n152), .Z(n153) );
  NAND U269 ( .A(n151), .B(n153), .Z(n750) );
  NAND U270 ( .A(sreg[84]), .B(n807), .Z(n154) );
  XOR U271 ( .A(n807), .B(sreg[84]), .Z(n155) );
  NANDN U272 ( .A(n808), .B(n155), .Z(n156) );
  NAND U273 ( .A(n154), .B(n156), .Z(n826) );
  NAND U274 ( .A(sreg[88]), .B(n883), .Z(n157) );
  XOR U275 ( .A(n883), .B(sreg[88]), .Z(n158) );
  NANDN U276 ( .A(n884), .B(n158), .Z(n159) );
  NAND U277 ( .A(n157), .B(n159), .Z(n902) );
  NAND U278 ( .A(sreg[92]), .B(n959), .Z(n160) );
  XOR U279 ( .A(n959), .B(sreg[92]), .Z(n161) );
  NANDN U280 ( .A(n960), .B(n161), .Z(n162) );
  NAND U281 ( .A(n160), .B(n162), .Z(n978) );
  NAND U282 ( .A(sreg[96]), .B(n1035), .Z(n163) );
  XOR U283 ( .A(n1035), .B(sreg[96]), .Z(n164) );
  NANDN U284 ( .A(n1036), .B(n164), .Z(n165) );
  NAND U285 ( .A(n163), .B(n165), .Z(n1054) );
  NAND U286 ( .A(sreg[100]), .B(n1111), .Z(n166) );
  XOR U287 ( .A(n1111), .B(sreg[100]), .Z(n167) );
  NANDN U288 ( .A(n1112), .B(n167), .Z(n168) );
  NAND U289 ( .A(n166), .B(n168), .Z(n1130) );
  NAND U290 ( .A(sreg[104]), .B(n1187), .Z(n169) );
  XOR U291 ( .A(n1187), .B(sreg[104]), .Z(n170) );
  NANDN U292 ( .A(n1188), .B(n170), .Z(n171) );
  NAND U293 ( .A(n169), .B(n171), .Z(n1206) );
  NAND U294 ( .A(sreg[108]), .B(n1263), .Z(n172) );
  XOR U295 ( .A(n1263), .B(sreg[108]), .Z(n173) );
  NANDN U296 ( .A(n1264), .B(n173), .Z(n174) );
  NAND U297 ( .A(n172), .B(n174), .Z(n1282) );
  NAND U298 ( .A(sreg[112]), .B(n1339), .Z(n175) );
  XOR U299 ( .A(n1339), .B(sreg[112]), .Z(n176) );
  NANDN U300 ( .A(n1340), .B(n176), .Z(n177) );
  NAND U301 ( .A(n175), .B(n177), .Z(n1358) );
  NAND U302 ( .A(sreg[116]), .B(n1415), .Z(n178) );
  XOR U303 ( .A(n1415), .B(sreg[116]), .Z(n179) );
  NANDN U304 ( .A(n1416), .B(n179), .Z(n180) );
  NAND U305 ( .A(n178), .B(n180), .Z(n1434) );
  NAND U306 ( .A(sreg[120]), .B(n1491), .Z(n181) );
  XOR U307 ( .A(n1491), .B(sreg[120]), .Z(n182) );
  NANDN U308 ( .A(n1492), .B(n182), .Z(n183) );
  NAND U309 ( .A(n181), .B(n183), .Z(n1510) );
  AND U310 ( .A(b[1]), .B(a[0]), .Z(n390) );
  NAND U311 ( .A(n463), .B(n461), .Z(n184) );
  XOR U312 ( .A(n461), .B(n463), .Z(n185) );
  NANDN U313 ( .A(n462), .B(n185), .Z(n186) );
  NAND U314 ( .A(n184), .B(n186), .Z(n477) );
  NAND U315 ( .A(n482), .B(n480), .Z(n187) );
  XOR U316 ( .A(n480), .B(n482), .Z(n188) );
  NANDN U317 ( .A(n481), .B(n188), .Z(n189) );
  NAND U318 ( .A(n187), .B(n189), .Z(n496) );
  NAND U319 ( .A(n520), .B(n518), .Z(n190) );
  XOR U320 ( .A(n518), .B(n520), .Z(n191) );
  NANDN U321 ( .A(n519), .B(n191), .Z(n192) );
  NAND U322 ( .A(n190), .B(n192), .Z(n534) );
  NAND U323 ( .A(n539), .B(n537), .Z(n193) );
  XOR U324 ( .A(n537), .B(n539), .Z(n194) );
  NANDN U325 ( .A(n538), .B(n194), .Z(n195) );
  NAND U326 ( .A(n193), .B(n195), .Z(n553) );
  NAND U327 ( .A(n558), .B(n556), .Z(n196) );
  XOR U328 ( .A(n556), .B(n558), .Z(n197) );
  NANDN U329 ( .A(n557), .B(n197), .Z(n198) );
  NAND U330 ( .A(n196), .B(n198), .Z(n572) );
  NAND U331 ( .A(n596), .B(n594), .Z(n199) );
  XOR U332 ( .A(n594), .B(n596), .Z(n200) );
  NANDN U333 ( .A(n595), .B(n200), .Z(n201) );
  NAND U334 ( .A(n199), .B(n201), .Z(n610) );
  NAND U335 ( .A(n615), .B(n613), .Z(n202) );
  XOR U336 ( .A(n613), .B(n615), .Z(n203) );
  NANDN U337 ( .A(n614), .B(n203), .Z(n204) );
  NAND U338 ( .A(n202), .B(n204), .Z(n629) );
  NAND U339 ( .A(n634), .B(n632), .Z(n205) );
  XOR U340 ( .A(n632), .B(n634), .Z(n206) );
  NANDN U341 ( .A(n633), .B(n206), .Z(n207) );
  NAND U342 ( .A(n205), .B(n207), .Z(n648) );
  NAND U343 ( .A(n672), .B(n670), .Z(n208) );
  XOR U344 ( .A(n670), .B(n672), .Z(n209) );
  NANDN U345 ( .A(n671), .B(n209), .Z(n210) );
  NAND U346 ( .A(n208), .B(n210), .Z(n686) );
  NAND U347 ( .A(n691), .B(n689), .Z(n211) );
  XOR U348 ( .A(n689), .B(n691), .Z(n212) );
  NANDN U349 ( .A(n690), .B(n212), .Z(n213) );
  NAND U350 ( .A(n211), .B(n213), .Z(n705) );
  NAND U351 ( .A(n710), .B(n708), .Z(n214) );
  XOR U352 ( .A(n708), .B(n710), .Z(n215) );
  NANDN U353 ( .A(n709), .B(n215), .Z(n216) );
  NAND U354 ( .A(n214), .B(n216), .Z(n724) );
  NAND U355 ( .A(n748), .B(n746), .Z(n217) );
  XOR U356 ( .A(n746), .B(n748), .Z(n218) );
  NANDN U357 ( .A(n747), .B(n218), .Z(n219) );
  NAND U358 ( .A(n217), .B(n219), .Z(n762) );
  NAND U359 ( .A(n767), .B(n765), .Z(n220) );
  XOR U360 ( .A(n765), .B(n767), .Z(n221) );
  NANDN U361 ( .A(n766), .B(n221), .Z(n222) );
  NAND U362 ( .A(n220), .B(n222), .Z(n781) );
  NAND U363 ( .A(n786), .B(n784), .Z(n223) );
  XOR U364 ( .A(n784), .B(n786), .Z(n224) );
  NANDN U365 ( .A(n785), .B(n224), .Z(n225) );
  NAND U366 ( .A(n223), .B(n225), .Z(n800) );
  NAND U367 ( .A(n824), .B(n822), .Z(n226) );
  XOR U368 ( .A(n822), .B(n824), .Z(n227) );
  NANDN U369 ( .A(n823), .B(n227), .Z(n228) );
  NAND U370 ( .A(n226), .B(n228), .Z(n838) );
  NAND U371 ( .A(n843), .B(n841), .Z(n229) );
  XOR U372 ( .A(n841), .B(n843), .Z(n230) );
  NANDN U373 ( .A(n842), .B(n230), .Z(n231) );
  NAND U374 ( .A(n229), .B(n231), .Z(n857) );
  NAND U375 ( .A(n862), .B(n860), .Z(n232) );
  XOR U376 ( .A(n860), .B(n862), .Z(n233) );
  NANDN U377 ( .A(n861), .B(n233), .Z(n234) );
  NAND U378 ( .A(n232), .B(n234), .Z(n876) );
  NAND U379 ( .A(n900), .B(n898), .Z(n235) );
  XOR U380 ( .A(n898), .B(n900), .Z(n236) );
  NANDN U381 ( .A(n899), .B(n236), .Z(n237) );
  NAND U382 ( .A(n235), .B(n237), .Z(n914) );
  NAND U383 ( .A(n919), .B(n917), .Z(n238) );
  XOR U384 ( .A(n917), .B(n919), .Z(n239) );
  NANDN U385 ( .A(n918), .B(n239), .Z(n240) );
  NAND U386 ( .A(n238), .B(n240), .Z(n933) );
  NAND U387 ( .A(n938), .B(n936), .Z(n241) );
  XOR U388 ( .A(n936), .B(n938), .Z(n242) );
  NANDN U389 ( .A(n937), .B(n242), .Z(n243) );
  NAND U390 ( .A(n241), .B(n243), .Z(n952) );
  NAND U391 ( .A(n976), .B(n974), .Z(n244) );
  XOR U392 ( .A(n974), .B(n976), .Z(n245) );
  NANDN U393 ( .A(n975), .B(n245), .Z(n246) );
  NAND U394 ( .A(n244), .B(n246), .Z(n990) );
  NAND U395 ( .A(n995), .B(n993), .Z(n247) );
  XOR U396 ( .A(n993), .B(n995), .Z(n248) );
  NANDN U397 ( .A(n994), .B(n248), .Z(n249) );
  NAND U398 ( .A(n247), .B(n249), .Z(n1009) );
  NAND U399 ( .A(n1014), .B(n1012), .Z(n250) );
  XOR U400 ( .A(n1012), .B(n1014), .Z(n251) );
  NANDN U401 ( .A(n1013), .B(n251), .Z(n252) );
  NAND U402 ( .A(n250), .B(n252), .Z(n1028) );
  NAND U403 ( .A(n1052), .B(n1050), .Z(n253) );
  XOR U404 ( .A(n1050), .B(n1052), .Z(n254) );
  NANDN U405 ( .A(n1051), .B(n254), .Z(n255) );
  NAND U406 ( .A(n253), .B(n255), .Z(n1066) );
  NAND U407 ( .A(n1071), .B(n1069), .Z(n256) );
  XOR U408 ( .A(n1069), .B(n1071), .Z(n257) );
  NANDN U409 ( .A(n1070), .B(n257), .Z(n258) );
  NAND U410 ( .A(n256), .B(n258), .Z(n1085) );
  NAND U411 ( .A(n1090), .B(n1088), .Z(n259) );
  XOR U412 ( .A(n1088), .B(n1090), .Z(n260) );
  NANDN U413 ( .A(n1089), .B(n260), .Z(n261) );
  NAND U414 ( .A(n259), .B(n261), .Z(n1104) );
  NAND U415 ( .A(n1128), .B(n1126), .Z(n262) );
  XOR U416 ( .A(n1126), .B(n1128), .Z(n263) );
  NANDN U417 ( .A(n1127), .B(n263), .Z(n264) );
  NAND U418 ( .A(n262), .B(n264), .Z(n1142) );
  NAND U419 ( .A(n1147), .B(n1145), .Z(n265) );
  XOR U420 ( .A(n1145), .B(n1147), .Z(n266) );
  NANDN U421 ( .A(n1146), .B(n266), .Z(n267) );
  NAND U422 ( .A(n265), .B(n267), .Z(n1161) );
  NAND U423 ( .A(n1166), .B(n1164), .Z(n268) );
  XOR U424 ( .A(n1164), .B(n1166), .Z(n269) );
  NANDN U425 ( .A(n1165), .B(n269), .Z(n270) );
  NAND U426 ( .A(n268), .B(n270), .Z(n1180) );
  NAND U427 ( .A(n1204), .B(n1202), .Z(n271) );
  XOR U428 ( .A(n1202), .B(n1204), .Z(n272) );
  NANDN U429 ( .A(n1203), .B(n272), .Z(n273) );
  NAND U430 ( .A(n271), .B(n273), .Z(n1218) );
  NAND U431 ( .A(n1223), .B(n1221), .Z(n274) );
  XOR U432 ( .A(n1221), .B(n1223), .Z(n275) );
  NANDN U433 ( .A(n1222), .B(n275), .Z(n276) );
  NAND U434 ( .A(n274), .B(n276), .Z(n1237) );
  NAND U435 ( .A(n1242), .B(n1240), .Z(n277) );
  XOR U436 ( .A(n1240), .B(n1242), .Z(n278) );
  NANDN U437 ( .A(n1241), .B(n278), .Z(n279) );
  NAND U438 ( .A(n277), .B(n279), .Z(n1256) );
  NAND U439 ( .A(n1280), .B(n1278), .Z(n280) );
  XOR U440 ( .A(n1278), .B(n1280), .Z(n281) );
  NANDN U441 ( .A(n1279), .B(n281), .Z(n282) );
  NAND U442 ( .A(n280), .B(n282), .Z(n1294) );
  NAND U443 ( .A(n1299), .B(n1297), .Z(n283) );
  XOR U444 ( .A(n1297), .B(n1299), .Z(n284) );
  NANDN U445 ( .A(n1298), .B(n284), .Z(n285) );
  NAND U446 ( .A(n283), .B(n285), .Z(n1313) );
  NAND U447 ( .A(n1318), .B(n1316), .Z(n286) );
  XOR U448 ( .A(n1316), .B(n1318), .Z(n287) );
  NANDN U449 ( .A(n1317), .B(n287), .Z(n288) );
  NAND U450 ( .A(n286), .B(n288), .Z(n1332) );
  NAND U451 ( .A(n1356), .B(n1354), .Z(n289) );
  XOR U452 ( .A(n1354), .B(n1356), .Z(n290) );
  NANDN U453 ( .A(n1355), .B(n290), .Z(n291) );
  NAND U454 ( .A(n289), .B(n291), .Z(n1370) );
  NAND U455 ( .A(n1375), .B(n1373), .Z(n292) );
  XOR U456 ( .A(n1373), .B(n1375), .Z(n293) );
  NANDN U457 ( .A(n1374), .B(n293), .Z(n294) );
  NAND U458 ( .A(n292), .B(n294), .Z(n1389) );
  NAND U459 ( .A(n1394), .B(n1392), .Z(n295) );
  XOR U460 ( .A(n1392), .B(n1394), .Z(n296) );
  NANDN U461 ( .A(n1393), .B(n296), .Z(n297) );
  NAND U462 ( .A(n295), .B(n297), .Z(n1408) );
  NAND U463 ( .A(n1432), .B(n1430), .Z(n298) );
  XOR U464 ( .A(n1430), .B(n1432), .Z(n299) );
  NANDN U465 ( .A(n1431), .B(n299), .Z(n300) );
  NAND U466 ( .A(n298), .B(n300), .Z(n1446) );
  NAND U467 ( .A(n1451), .B(n1449), .Z(n301) );
  XOR U468 ( .A(n1449), .B(n1451), .Z(n302) );
  NANDN U469 ( .A(n1450), .B(n302), .Z(n303) );
  NAND U470 ( .A(n301), .B(n303), .Z(n1465) );
  NAND U471 ( .A(n1470), .B(n1468), .Z(n304) );
  XOR U472 ( .A(n1468), .B(n1470), .Z(n305) );
  NANDN U473 ( .A(n1469), .B(n305), .Z(n306) );
  NAND U474 ( .A(n304), .B(n306), .Z(n1484) );
  NAND U475 ( .A(n1508), .B(n1506), .Z(n307) );
  XOR U476 ( .A(n1506), .B(n1508), .Z(n308) );
  NANDN U477 ( .A(n1507), .B(n308), .Z(n309) );
  NAND U478 ( .A(n307), .B(n309), .Z(n1524) );
  XOR U479 ( .A(n1538), .B(n1536), .Z(n310) );
  NANDN U480 ( .A(n1537), .B(n310), .Z(n311) );
  NAND U481 ( .A(n1538), .B(n1536), .Z(n312) );
  AND U482 ( .A(n311), .B(n312), .Z(n1555) );
  AND U483 ( .A(a[0]), .B(b[3]), .Z(n313) );
  NAND U484 ( .A(a[2]), .B(b[1]), .Z(n314) );
  XNOR U485 ( .A(n313), .B(n314), .Z(n315) );
  XNOR U486 ( .A(n315), .B(n391), .Z(n396) );
  XNOR U487 ( .A(n423), .B(n424), .Z(n417) );
  NAND U488 ( .A(sreg[65]), .B(n446), .Z(n316) );
  XOR U489 ( .A(n446), .B(sreg[65]), .Z(n317) );
  NANDN U490 ( .A(n447), .B(n317), .Z(n318) );
  NAND U491 ( .A(n316), .B(n318), .Z(n465) );
  NAND U492 ( .A(sreg[69]), .B(n522), .Z(n319) );
  XOR U493 ( .A(n522), .B(sreg[69]), .Z(n320) );
  NANDN U494 ( .A(n523), .B(n320), .Z(n321) );
  NAND U495 ( .A(n319), .B(n321), .Z(n541) );
  NAND U496 ( .A(sreg[73]), .B(n598), .Z(n322) );
  XOR U497 ( .A(n598), .B(sreg[73]), .Z(n323) );
  NANDN U498 ( .A(n599), .B(n323), .Z(n324) );
  NAND U499 ( .A(n322), .B(n324), .Z(n617) );
  NAND U500 ( .A(sreg[77]), .B(n674), .Z(n325) );
  XOR U501 ( .A(n674), .B(sreg[77]), .Z(n326) );
  NANDN U502 ( .A(n675), .B(n326), .Z(n327) );
  NAND U503 ( .A(n325), .B(n327), .Z(n693) );
  NAND U504 ( .A(sreg[81]), .B(n750), .Z(n328) );
  XOR U505 ( .A(n750), .B(sreg[81]), .Z(n329) );
  NANDN U506 ( .A(n751), .B(n329), .Z(n330) );
  NAND U507 ( .A(n328), .B(n330), .Z(n769) );
  NAND U508 ( .A(sreg[85]), .B(n826), .Z(n331) );
  XOR U509 ( .A(n826), .B(sreg[85]), .Z(n332) );
  NANDN U510 ( .A(n827), .B(n332), .Z(n333) );
  NAND U511 ( .A(n331), .B(n333), .Z(n845) );
  NAND U512 ( .A(sreg[89]), .B(n902), .Z(n334) );
  XOR U513 ( .A(n902), .B(sreg[89]), .Z(n335) );
  NANDN U514 ( .A(n903), .B(n335), .Z(n336) );
  NAND U515 ( .A(n334), .B(n336), .Z(n921) );
  NAND U516 ( .A(sreg[93]), .B(n978), .Z(n337) );
  XOR U517 ( .A(n978), .B(sreg[93]), .Z(n338) );
  NANDN U518 ( .A(n979), .B(n338), .Z(n339) );
  NAND U519 ( .A(n337), .B(n339), .Z(n997) );
  NAND U520 ( .A(sreg[97]), .B(n1054), .Z(n340) );
  XOR U521 ( .A(n1054), .B(sreg[97]), .Z(n341) );
  NANDN U522 ( .A(n1055), .B(n341), .Z(n342) );
  NAND U523 ( .A(n340), .B(n342), .Z(n1073) );
  NAND U524 ( .A(sreg[101]), .B(n1130), .Z(n343) );
  XOR U525 ( .A(n1130), .B(sreg[101]), .Z(n344) );
  NANDN U526 ( .A(n1131), .B(n344), .Z(n345) );
  NAND U527 ( .A(n343), .B(n345), .Z(n1149) );
  NAND U528 ( .A(sreg[105]), .B(n1206), .Z(n346) );
  XOR U529 ( .A(n1206), .B(sreg[105]), .Z(n347) );
  NANDN U530 ( .A(n1207), .B(n347), .Z(n348) );
  NAND U531 ( .A(n346), .B(n348), .Z(n1225) );
  NAND U532 ( .A(sreg[109]), .B(n1282), .Z(n349) );
  XOR U533 ( .A(n1282), .B(sreg[109]), .Z(n350) );
  NANDN U534 ( .A(n1283), .B(n350), .Z(n351) );
  NAND U535 ( .A(n349), .B(n351), .Z(n1301) );
  NAND U536 ( .A(sreg[113]), .B(n1358), .Z(n352) );
  XOR U537 ( .A(n1358), .B(sreg[113]), .Z(n353) );
  NANDN U538 ( .A(n1359), .B(n353), .Z(n354) );
  NAND U539 ( .A(n352), .B(n354), .Z(n1377) );
  NAND U540 ( .A(sreg[117]), .B(n1434), .Z(n355) );
  XOR U541 ( .A(n1434), .B(sreg[117]), .Z(n356) );
  NANDN U542 ( .A(n1435), .B(n356), .Z(n357) );
  NAND U543 ( .A(n355), .B(n357), .Z(n1453) );
  NAND U544 ( .A(sreg[121]), .B(n1510), .Z(n358) );
  XOR U545 ( .A(n1510), .B(sreg[121]), .Z(n359) );
  NANDN U546 ( .A(n1511), .B(n359), .Z(n360) );
  NAND U547 ( .A(n358), .B(n360), .Z(n1513) );
  NANDN U548 ( .A(n1585), .B(n1586), .Z(n361) );
  XNOR U549 ( .A(n1585), .B(n1586), .Z(n362) );
  NAND U550 ( .A(n362), .B(n1587), .Z(n363) );
  AND U551 ( .A(n361), .B(n363), .Z(n364) );
  XOR U552 ( .A(n1587), .B(n362), .Z(n365) );
  NANDN U553 ( .A(n1584), .B(n365), .Z(n366) );
  NAND U554 ( .A(n364), .B(n366), .Z(c[127]) );
  IV U555 ( .A(b[3]), .Z(n367) );
  NAND U556 ( .A(a[0]), .B(b[0]), .Z(n368) );
  XNOR U557 ( .A(n368), .B(sreg[60]), .Z(c[60]) );
  IV U558 ( .A(n390), .Z(n370) );
  NAND U559 ( .A(b[0]), .B(a[1]), .Z(n369) );
  XNOR U560 ( .A(n370), .B(n369), .Z(n371) );
  XOR U561 ( .A(sreg[61]), .B(n371), .Z(n373) );
  NANDN U562 ( .A(n368), .B(sreg[60]), .Z(n372) );
  XOR U563 ( .A(n373), .B(n372), .Z(c[61]) );
  NOR U564 ( .A(n370), .B(n369), .Z(n384) );
  AND U565 ( .A(b[2]), .B(a[0]), .Z(n381) );
  NAND U566 ( .A(b[1]), .B(a[1]), .Z(n380) );
  NAND U567 ( .A(a[2]), .B(b[0]), .Z(n379) );
  XOR U568 ( .A(n380), .B(n379), .Z(n382) );
  XOR U569 ( .A(n381), .B(n382), .Z(n383) );
  XOR U570 ( .A(n384), .B(n383), .Z(n377) );
  NANDN U571 ( .A(n371), .B(sreg[61]), .Z(n375) );
  OR U572 ( .A(n373), .B(n372), .Z(n374) );
  AND U573 ( .A(n375), .B(n374), .Z(n378) );
  XOR U574 ( .A(n377), .B(n378), .Z(n376) );
  XNOR U575 ( .A(sreg[62]), .B(n376), .Z(c[62]) );
  XNOR U576 ( .A(n400), .B(sreg[63]), .Z(n402) );
  OR U577 ( .A(n380), .B(n379), .Z(n391) );
  OR U578 ( .A(n382), .B(n381), .Z(n386) );
  NANDN U579 ( .A(n384), .B(n383), .Z(n385) );
  NAND U580 ( .A(n386), .B(n385), .Z(n393) );
  NAND U581 ( .A(a[3]), .B(b[0]), .Z(n388) );
  NAND U582 ( .A(b[2]), .B(a[1]), .Z(n387) );
  XOR U583 ( .A(n388), .B(n387), .Z(n394) );
  XNOR U584 ( .A(n393), .B(n394), .Z(n395) );
  XNOR U585 ( .A(n396), .B(n395), .Z(n401) );
  XOR U586 ( .A(n402), .B(n401), .Z(c[63]) );
  NAND U587 ( .A(b[2]), .B(a[2]), .Z(n409) );
  OR U588 ( .A(n388), .B(n387), .Z(n406) );
  IV U589 ( .A(n406), .Z(n407) );
  AND U590 ( .A(a[1]), .B(b[3]), .Z(n408) );
  XNOR U591 ( .A(n407), .B(n408), .Z(n389) );
  XNOR U592 ( .A(n409), .B(n389), .Z(n424) );
  NAND U593 ( .A(a[4]), .B(b[0]), .Z(n422) );
  AND U594 ( .A(a[3]), .B(b[1]), .Z(n421) );
  XNOR U595 ( .A(n422), .B(n421), .Z(n423) );
  ANDN U596 ( .B(a[2]), .A(n367), .Z(n442) );
  NAND U597 ( .A(n390), .B(n442), .Z(n392) );
  AND U598 ( .A(n392), .B(n391), .Z(n416) );
  IV U599 ( .A(n416), .Z(n414) );
  NANDN U600 ( .A(n394), .B(n393), .Z(n398) );
  NANDN U601 ( .A(n396), .B(n395), .Z(n397) );
  AND U602 ( .A(n398), .B(n397), .Z(n415) );
  XOR U603 ( .A(n414), .B(n415), .Z(n399) );
  XNOR U604 ( .A(n417), .B(n399), .Z(n428) );
  NAND U605 ( .A(sreg[63]), .B(n400), .Z(n404) );
  OR U606 ( .A(n402), .B(n401), .Z(n403) );
  AND U607 ( .A(n404), .B(n403), .Z(n427) );
  XNOR U608 ( .A(n427), .B(sreg[64]), .Z(n405) );
  XNOR U609 ( .A(n428), .B(n405), .Z(c[64]) );
  NANDN U610 ( .A(n408), .B(n406), .Z(n412) );
  AND U611 ( .A(n408), .B(n407), .Z(n410) );
  NANDN U612 ( .A(n410), .B(n409), .Z(n411) );
  NAND U613 ( .A(n412), .B(n411), .Z(n439) );
  AND U614 ( .A(a[4]), .B(b[1]), .Z(n443) );
  NAND U615 ( .A(b[2]), .B(a[3]), .Z(n444) );
  XOR U616 ( .A(n442), .B(n444), .Z(n413) );
  XNOR U617 ( .A(n443), .B(n413), .Z(n436) );
  NAND U618 ( .A(a[5]), .B(b[0]), .Z(n437) );
  XOR U619 ( .A(n439), .B(n438), .Z(n432) );
  NAND U620 ( .A(n414), .B(n415), .Z(n420) );
  ANDN U621 ( .B(n416), .A(n415), .Z(n418) );
  NANDN U622 ( .A(n418), .B(n417), .Z(n419) );
  NAND U623 ( .A(n420), .B(n419), .Z(n430) );
  NANDN U624 ( .A(n422), .B(n421), .Z(n426) );
  NANDN U625 ( .A(n424), .B(n423), .Z(n425) );
  AND U626 ( .A(n426), .B(n425), .Z(n431) );
  XOR U627 ( .A(n430), .B(n431), .Z(n433) );
  XNOR U628 ( .A(n432), .B(n433), .Z(n447) );
  XOR U629 ( .A(n446), .B(sreg[65]), .Z(n429) );
  XNOR U630 ( .A(n447), .B(n429), .Z(c[65]) );
  NANDN U631 ( .A(n431), .B(n430), .Z(n435) );
  OR U632 ( .A(n433), .B(n432), .Z(n434) );
  NAND U633 ( .A(n435), .B(n434), .Z(n449) );
  NANDN U634 ( .A(n437), .B(n436), .Z(n441) );
  NANDN U635 ( .A(n439), .B(n438), .Z(n440) );
  AND U636 ( .A(n441), .B(n440), .Z(n450) );
  XNOR U637 ( .A(n449), .B(n450), .Z(n451) );
  AND U638 ( .A(a[5]), .B(b[1]), .Z(n462) );
  NAND U639 ( .A(b[2]), .B(a[4]), .Z(n463) );
  NAND U640 ( .A(b[3]), .B(a[3]), .Z(n461) );
  XNOR U641 ( .A(n463), .B(n461), .Z(n445) );
  XNOR U642 ( .A(n462), .B(n445), .Z(n455) );
  NAND U643 ( .A(a[6]), .B(b[0]), .Z(n456) );
  XOR U644 ( .A(n458), .B(n457), .Z(n452) );
  XOR U645 ( .A(n451), .B(n452), .Z(n466) );
  XOR U646 ( .A(n465), .B(sreg[66]), .Z(n448) );
  XNOR U647 ( .A(n466), .B(n448), .Z(c[66]) );
  NANDN U648 ( .A(n450), .B(n449), .Z(n454) );
  NANDN U649 ( .A(n452), .B(n451), .Z(n453) );
  NAND U650 ( .A(n454), .B(n453), .Z(n468) );
  NANDN U651 ( .A(n456), .B(n455), .Z(n460) );
  NANDN U652 ( .A(n458), .B(n457), .Z(n459) );
  AND U653 ( .A(n460), .B(n459), .Z(n469) );
  XNOR U654 ( .A(n468), .B(n469), .Z(n470) );
  AND U655 ( .A(a[6]), .B(b[1]), .Z(n481) );
  NAND U656 ( .A(b[2]), .B(a[5]), .Z(n482) );
  NAND U657 ( .A(b[3]), .B(a[4]), .Z(n480) );
  XNOR U658 ( .A(n482), .B(n480), .Z(n464) );
  XNOR U659 ( .A(n481), .B(n464), .Z(n474) );
  NAND U660 ( .A(a[7]), .B(b[0]), .Z(n475) );
  XOR U661 ( .A(n477), .B(n476), .Z(n471) );
  XOR U662 ( .A(n470), .B(n471), .Z(n485) );
  XOR U663 ( .A(n484), .B(sreg[67]), .Z(n467) );
  XNOR U664 ( .A(n485), .B(n467), .Z(c[67]) );
  NANDN U665 ( .A(n469), .B(n468), .Z(n473) );
  NANDN U666 ( .A(n471), .B(n470), .Z(n472) );
  NAND U667 ( .A(n473), .B(n472), .Z(n487) );
  NANDN U668 ( .A(n475), .B(n474), .Z(n479) );
  NANDN U669 ( .A(n477), .B(n476), .Z(n478) );
  AND U670 ( .A(n479), .B(n478), .Z(n488) );
  XNOR U671 ( .A(n487), .B(n488), .Z(n489) );
  AND U672 ( .A(a[7]), .B(b[1]), .Z(n500) );
  NAND U673 ( .A(b[2]), .B(a[6]), .Z(n501) );
  NAND U674 ( .A(b[3]), .B(a[5]), .Z(n499) );
  XNOR U675 ( .A(n501), .B(n499), .Z(n483) );
  XNOR U676 ( .A(n500), .B(n483), .Z(n493) );
  NAND U677 ( .A(a[8]), .B(b[0]), .Z(n494) );
  XOR U678 ( .A(n496), .B(n495), .Z(n490) );
  XOR U679 ( .A(n489), .B(n490), .Z(n504) );
  XOR U680 ( .A(n503), .B(sreg[68]), .Z(n486) );
  XNOR U681 ( .A(n504), .B(n486), .Z(c[68]) );
  NANDN U682 ( .A(n488), .B(n487), .Z(n492) );
  NANDN U683 ( .A(n490), .B(n489), .Z(n491) );
  NAND U684 ( .A(n492), .B(n491), .Z(n506) );
  NANDN U685 ( .A(n494), .B(n493), .Z(n498) );
  NANDN U686 ( .A(n496), .B(n495), .Z(n497) );
  AND U687 ( .A(n498), .B(n497), .Z(n507) );
  XNOR U688 ( .A(n506), .B(n507), .Z(n508) );
  AND U689 ( .A(a[8]), .B(b[1]), .Z(n519) );
  NAND U690 ( .A(b[2]), .B(a[7]), .Z(n520) );
  NAND U691 ( .A(b[3]), .B(a[6]), .Z(n518) );
  XNOR U692 ( .A(n520), .B(n518), .Z(n502) );
  XNOR U693 ( .A(n519), .B(n502), .Z(n512) );
  NAND U694 ( .A(a[9]), .B(b[0]), .Z(n513) );
  XOR U695 ( .A(n515), .B(n514), .Z(n509) );
  XOR U696 ( .A(n508), .B(n509), .Z(n523) );
  XOR U697 ( .A(n522), .B(sreg[69]), .Z(n505) );
  XNOR U698 ( .A(n523), .B(n505), .Z(c[69]) );
  NANDN U699 ( .A(n507), .B(n506), .Z(n511) );
  NANDN U700 ( .A(n509), .B(n508), .Z(n510) );
  NAND U701 ( .A(n511), .B(n510), .Z(n525) );
  NANDN U702 ( .A(n513), .B(n512), .Z(n517) );
  NANDN U703 ( .A(n515), .B(n514), .Z(n516) );
  AND U704 ( .A(n517), .B(n516), .Z(n526) );
  XNOR U705 ( .A(n525), .B(n526), .Z(n527) );
  AND U706 ( .A(a[9]), .B(b[1]), .Z(n538) );
  NAND U707 ( .A(b[2]), .B(a[8]), .Z(n539) );
  NAND U708 ( .A(b[3]), .B(a[7]), .Z(n537) );
  XNOR U709 ( .A(n539), .B(n537), .Z(n521) );
  XNOR U710 ( .A(n538), .B(n521), .Z(n531) );
  NAND U711 ( .A(a[10]), .B(b[0]), .Z(n532) );
  XOR U712 ( .A(n534), .B(n533), .Z(n528) );
  XOR U713 ( .A(n527), .B(n528), .Z(n542) );
  XOR U714 ( .A(n541), .B(sreg[70]), .Z(n524) );
  XNOR U715 ( .A(n542), .B(n524), .Z(c[70]) );
  NANDN U716 ( .A(n526), .B(n525), .Z(n530) );
  NANDN U717 ( .A(n528), .B(n527), .Z(n529) );
  NAND U718 ( .A(n530), .B(n529), .Z(n544) );
  NANDN U719 ( .A(n532), .B(n531), .Z(n536) );
  NANDN U720 ( .A(n534), .B(n533), .Z(n535) );
  AND U721 ( .A(n536), .B(n535), .Z(n545) );
  XNOR U722 ( .A(n544), .B(n545), .Z(n546) );
  AND U723 ( .A(a[10]), .B(b[1]), .Z(n557) );
  NAND U724 ( .A(b[2]), .B(a[9]), .Z(n558) );
  NAND U725 ( .A(b[3]), .B(a[8]), .Z(n556) );
  XNOR U726 ( .A(n558), .B(n556), .Z(n540) );
  XNOR U727 ( .A(n557), .B(n540), .Z(n550) );
  NAND U728 ( .A(a[11]), .B(b[0]), .Z(n551) );
  XOR U729 ( .A(n553), .B(n552), .Z(n547) );
  XOR U730 ( .A(n546), .B(n547), .Z(n561) );
  XOR U731 ( .A(n560), .B(sreg[71]), .Z(n543) );
  XNOR U732 ( .A(n561), .B(n543), .Z(c[71]) );
  NANDN U733 ( .A(n545), .B(n544), .Z(n549) );
  NANDN U734 ( .A(n547), .B(n546), .Z(n548) );
  NAND U735 ( .A(n549), .B(n548), .Z(n563) );
  NANDN U736 ( .A(n551), .B(n550), .Z(n555) );
  NANDN U737 ( .A(n553), .B(n552), .Z(n554) );
  AND U738 ( .A(n555), .B(n554), .Z(n564) );
  XNOR U739 ( .A(n563), .B(n564), .Z(n565) );
  AND U740 ( .A(a[11]), .B(b[1]), .Z(n576) );
  NAND U741 ( .A(b[2]), .B(a[10]), .Z(n577) );
  NAND U742 ( .A(b[3]), .B(a[9]), .Z(n575) );
  XNOR U743 ( .A(n577), .B(n575), .Z(n559) );
  XNOR U744 ( .A(n576), .B(n559), .Z(n569) );
  NAND U745 ( .A(a[12]), .B(b[0]), .Z(n570) );
  XOR U746 ( .A(n572), .B(n571), .Z(n566) );
  XOR U747 ( .A(n565), .B(n566), .Z(n580) );
  XOR U748 ( .A(n579), .B(sreg[72]), .Z(n562) );
  XNOR U749 ( .A(n580), .B(n562), .Z(c[72]) );
  NANDN U750 ( .A(n564), .B(n563), .Z(n568) );
  NANDN U751 ( .A(n566), .B(n565), .Z(n567) );
  NAND U752 ( .A(n568), .B(n567), .Z(n582) );
  NANDN U753 ( .A(n570), .B(n569), .Z(n574) );
  NANDN U754 ( .A(n572), .B(n571), .Z(n573) );
  AND U755 ( .A(n574), .B(n573), .Z(n583) );
  XNOR U756 ( .A(n582), .B(n583), .Z(n584) );
  AND U757 ( .A(a[12]), .B(b[1]), .Z(n595) );
  NAND U758 ( .A(b[2]), .B(a[11]), .Z(n596) );
  NAND U759 ( .A(b[3]), .B(a[10]), .Z(n594) );
  XNOR U760 ( .A(n596), .B(n594), .Z(n578) );
  XNOR U761 ( .A(n595), .B(n578), .Z(n588) );
  NAND U762 ( .A(a[13]), .B(b[0]), .Z(n589) );
  XOR U763 ( .A(n591), .B(n590), .Z(n585) );
  XOR U764 ( .A(n584), .B(n585), .Z(n599) );
  XOR U765 ( .A(n598), .B(sreg[73]), .Z(n581) );
  XNOR U766 ( .A(n599), .B(n581), .Z(c[73]) );
  NANDN U767 ( .A(n583), .B(n582), .Z(n587) );
  NANDN U768 ( .A(n585), .B(n584), .Z(n586) );
  NAND U769 ( .A(n587), .B(n586), .Z(n601) );
  NANDN U770 ( .A(n589), .B(n588), .Z(n593) );
  NANDN U771 ( .A(n591), .B(n590), .Z(n592) );
  AND U772 ( .A(n593), .B(n592), .Z(n602) );
  XNOR U773 ( .A(n601), .B(n602), .Z(n603) );
  AND U774 ( .A(a[13]), .B(b[1]), .Z(n614) );
  NAND U775 ( .A(b[2]), .B(a[12]), .Z(n615) );
  NAND U776 ( .A(b[3]), .B(a[11]), .Z(n613) );
  XNOR U777 ( .A(n615), .B(n613), .Z(n597) );
  XNOR U778 ( .A(n614), .B(n597), .Z(n607) );
  NAND U779 ( .A(a[14]), .B(b[0]), .Z(n608) );
  XOR U780 ( .A(n610), .B(n609), .Z(n604) );
  XOR U781 ( .A(n603), .B(n604), .Z(n618) );
  XOR U782 ( .A(n617), .B(sreg[74]), .Z(n600) );
  XNOR U783 ( .A(n618), .B(n600), .Z(c[74]) );
  NANDN U784 ( .A(n602), .B(n601), .Z(n606) );
  NANDN U785 ( .A(n604), .B(n603), .Z(n605) );
  NAND U786 ( .A(n606), .B(n605), .Z(n620) );
  NANDN U787 ( .A(n608), .B(n607), .Z(n612) );
  NANDN U788 ( .A(n610), .B(n609), .Z(n611) );
  AND U789 ( .A(n612), .B(n611), .Z(n621) );
  XNOR U790 ( .A(n620), .B(n621), .Z(n622) );
  AND U791 ( .A(a[14]), .B(b[1]), .Z(n633) );
  NAND U792 ( .A(b[2]), .B(a[13]), .Z(n634) );
  NAND U793 ( .A(b[3]), .B(a[12]), .Z(n632) );
  XNOR U794 ( .A(n634), .B(n632), .Z(n616) );
  XNOR U795 ( .A(n633), .B(n616), .Z(n626) );
  NAND U796 ( .A(a[15]), .B(b[0]), .Z(n627) );
  XOR U797 ( .A(n629), .B(n628), .Z(n623) );
  XOR U798 ( .A(n622), .B(n623), .Z(n637) );
  XOR U799 ( .A(n636), .B(sreg[75]), .Z(n619) );
  XNOR U800 ( .A(n637), .B(n619), .Z(c[75]) );
  NANDN U801 ( .A(n621), .B(n620), .Z(n625) );
  NANDN U802 ( .A(n623), .B(n622), .Z(n624) );
  NAND U803 ( .A(n625), .B(n624), .Z(n639) );
  NANDN U804 ( .A(n627), .B(n626), .Z(n631) );
  NANDN U805 ( .A(n629), .B(n628), .Z(n630) );
  AND U806 ( .A(n631), .B(n630), .Z(n640) );
  XNOR U807 ( .A(n639), .B(n640), .Z(n641) );
  AND U808 ( .A(a[15]), .B(b[1]), .Z(n652) );
  NAND U809 ( .A(b[2]), .B(a[14]), .Z(n653) );
  NAND U810 ( .A(b[3]), .B(a[13]), .Z(n651) );
  XNOR U811 ( .A(n653), .B(n651), .Z(n635) );
  XNOR U812 ( .A(n652), .B(n635), .Z(n645) );
  NAND U813 ( .A(a[16]), .B(b[0]), .Z(n646) );
  XOR U814 ( .A(n648), .B(n647), .Z(n642) );
  XOR U815 ( .A(n641), .B(n642), .Z(n656) );
  XOR U816 ( .A(n655), .B(sreg[76]), .Z(n638) );
  XNOR U817 ( .A(n656), .B(n638), .Z(c[76]) );
  NANDN U818 ( .A(n640), .B(n639), .Z(n644) );
  NANDN U819 ( .A(n642), .B(n641), .Z(n643) );
  NAND U820 ( .A(n644), .B(n643), .Z(n658) );
  NANDN U821 ( .A(n646), .B(n645), .Z(n650) );
  NANDN U822 ( .A(n648), .B(n647), .Z(n649) );
  AND U823 ( .A(n650), .B(n649), .Z(n659) );
  XNOR U824 ( .A(n658), .B(n659), .Z(n660) );
  AND U825 ( .A(a[16]), .B(b[1]), .Z(n671) );
  NAND U826 ( .A(b[2]), .B(a[15]), .Z(n672) );
  NAND U827 ( .A(b[3]), .B(a[14]), .Z(n670) );
  XNOR U828 ( .A(n672), .B(n670), .Z(n654) );
  XNOR U829 ( .A(n671), .B(n654), .Z(n664) );
  NAND U830 ( .A(a[17]), .B(b[0]), .Z(n665) );
  XOR U831 ( .A(n667), .B(n666), .Z(n661) );
  XOR U832 ( .A(n660), .B(n661), .Z(n675) );
  XOR U833 ( .A(n674), .B(sreg[77]), .Z(n657) );
  XNOR U834 ( .A(n675), .B(n657), .Z(c[77]) );
  NANDN U835 ( .A(n659), .B(n658), .Z(n663) );
  NANDN U836 ( .A(n661), .B(n660), .Z(n662) );
  NAND U837 ( .A(n663), .B(n662), .Z(n677) );
  NANDN U838 ( .A(n665), .B(n664), .Z(n669) );
  NANDN U839 ( .A(n667), .B(n666), .Z(n668) );
  AND U840 ( .A(n669), .B(n668), .Z(n678) );
  XNOR U841 ( .A(n677), .B(n678), .Z(n679) );
  AND U842 ( .A(a[17]), .B(b[1]), .Z(n690) );
  NAND U843 ( .A(b[2]), .B(a[16]), .Z(n691) );
  NAND U844 ( .A(b[3]), .B(a[15]), .Z(n689) );
  XNOR U845 ( .A(n691), .B(n689), .Z(n673) );
  XNOR U846 ( .A(n690), .B(n673), .Z(n683) );
  NAND U847 ( .A(a[18]), .B(b[0]), .Z(n684) );
  XOR U848 ( .A(n686), .B(n685), .Z(n680) );
  XOR U849 ( .A(n679), .B(n680), .Z(n694) );
  XOR U850 ( .A(n693), .B(sreg[78]), .Z(n676) );
  XNOR U851 ( .A(n694), .B(n676), .Z(c[78]) );
  NANDN U852 ( .A(n678), .B(n677), .Z(n682) );
  NANDN U853 ( .A(n680), .B(n679), .Z(n681) );
  NAND U854 ( .A(n682), .B(n681), .Z(n696) );
  NANDN U855 ( .A(n684), .B(n683), .Z(n688) );
  NANDN U856 ( .A(n686), .B(n685), .Z(n687) );
  AND U857 ( .A(n688), .B(n687), .Z(n697) );
  XNOR U858 ( .A(n696), .B(n697), .Z(n698) );
  AND U859 ( .A(a[18]), .B(b[1]), .Z(n709) );
  NAND U860 ( .A(b[2]), .B(a[17]), .Z(n710) );
  NAND U861 ( .A(b[3]), .B(a[16]), .Z(n708) );
  XNOR U862 ( .A(n710), .B(n708), .Z(n692) );
  XNOR U863 ( .A(n709), .B(n692), .Z(n702) );
  NAND U864 ( .A(a[19]), .B(b[0]), .Z(n703) );
  XOR U865 ( .A(n705), .B(n704), .Z(n699) );
  XOR U866 ( .A(n698), .B(n699), .Z(n713) );
  XOR U867 ( .A(n712), .B(sreg[79]), .Z(n695) );
  XNOR U868 ( .A(n713), .B(n695), .Z(c[79]) );
  NANDN U869 ( .A(n697), .B(n696), .Z(n701) );
  NANDN U870 ( .A(n699), .B(n698), .Z(n700) );
  NAND U871 ( .A(n701), .B(n700), .Z(n715) );
  NANDN U872 ( .A(n703), .B(n702), .Z(n707) );
  NANDN U873 ( .A(n705), .B(n704), .Z(n706) );
  AND U874 ( .A(n707), .B(n706), .Z(n716) );
  XNOR U875 ( .A(n715), .B(n716), .Z(n717) );
  AND U876 ( .A(a[19]), .B(b[1]), .Z(n728) );
  NAND U877 ( .A(b[2]), .B(a[18]), .Z(n729) );
  NAND U878 ( .A(b[3]), .B(a[17]), .Z(n727) );
  XNOR U879 ( .A(n729), .B(n727), .Z(n711) );
  XNOR U880 ( .A(n728), .B(n711), .Z(n721) );
  NAND U881 ( .A(a[20]), .B(b[0]), .Z(n722) );
  XOR U882 ( .A(n724), .B(n723), .Z(n718) );
  XOR U883 ( .A(n717), .B(n718), .Z(n732) );
  XOR U884 ( .A(n731), .B(sreg[80]), .Z(n714) );
  XNOR U885 ( .A(n732), .B(n714), .Z(c[80]) );
  NANDN U886 ( .A(n716), .B(n715), .Z(n720) );
  NANDN U887 ( .A(n718), .B(n717), .Z(n719) );
  NAND U888 ( .A(n720), .B(n719), .Z(n734) );
  NANDN U889 ( .A(n722), .B(n721), .Z(n726) );
  NANDN U890 ( .A(n724), .B(n723), .Z(n725) );
  AND U891 ( .A(n726), .B(n725), .Z(n735) );
  XNOR U892 ( .A(n734), .B(n735), .Z(n736) );
  AND U893 ( .A(a[20]), .B(b[1]), .Z(n747) );
  NAND U894 ( .A(b[2]), .B(a[19]), .Z(n748) );
  NAND U895 ( .A(b[3]), .B(a[18]), .Z(n746) );
  XNOR U896 ( .A(n748), .B(n746), .Z(n730) );
  XNOR U897 ( .A(n747), .B(n730), .Z(n740) );
  NAND U898 ( .A(a[21]), .B(b[0]), .Z(n741) );
  XOR U899 ( .A(n743), .B(n742), .Z(n737) );
  XOR U900 ( .A(n736), .B(n737), .Z(n751) );
  XOR U901 ( .A(n750), .B(sreg[81]), .Z(n733) );
  XNOR U902 ( .A(n751), .B(n733), .Z(c[81]) );
  NANDN U903 ( .A(n735), .B(n734), .Z(n739) );
  NANDN U904 ( .A(n737), .B(n736), .Z(n738) );
  NAND U905 ( .A(n739), .B(n738), .Z(n753) );
  NANDN U906 ( .A(n741), .B(n740), .Z(n745) );
  NANDN U907 ( .A(n743), .B(n742), .Z(n744) );
  AND U908 ( .A(n745), .B(n744), .Z(n754) );
  XNOR U909 ( .A(n753), .B(n754), .Z(n755) );
  AND U910 ( .A(a[21]), .B(b[1]), .Z(n766) );
  NAND U911 ( .A(b[2]), .B(a[20]), .Z(n767) );
  NAND U912 ( .A(b[3]), .B(a[19]), .Z(n765) );
  XNOR U913 ( .A(n767), .B(n765), .Z(n749) );
  XNOR U914 ( .A(n766), .B(n749), .Z(n759) );
  NAND U915 ( .A(a[22]), .B(b[0]), .Z(n760) );
  XOR U916 ( .A(n762), .B(n761), .Z(n756) );
  XOR U917 ( .A(n755), .B(n756), .Z(n770) );
  XOR U918 ( .A(n769), .B(sreg[82]), .Z(n752) );
  XNOR U919 ( .A(n770), .B(n752), .Z(c[82]) );
  NANDN U920 ( .A(n754), .B(n753), .Z(n758) );
  NANDN U921 ( .A(n756), .B(n755), .Z(n757) );
  NAND U922 ( .A(n758), .B(n757), .Z(n772) );
  NANDN U923 ( .A(n760), .B(n759), .Z(n764) );
  NANDN U924 ( .A(n762), .B(n761), .Z(n763) );
  AND U925 ( .A(n764), .B(n763), .Z(n773) );
  XNOR U926 ( .A(n772), .B(n773), .Z(n774) );
  AND U927 ( .A(a[22]), .B(b[1]), .Z(n785) );
  NAND U928 ( .A(b[2]), .B(a[21]), .Z(n786) );
  NAND U929 ( .A(b[3]), .B(a[20]), .Z(n784) );
  XNOR U930 ( .A(n786), .B(n784), .Z(n768) );
  XNOR U931 ( .A(n785), .B(n768), .Z(n778) );
  NAND U932 ( .A(a[23]), .B(b[0]), .Z(n779) );
  XOR U933 ( .A(n781), .B(n780), .Z(n775) );
  XOR U934 ( .A(n774), .B(n775), .Z(n789) );
  XOR U935 ( .A(n788), .B(sreg[83]), .Z(n771) );
  XNOR U936 ( .A(n789), .B(n771), .Z(c[83]) );
  NANDN U937 ( .A(n773), .B(n772), .Z(n777) );
  NANDN U938 ( .A(n775), .B(n774), .Z(n776) );
  NAND U939 ( .A(n777), .B(n776), .Z(n791) );
  NANDN U940 ( .A(n779), .B(n778), .Z(n783) );
  NANDN U941 ( .A(n781), .B(n780), .Z(n782) );
  AND U942 ( .A(n783), .B(n782), .Z(n792) );
  XNOR U943 ( .A(n791), .B(n792), .Z(n793) );
  AND U944 ( .A(a[23]), .B(b[1]), .Z(n804) );
  NAND U945 ( .A(b[2]), .B(a[22]), .Z(n805) );
  NAND U946 ( .A(b[3]), .B(a[21]), .Z(n803) );
  XNOR U947 ( .A(n805), .B(n803), .Z(n787) );
  XNOR U948 ( .A(n804), .B(n787), .Z(n797) );
  NAND U949 ( .A(a[24]), .B(b[0]), .Z(n798) );
  XOR U950 ( .A(n800), .B(n799), .Z(n794) );
  XOR U951 ( .A(n793), .B(n794), .Z(n808) );
  XOR U952 ( .A(n807), .B(sreg[84]), .Z(n790) );
  XNOR U953 ( .A(n808), .B(n790), .Z(c[84]) );
  NANDN U954 ( .A(n792), .B(n791), .Z(n796) );
  NANDN U955 ( .A(n794), .B(n793), .Z(n795) );
  NAND U956 ( .A(n796), .B(n795), .Z(n810) );
  NANDN U957 ( .A(n798), .B(n797), .Z(n802) );
  NANDN U958 ( .A(n800), .B(n799), .Z(n801) );
  AND U959 ( .A(n802), .B(n801), .Z(n811) );
  XNOR U960 ( .A(n810), .B(n811), .Z(n812) );
  AND U961 ( .A(a[24]), .B(b[1]), .Z(n823) );
  NAND U962 ( .A(b[2]), .B(a[23]), .Z(n824) );
  NAND U963 ( .A(b[3]), .B(a[22]), .Z(n822) );
  XNOR U964 ( .A(n824), .B(n822), .Z(n806) );
  XNOR U965 ( .A(n823), .B(n806), .Z(n816) );
  NAND U966 ( .A(a[25]), .B(b[0]), .Z(n817) );
  XOR U967 ( .A(n819), .B(n818), .Z(n813) );
  XOR U968 ( .A(n812), .B(n813), .Z(n827) );
  XOR U969 ( .A(n826), .B(sreg[85]), .Z(n809) );
  XNOR U970 ( .A(n827), .B(n809), .Z(c[85]) );
  NANDN U971 ( .A(n811), .B(n810), .Z(n815) );
  NANDN U972 ( .A(n813), .B(n812), .Z(n814) );
  NAND U973 ( .A(n815), .B(n814), .Z(n829) );
  NANDN U974 ( .A(n817), .B(n816), .Z(n821) );
  NANDN U975 ( .A(n819), .B(n818), .Z(n820) );
  AND U976 ( .A(n821), .B(n820), .Z(n830) );
  XNOR U977 ( .A(n829), .B(n830), .Z(n831) );
  AND U978 ( .A(a[25]), .B(b[1]), .Z(n842) );
  NAND U979 ( .A(b[2]), .B(a[24]), .Z(n843) );
  NAND U980 ( .A(b[3]), .B(a[23]), .Z(n841) );
  XNOR U981 ( .A(n843), .B(n841), .Z(n825) );
  XNOR U982 ( .A(n842), .B(n825), .Z(n835) );
  NAND U983 ( .A(a[26]), .B(b[0]), .Z(n836) );
  XOR U984 ( .A(n838), .B(n837), .Z(n832) );
  XOR U985 ( .A(n831), .B(n832), .Z(n846) );
  XOR U986 ( .A(n845), .B(sreg[86]), .Z(n828) );
  XNOR U987 ( .A(n846), .B(n828), .Z(c[86]) );
  NANDN U988 ( .A(n830), .B(n829), .Z(n834) );
  NANDN U989 ( .A(n832), .B(n831), .Z(n833) );
  NAND U990 ( .A(n834), .B(n833), .Z(n848) );
  NANDN U991 ( .A(n836), .B(n835), .Z(n840) );
  NANDN U992 ( .A(n838), .B(n837), .Z(n839) );
  AND U993 ( .A(n840), .B(n839), .Z(n849) );
  XNOR U994 ( .A(n848), .B(n849), .Z(n850) );
  AND U995 ( .A(a[26]), .B(b[1]), .Z(n861) );
  NAND U996 ( .A(b[2]), .B(a[25]), .Z(n862) );
  NAND U997 ( .A(b[3]), .B(a[24]), .Z(n860) );
  XNOR U998 ( .A(n862), .B(n860), .Z(n844) );
  XNOR U999 ( .A(n861), .B(n844), .Z(n854) );
  NAND U1000 ( .A(a[27]), .B(b[0]), .Z(n855) );
  XOR U1001 ( .A(n857), .B(n856), .Z(n851) );
  XOR U1002 ( .A(n850), .B(n851), .Z(n865) );
  XOR U1003 ( .A(n864), .B(sreg[87]), .Z(n847) );
  XNOR U1004 ( .A(n865), .B(n847), .Z(c[87]) );
  NANDN U1005 ( .A(n849), .B(n848), .Z(n853) );
  NANDN U1006 ( .A(n851), .B(n850), .Z(n852) );
  NAND U1007 ( .A(n853), .B(n852), .Z(n867) );
  NANDN U1008 ( .A(n855), .B(n854), .Z(n859) );
  NANDN U1009 ( .A(n857), .B(n856), .Z(n858) );
  AND U1010 ( .A(n859), .B(n858), .Z(n868) );
  XNOR U1011 ( .A(n867), .B(n868), .Z(n869) );
  AND U1012 ( .A(a[27]), .B(b[1]), .Z(n880) );
  NAND U1013 ( .A(b[2]), .B(a[26]), .Z(n881) );
  NAND U1014 ( .A(b[3]), .B(a[25]), .Z(n879) );
  XNOR U1015 ( .A(n881), .B(n879), .Z(n863) );
  XNOR U1016 ( .A(n880), .B(n863), .Z(n873) );
  NAND U1017 ( .A(a[28]), .B(b[0]), .Z(n874) );
  XOR U1018 ( .A(n876), .B(n875), .Z(n870) );
  XOR U1019 ( .A(n869), .B(n870), .Z(n884) );
  XOR U1020 ( .A(n883), .B(sreg[88]), .Z(n866) );
  XNOR U1021 ( .A(n884), .B(n866), .Z(c[88]) );
  NANDN U1022 ( .A(n868), .B(n867), .Z(n872) );
  NANDN U1023 ( .A(n870), .B(n869), .Z(n871) );
  NAND U1024 ( .A(n872), .B(n871), .Z(n886) );
  NANDN U1025 ( .A(n874), .B(n873), .Z(n878) );
  NANDN U1026 ( .A(n876), .B(n875), .Z(n877) );
  AND U1027 ( .A(n878), .B(n877), .Z(n887) );
  XNOR U1028 ( .A(n886), .B(n887), .Z(n888) );
  AND U1029 ( .A(a[28]), .B(b[1]), .Z(n899) );
  NAND U1030 ( .A(b[2]), .B(a[27]), .Z(n900) );
  NAND U1031 ( .A(b[3]), .B(a[26]), .Z(n898) );
  XNOR U1032 ( .A(n900), .B(n898), .Z(n882) );
  XNOR U1033 ( .A(n899), .B(n882), .Z(n892) );
  NAND U1034 ( .A(a[29]), .B(b[0]), .Z(n893) );
  XOR U1035 ( .A(n895), .B(n894), .Z(n889) );
  XOR U1036 ( .A(n888), .B(n889), .Z(n903) );
  XOR U1037 ( .A(n902), .B(sreg[89]), .Z(n885) );
  XNOR U1038 ( .A(n903), .B(n885), .Z(c[89]) );
  NANDN U1039 ( .A(n887), .B(n886), .Z(n891) );
  NANDN U1040 ( .A(n889), .B(n888), .Z(n890) );
  NAND U1041 ( .A(n891), .B(n890), .Z(n905) );
  NANDN U1042 ( .A(n893), .B(n892), .Z(n897) );
  NANDN U1043 ( .A(n895), .B(n894), .Z(n896) );
  AND U1044 ( .A(n897), .B(n896), .Z(n906) );
  XNOR U1045 ( .A(n905), .B(n906), .Z(n907) );
  AND U1046 ( .A(a[29]), .B(b[1]), .Z(n918) );
  NAND U1047 ( .A(b[2]), .B(a[28]), .Z(n919) );
  NAND U1048 ( .A(b[3]), .B(a[27]), .Z(n917) );
  XNOR U1049 ( .A(n919), .B(n917), .Z(n901) );
  XNOR U1050 ( .A(n918), .B(n901), .Z(n911) );
  NAND U1051 ( .A(a[30]), .B(b[0]), .Z(n912) );
  XOR U1052 ( .A(n914), .B(n913), .Z(n908) );
  XOR U1053 ( .A(n907), .B(n908), .Z(n922) );
  XOR U1054 ( .A(n921), .B(sreg[90]), .Z(n904) );
  XNOR U1055 ( .A(n922), .B(n904), .Z(c[90]) );
  NANDN U1056 ( .A(n906), .B(n905), .Z(n910) );
  NANDN U1057 ( .A(n908), .B(n907), .Z(n909) );
  NAND U1058 ( .A(n910), .B(n909), .Z(n924) );
  NANDN U1059 ( .A(n912), .B(n911), .Z(n916) );
  NANDN U1060 ( .A(n914), .B(n913), .Z(n915) );
  AND U1061 ( .A(n916), .B(n915), .Z(n925) );
  XNOR U1062 ( .A(n924), .B(n925), .Z(n926) );
  AND U1063 ( .A(a[30]), .B(b[1]), .Z(n937) );
  NAND U1064 ( .A(b[2]), .B(a[29]), .Z(n938) );
  NAND U1065 ( .A(b[3]), .B(a[28]), .Z(n936) );
  XNOR U1066 ( .A(n938), .B(n936), .Z(n920) );
  XNOR U1067 ( .A(n937), .B(n920), .Z(n930) );
  NAND U1068 ( .A(a[31]), .B(b[0]), .Z(n931) );
  XOR U1069 ( .A(n933), .B(n932), .Z(n927) );
  XOR U1070 ( .A(n926), .B(n927), .Z(n941) );
  XOR U1071 ( .A(n940), .B(sreg[91]), .Z(n923) );
  XNOR U1072 ( .A(n941), .B(n923), .Z(c[91]) );
  NANDN U1073 ( .A(n925), .B(n924), .Z(n929) );
  NANDN U1074 ( .A(n927), .B(n926), .Z(n928) );
  NAND U1075 ( .A(n929), .B(n928), .Z(n943) );
  NANDN U1076 ( .A(n931), .B(n930), .Z(n935) );
  NANDN U1077 ( .A(n933), .B(n932), .Z(n934) );
  AND U1078 ( .A(n935), .B(n934), .Z(n944) );
  XNOR U1079 ( .A(n943), .B(n944), .Z(n945) );
  AND U1080 ( .A(a[31]), .B(b[1]), .Z(n956) );
  NAND U1081 ( .A(b[2]), .B(a[30]), .Z(n957) );
  NAND U1082 ( .A(b[3]), .B(a[29]), .Z(n955) );
  XNOR U1083 ( .A(n957), .B(n955), .Z(n939) );
  XNOR U1084 ( .A(n956), .B(n939), .Z(n949) );
  NAND U1085 ( .A(a[32]), .B(b[0]), .Z(n950) );
  XOR U1086 ( .A(n952), .B(n951), .Z(n946) );
  XOR U1087 ( .A(n945), .B(n946), .Z(n960) );
  XOR U1088 ( .A(n959), .B(sreg[92]), .Z(n942) );
  XNOR U1089 ( .A(n960), .B(n942), .Z(c[92]) );
  NANDN U1090 ( .A(n944), .B(n943), .Z(n948) );
  NANDN U1091 ( .A(n946), .B(n945), .Z(n947) );
  NAND U1092 ( .A(n948), .B(n947), .Z(n962) );
  NANDN U1093 ( .A(n950), .B(n949), .Z(n954) );
  NANDN U1094 ( .A(n952), .B(n951), .Z(n953) );
  AND U1095 ( .A(n954), .B(n953), .Z(n963) );
  XNOR U1096 ( .A(n962), .B(n963), .Z(n964) );
  AND U1097 ( .A(a[32]), .B(b[1]), .Z(n975) );
  NAND U1098 ( .A(b[2]), .B(a[31]), .Z(n976) );
  NAND U1099 ( .A(b[3]), .B(a[30]), .Z(n974) );
  XNOR U1100 ( .A(n976), .B(n974), .Z(n958) );
  XNOR U1101 ( .A(n975), .B(n958), .Z(n968) );
  NAND U1102 ( .A(a[33]), .B(b[0]), .Z(n969) );
  XOR U1103 ( .A(n971), .B(n970), .Z(n965) );
  XOR U1104 ( .A(n964), .B(n965), .Z(n979) );
  XOR U1105 ( .A(n978), .B(sreg[93]), .Z(n961) );
  XNOR U1106 ( .A(n979), .B(n961), .Z(c[93]) );
  NANDN U1107 ( .A(n963), .B(n962), .Z(n967) );
  NANDN U1108 ( .A(n965), .B(n964), .Z(n966) );
  NAND U1109 ( .A(n967), .B(n966), .Z(n981) );
  NANDN U1110 ( .A(n969), .B(n968), .Z(n973) );
  NANDN U1111 ( .A(n971), .B(n970), .Z(n972) );
  AND U1112 ( .A(n973), .B(n972), .Z(n982) );
  XNOR U1113 ( .A(n981), .B(n982), .Z(n983) );
  AND U1114 ( .A(a[33]), .B(b[1]), .Z(n994) );
  NAND U1115 ( .A(b[2]), .B(a[32]), .Z(n995) );
  NAND U1116 ( .A(b[3]), .B(a[31]), .Z(n993) );
  XNOR U1117 ( .A(n995), .B(n993), .Z(n977) );
  XNOR U1118 ( .A(n994), .B(n977), .Z(n987) );
  NAND U1119 ( .A(a[34]), .B(b[0]), .Z(n988) );
  XOR U1120 ( .A(n990), .B(n989), .Z(n984) );
  XOR U1121 ( .A(n983), .B(n984), .Z(n998) );
  XOR U1122 ( .A(n997), .B(sreg[94]), .Z(n980) );
  XNOR U1123 ( .A(n998), .B(n980), .Z(c[94]) );
  NANDN U1124 ( .A(n982), .B(n981), .Z(n986) );
  NANDN U1125 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1126 ( .A(n986), .B(n985), .Z(n1000) );
  NANDN U1127 ( .A(n988), .B(n987), .Z(n992) );
  NANDN U1128 ( .A(n990), .B(n989), .Z(n991) );
  AND U1129 ( .A(n992), .B(n991), .Z(n1001) );
  XNOR U1130 ( .A(n1000), .B(n1001), .Z(n1002) );
  AND U1131 ( .A(a[34]), .B(b[1]), .Z(n1013) );
  NAND U1132 ( .A(b[2]), .B(a[33]), .Z(n1014) );
  NAND U1133 ( .A(b[3]), .B(a[32]), .Z(n1012) );
  XNOR U1134 ( .A(n1014), .B(n1012), .Z(n996) );
  XNOR U1135 ( .A(n1013), .B(n996), .Z(n1006) );
  NAND U1136 ( .A(a[35]), .B(b[0]), .Z(n1007) );
  XOR U1137 ( .A(n1009), .B(n1008), .Z(n1003) );
  XOR U1138 ( .A(n1002), .B(n1003), .Z(n1017) );
  XOR U1139 ( .A(n1016), .B(sreg[95]), .Z(n999) );
  XNOR U1140 ( .A(n1017), .B(n999), .Z(c[95]) );
  NANDN U1141 ( .A(n1001), .B(n1000), .Z(n1005) );
  NANDN U1142 ( .A(n1003), .B(n1002), .Z(n1004) );
  NAND U1143 ( .A(n1005), .B(n1004), .Z(n1019) );
  NANDN U1144 ( .A(n1007), .B(n1006), .Z(n1011) );
  NANDN U1145 ( .A(n1009), .B(n1008), .Z(n1010) );
  AND U1146 ( .A(n1011), .B(n1010), .Z(n1020) );
  XNOR U1147 ( .A(n1019), .B(n1020), .Z(n1021) );
  AND U1148 ( .A(a[35]), .B(b[1]), .Z(n1032) );
  NAND U1149 ( .A(b[2]), .B(a[34]), .Z(n1033) );
  NAND U1150 ( .A(b[3]), .B(a[33]), .Z(n1031) );
  XNOR U1151 ( .A(n1033), .B(n1031), .Z(n1015) );
  XNOR U1152 ( .A(n1032), .B(n1015), .Z(n1025) );
  NAND U1153 ( .A(a[36]), .B(b[0]), .Z(n1026) );
  XOR U1154 ( .A(n1028), .B(n1027), .Z(n1022) );
  XOR U1155 ( .A(n1021), .B(n1022), .Z(n1036) );
  XOR U1156 ( .A(n1035), .B(sreg[96]), .Z(n1018) );
  XNOR U1157 ( .A(n1036), .B(n1018), .Z(c[96]) );
  NANDN U1158 ( .A(n1020), .B(n1019), .Z(n1024) );
  NANDN U1159 ( .A(n1022), .B(n1021), .Z(n1023) );
  NAND U1160 ( .A(n1024), .B(n1023), .Z(n1038) );
  NANDN U1161 ( .A(n1026), .B(n1025), .Z(n1030) );
  NANDN U1162 ( .A(n1028), .B(n1027), .Z(n1029) );
  AND U1163 ( .A(n1030), .B(n1029), .Z(n1039) );
  XNOR U1164 ( .A(n1038), .B(n1039), .Z(n1040) );
  AND U1165 ( .A(a[36]), .B(b[1]), .Z(n1051) );
  NAND U1166 ( .A(b[2]), .B(a[35]), .Z(n1052) );
  NAND U1167 ( .A(b[3]), .B(a[34]), .Z(n1050) );
  XNOR U1168 ( .A(n1052), .B(n1050), .Z(n1034) );
  XNOR U1169 ( .A(n1051), .B(n1034), .Z(n1044) );
  NAND U1170 ( .A(a[37]), .B(b[0]), .Z(n1045) );
  XOR U1171 ( .A(n1047), .B(n1046), .Z(n1041) );
  XOR U1172 ( .A(n1040), .B(n1041), .Z(n1055) );
  XOR U1173 ( .A(n1054), .B(sreg[97]), .Z(n1037) );
  XNOR U1174 ( .A(n1055), .B(n1037), .Z(c[97]) );
  NANDN U1175 ( .A(n1039), .B(n1038), .Z(n1043) );
  NANDN U1176 ( .A(n1041), .B(n1040), .Z(n1042) );
  NAND U1177 ( .A(n1043), .B(n1042), .Z(n1057) );
  NANDN U1178 ( .A(n1045), .B(n1044), .Z(n1049) );
  NANDN U1179 ( .A(n1047), .B(n1046), .Z(n1048) );
  AND U1180 ( .A(n1049), .B(n1048), .Z(n1058) );
  XNOR U1181 ( .A(n1057), .B(n1058), .Z(n1059) );
  AND U1182 ( .A(a[37]), .B(b[1]), .Z(n1070) );
  NAND U1183 ( .A(b[2]), .B(a[36]), .Z(n1071) );
  NAND U1184 ( .A(b[3]), .B(a[35]), .Z(n1069) );
  XNOR U1185 ( .A(n1071), .B(n1069), .Z(n1053) );
  XNOR U1186 ( .A(n1070), .B(n1053), .Z(n1063) );
  NAND U1187 ( .A(a[38]), .B(b[0]), .Z(n1064) );
  XOR U1188 ( .A(n1066), .B(n1065), .Z(n1060) );
  XOR U1189 ( .A(n1059), .B(n1060), .Z(n1074) );
  XOR U1190 ( .A(n1073), .B(sreg[98]), .Z(n1056) );
  XNOR U1191 ( .A(n1074), .B(n1056), .Z(c[98]) );
  NANDN U1192 ( .A(n1058), .B(n1057), .Z(n1062) );
  NANDN U1193 ( .A(n1060), .B(n1059), .Z(n1061) );
  NAND U1194 ( .A(n1062), .B(n1061), .Z(n1076) );
  NANDN U1195 ( .A(n1064), .B(n1063), .Z(n1068) );
  NANDN U1196 ( .A(n1066), .B(n1065), .Z(n1067) );
  AND U1197 ( .A(n1068), .B(n1067), .Z(n1077) );
  XNOR U1198 ( .A(n1076), .B(n1077), .Z(n1078) );
  AND U1199 ( .A(a[38]), .B(b[1]), .Z(n1089) );
  NAND U1200 ( .A(b[2]), .B(a[37]), .Z(n1090) );
  NAND U1201 ( .A(b[3]), .B(a[36]), .Z(n1088) );
  XNOR U1202 ( .A(n1090), .B(n1088), .Z(n1072) );
  XNOR U1203 ( .A(n1089), .B(n1072), .Z(n1082) );
  NAND U1204 ( .A(a[39]), .B(b[0]), .Z(n1083) );
  XOR U1205 ( .A(n1085), .B(n1084), .Z(n1079) );
  XOR U1206 ( .A(n1078), .B(n1079), .Z(n1093) );
  XOR U1207 ( .A(n1092), .B(sreg[99]), .Z(n1075) );
  XNOR U1208 ( .A(n1093), .B(n1075), .Z(c[99]) );
  NANDN U1209 ( .A(n1077), .B(n1076), .Z(n1081) );
  NANDN U1210 ( .A(n1079), .B(n1078), .Z(n1080) );
  NAND U1211 ( .A(n1081), .B(n1080), .Z(n1095) );
  NANDN U1212 ( .A(n1083), .B(n1082), .Z(n1087) );
  NANDN U1213 ( .A(n1085), .B(n1084), .Z(n1086) );
  AND U1214 ( .A(n1087), .B(n1086), .Z(n1096) );
  XNOR U1215 ( .A(n1095), .B(n1096), .Z(n1097) );
  AND U1216 ( .A(a[39]), .B(b[1]), .Z(n1108) );
  NAND U1217 ( .A(b[2]), .B(a[38]), .Z(n1109) );
  NAND U1218 ( .A(b[3]), .B(a[37]), .Z(n1107) );
  XNOR U1219 ( .A(n1109), .B(n1107), .Z(n1091) );
  XNOR U1220 ( .A(n1108), .B(n1091), .Z(n1101) );
  NAND U1221 ( .A(a[40]), .B(b[0]), .Z(n1102) );
  XOR U1222 ( .A(n1104), .B(n1103), .Z(n1098) );
  XOR U1223 ( .A(n1097), .B(n1098), .Z(n1112) );
  XOR U1224 ( .A(n1111), .B(sreg[100]), .Z(n1094) );
  XNOR U1225 ( .A(n1112), .B(n1094), .Z(c[100]) );
  NANDN U1226 ( .A(n1096), .B(n1095), .Z(n1100) );
  NANDN U1227 ( .A(n1098), .B(n1097), .Z(n1099) );
  NAND U1228 ( .A(n1100), .B(n1099), .Z(n1114) );
  NANDN U1229 ( .A(n1102), .B(n1101), .Z(n1106) );
  NANDN U1230 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U1231 ( .A(n1106), .B(n1105), .Z(n1115) );
  XNOR U1232 ( .A(n1114), .B(n1115), .Z(n1116) );
  AND U1233 ( .A(a[40]), .B(b[1]), .Z(n1127) );
  NAND U1234 ( .A(b[2]), .B(a[39]), .Z(n1128) );
  NAND U1235 ( .A(b[3]), .B(a[38]), .Z(n1126) );
  XNOR U1236 ( .A(n1128), .B(n1126), .Z(n1110) );
  XNOR U1237 ( .A(n1127), .B(n1110), .Z(n1120) );
  NAND U1238 ( .A(a[41]), .B(b[0]), .Z(n1121) );
  XOR U1239 ( .A(n1123), .B(n1122), .Z(n1117) );
  XOR U1240 ( .A(n1116), .B(n1117), .Z(n1131) );
  XOR U1241 ( .A(n1130), .B(sreg[101]), .Z(n1113) );
  XNOR U1242 ( .A(n1131), .B(n1113), .Z(c[101]) );
  NANDN U1243 ( .A(n1115), .B(n1114), .Z(n1119) );
  NANDN U1244 ( .A(n1117), .B(n1116), .Z(n1118) );
  NAND U1245 ( .A(n1119), .B(n1118), .Z(n1133) );
  NANDN U1246 ( .A(n1121), .B(n1120), .Z(n1125) );
  NANDN U1247 ( .A(n1123), .B(n1122), .Z(n1124) );
  AND U1248 ( .A(n1125), .B(n1124), .Z(n1134) );
  XNOR U1249 ( .A(n1133), .B(n1134), .Z(n1135) );
  AND U1250 ( .A(a[41]), .B(b[1]), .Z(n1146) );
  NAND U1251 ( .A(b[2]), .B(a[40]), .Z(n1147) );
  NAND U1252 ( .A(b[3]), .B(a[39]), .Z(n1145) );
  XNOR U1253 ( .A(n1147), .B(n1145), .Z(n1129) );
  XNOR U1254 ( .A(n1146), .B(n1129), .Z(n1139) );
  NAND U1255 ( .A(a[42]), .B(b[0]), .Z(n1140) );
  XOR U1256 ( .A(n1142), .B(n1141), .Z(n1136) );
  XOR U1257 ( .A(n1135), .B(n1136), .Z(n1150) );
  XOR U1258 ( .A(n1149), .B(sreg[102]), .Z(n1132) );
  XNOR U1259 ( .A(n1150), .B(n1132), .Z(c[102]) );
  NANDN U1260 ( .A(n1134), .B(n1133), .Z(n1138) );
  NANDN U1261 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1262 ( .A(n1138), .B(n1137), .Z(n1152) );
  NANDN U1263 ( .A(n1140), .B(n1139), .Z(n1144) );
  NANDN U1264 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U1265 ( .A(n1144), .B(n1143), .Z(n1153) );
  XNOR U1266 ( .A(n1152), .B(n1153), .Z(n1154) );
  AND U1267 ( .A(a[42]), .B(b[1]), .Z(n1165) );
  NAND U1268 ( .A(b[2]), .B(a[41]), .Z(n1166) );
  NAND U1269 ( .A(b[3]), .B(a[40]), .Z(n1164) );
  XNOR U1270 ( .A(n1166), .B(n1164), .Z(n1148) );
  XNOR U1271 ( .A(n1165), .B(n1148), .Z(n1158) );
  NAND U1272 ( .A(a[43]), .B(b[0]), .Z(n1159) );
  XOR U1273 ( .A(n1161), .B(n1160), .Z(n1155) );
  XOR U1274 ( .A(n1154), .B(n1155), .Z(n1169) );
  XOR U1275 ( .A(n1168), .B(sreg[103]), .Z(n1151) );
  XNOR U1276 ( .A(n1169), .B(n1151), .Z(c[103]) );
  NANDN U1277 ( .A(n1153), .B(n1152), .Z(n1157) );
  NANDN U1278 ( .A(n1155), .B(n1154), .Z(n1156) );
  NAND U1279 ( .A(n1157), .B(n1156), .Z(n1171) );
  NANDN U1280 ( .A(n1159), .B(n1158), .Z(n1163) );
  NANDN U1281 ( .A(n1161), .B(n1160), .Z(n1162) );
  AND U1282 ( .A(n1163), .B(n1162), .Z(n1172) );
  XNOR U1283 ( .A(n1171), .B(n1172), .Z(n1173) );
  AND U1284 ( .A(a[43]), .B(b[1]), .Z(n1184) );
  NAND U1285 ( .A(b[2]), .B(a[42]), .Z(n1185) );
  NAND U1286 ( .A(b[3]), .B(a[41]), .Z(n1183) );
  XNOR U1287 ( .A(n1185), .B(n1183), .Z(n1167) );
  XNOR U1288 ( .A(n1184), .B(n1167), .Z(n1177) );
  NAND U1289 ( .A(a[44]), .B(b[0]), .Z(n1178) );
  XOR U1290 ( .A(n1180), .B(n1179), .Z(n1174) );
  XOR U1291 ( .A(n1173), .B(n1174), .Z(n1188) );
  XOR U1292 ( .A(n1187), .B(sreg[104]), .Z(n1170) );
  XNOR U1293 ( .A(n1188), .B(n1170), .Z(c[104]) );
  NANDN U1294 ( .A(n1172), .B(n1171), .Z(n1176) );
  NANDN U1295 ( .A(n1174), .B(n1173), .Z(n1175) );
  NAND U1296 ( .A(n1176), .B(n1175), .Z(n1190) );
  NANDN U1297 ( .A(n1178), .B(n1177), .Z(n1182) );
  NANDN U1298 ( .A(n1180), .B(n1179), .Z(n1181) );
  AND U1299 ( .A(n1182), .B(n1181), .Z(n1191) );
  XNOR U1300 ( .A(n1190), .B(n1191), .Z(n1192) );
  AND U1301 ( .A(a[44]), .B(b[1]), .Z(n1203) );
  NAND U1302 ( .A(b[2]), .B(a[43]), .Z(n1204) );
  NAND U1303 ( .A(b[3]), .B(a[42]), .Z(n1202) );
  XNOR U1304 ( .A(n1204), .B(n1202), .Z(n1186) );
  XNOR U1305 ( .A(n1203), .B(n1186), .Z(n1196) );
  NAND U1306 ( .A(a[45]), .B(b[0]), .Z(n1197) );
  XOR U1307 ( .A(n1199), .B(n1198), .Z(n1193) );
  XOR U1308 ( .A(n1192), .B(n1193), .Z(n1207) );
  XOR U1309 ( .A(n1206), .B(sreg[105]), .Z(n1189) );
  XNOR U1310 ( .A(n1207), .B(n1189), .Z(c[105]) );
  NANDN U1311 ( .A(n1191), .B(n1190), .Z(n1195) );
  NANDN U1312 ( .A(n1193), .B(n1192), .Z(n1194) );
  NAND U1313 ( .A(n1195), .B(n1194), .Z(n1209) );
  NANDN U1314 ( .A(n1197), .B(n1196), .Z(n1201) );
  NANDN U1315 ( .A(n1199), .B(n1198), .Z(n1200) );
  AND U1316 ( .A(n1201), .B(n1200), .Z(n1210) );
  XNOR U1317 ( .A(n1209), .B(n1210), .Z(n1211) );
  AND U1318 ( .A(a[45]), .B(b[1]), .Z(n1222) );
  NAND U1319 ( .A(b[2]), .B(a[44]), .Z(n1223) );
  NAND U1320 ( .A(b[3]), .B(a[43]), .Z(n1221) );
  XNOR U1321 ( .A(n1223), .B(n1221), .Z(n1205) );
  XNOR U1322 ( .A(n1222), .B(n1205), .Z(n1215) );
  NAND U1323 ( .A(a[46]), .B(b[0]), .Z(n1216) );
  XOR U1324 ( .A(n1218), .B(n1217), .Z(n1212) );
  XOR U1325 ( .A(n1211), .B(n1212), .Z(n1226) );
  XOR U1326 ( .A(n1225), .B(sreg[106]), .Z(n1208) );
  XNOR U1327 ( .A(n1226), .B(n1208), .Z(c[106]) );
  NANDN U1328 ( .A(n1210), .B(n1209), .Z(n1214) );
  NANDN U1329 ( .A(n1212), .B(n1211), .Z(n1213) );
  NAND U1330 ( .A(n1214), .B(n1213), .Z(n1228) );
  NANDN U1331 ( .A(n1216), .B(n1215), .Z(n1220) );
  NANDN U1332 ( .A(n1218), .B(n1217), .Z(n1219) );
  AND U1333 ( .A(n1220), .B(n1219), .Z(n1229) );
  XNOR U1334 ( .A(n1228), .B(n1229), .Z(n1230) );
  AND U1335 ( .A(a[46]), .B(b[1]), .Z(n1241) );
  NAND U1336 ( .A(b[2]), .B(a[45]), .Z(n1242) );
  NAND U1337 ( .A(b[3]), .B(a[44]), .Z(n1240) );
  XNOR U1338 ( .A(n1242), .B(n1240), .Z(n1224) );
  XNOR U1339 ( .A(n1241), .B(n1224), .Z(n1234) );
  NAND U1340 ( .A(a[47]), .B(b[0]), .Z(n1235) );
  XOR U1341 ( .A(n1237), .B(n1236), .Z(n1231) );
  XOR U1342 ( .A(n1230), .B(n1231), .Z(n1245) );
  XOR U1343 ( .A(n1244), .B(sreg[107]), .Z(n1227) );
  XNOR U1344 ( .A(n1245), .B(n1227), .Z(c[107]) );
  NANDN U1345 ( .A(n1229), .B(n1228), .Z(n1233) );
  NANDN U1346 ( .A(n1231), .B(n1230), .Z(n1232) );
  NAND U1347 ( .A(n1233), .B(n1232), .Z(n1247) );
  NANDN U1348 ( .A(n1235), .B(n1234), .Z(n1239) );
  NANDN U1349 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U1350 ( .A(n1239), .B(n1238), .Z(n1248) );
  XNOR U1351 ( .A(n1247), .B(n1248), .Z(n1249) );
  AND U1352 ( .A(a[47]), .B(b[1]), .Z(n1260) );
  NAND U1353 ( .A(b[2]), .B(a[46]), .Z(n1261) );
  NAND U1354 ( .A(b[3]), .B(a[45]), .Z(n1259) );
  XNOR U1355 ( .A(n1261), .B(n1259), .Z(n1243) );
  XNOR U1356 ( .A(n1260), .B(n1243), .Z(n1253) );
  NAND U1357 ( .A(a[48]), .B(b[0]), .Z(n1254) );
  XOR U1358 ( .A(n1256), .B(n1255), .Z(n1250) );
  XOR U1359 ( .A(n1249), .B(n1250), .Z(n1264) );
  XOR U1360 ( .A(n1263), .B(sreg[108]), .Z(n1246) );
  XNOR U1361 ( .A(n1264), .B(n1246), .Z(c[108]) );
  NANDN U1362 ( .A(n1248), .B(n1247), .Z(n1252) );
  NANDN U1363 ( .A(n1250), .B(n1249), .Z(n1251) );
  NAND U1364 ( .A(n1252), .B(n1251), .Z(n1266) );
  NANDN U1365 ( .A(n1254), .B(n1253), .Z(n1258) );
  NANDN U1366 ( .A(n1256), .B(n1255), .Z(n1257) );
  AND U1367 ( .A(n1258), .B(n1257), .Z(n1267) );
  XNOR U1368 ( .A(n1266), .B(n1267), .Z(n1268) );
  AND U1369 ( .A(a[48]), .B(b[1]), .Z(n1279) );
  NAND U1370 ( .A(b[2]), .B(a[47]), .Z(n1280) );
  NAND U1371 ( .A(b[3]), .B(a[46]), .Z(n1278) );
  XNOR U1372 ( .A(n1280), .B(n1278), .Z(n1262) );
  XNOR U1373 ( .A(n1279), .B(n1262), .Z(n1272) );
  NAND U1374 ( .A(a[49]), .B(b[0]), .Z(n1273) );
  XOR U1375 ( .A(n1275), .B(n1274), .Z(n1269) );
  XOR U1376 ( .A(n1268), .B(n1269), .Z(n1283) );
  XOR U1377 ( .A(n1282), .B(sreg[109]), .Z(n1265) );
  XNOR U1378 ( .A(n1283), .B(n1265), .Z(c[109]) );
  NANDN U1379 ( .A(n1267), .B(n1266), .Z(n1271) );
  NANDN U1380 ( .A(n1269), .B(n1268), .Z(n1270) );
  NAND U1381 ( .A(n1271), .B(n1270), .Z(n1285) );
  NANDN U1382 ( .A(n1273), .B(n1272), .Z(n1277) );
  NANDN U1383 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U1384 ( .A(n1277), .B(n1276), .Z(n1286) );
  XNOR U1385 ( .A(n1285), .B(n1286), .Z(n1287) );
  AND U1386 ( .A(a[49]), .B(b[1]), .Z(n1298) );
  NAND U1387 ( .A(b[2]), .B(a[48]), .Z(n1299) );
  NAND U1388 ( .A(b[3]), .B(a[47]), .Z(n1297) );
  XNOR U1389 ( .A(n1299), .B(n1297), .Z(n1281) );
  XNOR U1390 ( .A(n1298), .B(n1281), .Z(n1291) );
  NAND U1391 ( .A(a[50]), .B(b[0]), .Z(n1292) );
  XOR U1392 ( .A(n1294), .B(n1293), .Z(n1288) );
  XOR U1393 ( .A(n1287), .B(n1288), .Z(n1302) );
  XOR U1394 ( .A(n1301), .B(sreg[110]), .Z(n1284) );
  XNOR U1395 ( .A(n1302), .B(n1284), .Z(c[110]) );
  NANDN U1396 ( .A(n1286), .B(n1285), .Z(n1290) );
  NANDN U1397 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U1398 ( .A(n1290), .B(n1289), .Z(n1304) );
  NANDN U1399 ( .A(n1292), .B(n1291), .Z(n1296) );
  NANDN U1400 ( .A(n1294), .B(n1293), .Z(n1295) );
  AND U1401 ( .A(n1296), .B(n1295), .Z(n1305) );
  XNOR U1402 ( .A(n1304), .B(n1305), .Z(n1306) );
  AND U1403 ( .A(a[50]), .B(b[1]), .Z(n1317) );
  NAND U1404 ( .A(b[2]), .B(a[49]), .Z(n1318) );
  NAND U1405 ( .A(b[3]), .B(a[48]), .Z(n1316) );
  XNOR U1406 ( .A(n1318), .B(n1316), .Z(n1300) );
  XNOR U1407 ( .A(n1317), .B(n1300), .Z(n1310) );
  NAND U1408 ( .A(a[51]), .B(b[0]), .Z(n1311) );
  XOR U1409 ( .A(n1313), .B(n1312), .Z(n1307) );
  XOR U1410 ( .A(n1306), .B(n1307), .Z(n1321) );
  XOR U1411 ( .A(n1320), .B(sreg[111]), .Z(n1303) );
  XNOR U1412 ( .A(n1321), .B(n1303), .Z(c[111]) );
  NANDN U1413 ( .A(n1305), .B(n1304), .Z(n1309) );
  NANDN U1414 ( .A(n1307), .B(n1306), .Z(n1308) );
  NAND U1415 ( .A(n1309), .B(n1308), .Z(n1323) );
  NANDN U1416 ( .A(n1311), .B(n1310), .Z(n1315) );
  NANDN U1417 ( .A(n1313), .B(n1312), .Z(n1314) );
  AND U1418 ( .A(n1315), .B(n1314), .Z(n1324) );
  XNOR U1419 ( .A(n1323), .B(n1324), .Z(n1325) );
  AND U1420 ( .A(a[51]), .B(b[1]), .Z(n1336) );
  NAND U1421 ( .A(b[2]), .B(a[50]), .Z(n1337) );
  NAND U1422 ( .A(b[3]), .B(a[49]), .Z(n1335) );
  XNOR U1423 ( .A(n1337), .B(n1335), .Z(n1319) );
  XNOR U1424 ( .A(n1336), .B(n1319), .Z(n1329) );
  NAND U1425 ( .A(a[52]), .B(b[0]), .Z(n1330) );
  XOR U1426 ( .A(n1332), .B(n1331), .Z(n1326) );
  XOR U1427 ( .A(n1325), .B(n1326), .Z(n1340) );
  XOR U1428 ( .A(n1339), .B(sreg[112]), .Z(n1322) );
  XNOR U1429 ( .A(n1340), .B(n1322), .Z(c[112]) );
  NANDN U1430 ( .A(n1324), .B(n1323), .Z(n1328) );
  NANDN U1431 ( .A(n1326), .B(n1325), .Z(n1327) );
  NAND U1432 ( .A(n1328), .B(n1327), .Z(n1342) );
  NANDN U1433 ( .A(n1330), .B(n1329), .Z(n1334) );
  NANDN U1434 ( .A(n1332), .B(n1331), .Z(n1333) );
  AND U1435 ( .A(n1334), .B(n1333), .Z(n1343) );
  XNOR U1436 ( .A(n1342), .B(n1343), .Z(n1344) );
  AND U1437 ( .A(a[52]), .B(b[1]), .Z(n1355) );
  NAND U1438 ( .A(b[2]), .B(a[51]), .Z(n1356) );
  NAND U1439 ( .A(b[3]), .B(a[50]), .Z(n1354) );
  XNOR U1440 ( .A(n1356), .B(n1354), .Z(n1338) );
  XNOR U1441 ( .A(n1355), .B(n1338), .Z(n1348) );
  NAND U1442 ( .A(a[53]), .B(b[0]), .Z(n1349) );
  XOR U1443 ( .A(n1351), .B(n1350), .Z(n1345) );
  XOR U1444 ( .A(n1344), .B(n1345), .Z(n1359) );
  XOR U1445 ( .A(n1358), .B(sreg[113]), .Z(n1341) );
  XNOR U1446 ( .A(n1359), .B(n1341), .Z(c[113]) );
  NANDN U1447 ( .A(n1343), .B(n1342), .Z(n1347) );
  NANDN U1448 ( .A(n1345), .B(n1344), .Z(n1346) );
  NAND U1449 ( .A(n1347), .B(n1346), .Z(n1361) );
  NANDN U1450 ( .A(n1349), .B(n1348), .Z(n1353) );
  NANDN U1451 ( .A(n1351), .B(n1350), .Z(n1352) );
  AND U1452 ( .A(n1353), .B(n1352), .Z(n1362) );
  XNOR U1453 ( .A(n1361), .B(n1362), .Z(n1363) );
  AND U1454 ( .A(a[53]), .B(b[1]), .Z(n1374) );
  NAND U1455 ( .A(b[2]), .B(a[52]), .Z(n1375) );
  NAND U1456 ( .A(b[3]), .B(a[51]), .Z(n1373) );
  XNOR U1457 ( .A(n1375), .B(n1373), .Z(n1357) );
  XNOR U1458 ( .A(n1374), .B(n1357), .Z(n1367) );
  NAND U1459 ( .A(a[54]), .B(b[0]), .Z(n1368) );
  XOR U1460 ( .A(n1370), .B(n1369), .Z(n1364) );
  XOR U1461 ( .A(n1363), .B(n1364), .Z(n1378) );
  XOR U1462 ( .A(n1377), .B(sreg[114]), .Z(n1360) );
  XNOR U1463 ( .A(n1378), .B(n1360), .Z(c[114]) );
  NANDN U1464 ( .A(n1362), .B(n1361), .Z(n1366) );
  NANDN U1465 ( .A(n1364), .B(n1363), .Z(n1365) );
  NAND U1466 ( .A(n1366), .B(n1365), .Z(n1380) );
  NANDN U1467 ( .A(n1368), .B(n1367), .Z(n1372) );
  NANDN U1468 ( .A(n1370), .B(n1369), .Z(n1371) );
  AND U1469 ( .A(n1372), .B(n1371), .Z(n1381) );
  XNOR U1470 ( .A(n1380), .B(n1381), .Z(n1382) );
  AND U1471 ( .A(a[54]), .B(b[1]), .Z(n1393) );
  NAND U1472 ( .A(b[2]), .B(a[53]), .Z(n1394) );
  NAND U1473 ( .A(b[3]), .B(a[52]), .Z(n1392) );
  XNOR U1474 ( .A(n1394), .B(n1392), .Z(n1376) );
  XNOR U1475 ( .A(n1393), .B(n1376), .Z(n1386) );
  NAND U1476 ( .A(a[55]), .B(b[0]), .Z(n1387) );
  XOR U1477 ( .A(n1389), .B(n1388), .Z(n1383) );
  XOR U1478 ( .A(n1382), .B(n1383), .Z(n1397) );
  XOR U1479 ( .A(n1396), .B(sreg[115]), .Z(n1379) );
  XNOR U1480 ( .A(n1397), .B(n1379), .Z(c[115]) );
  NANDN U1481 ( .A(n1381), .B(n1380), .Z(n1385) );
  NANDN U1482 ( .A(n1383), .B(n1382), .Z(n1384) );
  NAND U1483 ( .A(n1385), .B(n1384), .Z(n1399) );
  NANDN U1484 ( .A(n1387), .B(n1386), .Z(n1391) );
  NANDN U1485 ( .A(n1389), .B(n1388), .Z(n1390) );
  AND U1486 ( .A(n1391), .B(n1390), .Z(n1400) );
  XNOR U1487 ( .A(n1399), .B(n1400), .Z(n1401) );
  AND U1488 ( .A(a[55]), .B(b[1]), .Z(n1412) );
  NAND U1489 ( .A(b[2]), .B(a[54]), .Z(n1413) );
  NAND U1490 ( .A(b[3]), .B(a[53]), .Z(n1411) );
  XNOR U1491 ( .A(n1413), .B(n1411), .Z(n1395) );
  XNOR U1492 ( .A(n1412), .B(n1395), .Z(n1405) );
  NAND U1493 ( .A(a[56]), .B(b[0]), .Z(n1406) );
  XOR U1494 ( .A(n1408), .B(n1407), .Z(n1402) );
  XOR U1495 ( .A(n1401), .B(n1402), .Z(n1416) );
  XOR U1496 ( .A(n1415), .B(sreg[116]), .Z(n1398) );
  XNOR U1497 ( .A(n1416), .B(n1398), .Z(c[116]) );
  NANDN U1498 ( .A(n1400), .B(n1399), .Z(n1404) );
  NANDN U1499 ( .A(n1402), .B(n1401), .Z(n1403) );
  NAND U1500 ( .A(n1404), .B(n1403), .Z(n1418) );
  NANDN U1501 ( .A(n1406), .B(n1405), .Z(n1410) );
  NANDN U1502 ( .A(n1408), .B(n1407), .Z(n1409) );
  AND U1503 ( .A(n1410), .B(n1409), .Z(n1419) );
  XNOR U1504 ( .A(n1418), .B(n1419), .Z(n1420) );
  AND U1505 ( .A(a[56]), .B(b[1]), .Z(n1431) );
  NAND U1506 ( .A(b[2]), .B(a[55]), .Z(n1432) );
  NAND U1507 ( .A(b[3]), .B(a[54]), .Z(n1430) );
  XNOR U1508 ( .A(n1432), .B(n1430), .Z(n1414) );
  XNOR U1509 ( .A(n1431), .B(n1414), .Z(n1424) );
  NAND U1510 ( .A(a[57]), .B(b[0]), .Z(n1425) );
  XOR U1511 ( .A(n1427), .B(n1426), .Z(n1421) );
  XOR U1512 ( .A(n1420), .B(n1421), .Z(n1435) );
  XOR U1513 ( .A(n1434), .B(sreg[117]), .Z(n1417) );
  XNOR U1514 ( .A(n1435), .B(n1417), .Z(c[117]) );
  NANDN U1515 ( .A(n1419), .B(n1418), .Z(n1423) );
  NANDN U1516 ( .A(n1421), .B(n1420), .Z(n1422) );
  NAND U1517 ( .A(n1423), .B(n1422), .Z(n1437) );
  NANDN U1518 ( .A(n1425), .B(n1424), .Z(n1429) );
  NANDN U1519 ( .A(n1427), .B(n1426), .Z(n1428) );
  AND U1520 ( .A(n1429), .B(n1428), .Z(n1438) );
  XNOR U1521 ( .A(n1437), .B(n1438), .Z(n1439) );
  AND U1522 ( .A(a[57]), .B(b[1]), .Z(n1450) );
  NAND U1523 ( .A(b[2]), .B(a[56]), .Z(n1451) );
  NAND U1524 ( .A(b[3]), .B(a[55]), .Z(n1449) );
  XNOR U1525 ( .A(n1451), .B(n1449), .Z(n1433) );
  XNOR U1526 ( .A(n1450), .B(n1433), .Z(n1443) );
  NAND U1527 ( .A(a[58]), .B(b[0]), .Z(n1444) );
  XOR U1528 ( .A(n1446), .B(n1445), .Z(n1440) );
  XOR U1529 ( .A(n1439), .B(n1440), .Z(n1454) );
  XOR U1530 ( .A(n1453), .B(sreg[118]), .Z(n1436) );
  XNOR U1531 ( .A(n1454), .B(n1436), .Z(c[118]) );
  NANDN U1532 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U1533 ( .A(n1440), .B(n1439), .Z(n1441) );
  NAND U1534 ( .A(n1442), .B(n1441), .Z(n1456) );
  NANDN U1535 ( .A(n1444), .B(n1443), .Z(n1448) );
  NANDN U1536 ( .A(n1446), .B(n1445), .Z(n1447) );
  AND U1537 ( .A(n1448), .B(n1447), .Z(n1457) );
  XNOR U1538 ( .A(n1456), .B(n1457), .Z(n1458) );
  AND U1539 ( .A(a[58]), .B(b[1]), .Z(n1469) );
  NAND U1540 ( .A(b[2]), .B(a[57]), .Z(n1470) );
  NAND U1541 ( .A(b[3]), .B(a[56]), .Z(n1468) );
  XNOR U1542 ( .A(n1470), .B(n1468), .Z(n1452) );
  XNOR U1543 ( .A(n1469), .B(n1452), .Z(n1462) );
  NAND U1544 ( .A(a[59]), .B(b[0]), .Z(n1463) );
  XOR U1545 ( .A(n1465), .B(n1464), .Z(n1459) );
  XOR U1546 ( .A(n1458), .B(n1459), .Z(n1473) );
  XOR U1547 ( .A(n1472), .B(sreg[119]), .Z(n1455) );
  XNOR U1548 ( .A(n1473), .B(n1455), .Z(c[119]) );
  NANDN U1549 ( .A(n1457), .B(n1456), .Z(n1461) );
  NANDN U1550 ( .A(n1459), .B(n1458), .Z(n1460) );
  NAND U1551 ( .A(n1461), .B(n1460), .Z(n1475) );
  NANDN U1552 ( .A(n1463), .B(n1462), .Z(n1467) );
  NANDN U1553 ( .A(n1465), .B(n1464), .Z(n1466) );
  AND U1554 ( .A(n1467), .B(n1466), .Z(n1476) );
  XNOR U1555 ( .A(n1475), .B(n1476), .Z(n1477) );
  AND U1556 ( .A(a[59]), .B(b[1]), .Z(n1488) );
  NAND U1557 ( .A(b[2]), .B(a[58]), .Z(n1489) );
  NAND U1558 ( .A(b[3]), .B(a[57]), .Z(n1487) );
  XNOR U1559 ( .A(n1489), .B(n1487), .Z(n1471) );
  XNOR U1560 ( .A(n1488), .B(n1471), .Z(n1481) );
  NAND U1561 ( .A(a[60]), .B(b[0]), .Z(n1482) );
  XOR U1562 ( .A(n1484), .B(n1483), .Z(n1478) );
  XOR U1563 ( .A(n1477), .B(n1478), .Z(n1492) );
  XOR U1564 ( .A(n1491), .B(sreg[120]), .Z(n1474) );
  XNOR U1565 ( .A(n1492), .B(n1474), .Z(c[120]) );
  NANDN U1566 ( .A(n1476), .B(n1475), .Z(n1480) );
  NANDN U1567 ( .A(n1478), .B(n1477), .Z(n1479) );
  NAND U1568 ( .A(n1480), .B(n1479), .Z(n1494) );
  NANDN U1569 ( .A(n1482), .B(n1481), .Z(n1486) );
  NANDN U1570 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1571 ( .A(n1486), .B(n1485), .Z(n1495) );
  XNOR U1572 ( .A(n1494), .B(n1495), .Z(n1496) );
  AND U1573 ( .A(a[60]), .B(b[1]), .Z(n1507) );
  NAND U1574 ( .A(b[2]), .B(a[59]), .Z(n1508) );
  NAND U1575 ( .A(b[3]), .B(a[58]), .Z(n1506) );
  XNOR U1576 ( .A(n1508), .B(n1506), .Z(n1490) );
  XNOR U1577 ( .A(n1507), .B(n1490), .Z(n1500) );
  NAND U1578 ( .A(a[61]), .B(b[0]), .Z(n1501) );
  XOR U1579 ( .A(n1503), .B(n1502), .Z(n1497) );
  XOR U1580 ( .A(n1496), .B(n1497), .Z(n1511) );
  XOR U1581 ( .A(n1510), .B(sreg[121]), .Z(n1493) );
  XNOR U1582 ( .A(n1511), .B(n1493), .Z(c[121]) );
  NANDN U1583 ( .A(n1495), .B(n1494), .Z(n1499) );
  NANDN U1584 ( .A(n1497), .B(n1496), .Z(n1498) );
  NAND U1585 ( .A(n1499), .B(n1498), .Z(n1515) );
  NANDN U1586 ( .A(n1501), .B(n1500), .Z(n1505) );
  NANDN U1587 ( .A(n1503), .B(n1502), .Z(n1504) );
  AND U1588 ( .A(n1505), .B(n1504), .Z(n1516) );
  XNOR U1589 ( .A(n1515), .B(n1516), .Z(n1517) );
  AND U1590 ( .A(a[61]), .B(b[1]), .Z(n1529) );
  AND U1591 ( .A(a[60]), .B(b[2]), .Z(n1531) );
  AND U1592 ( .A(a[59]), .B(b[3]), .Z(n1528) );
  IV U1593 ( .A(n1528), .Z(n1527) );
  XOR U1594 ( .A(n1531), .B(n1527), .Z(n1509) );
  XNOR U1595 ( .A(n1529), .B(n1509), .Z(n1521) );
  NAND U1596 ( .A(a[62]), .B(b[0]), .Z(n1522) );
  XOR U1597 ( .A(n1524), .B(n1523), .Z(n1518) );
  XOR U1598 ( .A(n1517), .B(n1518), .Z(n1514) );
  XOR U1599 ( .A(n1513), .B(sreg[122]), .Z(n1512) );
  XNOR U1600 ( .A(n1514), .B(n1512), .Z(c[122]) );
  XNOR U1601 ( .A(n1548), .B(sreg[123]), .Z(n1550) );
  NANDN U1602 ( .A(n1516), .B(n1515), .Z(n1520) );
  NANDN U1603 ( .A(n1518), .B(n1517), .Z(n1519) );
  NAND U1604 ( .A(n1520), .B(n1519), .Z(n1539) );
  NANDN U1605 ( .A(n1522), .B(n1521), .Z(n1526) );
  NANDN U1606 ( .A(n1524), .B(n1523), .Z(n1525) );
  AND U1607 ( .A(n1526), .B(n1525), .Z(n1540) );
  XNOR U1608 ( .A(n1539), .B(n1540), .Z(n1541) );
  NANDN U1609 ( .A(n1529), .B(n1527), .Z(n1533) );
  AND U1610 ( .A(n1529), .B(n1528), .Z(n1530) );
  OR U1611 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U1612 ( .A(n1533), .B(n1532), .Z(n1538) );
  AND U1613 ( .A(a[61]), .B(b[2]), .Z(n1547) );
  ANDN U1614 ( .B(a[60]), .A(n367), .Z(n1546) );
  XNOR U1615 ( .A(n1545), .B(n1546), .Z(n1534) );
  XNOR U1616 ( .A(n1547), .B(n1534), .Z(n1537) );
  NAND U1617 ( .A(b[0]), .B(a[63]), .Z(n1536) );
  XOR U1618 ( .A(n1537), .B(n1536), .Z(n1535) );
  XOR U1619 ( .A(n1538), .B(n1535), .Z(n1542) );
  XNOR U1620 ( .A(n1541), .B(n1542), .Z(n1549) );
  XOR U1621 ( .A(n1550), .B(n1549), .Z(c[123]) );
  NANDN U1622 ( .A(n1540), .B(n1539), .Z(n1544) );
  NAND U1623 ( .A(n1542), .B(n1541), .Z(n1543) );
  AND U1624 ( .A(n1544), .B(n1543), .Z(n1556) );
  XOR U1625 ( .A(n1555), .B(n1556), .Z(n1558) );
  NAND U1626 ( .A(b[3]), .B(a[61]), .Z(n1566) );
  NAND U1627 ( .A(a[62]), .B(b[2]), .Z(n1573) );
  AND U1628 ( .A(a[63]), .B(b[1]), .Z(n1571) );
  XOR U1629 ( .A(n1573), .B(n1571), .Z(n1565) );
  XNOR U1630 ( .A(n1566), .B(n1565), .Z(n1568) );
  XOR U1631 ( .A(n1567), .B(n1568), .Z(n1557) );
  XOR U1632 ( .A(n1558), .B(n1557), .Z(n1553) );
  NAND U1633 ( .A(sreg[123]), .B(n1548), .Z(n1552) );
  OR U1634 ( .A(n1550), .B(n1549), .Z(n1551) );
  AND U1635 ( .A(n1552), .B(n1551), .Z(n1554) );
  XNOR U1636 ( .A(n1553), .B(n1554), .Z(c[124]) );
  NANDN U1637 ( .A(n1554), .B(n1553), .Z(n1581) );
  NANDN U1638 ( .A(n1556), .B(n1555), .Z(n1560) );
  OR U1639 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U1640 ( .A(n1560), .B(n1559), .Z(n1576) );
  ANDN U1641 ( .B(n1571), .A(n1573), .Z(n1564) );
  AND U1642 ( .A(a[62]), .B(b[3]), .Z(n1562) );
  AND U1643 ( .A(a[63]), .B(b[2]), .Z(n1561) );
  XNOR U1644 ( .A(n1562), .B(n1561), .Z(n1563) );
  XOR U1645 ( .A(n1564), .B(n1563), .Z(n1575) );
  OR U1646 ( .A(n1566), .B(n1565), .Z(n1570) );
  NANDN U1647 ( .A(n1568), .B(n1567), .Z(n1569) );
  AND U1648 ( .A(n1570), .B(n1569), .Z(n1574) );
  XNOR U1649 ( .A(n1575), .B(n1574), .Z(n1577) );
  XNOR U1650 ( .A(n1576), .B(n1577), .Z(n1580) );
  XOR U1651 ( .A(n1581), .B(n1580), .Z(c[125]) );
  ANDN U1652 ( .B(a[63]), .A(n367), .Z(n1586) );
  OR U1653 ( .A(n1586), .B(n1571), .Z(n1572) );
  NANDN U1654 ( .A(n1573), .B(n1572), .Z(n1584) );
  OR U1655 ( .A(n1575), .B(n1574), .Z(n1579) );
  OR U1656 ( .A(n1577), .B(n1576), .Z(n1578) );
  NAND U1657 ( .A(n1579), .B(n1578), .Z(n1587) );
  XOR U1658 ( .A(n1586), .B(n1587), .Z(n1582) );
  OR U1659 ( .A(n1581), .B(n1580), .Z(n1585) );
  XOR U1660 ( .A(n1582), .B(n1585), .Z(n1583) );
  XOR U1661 ( .A(n1584), .B(n1583), .Z(c[126]) );
endmodule

