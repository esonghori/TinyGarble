
module hamming_N16000_CC128 ( clk, rst, x, y, o );
  input [124:0] x;
  input [124:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[13]) );
  XOR U142 ( .A(n89), .B(n78), .Z(n124) );
  XOR U143 ( .A(n186), .B(n188), .Z(n194) );
  XOR U144 ( .A(n254), .B(n256), .Z(n262) );
  XNOR U145 ( .A(n156), .B(n223), .Z(n128) );
  XNOR U146 ( .A(oglobal[4]), .B(n63), .Z(n19) );
  XOR U147 ( .A(n370), .B(n369), .Z(n367) );
  XOR U148 ( .A(n326), .B(n325), .Z(n323) );
  XNOR U149 ( .A(n288), .B(n423), .Z(n260) );
  XNOR U150 ( .A(n55), .B(n75), .Z(n60) );
  XOR U151 ( .A(n192), .B(n194), .Z(n228) );
  XNOR U152 ( .A(oglobal[6]), .B(n36), .Z(n15) );
  XNOR U153 ( .A(oglobal[3]), .B(n94), .Z(n21) );
  XOR U154 ( .A(n412), .B(n411), .Z(n409) );
  XOR U155 ( .A(n458), .B(n457), .Z(n455) );
  XNOR U156 ( .A(n220), .B(n335), .Z(n192) );
  XNOR U157 ( .A(n39), .B(n51), .Z(n41) );
  XOR U158 ( .A(n122), .B(n123), .Z(n129) );
  XNOR U159 ( .A(n260), .B(n379), .Z(n226) );
  XNOR U160 ( .A(oglobal[5]), .B(n44), .Z(n17) );
  XNOR U161 ( .A(oglobal[2]), .B(n159), .Z(n23) );
  XOR U162 ( .A(n390), .B(n389), .Z(n408) );
  XOR U163 ( .A(n434), .B(n433), .Z(n454) );
  XOR U164 ( .A(n346), .B(n345), .Z(n366) );
  XOR U165 ( .A(n304), .B(n303), .Z(n322) );
  XOR U166 ( .A(n41), .B(n42), .Z(n18) );
  XOR U167 ( .A(n60), .B(n61), .Z(n20) );
  XOR U168 ( .A(n80), .B(n81), .Z(n22) );
  XOR U169 ( .A(n128), .B(n129), .Z(n24) );
  XOR U170 ( .A(n226), .B(n228), .Z(n26) );
  XNOR U171 ( .A(n15), .B(n16), .Z(o[6]) );
  XOR U172 ( .A(n17), .B(n18), .Z(o[5]) );
  XOR U173 ( .A(n19), .B(n20), .Z(o[4]) );
  XOR U174 ( .A(n21), .B(n22), .Z(o[3]) );
  XOR U175 ( .A(n23), .B(n24), .Z(o[2]) );
  XOR U176 ( .A(n25), .B(n26), .Z(o[1]) );
  XOR U177 ( .A(n27), .B(n28), .Z(o[13]) );
  XOR U178 ( .A(oglobal[13]), .B(n29), .Z(n28) );
  AND U179 ( .A(n27), .B(o[12]), .Z(n29) );
  XOR U180 ( .A(oglobal[12]), .B(n27), .Z(o[12]) );
  ANDN U181 ( .B(n30), .A(o[11]), .Z(n27) );
  XOR U182 ( .A(oglobal[11]), .B(n30), .Z(o[11]) );
  ANDN U183 ( .B(n31), .A(o[10]), .Z(n30) );
  XOR U184 ( .A(oglobal[10]), .B(n31), .Z(o[10]) );
  ANDN U185 ( .B(n32), .A(o[9]), .Z(n31) );
  XOR U186 ( .A(oglobal[9]), .B(n32), .Z(o[9]) );
  ANDN U187 ( .B(n33), .A(o[8]), .Z(n32) );
  XOR U188 ( .A(oglobal[8]), .B(n33), .Z(o[8]) );
  ANDN U189 ( .B(n34), .A(o[7]), .Z(n33) );
  XOR U190 ( .A(oglobal[7]), .B(n34), .Z(o[7]) );
  XOR U191 ( .A(n35), .B(n36), .Z(n34) );
  ANDN U192 ( .B(n37), .A(n15), .Z(n35) );
  XOR U193 ( .A(n36), .B(n16), .Z(n37) );
  XOR U194 ( .A(n38), .B(n39), .Z(n16) );
  AND U195 ( .A(n40), .B(n41), .Z(n38) );
  XNOR U196 ( .A(n39), .B(n42), .Z(n40) );
  XOR U197 ( .A(n43), .B(n44), .Z(n36) );
  ANDN U198 ( .B(n45), .A(n17), .Z(n43) );
  XNOR U199 ( .A(n44), .B(n18), .Z(n45) );
  XNOR U200 ( .A(n46), .B(n47), .Z(n42) );
  ANDN U201 ( .B(n48), .A(n49), .Z(n46) );
  XNOR U202 ( .A(n50), .B(n47), .Z(n48) );
  XNOR U203 ( .A(n52), .B(n53), .Z(n51) );
  AND U204 ( .A(n54), .B(n55), .Z(n52) );
  XNOR U205 ( .A(n56), .B(n53), .Z(n54) );
  XOR U206 ( .A(n57), .B(n58), .Z(n39) );
  AND U207 ( .A(n59), .B(n60), .Z(n57) );
  XNOR U208 ( .A(n58), .B(n61), .Z(n59) );
  XOR U209 ( .A(n62), .B(n63), .Z(n44) );
  ANDN U210 ( .B(n64), .A(n19), .Z(n62) );
  XNOR U211 ( .A(n63), .B(n20), .Z(n64) );
  XNOR U212 ( .A(n50), .B(n49), .Z(n61) );
  XNOR U213 ( .A(n65), .B(n47), .Z(n49) );
  XNOR U214 ( .A(n66), .B(n67), .Z(n47) );
  AND U215 ( .A(n68), .B(n69), .Z(n66) );
  XOR U216 ( .A(n67), .B(n70), .Z(n69) );
  NOR U217 ( .A(n71), .B(n72), .Z(n65) );
  OR U218 ( .A(n73), .B(n74), .Z(n50) );
  XNOR U219 ( .A(n56), .B(n76), .Z(n75) );
  IV U220 ( .A(n58), .Z(n76) );
  XOR U221 ( .A(n77), .B(n78), .Z(n58) );
  AND U222 ( .A(n79), .B(n80), .Z(n77) );
  XNOR U223 ( .A(n78), .B(n81), .Z(n79) );
  OR U224 ( .A(n82), .B(n83), .Z(n56) );
  XOR U225 ( .A(n84), .B(n53), .Z(n55) );
  XOR U226 ( .A(n85), .B(n86), .Z(n53) );
  AND U227 ( .A(n87), .B(n88), .Z(n85) );
  XNOR U228 ( .A(n89), .B(n90), .Z(n88) );
  IV U229 ( .A(n86), .Z(n90) );
  NOR U230 ( .A(n91), .B(n92), .Z(n84) );
  XOR U231 ( .A(n93), .B(n94), .Z(n63) );
  ANDN U232 ( .B(n95), .A(n21), .Z(n93) );
  XNOR U233 ( .A(n94), .B(n22), .Z(n95) );
  XOR U234 ( .A(n68), .B(n70), .Z(n81) );
  XNOR U235 ( .A(n73), .B(n74), .Z(n70) );
  AND U236 ( .A(n96), .B(n97), .Z(n74) );
  OR U237 ( .A(n98), .B(n99), .Z(n97) );
  XOR U238 ( .A(n100), .B(n101), .Z(n96) );
  AND U239 ( .A(n102), .B(n103), .Z(n100) );
  XOR U240 ( .A(n101), .B(n104), .Z(n103) );
  OR U241 ( .A(n105), .B(n106), .Z(n73) );
  XNOR U242 ( .A(n67), .B(n107), .Z(n68) );
  XOR U243 ( .A(n71), .B(n72), .Z(n107) );
  AND U244 ( .A(n108), .B(n109), .Z(n72) );
  OR U245 ( .A(n110), .B(n111), .Z(n109) );
  XOR U246 ( .A(n112), .B(n113), .Z(n108) );
  AND U247 ( .A(n114), .B(n115), .Z(n112) );
  XNOR U248 ( .A(n116), .B(n113), .Z(n115) );
  OR U249 ( .A(n117), .B(n118), .Z(n71) );
  XOR U250 ( .A(n119), .B(n120), .Z(n67) );
  AND U251 ( .A(n121), .B(n122), .Z(n119) );
  XOR U252 ( .A(n120), .B(n123), .Z(n121) );
  XOR U253 ( .A(n87), .B(n124), .Z(n80) );
  XNOR U254 ( .A(n125), .B(n126), .Z(n78) );
  AND U255 ( .A(n127), .B(n128), .Z(n125) );
  XOR U256 ( .A(n126), .B(n129), .Z(n127) );
  XOR U257 ( .A(n82), .B(n83), .Z(n89) );
  AND U258 ( .A(n130), .B(n131), .Z(n83) );
  OR U259 ( .A(n132), .B(n133), .Z(n131) );
  XOR U260 ( .A(n134), .B(n135), .Z(n130) );
  ANDN U261 ( .B(n136), .A(n137), .Z(n134) );
  XOR U262 ( .A(n135), .B(n138), .Z(n136) );
  OR U263 ( .A(n139), .B(n140), .Z(n82) );
  XOR U264 ( .A(n86), .B(n141), .Z(n87) );
  XOR U265 ( .A(n91), .B(n92), .Z(n141) );
  AND U266 ( .A(n142), .B(n143), .Z(n92) );
  OR U267 ( .A(n144), .B(n145), .Z(n143) );
  XOR U268 ( .A(n146), .B(n147), .Z(n142) );
  AND U269 ( .A(n148), .B(n149), .Z(n146) );
  XNOR U270 ( .A(n150), .B(n147), .Z(n149) );
  OR U271 ( .A(n151), .B(n152), .Z(n91) );
  XNOR U272 ( .A(n153), .B(n154), .Z(n86) );
  AND U273 ( .A(n155), .B(n156), .Z(n153) );
  XOR U274 ( .A(n157), .B(n154), .Z(n155) );
  XOR U275 ( .A(n158), .B(n159), .Z(n94) );
  ANDN U276 ( .B(n160), .A(n23), .Z(n158) );
  XNOR U277 ( .A(n159), .B(n24), .Z(n160) );
  XOR U278 ( .A(n102), .B(n104), .Z(n123) );
  XNOR U279 ( .A(n105), .B(n106), .Z(n104) );
  AND U280 ( .A(n161), .B(n162), .Z(n106) );
  OR U281 ( .A(n163), .B(n164), .Z(n162) );
  XOR U282 ( .A(n165), .B(n166), .Z(n161) );
  NAND U283 ( .A(n167), .B(n168), .Z(n166) );
  XNOR U284 ( .A(n165), .B(n169), .Z(n167) );
  OR U285 ( .A(n170), .B(n171), .Z(n105) );
  XNOR U286 ( .A(n101), .B(n172), .Z(n102) );
  XOR U287 ( .A(n98), .B(n99), .Z(n172) );
  AND U288 ( .A(n173), .B(n174), .Z(n99) );
  OR U289 ( .A(n175), .B(n176), .Z(n174) );
  XOR U290 ( .A(n177), .B(n178), .Z(n173) );
  NAND U291 ( .A(n179), .B(n180), .Z(n178) );
  XNOR U292 ( .A(n177), .B(n181), .Z(n179) );
  OR U293 ( .A(n182), .B(n183), .Z(n98) );
  XNOR U294 ( .A(n184), .B(n185), .Z(n101) );
  NAND U295 ( .A(n186), .B(n187), .Z(n185) );
  XOR U296 ( .A(n184), .B(n188), .Z(n187) );
  XOR U297 ( .A(n114), .B(n189), .Z(n122) );
  XNOR U298 ( .A(n116), .B(n120), .Z(n189) );
  XNOR U299 ( .A(n190), .B(n191), .Z(n120) );
  NAND U300 ( .A(n192), .B(n193), .Z(n191) );
  XOR U301 ( .A(n190), .B(n194), .Z(n193) );
  XOR U302 ( .A(n117), .B(n118), .Z(n116) );
  AND U303 ( .A(n195), .B(n196), .Z(n118) );
  OR U304 ( .A(n197), .B(n198), .Z(n196) );
  XOR U305 ( .A(n199), .B(n200), .Z(n195) );
  NAND U306 ( .A(n201), .B(n202), .Z(n200) );
  XNOR U307 ( .A(n199), .B(n203), .Z(n201) );
  OR U308 ( .A(n204), .B(n205), .Z(n117) );
  XNOR U309 ( .A(n113), .B(n206), .Z(n114) );
  XOR U310 ( .A(n110), .B(n111), .Z(n206) );
  AND U311 ( .A(n207), .B(n208), .Z(n111) );
  OR U312 ( .A(n209), .B(n210), .Z(n208) );
  XOR U313 ( .A(n211), .B(n212), .Z(n207) );
  NAND U314 ( .A(n213), .B(n214), .Z(n212) );
  XNOR U315 ( .A(n211), .B(n215), .Z(n213) );
  OR U316 ( .A(n216), .B(n217), .Z(n110) );
  XNOR U317 ( .A(n218), .B(n219), .Z(n113) );
  NAND U318 ( .A(n220), .B(n221), .Z(n219) );
  XOR U319 ( .A(n218), .B(n222), .Z(n221) );
  XNOR U320 ( .A(n157), .B(n126), .Z(n223) );
  XNOR U321 ( .A(n224), .B(n225), .Z(n126) );
  NAND U322 ( .A(n226), .B(n227), .Z(n225) );
  XOR U323 ( .A(n224), .B(n228), .Z(n227) );
  XNOR U324 ( .A(n137), .B(n138), .Z(n157) );
  XNOR U325 ( .A(n139), .B(n140), .Z(n138) );
  AND U326 ( .A(n229), .B(n230), .Z(n140) );
  OR U327 ( .A(n231), .B(n232), .Z(n230) );
  XOR U328 ( .A(n233), .B(n234), .Z(n229) );
  NAND U329 ( .A(n235), .B(n236), .Z(n234) );
  XNOR U330 ( .A(n233), .B(n237), .Z(n235) );
  OR U331 ( .A(n238), .B(n239), .Z(n139) );
  XOR U332 ( .A(n135), .B(n240), .Z(n137) );
  XOR U333 ( .A(n132), .B(n133), .Z(n240) );
  AND U334 ( .A(n241), .B(n242), .Z(n133) );
  OR U335 ( .A(n243), .B(n244), .Z(n242) );
  XOR U336 ( .A(n245), .B(n246), .Z(n241) );
  NAND U337 ( .A(n247), .B(n248), .Z(n246) );
  XNOR U338 ( .A(n245), .B(n249), .Z(n247) );
  OR U339 ( .A(n250), .B(n251), .Z(n132) );
  XNOR U340 ( .A(n252), .B(n253), .Z(n135) );
  NAND U341 ( .A(n254), .B(n255), .Z(n253) );
  XOR U342 ( .A(n252), .B(n256), .Z(n255) );
  XOR U343 ( .A(n148), .B(n257), .Z(n156) );
  XNOR U344 ( .A(n150), .B(n154), .Z(n257) );
  XNOR U345 ( .A(n258), .B(n259), .Z(n154) );
  NAND U346 ( .A(n260), .B(n261), .Z(n259) );
  XOR U347 ( .A(n258), .B(n262), .Z(n261) );
  XOR U348 ( .A(n151), .B(n152), .Z(n150) );
  AND U349 ( .A(n263), .B(n264), .Z(n152) );
  OR U350 ( .A(n265), .B(n266), .Z(n264) );
  XOR U351 ( .A(n267), .B(n268), .Z(n263) );
  NAND U352 ( .A(n269), .B(n270), .Z(n268) );
  XNOR U353 ( .A(n267), .B(n271), .Z(n269) );
  OR U354 ( .A(n272), .B(n273), .Z(n151) );
  XNOR U355 ( .A(n147), .B(n274), .Z(n148) );
  XOR U356 ( .A(n144), .B(n145), .Z(n274) );
  AND U357 ( .A(n275), .B(n276), .Z(n145) );
  OR U358 ( .A(n277), .B(n278), .Z(n276) );
  XOR U359 ( .A(n279), .B(n280), .Z(n275) );
  NAND U360 ( .A(n281), .B(n282), .Z(n280) );
  XNOR U361 ( .A(n279), .B(n283), .Z(n281) );
  OR U362 ( .A(n284), .B(n285), .Z(n144) );
  XNOR U363 ( .A(n286), .B(n287), .Z(n147) );
  NAND U364 ( .A(n288), .B(n289), .Z(n287) );
  XOR U365 ( .A(n286), .B(n290), .Z(n289) );
  XNOR U366 ( .A(n291), .B(n292), .Z(n159) );
  NANDN U367 ( .A(n25), .B(n293), .Z(n292) );
  XNOR U368 ( .A(n291), .B(n26), .Z(n293) );
  XOR U369 ( .A(n168), .B(n169), .Z(n188) );
  XNOR U370 ( .A(n170), .B(n171), .Z(n169) );
  AND U371 ( .A(n294), .B(n295), .Z(n171) );
  OR U372 ( .A(n296), .B(n297), .Z(n295) );
  OR U373 ( .A(n298), .B(n299), .Z(n294) );
  OR U374 ( .A(n300), .B(n301), .Z(n170) );
  XOR U375 ( .A(n164), .B(n302), .Z(n168) );
  XOR U376 ( .A(n163), .B(n165), .Z(n302) );
  ANDN U377 ( .B(n303), .A(n304), .Z(n165) );
  OR U378 ( .A(n305), .B(n306), .Z(n163) );
  AND U379 ( .A(n307), .B(n308), .Z(n164) );
  OR U380 ( .A(n309), .B(n310), .Z(n308) );
  OR U381 ( .A(n311), .B(n312), .Z(n307) );
  XOR U382 ( .A(n180), .B(n313), .Z(n186) );
  XOR U383 ( .A(n184), .B(n181), .Z(n313) );
  XNOR U384 ( .A(n182), .B(n183), .Z(n181) );
  AND U385 ( .A(n314), .B(n315), .Z(n183) );
  OR U386 ( .A(n316), .B(n317), .Z(n315) );
  OR U387 ( .A(n318), .B(n319), .Z(n314) );
  OR U388 ( .A(n320), .B(n321), .Z(n182) );
  OR U389 ( .A(n322), .B(n323), .Z(n184) );
  XOR U390 ( .A(n176), .B(n324), .Z(n180) );
  XOR U391 ( .A(n175), .B(n177), .Z(n324) );
  ANDN U392 ( .B(n325), .A(n326), .Z(n177) );
  OR U393 ( .A(n327), .B(n328), .Z(n175) );
  AND U394 ( .A(n329), .B(n330), .Z(n176) );
  OR U395 ( .A(n331), .B(n332), .Z(n330) );
  OR U396 ( .A(n333), .B(n334), .Z(n329) );
  XNOR U397 ( .A(n190), .B(n222), .Z(n335) );
  XOR U398 ( .A(n202), .B(n203), .Z(n222) );
  XNOR U399 ( .A(n204), .B(n205), .Z(n203) );
  AND U400 ( .A(n336), .B(n337), .Z(n205) );
  OR U401 ( .A(n338), .B(n339), .Z(n337) );
  OR U402 ( .A(n340), .B(n341), .Z(n336) );
  OR U403 ( .A(n342), .B(n343), .Z(n204) );
  XOR U404 ( .A(n198), .B(n344), .Z(n202) );
  XOR U405 ( .A(n197), .B(n199), .Z(n344) );
  ANDN U406 ( .B(n345), .A(n346), .Z(n199) );
  OR U407 ( .A(n347), .B(n348), .Z(n197) );
  AND U408 ( .A(n349), .B(n350), .Z(n198) );
  OR U409 ( .A(n351), .B(n352), .Z(n350) );
  OR U410 ( .A(n353), .B(n354), .Z(n349) );
  OR U411 ( .A(n355), .B(n356), .Z(n190) );
  XOR U412 ( .A(n214), .B(n357), .Z(n220) );
  XOR U413 ( .A(n218), .B(n215), .Z(n357) );
  XNOR U414 ( .A(n216), .B(n217), .Z(n215) );
  AND U415 ( .A(n358), .B(n359), .Z(n217) );
  OR U416 ( .A(n360), .B(n361), .Z(n359) );
  OR U417 ( .A(n362), .B(n363), .Z(n358) );
  OR U418 ( .A(n364), .B(n365), .Z(n216) );
  OR U419 ( .A(n366), .B(n367), .Z(n218) );
  XOR U420 ( .A(n210), .B(n368), .Z(n214) );
  XOR U421 ( .A(n209), .B(n211), .Z(n368) );
  ANDN U422 ( .B(n369), .A(n370), .Z(n211) );
  OR U423 ( .A(n371), .B(n372), .Z(n209) );
  AND U424 ( .A(n373), .B(n374), .Z(n210) );
  OR U425 ( .A(n375), .B(n376), .Z(n374) );
  OR U426 ( .A(n377), .B(n378), .Z(n373) );
  XNOR U427 ( .A(n224), .B(n262), .Z(n379) );
  XOR U428 ( .A(n236), .B(n237), .Z(n256) );
  XNOR U429 ( .A(n238), .B(n239), .Z(n237) );
  AND U430 ( .A(n380), .B(n381), .Z(n239) );
  OR U431 ( .A(n382), .B(n383), .Z(n381) );
  OR U432 ( .A(n384), .B(n385), .Z(n380) );
  OR U433 ( .A(n386), .B(n387), .Z(n238) );
  XOR U434 ( .A(n232), .B(n388), .Z(n236) );
  XOR U435 ( .A(n231), .B(n233), .Z(n388) );
  ANDN U436 ( .B(n389), .A(n390), .Z(n233) );
  OR U437 ( .A(n391), .B(n392), .Z(n231) );
  AND U438 ( .A(n393), .B(n394), .Z(n232) );
  OR U439 ( .A(n395), .B(n396), .Z(n394) );
  OR U440 ( .A(n397), .B(n398), .Z(n393) );
  XOR U441 ( .A(n248), .B(n399), .Z(n254) );
  XOR U442 ( .A(n252), .B(n249), .Z(n399) );
  XNOR U443 ( .A(n250), .B(n251), .Z(n249) );
  AND U444 ( .A(n400), .B(n401), .Z(n251) );
  OR U445 ( .A(n402), .B(n403), .Z(n401) );
  OR U446 ( .A(n404), .B(n405), .Z(n400) );
  OR U447 ( .A(n406), .B(n407), .Z(n250) );
  OR U448 ( .A(n408), .B(n409), .Z(n252) );
  XOR U449 ( .A(n244), .B(n410), .Z(n248) );
  XOR U450 ( .A(n243), .B(n245), .Z(n410) );
  ANDN U451 ( .B(n411), .A(n412), .Z(n245) );
  OR U452 ( .A(n413), .B(n414), .Z(n243) );
  AND U453 ( .A(n415), .B(n416), .Z(n244) );
  OR U454 ( .A(n417), .B(n418), .Z(n416) );
  OR U455 ( .A(n419), .B(n420), .Z(n415) );
  OR U456 ( .A(n421), .B(n422), .Z(n224) );
  XNOR U457 ( .A(n258), .B(n290), .Z(n423) );
  XOR U458 ( .A(n270), .B(n271), .Z(n290) );
  XNOR U459 ( .A(n272), .B(n273), .Z(n271) );
  AND U460 ( .A(n424), .B(n425), .Z(n273) );
  OR U461 ( .A(n426), .B(n427), .Z(n425) );
  OR U462 ( .A(n428), .B(n429), .Z(n424) );
  OR U463 ( .A(n430), .B(n431), .Z(n272) );
  XOR U464 ( .A(n266), .B(n432), .Z(n270) );
  XOR U465 ( .A(n265), .B(n267), .Z(n432) );
  ANDN U466 ( .B(n433), .A(n434), .Z(n267) );
  OR U467 ( .A(n435), .B(n436), .Z(n265) );
  AND U468 ( .A(n437), .B(n438), .Z(n266) );
  OR U469 ( .A(n439), .B(n440), .Z(n438) );
  OR U470 ( .A(n441), .B(n442), .Z(n437) );
  OR U471 ( .A(n443), .B(n444), .Z(n258) );
  XOR U472 ( .A(n282), .B(n445), .Z(n288) );
  XOR U473 ( .A(n286), .B(n283), .Z(n445) );
  XNOR U474 ( .A(n284), .B(n285), .Z(n283) );
  AND U475 ( .A(n446), .B(n447), .Z(n285) );
  OR U476 ( .A(n448), .B(n449), .Z(n447) );
  OR U477 ( .A(n450), .B(n451), .Z(n446) );
  OR U478 ( .A(n452), .B(n453), .Z(n284) );
  OR U479 ( .A(n454), .B(n455), .Z(n286) );
  XOR U480 ( .A(n278), .B(n456), .Z(n282) );
  XOR U481 ( .A(n277), .B(n279), .Z(n456) );
  ANDN U482 ( .B(n457), .A(n458), .Z(n279) );
  OR U483 ( .A(n459), .B(n460), .Z(n277) );
  AND U484 ( .A(n461), .B(n462), .Z(n278) );
  OR U485 ( .A(n463), .B(n464), .Z(n462) );
  OR U486 ( .A(n465), .B(n466), .Z(n461) );
  XNOR U487 ( .A(oglobal[1]), .B(n291), .Z(n25) );
  ANDN U488 ( .B(oglobal[0]), .A(n467), .Z(n291) );
  XNOR U489 ( .A(oglobal[0]), .B(n467), .Z(o[0]) );
  XNOR U490 ( .A(n422), .B(n421), .Z(n467) );
  XNOR U491 ( .A(n356), .B(n355), .Z(n421) );
  XNOR U492 ( .A(n323), .B(n322), .Z(n355) );
  XOR U493 ( .A(n298), .B(n299), .Z(n303) );
  XNOR U494 ( .A(n301), .B(n300), .Z(n299) );
  XNOR U495 ( .A(y[63]), .B(x[63]), .Z(n300) );
  XNOR U496 ( .A(y[62]), .B(x[62]), .Z(n301) );
  XNOR U497 ( .A(n296), .B(n297), .Z(n298) );
  XNOR U498 ( .A(y[61]), .B(x[61]), .Z(n297) );
  XNOR U499 ( .A(y[60]), .B(x[60]), .Z(n296) );
  XNOR U500 ( .A(n311), .B(n312), .Z(n304) );
  XNOR U501 ( .A(n306), .B(n305), .Z(n312) );
  XNOR U502 ( .A(y[59]), .B(x[59]), .Z(n305) );
  XNOR U503 ( .A(y[58]), .B(x[58]), .Z(n306) );
  XNOR U504 ( .A(n309), .B(n310), .Z(n311) );
  XNOR U505 ( .A(y[57]), .B(x[57]), .Z(n310) );
  XNOR U506 ( .A(y[56]), .B(x[56]), .Z(n309) );
  XOR U507 ( .A(n318), .B(n319), .Z(n325) );
  XNOR U508 ( .A(n321), .B(n320), .Z(n319) );
  XNOR U509 ( .A(y[55]), .B(x[55]), .Z(n320) );
  XNOR U510 ( .A(y[54]), .B(x[54]), .Z(n321) );
  XNOR U511 ( .A(n316), .B(n317), .Z(n318) );
  XNOR U512 ( .A(y[53]), .B(x[53]), .Z(n317) );
  XNOR U513 ( .A(y[52]), .B(x[52]), .Z(n316) );
  XNOR U514 ( .A(n333), .B(n334), .Z(n326) );
  XNOR U515 ( .A(n328), .B(n327), .Z(n334) );
  XNOR U516 ( .A(y[51]), .B(x[51]), .Z(n327) );
  XNOR U517 ( .A(y[50]), .B(x[50]), .Z(n328) );
  XNOR U518 ( .A(n331), .B(n332), .Z(n333) );
  XNOR U519 ( .A(y[49]), .B(x[49]), .Z(n332) );
  XNOR U520 ( .A(y[48]), .B(x[48]), .Z(n331) );
  XNOR U521 ( .A(n367), .B(n366), .Z(n356) );
  XOR U522 ( .A(n340), .B(n341), .Z(n345) );
  XNOR U523 ( .A(n343), .B(n342), .Z(n341) );
  XNOR U524 ( .A(y[47]), .B(x[47]), .Z(n342) );
  XNOR U525 ( .A(y[46]), .B(x[46]), .Z(n343) );
  XNOR U526 ( .A(n338), .B(n339), .Z(n340) );
  XNOR U527 ( .A(y[45]), .B(x[45]), .Z(n339) );
  XNOR U528 ( .A(y[44]), .B(x[44]), .Z(n338) );
  XNOR U529 ( .A(n353), .B(n354), .Z(n346) );
  XNOR U530 ( .A(n348), .B(n347), .Z(n354) );
  XNOR U531 ( .A(y[43]), .B(x[43]), .Z(n347) );
  XNOR U532 ( .A(y[42]), .B(x[42]), .Z(n348) );
  XNOR U533 ( .A(n351), .B(n352), .Z(n353) );
  XNOR U534 ( .A(y[41]), .B(x[41]), .Z(n352) );
  XNOR U535 ( .A(y[40]), .B(x[40]), .Z(n351) );
  XOR U536 ( .A(n362), .B(n363), .Z(n369) );
  XNOR U537 ( .A(n365), .B(n364), .Z(n363) );
  XNOR U538 ( .A(y[39]), .B(x[39]), .Z(n364) );
  XNOR U539 ( .A(y[38]), .B(x[38]), .Z(n365) );
  XNOR U540 ( .A(n360), .B(n361), .Z(n362) );
  XNOR U541 ( .A(y[37]), .B(x[37]), .Z(n361) );
  XNOR U542 ( .A(y[36]), .B(x[36]), .Z(n360) );
  XNOR U543 ( .A(n377), .B(n378), .Z(n370) );
  XNOR U544 ( .A(n372), .B(n371), .Z(n378) );
  XNOR U545 ( .A(y[35]), .B(x[35]), .Z(n371) );
  XNOR U546 ( .A(y[34]), .B(x[34]), .Z(n372) );
  XNOR U547 ( .A(n375), .B(n376), .Z(n377) );
  XNOR U548 ( .A(y[33]), .B(x[33]), .Z(n376) );
  XNOR U549 ( .A(y[32]), .B(x[32]), .Z(n375) );
  XNOR U550 ( .A(n444), .B(n443), .Z(n422) );
  XNOR U551 ( .A(n409), .B(n408), .Z(n443) );
  XOR U552 ( .A(n384), .B(n385), .Z(n389) );
  XNOR U553 ( .A(n387), .B(n386), .Z(n385) );
  XNOR U554 ( .A(y[31]), .B(x[31]), .Z(n386) );
  XNOR U555 ( .A(y[30]), .B(x[30]), .Z(n387) );
  XNOR U556 ( .A(n382), .B(n383), .Z(n384) );
  XNOR U557 ( .A(y[29]), .B(x[29]), .Z(n383) );
  XNOR U558 ( .A(y[28]), .B(x[28]), .Z(n382) );
  XNOR U559 ( .A(n397), .B(n398), .Z(n390) );
  XNOR U560 ( .A(n392), .B(n391), .Z(n398) );
  XNOR U561 ( .A(y[27]), .B(x[27]), .Z(n391) );
  XNOR U562 ( .A(y[26]), .B(x[26]), .Z(n392) );
  XNOR U563 ( .A(n395), .B(n396), .Z(n397) );
  XNOR U564 ( .A(y[25]), .B(x[25]), .Z(n396) );
  XNOR U565 ( .A(y[24]), .B(x[24]), .Z(n395) );
  XOR U566 ( .A(n404), .B(n405), .Z(n411) );
  XNOR U567 ( .A(n407), .B(n406), .Z(n405) );
  XNOR U568 ( .A(y[23]), .B(x[23]), .Z(n406) );
  XNOR U569 ( .A(y[22]), .B(x[22]), .Z(n407) );
  XNOR U570 ( .A(n402), .B(n403), .Z(n404) );
  XNOR U571 ( .A(y[21]), .B(x[21]), .Z(n403) );
  XNOR U572 ( .A(y[20]), .B(x[20]), .Z(n402) );
  XNOR U573 ( .A(n419), .B(n420), .Z(n412) );
  XNOR U574 ( .A(n414), .B(n413), .Z(n420) );
  XNOR U575 ( .A(y[19]), .B(x[19]), .Z(n413) );
  XNOR U576 ( .A(y[18]), .B(x[18]), .Z(n414) );
  XNOR U577 ( .A(n417), .B(n418), .Z(n419) );
  XNOR U578 ( .A(y[17]), .B(x[17]), .Z(n418) );
  XNOR U579 ( .A(y[16]), .B(x[16]), .Z(n417) );
  XNOR U580 ( .A(n455), .B(n454), .Z(n444) );
  XOR U581 ( .A(n428), .B(n429), .Z(n433) );
  XNOR U582 ( .A(n431), .B(n430), .Z(n429) );
  XNOR U583 ( .A(y[15]), .B(x[15]), .Z(n430) );
  XNOR U584 ( .A(y[14]), .B(x[14]), .Z(n431) );
  XNOR U585 ( .A(n426), .B(n427), .Z(n428) );
  XNOR U586 ( .A(y[13]), .B(x[13]), .Z(n427) );
  XNOR U587 ( .A(y[12]), .B(x[12]), .Z(n426) );
  XNOR U588 ( .A(n441), .B(n442), .Z(n434) );
  XNOR U589 ( .A(n436), .B(n435), .Z(n442) );
  XNOR U590 ( .A(y[11]), .B(x[11]), .Z(n435) );
  XNOR U591 ( .A(y[10]), .B(x[10]), .Z(n436) );
  XNOR U592 ( .A(n439), .B(n440), .Z(n441) );
  XNOR U593 ( .A(y[9]), .B(x[9]), .Z(n440) );
  XNOR U594 ( .A(y[8]), .B(x[8]), .Z(n439) );
  XOR U595 ( .A(n450), .B(n451), .Z(n457) );
  XNOR U596 ( .A(n453), .B(n452), .Z(n451) );
  XNOR U597 ( .A(y[7]), .B(x[7]), .Z(n452) );
  XNOR U598 ( .A(y[6]), .B(x[6]), .Z(n453) );
  XNOR U599 ( .A(n448), .B(n449), .Z(n450) );
  XNOR U600 ( .A(y[5]), .B(x[5]), .Z(n449) );
  XNOR U601 ( .A(y[4]), .B(x[4]), .Z(n448) );
  XNOR U602 ( .A(n465), .B(n466), .Z(n458) );
  XNOR U603 ( .A(n460), .B(n459), .Z(n466) );
  XNOR U604 ( .A(y[3]), .B(x[3]), .Z(n459) );
  XNOR U605 ( .A(y[2]), .B(x[2]), .Z(n460) );
  XNOR U606 ( .A(n463), .B(n464), .Z(n465) );
  XNOR U607 ( .A(y[1]), .B(x[1]), .Z(n464) );
  XNOR U608 ( .A(y[0]), .B(x[0]), .Z(n463) );
endmodule

