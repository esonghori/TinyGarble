
module knns_seq_W32_K4 ( clk, rst, g_input, e_input, o );
  input [63:0] g_input;
  input [63:0] e_input;
  output [255:0] o;
  input clk, rst;
  wire   \min_dist_reg[3][33] , \min_dist_reg[3][32] , \min_dist_reg[3][31] ,
         \min_dist_reg[3][30] , \min_dist_reg[3][29] , \min_dist_reg[3][28] ,
         \min_dist_reg[3][27] , \min_dist_reg[3][26] , \min_dist_reg[3][25] ,
         \min_dist_reg[3][24] , \min_dist_reg[3][23] , \min_dist_reg[3][22] ,
         \min_dist_reg[3][21] , \min_dist_reg[3][20] , \min_dist_reg[3][19] ,
         \min_dist_reg[3][18] , \min_dist_reg[3][17] , \min_dist_reg[3][16] ,
         \min_dist_reg[3][15] , \min_dist_reg[3][14] , \min_dist_reg[3][13] ,
         \min_dist_reg[3][12] , \min_dist_reg[3][11] , \min_dist_reg[3][10] ,
         \min_dist_reg[3][9] , \min_dist_reg[3][8] , \min_dist_reg[3][7] ,
         \min_dist_reg[3][6] , \min_dist_reg[3][5] , \min_dist_reg[3][4] ,
         \min_dist_reg[3][3] , \min_dist_reg[3][2] , \min_dist_reg[3][1] ,
         \min_dist_reg[3][0] , \min_dist_reg[2][33] , \min_dist_reg[2][32] ,
         \min_dist_reg[2][31] , \min_dist_reg[2][30] , \min_dist_reg[2][29] ,
         \min_dist_reg[2][28] , \min_dist_reg[2][27] , \min_dist_reg[2][26] ,
         \min_dist_reg[2][25] , \min_dist_reg[2][24] , \min_dist_reg[2][23] ,
         \min_dist_reg[2][22] , \min_dist_reg[2][21] , \min_dist_reg[2][20] ,
         \min_dist_reg[2][19] , \min_dist_reg[2][18] , \min_dist_reg[2][17] ,
         \min_dist_reg[2][16] , \min_dist_reg[2][15] , \min_dist_reg[2][14] ,
         \min_dist_reg[2][13] , \min_dist_reg[2][12] , \min_dist_reg[2][11] ,
         \min_dist_reg[2][10] , \min_dist_reg[2][9] , \min_dist_reg[2][8] ,
         \min_dist_reg[2][7] , \min_dist_reg[2][6] , \min_dist_reg[2][5] ,
         \min_dist_reg[2][4] , \min_dist_reg[2][3] , \min_dist_reg[2][2] ,
         \min_dist_reg[2][1] , \min_dist_reg[2][0] , \min_dist_reg[1][33] ,
         \min_dist_reg[1][32] , \min_dist_reg[1][31] , \min_dist_reg[1][30] ,
         \min_dist_reg[1][29] , \min_dist_reg[1][28] , \min_dist_reg[1][27] ,
         \min_dist_reg[1][26] , \min_dist_reg[1][25] , \min_dist_reg[1][24] ,
         \min_dist_reg[1][23] , \min_dist_reg[1][22] , \min_dist_reg[1][21] ,
         \min_dist_reg[1][20] , \min_dist_reg[1][19] , \min_dist_reg[1][18] ,
         \min_dist_reg[1][17] , \min_dist_reg[1][16] , \min_dist_reg[1][15] ,
         \min_dist_reg[1][14] , \min_dist_reg[1][13] , \min_dist_reg[1][12] ,
         \min_dist_reg[1][11] , \min_dist_reg[1][10] , \min_dist_reg[1][9] ,
         \min_dist_reg[1][8] , \min_dist_reg[1][7] , \min_dist_reg[1][6] ,
         \min_dist_reg[1][5] , \min_dist_reg[1][4] , \min_dist_reg[1][3] ,
         \min_dist_reg[1][2] , \min_dist_reg[1][1] , \min_dist_reg[1][0] ,
         \min_dist_reg[0][33] , \min_dist_reg[0][32] , \min_dist_reg[0][31] ,
         \min_dist_reg[0][30] , \min_dist_reg[0][29] , \min_dist_reg[0][28] ,
         \min_dist_reg[0][27] , \min_dist_reg[0][26] , \min_dist_reg[0][25] ,
         \min_dist_reg[0][24] , \min_dist_reg[0][23] , \min_dist_reg[0][22] ,
         \min_dist_reg[0][21] , \min_dist_reg[0][20] , \min_dist_reg[0][19] ,
         \min_dist_reg[0][18] , \min_dist_reg[0][17] , \min_dist_reg[0][16] ,
         \min_dist_reg[0][15] , \min_dist_reg[0][14] , \min_dist_reg[0][13] ,
         \min_dist_reg[0][12] , \min_dist_reg[0][11] , \min_dist_reg[0][10] ,
         \min_dist_reg[0][9] , \min_dist_reg[0][8] , \min_dist_reg[0][7] ,
         \min_dist_reg[0][6] , \min_dist_reg[0][5] , \min_dist_reg[0][4] ,
         \min_dist_reg[0][3] , \min_dist_reg[0][2] , \min_dist_reg[0][1] ,
         \min_dist_reg[0][0] , \local_min_dist[0][33] ,
         \local_min_dist[0][32] , \local_min_dist[0][31] ,
         \local_min_dist[0][30] , \local_min_dist[0][29] ,
         \local_min_dist[0][28] , \local_min_dist[0][27] ,
         \local_min_dist[0][26] , \local_min_dist[0][25] ,
         \local_min_dist[0][24] , \local_min_dist[0][23] ,
         \local_min_dist[0][22] , \local_min_dist[0][21] ,
         \local_min_dist[0][20] , \local_min_dist[0][19] ,
         \local_min_dist[0][18] , \local_min_dist[0][17] ,
         \local_min_dist[0][16] , \local_min_dist[0][15] ,
         \local_min_dist[0][14] , \local_min_dist[0][13] ,
         \local_min_dist[0][12] , \local_min_dist[0][11] ,
         \local_min_dist[0][10] , \local_min_dist[0][9] ,
         \local_min_dist[0][8] , \local_min_dist[0][7] ,
         \local_min_dist[0][6] , \local_min_dist[0][5] ,
         \local_min_dist[0][4] , \local_min_dist[0][3] ,
         \local_min_dist[0][2] , \local_min_dist[0][1] ,
         \local_min_dist[0][0] , \min_dist[3][33] , \min_dist[3][32] ,
         \min_dist[3][31] , \min_dist[3][30] , \min_dist[3][29] ,
         \min_dist[3][28] , \min_dist[3][27] , \min_dist[3][26] ,
         \min_dist[3][25] , \min_dist[3][24] , \min_dist[3][23] ,
         \min_dist[3][22] , \min_dist[3][21] , \min_dist[3][20] ,
         \min_dist[3][19] , \min_dist[3][18] , \min_dist[3][17] ,
         \min_dist[3][16] , \min_dist[3][15] , \min_dist[3][14] ,
         \min_dist[3][13] , \min_dist[3][12] , \min_dist[3][11] ,
         \min_dist[3][10] , \min_dist[3][9] , \min_dist[3][8] ,
         \min_dist[3][7] , \min_dist[3][6] , \min_dist[3][5] ,
         \min_dist[3][4] , \min_dist[3][3] , \min_dist[3][2] ,
         \min_dist[3][1] , \min_dist[3][0] , \min_dist[2][33] ,
         \min_dist[2][32] , \min_dist[2][31] , \min_dist[2][30] ,
         \min_dist[2][29] , \min_dist[2][28] , \min_dist[2][27] ,
         \min_dist[2][26] , \min_dist[2][25] , \min_dist[2][24] ,
         \min_dist[2][23] , \min_dist[2][22] , \min_dist[2][21] ,
         \min_dist[2][20] , \min_dist[2][19] , \min_dist[2][18] ,
         \min_dist[2][17] , \min_dist[2][16] , \min_dist[2][15] ,
         \min_dist[2][14] , \min_dist[2][13] , \min_dist[2][12] ,
         \min_dist[2][11] , \min_dist[2][10] , \min_dist[2][9] ,
         \min_dist[2][8] , \min_dist[2][7] , \min_dist[2][6] ,
         \min_dist[2][5] , \min_dist[2][4] , \min_dist[2][3] ,
         \min_dist[2][2] , \min_dist[2][1] , \min_dist[2][0] ,
         \min_dist[1][33] , \min_dist[1][32] , \min_dist[1][31] ,
         \min_dist[1][30] , \min_dist[1][29] , \min_dist[1][28] ,
         \min_dist[1][27] , \min_dist[1][26] , \min_dist[1][25] ,
         \min_dist[1][24] , \min_dist[1][23] , \min_dist[1][22] ,
         \min_dist[1][21] , \min_dist[1][20] , \min_dist[1][19] ,
         \min_dist[1][18] , \min_dist[1][17] , \min_dist[1][16] ,
         \min_dist[1][15] , \min_dist[1][14] , \min_dist[1][13] ,
         \min_dist[1][12] , \min_dist[1][11] , \min_dist[1][10] ,
         \min_dist[1][9] , \min_dist[1][8] , \min_dist[1][7] ,
         \min_dist[1][6] , \min_dist[1][5] , \min_dist[1][4] ,
         \min_dist[1][3] , \min_dist[1][2] , \min_dist[1][1] ,
         \min_dist[1][0] , \min_val_reg[3][63] , \min_val_reg[3][62] ,
         \min_val_reg[3][61] , \min_val_reg[3][60] , \min_val_reg[3][59] ,
         \min_val_reg[3][58] , \min_val_reg[3][57] , \min_val_reg[3][56] ,
         \min_val_reg[3][55] , \min_val_reg[3][54] , \min_val_reg[3][53] ,
         \min_val_reg[3][52] , \min_val_reg[3][51] , \min_val_reg[3][50] ,
         \min_val_reg[3][49] , \min_val_reg[3][48] , \min_val_reg[3][47] ,
         \min_val_reg[3][46] , \min_val_reg[3][45] , \min_val_reg[3][44] ,
         \min_val_reg[3][43] , \min_val_reg[3][42] , \min_val_reg[3][41] ,
         \min_val_reg[3][40] , \min_val_reg[3][39] , \min_val_reg[3][38] ,
         \min_val_reg[3][37] , \min_val_reg[3][36] , \min_val_reg[3][35] ,
         \min_val_reg[3][34] , \min_val_reg[3][33] , \min_val_reg[3][32] ,
         \min_val_reg[3][31] , \min_val_reg[3][30] , \min_val_reg[3][29] ,
         \min_val_reg[3][28] , \min_val_reg[3][27] , \min_val_reg[3][26] ,
         \min_val_reg[3][25] , \min_val_reg[3][24] , \min_val_reg[3][23] ,
         \min_val_reg[3][22] , \min_val_reg[3][21] , \min_val_reg[3][20] ,
         \min_val_reg[3][19] , \min_val_reg[3][18] , \min_val_reg[3][17] ,
         \min_val_reg[3][16] , \min_val_reg[3][15] , \min_val_reg[3][14] ,
         \min_val_reg[3][13] , \min_val_reg[3][12] , \min_val_reg[3][11] ,
         \min_val_reg[3][10] , \min_val_reg[3][9] , \min_val_reg[3][8] ,
         \min_val_reg[3][7] , \min_val_reg[3][6] , \min_val_reg[3][5] ,
         \min_val_reg[3][4] , \min_val_reg[3][3] , \min_val_reg[3][2] ,
         \min_val_reg[3][1] , \min_val_reg[3][0] , \min_val_reg[2][63] ,
         \min_val_reg[2][62] , \min_val_reg[2][61] , \min_val_reg[2][60] ,
         \min_val_reg[2][59] , \min_val_reg[2][58] , \min_val_reg[2][57] ,
         \min_val_reg[2][56] , \min_val_reg[2][55] , \min_val_reg[2][54] ,
         \min_val_reg[2][53] , \min_val_reg[2][52] , \min_val_reg[2][51] ,
         \min_val_reg[2][50] , \min_val_reg[2][49] , \min_val_reg[2][48] ,
         \min_val_reg[2][47] , \min_val_reg[2][46] , \min_val_reg[2][45] ,
         \min_val_reg[2][44] , \min_val_reg[2][43] , \min_val_reg[2][42] ,
         \min_val_reg[2][41] , \min_val_reg[2][40] , \min_val_reg[2][39] ,
         \min_val_reg[2][38] , \min_val_reg[2][37] , \min_val_reg[2][36] ,
         \min_val_reg[2][35] , \min_val_reg[2][34] , \min_val_reg[2][33] ,
         \min_val_reg[2][32] , \min_val_reg[2][31] , \min_val_reg[2][30] ,
         \min_val_reg[2][29] , \min_val_reg[2][28] , \min_val_reg[2][27] ,
         \min_val_reg[2][26] , \min_val_reg[2][25] , \min_val_reg[2][24] ,
         \min_val_reg[2][23] , \min_val_reg[2][22] , \min_val_reg[2][21] ,
         \min_val_reg[2][20] , \min_val_reg[2][19] , \min_val_reg[2][18] ,
         \min_val_reg[2][17] , \min_val_reg[2][16] , \min_val_reg[2][15] ,
         \min_val_reg[2][14] , \min_val_reg[2][13] , \min_val_reg[2][12] ,
         \min_val_reg[2][11] , \min_val_reg[2][10] , \min_val_reg[2][9] ,
         \min_val_reg[2][8] , \min_val_reg[2][7] , \min_val_reg[2][6] ,
         \min_val_reg[2][5] , \min_val_reg[2][4] , \min_val_reg[2][3] ,
         \min_val_reg[2][2] , \min_val_reg[2][1] , \min_val_reg[2][0] ,
         \min_val_reg[1][63] , \min_val_reg[1][62] , \min_val_reg[1][61] ,
         \min_val_reg[1][60] , \min_val_reg[1][59] , \min_val_reg[1][58] ,
         \min_val_reg[1][57] , \min_val_reg[1][56] , \min_val_reg[1][55] ,
         \min_val_reg[1][54] , \min_val_reg[1][53] , \min_val_reg[1][52] ,
         \min_val_reg[1][51] , \min_val_reg[1][50] , \min_val_reg[1][49] ,
         \min_val_reg[1][48] , \min_val_reg[1][47] , \min_val_reg[1][46] ,
         \min_val_reg[1][45] , \min_val_reg[1][44] , \min_val_reg[1][43] ,
         \min_val_reg[1][42] , \min_val_reg[1][41] , \min_val_reg[1][40] ,
         \min_val_reg[1][39] , \min_val_reg[1][38] , \min_val_reg[1][37] ,
         \min_val_reg[1][36] , \min_val_reg[1][35] , \min_val_reg[1][34] ,
         \min_val_reg[1][33] , \min_val_reg[1][32] , \min_val_reg[1][31] ,
         \min_val_reg[1][30] , \min_val_reg[1][29] , \min_val_reg[1][28] ,
         \min_val_reg[1][27] , \min_val_reg[1][26] , \min_val_reg[1][25] ,
         \min_val_reg[1][24] , \min_val_reg[1][23] , \min_val_reg[1][22] ,
         \min_val_reg[1][21] , \min_val_reg[1][20] , \min_val_reg[1][19] ,
         \min_val_reg[1][18] , \min_val_reg[1][17] , \min_val_reg[1][16] ,
         \min_val_reg[1][15] , \min_val_reg[1][14] , \min_val_reg[1][13] ,
         \min_val_reg[1][12] , \min_val_reg[1][11] , \min_val_reg[1][10] ,
         \min_val_reg[1][9] , \min_val_reg[1][8] , \min_val_reg[1][7] ,
         \min_val_reg[1][6] , \min_val_reg[1][5] , \min_val_reg[1][4] ,
         \min_val_reg[1][3] , \min_val_reg[1][2] , \min_val_reg[1][1] ,
         \min_val_reg[1][0] , \min_val_reg[0][63] , \min_val_reg[0][62] ,
         \min_val_reg[0][61] , \min_val_reg[0][60] , \min_val_reg[0][59] ,
         \min_val_reg[0][58] , \min_val_reg[0][57] , \min_val_reg[0][56] ,
         \min_val_reg[0][55] , \min_val_reg[0][54] , \min_val_reg[0][53] ,
         \min_val_reg[0][52] , \min_val_reg[0][51] , \min_val_reg[0][50] ,
         \min_val_reg[0][49] , \min_val_reg[0][48] , \min_val_reg[0][47] ,
         \min_val_reg[0][46] , \min_val_reg[0][45] , \min_val_reg[0][44] ,
         \min_val_reg[0][43] , \min_val_reg[0][42] , \min_val_reg[0][41] ,
         \min_val_reg[0][40] , \min_val_reg[0][39] , \min_val_reg[0][38] ,
         \min_val_reg[0][37] , \min_val_reg[0][36] , \min_val_reg[0][35] ,
         \min_val_reg[0][34] , \min_val_reg[0][33] , \min_val_reg[0][32] ,
         \min_val_reg[0][31] , \min_val_reg[0][30] , \min_val_reg[0][29] ,
         \min_val_reg[0][28] , \min_val_reg[0][27] , \min_val_reg[0][26] ,
         \min_val_reg[0][25] , \min_val_reg[0][24] , \min_val_reg[0][23] ,
         \min_val_reg[0][22] , \min_val_reg[0][21] , \min_val_reg[0][20] ,
         \min_val_reg[0][19] , \min_val_reg[0][18] , \min_val_reg[0][17] ,
         \min_val_reg[0][16] , \min_val_reg[0][15] , \min_val_reg[0][14] ,
         \min_val_reg[0][13] , \min_val_reg[0][12] , \min_val_reg[0][11] ,
         \min_val_reg[0][10] , \min_val_reg[0][9] , \min_val_reg[0][8] ,
         \min_val_reg[0][7] , \min_val_reg[0][6] , \min_val_reg[0][5] ,
         \min_val_reg[0][4] , \min_val_reg[0][3] , \min_val_reg[0][2] ,
         \min_val_reg[0][1] , \min_val_reg[0][0] , n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900;

  DFF \min_dist_reg_reg[0][0]  ( .D(\local_min_dist[0][0] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][0] ) );
  DFF \min_dist_reg_reg[0][1]  ( .D(\local_min_dist[0][1] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][1] ) );
  DFF \min_dist_reg_reg[0][2]  ( .D(\local_min_dist[0][2] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][2] ) );
  DFF \min_dist_reg_reg[0][3]  ( .D(\local_min_dist[0][3] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][3] ) );
  DFF \min_dist_reg_reg[0][4]  ( .D(\local_min_dist[0][4] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][4] ) );
  DFF \min_dist_reg_reg[0][5]  ( .D(\local_min_dist[0][5] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][5] ) );
  DFF \min_dist_reg_reg[0][6]  ( .D(\local_min_dist[0][6] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][6] ) );
  DFF \min_dist_reg_reg[0][7]  ( .D(\local_min_dist[0][7] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][7] ) );
  DFF \min_dist_reg_reg[0][8]  ( .D(\local_min_dist[0][8] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][8] ) );
  DFF \min_dist_reg_reg[0][9]  ( .D(\local_min_dist[0][9] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][9] ) );
  DFF \min_dist_reg_reg[0][10]  ( .D(\local_min_dist[0][10] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][10] ) );
  DFF \min_dist_reg_reg[0][11]  ( .D(\local_min_dist[0][11] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][11] ) );
  DFF \min_dist_reg_reg[0][12]  ( .D(\local_min_dist[0][12] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][12] ) );
  DFF \min_dist_reg_reg[0][13]  ( .D(\local_min_dist[0][13] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][13] ) );
  DFF \min_dist_reg_reg[0][14]  ( .D(\local_min_dist[0][14] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][14] ) );
  DFF \min_dist_reg_reg[0][15]  ( .D(\local_min_dist[0][15] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][15] ) );
  DFF \min_dist_reg_reg[0][16]  ( .D(\local_min_dist[0][16] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][16] ) );
  DFF \min_dist_reg_reg[0][17]  ( .D(\local_min_dist[0][17] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][17] ) );
  DFF \min_dist_reg_reg[0][18]  ( .D(\local_min_dist[0][18] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][18] ) );
  DFF \min_dist_reg_reg[0][19]  ( .D(\local_min_dist[0][19] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][19] ) );
  DFF \min_dist_reg_reg[0][20]  ( .D(\local_min_dist[0][20] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][20] ) );
  DFF \min_dist_reg_reg[0][21]  ( .D(\local_min_dist[0][21] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][21] ) );
  DFF \min_dist_reg_reg[0][22]  ( .D(\local_min_dist[0][22] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][22] ) );
  DFF \min_dist_reg_reg[0][23]  ( .D(\local_min_dist[0][23] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][23] ) );
  DFF \min_dist_reg_reg[0][24]  ( .D(\local_min_dist[0][24] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][24] ) );
  DFF \min_dist_reg_reg[0][25]  ( .D(\local_min_dist[0][25] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][25] ) );
  DFF \min_dist_reg_reg[0][26]  ( .D(\local_min_dist[0][26] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][26] ) );
  DFF \min_dist_reg_reg[0][27]  ( .D(\local_min_dist[0][27] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][27] ) );
  DFF \min_dist_reg_reg[0][28]  ( .D(\local_min_dist[0][28] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][28] ) );
  DFF \min_dist_reg_reg[0][29]  ( .D(\local_min_dist[0][29] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][29] ) );
  DFF \min_dist_reg_reg[0][30]  ( .D(\local_min_dist[0][30] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][30] ) );
  DFF \min_dist_reg_reg[0][31]  ( .D(\local_min_dist[0][31] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][31] ) );
  DFF \min_dist_reg_reg[0][32]  ( .D(\local_min_dist[0][32] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][32] ) );
  DFF \min_dist_reg_reg[0][33]  ( .D(\local_min_dist[0][33] ), .CLK(clk), 
        .RST(rst), .I(1'b1), .Q(\min_dist_reg[0][33] ) );
  DFF \min_dist_reg_reg[1][0]  ( .D(\min_dist[1][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][0] ) );
  DFF \min_dist_reg_reg[1][1]  ( .D(\min_dist[1][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][1] ) );
  DFF \min_dist_reg_reg[1][2]  ( .D(\min_dist[1][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][2] ) );
  DFF \min_dist_reg_reg[1][3]  ( .D(\min_dist[1][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][3] ) );
  DFF \min_dist_reg_reg[1][4]  ( .D(\min_dist[1][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][4] ) );
  DFF \min_dist_reg_reg[1][5]  ( .D(\min_dist[1][5] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][5] ) );
  DFF \min_dist_reg_reg[1][6]  ( .D(\min_dist[1][6] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][6] ) );
  DFF \min_dist_reg_reg[1][7]  ( .D(\min_dist[1][7] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][7] ) );
  DFF \min_dist_reg_reg[1][8]  ( .D(\min_dist[1][8] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][8] ) );
  DFF \min_dist_reg_reg[1][9]  ( .D(\min_dist[1][9] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][9] ) );
  DFF \min_dist_reg_reg[1][10]  ( .D(\min_dist[1][10] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][10] ) );
  DFF \min_dist_reg_reg[1][11]  ( .D(\min_dist[1][11] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][11] ) );
  DFF \min_dist_reg_reg[1][12]  ( .D(\min_dist[1][12] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][12] ) );
  DFF \min_dist_reg_reg[1][13]  ( .D(\min_dist[1][13] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][13] ) );
  DFF \min_dist_reg_reg[1][14]  ( .D(\min_dist[1][14] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][14] ) );
  DFF \min_dist_reg_reg[1][15]  ( .D(\min_dist[1][15] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][15] ) );
  DFF \min_dist_reg_reg[1][16]  ( .D(\min_dist[1][16] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][16] ) );
  DFF \min_dist_reg_reg[1][17]  ( .D(\min_dist[1][17] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][17] ) );
  DFF \min_dist_reg_reg[1][18]  ( .D(\min_dist[1][18] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][18] ) );
  DFF \min_dist_reg_reg[1][19]  ( .D(\min_dist[1][19] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][19] ) );
  DFF \min_dist_reg_reg[1][20]  ( .D(\min_dist[1][20] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][20] ) );
  DFF \min_dist_reg_reg[1][21]  ( .D(\min_dist[1][21] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][21] ) );
  DFF \min_dist_reg_reg[1][22]  ( .D(\min_dist[1][22] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][22] ) );
  DFF \min_dist_reg_reg[1][23]  ( .D(\min_dist[1][23] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][23] ) );
  DFF \min_dist_reg_reg[1][24]  ( .D(\min_dist[1][24] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][24] ) );
  DFF \min_dist_reg_reg[1][25]  ( .D(\min_dist[1][25] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][25] ) );
  DFF \min_dist_reg_reg[1][26]  ( .D(\min_dist[1][26] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][26] ) );
  DFF \min_dist_reg_reg[1][27]  ( .D(\min_dist[1][27] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][27] ) );
  DFF \min_dist_reg_reg[1][28]  ( .D(\min_dist[1][28] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][28] ) );
  DFF \min_dist_reg_reg[1][29]  ( .D(\min_dist[1][29] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][29] ) );
  DFF \min_dist_reg_reg[1][30]  ( .D(\min_dist[1][30] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][30] ) );
  DFF \min_dist_reg_reg[1][31]  ( .D(\min_dist[1][31] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][31] ) );
  DFF \min_dist_reg_reg[1][32]  ( .D(\min_dist[1][32] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][32] ) );
  DFF \min_dist_reg_reg[1][33]  ( .D(\min_dist[1][33] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][33] ) );
  DFF \min_dist_reg_reg[2][0]  ( .D(\min_dist[2][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][0] ) );
  DFF \min_dist_reg_reg[2][1]  ( .D(\min_dist[2][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][1] ) );
  DFF \min_dist_reg_reg[2][2]  ( .D(\min_dist[2][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][2] ) );
  DFF \min_dist_reg_reg[2][3]  ( .D(\min_dist[2][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][3] ) );
  DFF \min_dist_reg_reg[2][4]  ( .D(\min_dist[2][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][4] ) );
  DFF \min_dist_reg_reg[2][5]  ( .D(\min_dist[2][5] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][5] ) );
  DFF \min_dist_reg_reg[2][6]  ( .D(\min_dist[2][6] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][6] ) );
  DFF \min_dist_reg_reg[2][7]  ( .D(\min_dist[2][7] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][7] ) );
  DFF \min_dist_reg_reg[2][8]  ( .D(\min_dist[2][8] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][8] ) );
  DFF \min_dist_reg_reg[2][9]  ( .D(\min_dist[2][9] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][9] ) );
  DFF \min_dist_reg_reg[2][10]  ( .D(\min_dist[2][10] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][10] ) );
  DFF \min_dist_reg_reg[2][11]  ( .D(\min_dist[2][11] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][11] ) );
  DFF \min_dist_reg_reg[2][12]  ( .D(\min_dist[2][12] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][12] ) );
  DFF \min_dist_reg_reg[2][13]  ( .D(\min_dist[2][13] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][13] ) );
  DFF \min_dist_reg_reg[2][14]  ( .D(\min_dist[2][14] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][14] ) );
  DFF \min_dist_reg_reg[2][15]  ( .D(\min_dist[2][15] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][15] ) );
  DFF \min_dist_reg_reg[2][16]  ( .D(\min_dist[2][16] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][16] ) );
  DFF \min_dist_reg_reg[2][17]  ( .D(\min_dist[2][17] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][17] ) );
  DFF \min_dist_reg_reg[2][18]  ( .D(\min_dist[2][18] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][18] ) );
  DFF \min_dist_reg_reg[2][19]  ( .D(\min_dist[2][19] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][19] ) );
  DFF \min_dist_reg_reg[2][20]  ( .D(\min_dist[2][20] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][20] ) );
  DFF \min_dist_reg_reg[2][21]  ( .D(\min_dist[2][21] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][21] ) );
  DFF \min_dist_reg_reg[2][22]  ( .D(\min_dist[2][22] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][22] ) );
  DFF \min_dist_reg_reg[2][23]  ( .D(\min_dist[2][23] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][23] ) );
  DFF \min_dist_reg_reg[2][24]  ( .D(\min_dist[2][24] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][24] ) );
  DFF \min_dist_reg_reg[2][25]  ( .D(\min_dist[2][25] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][25] ) );
  DFF \min_dist_reg_reg[2][26]  ( .D(\min_dist[2][26] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][26] ) );
  DFF \min_dist_reg_reg[2][27]  ( .D(\min_dist[2][27] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][27] ) );
  DFF \min_dist_reg_reg[2][28]  ( .D(\min_dist[2][28] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][28] ) );
  DFF \min_dist_reg_reg[2][29]  ( .D(\min_dist[2][29] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][29] ) );
  DFF \min_dist_reg_reg[2][30]  ( .D(\min_dist[2][30] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][30] ) );
  DFF \min_dist_reg_reg[2][31]  ( .D(\min_dist[2][31] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][31] ) );
  DFF \min_dist_reg_reg[2][32]  ( .D(\min_dist[2][32] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][32] ) );
  DFF \min_dist_reg_reg[2][33]  ( .D(\min_dist[2][33] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][33] ) );
  DFF \min_dist_reg_reg[3][0]  ( .D(\min_dist[3][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][0] ) );
  DFF \min_dist_reg_reg[3][1]  ( .D(\min_dist[3][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][1] ) );
  DFF \min_dist_reg_reg[3][2]  ( .D(\min_dist[3][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][2] ) );
  DFF \min_dist_reg_reg[3][3]  ( .D(\min_dist[3][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][3] ) );
  DFF \min_dist_reg_reg[3][4]  ( .D(\min_dist[3][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][4] ) );
  DFF \min_dist_reg_reg[3][5]  ( .D(\min_dist[3][5] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][5] ) );
  DFF \min_dist_reg_reg[3][6]  ( .D(\min_dist[3][6] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][6] ) );
  DFF \min_dist_reg_reg[3][7]  ( .D(\min_dist[3][7] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][7] ) );
  DFF \min_dist_reg_reg[3][8]  ( .D(\min_dist[3][8] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][8] ) );
  DFF \min_dist_reg_reg[3][9]  ( .D(\min_dist[3][9] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][9] ) );
  DFF \min_dist_reg_reg[3][10]  ( .D(\min_dist[3][10] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][10] ) );
  DFF \min_dist_reg_reg[3][11]  ( .D(\min_dist[3][11] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][11] ) );
  DFF \min_dist_reg_reg[3][12]  ( .D(\min_dist[3][12] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][12] ) );
  DFF \min_dist_reg_reg[3][13]  ( .D(\min_dist[3][13] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][13] ) );
  DFF \min_dist_reg_reg[3][14]  ( .D(\min_dist[3][14] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][14] ) );
  DFF \min_dist_reg_reg[3][15]  ( .D(\min_dist[3][15] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][15] ) );
  DFF \min_dist_reg_reg[3][16]  ( .D(\min_dist[3][16] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][16] ) );
  DFF \min_dist_reg_reg[3][17]  ( .D(\min_dist[3][17] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][17] ) );
  DFF \min_dist_reg_reg[3][18]  ( .D(\min_dist[3][18] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][18] ) );
  DFF \min_dist_reg_reg[3][19]  ( .D(\min_dist[3][19] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][19] ) );
  DFF \min_dist_reg_reg[3][20]  ( .D(\min_dist[3][20] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][20] ) );
  DFF \min_dist_reg_reg[3][21]  ( .D(\min_dist[3][21] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][21] ) );
  DFF \min_dist_reg_reg[3][22]  ( .D(\min_dist[3][22] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][22] ) );
  DFF \min_dist_reg_reg[3][23]  ( .D(\min_dist[3][23] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][23] ) );
  DFF \min_dist_reg_reg[3][24]  ( .D(\min_dist[3][24] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][24] ) );
  DFF \min_dist_reg_reg[3][25]  ( .D(\min_dist[3][25] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][25] ) );
  DFF \min_dist_reg_reg[3][26]  ( .D(\min_dist[3][26] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][26] ) );
  DFF \min_dist_reg_reg[3][27]  ( .D(\min_dist[3][27] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][27] ) );
  DFF \min_dist_reg_reg[3][28]  ( .D(\min_dist[3][28] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][28] ) );
  DFF \min_dist_reg_reg[3][29]  ( .D(\min_dist[3][29] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][29] ) );
  DFF \min_dist_reg_reg[3][30]  ( .D(\min_dist[3][30] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][30] ) );
  DFF \min_dist_reg_reg[3][31]  ( .D(\min_dist[3][31] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][31] ) );
  DFF \min_dist_reg_reg[3][32]  ( .D(\min_dist[3][32] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][32] ) );
  DFF \min_dist_reg_reg[3][33]  ( .D(\min_dist[3][33] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][33] ) );
  DFF \min_val_reg_reg[0][0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][0] ) );
  DFF \min_val_reg_reg[0][1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][1] ) );
  DFF \min_val_reg_reg[0][2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][2] ) );
  DFF \min_val_reg_reg[0][3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][3] ) );
  DFF \min_val_reg_reg[0][4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][4] ) );
  DFF \min_val_reg_reg[0][5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][5] ) );
  DFF \min_val_reg_reg[0][6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][6] ) );
  DFF \min_val_reg_reg[0][7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][7] ) );
  DFF \min_val_reg_reg[0][8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][8] ) );
  DFF \min_val_reg_reg[0][9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][9] ) );
  DFF \min_val_reg_reg[0][10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][10] ) );
  DFF \min_val_reg_reg[0][11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][11] ) );
  DFF \min_val_reg_reg[0][12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][12] ) );
  DFF \min_val_reg_reg[0][13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][13] ) );
  DFF \min_val_reg_reg[0][14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][14] ) );
  DFF \min_val_reg_reg[0][15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][15] ) );
  DFF \min_val_reg_reg[0][16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][16] ) );
  DFF \min_val_reg_reg[0][17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][17] ) );
  DFF \min_val_reg_reg[0][18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][18] ) );
  DFF \min_val_reg_reg[0][19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][19] ) );
  DFF \min_val_reg_reg[0][20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][20] ) );
  DFF \min_val_reg_reg[0][21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][21] ) );
  DFF \min_val_reg_reg[0][22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][22] ) );
  DFF \min_val_reg_reg[0][23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][23] ) );
  DFF \min_val_reg_reg[0][24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][24] ) );
  DFF \min_val_reg_reg[0][25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][25] ) );
  DFF \min_val_reg_reg[0][26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][26] ) );
  DFF \min_val_reg_reg[0][27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][27] ) );
  DFF \min_val_reg_reg[0][28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][28] ) );
  DFF \min_val_reg_reg[0][29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][29] ) );
  DFF \min_val_reg_reg[0][30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][30] ) );
  DFF \min_val_reg_reg[0][31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][31] ) );
  DFF \min_val_reg_reg[0][32]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][32] ) );
  DFF \min_val_reg_reg[0][33]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][33] ) );
  DFF \min_val_reg_reg[0][34]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][34] ) );
  DFF \min_val_reg_reg[0][35]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][35] ) );
  DFF \min_val_reg_reg[0][36]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][36] ) );
  DFF \min_val_reg_reg[0][37]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][37] ) );
  DFF \min_val_reg_reg[0][38]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][38] ) );
  DFF \min_val_reg_reg[0][39]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][39] ) );
  DFF \min_val_reg_reg[0][40]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][40] ) );
  DFF \min_val_reg_reg[0][41]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][41] ) );
  DFF \min_val_reg_reg[0][42]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][42] ) );
  DFF \min_val_reg_reg[0][43]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][43] ) );
  DFF \min_val_reg_reg[0][44]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][44] ) );
  DFF \min_val_reg_reg[0][45]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][45] ) );
  DFF \min_val_reg_reg[0][46]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][46] ) );
  DFF \min_val_reg_reg[0][47]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][47] ) );
  DFF \min_val_reg_reg[0][48]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][48] ) );
  DFF \min_val_reg_reg[0][49]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][49] ) );
  DFF \min_val_reg_reg[0][50]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][50] ) );
  DFF \min_val_reg_reg[0][51]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][51] ) );
  DFF \min_val_reg_reg[0][52]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][52] ) );
  DFF \min_val_reg_reg[0][53]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][53] ) );
  DFF \min_val_reg_reg[0][54]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][54] ) );
  DFF \min_val_reg_reg[0][55]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][55] ) );
  DFF \min_val_reg_reg[0][56]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][56] ) );
  DFF \min_val_reg_reg[0][57]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][57] ) );
  DFF \min_val_reg_reg[0][58]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][58] ) );
  DFF \min_val_reg_reg[0][59]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][59] ) );
  DFF \min_val_reg_reg[0][60]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][60] ) );
  DFF \min_val_reg_reg[0][61]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][61] ) );
  DFF \min_val_reg_reg[0][62]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][62] ) );
  DFF \min_val_reg_reg[0][63]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][63] ) );
  DFF \min_val_reg_reg[1][0]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][0] ) );
  DFF \min_val_reg_reg[1][1]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][1] ) );
  DFF \min_val_reg_reg[1][2]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][2] ) );
  DFF \min_val_reg_reg[1][3]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][3] ) );
  DFF \min_val_reg_reg[1][4]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][4] ) );
  DFF \min_val_reg_reg[1][5]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][5] ) );
  DFF \min_val_reg_reg[1][6]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][6] ) );
  DFF \min_val_reg_reg[1][7]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][7] ) );
  DFF \min_val_reg_reg[1][8]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][8] ) );
  DFF \min_val_reg_reg[1][9]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][9] ) );
  DFF \min_val_reg_reg[1][10]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][10] ) );
  DFF \min_val_reg_reg[1][11]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][11] ) );
  DFF \min_val_reg_reg[1][12]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][12] ) );
  DFF \min_val_reg_reg[1][13]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][13] ) );
  DFF \min_val_reg_reg[1][14]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][14] ) );
  DFF \min_val_reg_reg[1][15]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][15] ) );
  DFF \min_val_reg_reg[1][16]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][16] ) );
  DFF \min_val_reg_reg[1][17]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][17] ) );
  DFF \min_val_reg_reg[1][18]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][18] ) );
  DFF \min_val_reg_reg[1][19]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][19] ) );
  DFF \min_val_reg_reg[1][20]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][20] ) );
  DFF \min_val_reg_reg[1][21]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][21] ) );
  DFF \min_val_reg_reg[1][22]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][22] ) );
  DFF \min_val_reg_reg[1][23]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][23] ) );
  DFF \min_val_reg_reg[1][24]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][24] ) );
  DFF \min_val_reg_reg[1][25]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][25] ) );
  DFF \min_val_reg_reg[1][26]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][26] ) );
  DFF \min_val_reg_reg[1][27]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][27] ) );
  DFF \min_val_reg_reg[1][28]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][28] ) );
  DFF \min_val_reg_reg[1][29]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][29] ) );
  DFF \min_val_reg_reg[1][30]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][30] ) );
  DFF \min_val_reg_reg[1][31]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][31] ) );
  DFF \min_val_reg_reg[1][32]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][32] ) );
  DFF \min_val_reg_reg[1][33]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][33] ) );
  DFF \min_val_reg_reg[1][34]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][34] ) );
  DFF \min_val_reg_reg[1][35]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][35] ) );
  DFF \min_val_reg_reg[1][36]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][36] ) );
  DFF \min_val_reg_reg[1][37]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][37] ) );
  DFF \min_val_reg_reg[1][38]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][38] ) );
  DFF \min_val_reg_reg[1][39]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][39] ) );
  DFF \min_val_reg_reg[1][40]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][40] ) );
  DFF \min_val_reg_reg[1][41]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][41] ) );
  DFF \min_val_reg_reg[1][42]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][42] ) );
  DFF \min_val_reg_reg[1][43]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][43] ) );
  DFF \min_val_reg_reg[1][44]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][44] ) );
  DFF \min_val_reg_reg[1][45]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][45] ) );
  DFF \min_val_reg_reg[1][46]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][46] ) );
  DFF \min_val_reg_reg[1][47]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][47] ) );
  DFF \min_val_reg_reg[1][48]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][48] ) );
  DFF \min_val_reg_reg[1][49]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][49] ) );
  DFF \min_val_reg_reg[1][50]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][50] ) );
  DFF \min_val_reg_reg[1][51]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][51] ) );
  DFF \min_val_reg_reg[1][52]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][52] ) );
  DFF \min_val_reg_reg[1][53]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][53] ) );
  DFF \min_val_reg_reg[1][54]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][54] ) );
  DFF \min_val_reg_reg[1][55]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][55] ) );
  DFF \min_val_reg_reg[1][56]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][56] ) );
  DFF \min_val_reg_reg[1][57]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][57] ) );
  DFF \min_val_reg_reg[1][58]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][58] ) );
  DFF \min_val_reg_reg[1][59]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][59] ) );
  DFF \min_val_reg_reg[1][60]  ( .D(o[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][60] ) );
  DFF \min_val_reg_reg[1][61]  ( .D(o[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][61] ) );
  DFF \min_val_reg_reg[1][62]  ( .D(o[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][62] ) );
  DFF \min_val_reg_reg[1][63]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][63] ) );
  DFF \min_val_reg_reg[2][0]  ( .D(o[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][0] ) );
  DFF \min_val_reg_reg[2][1]  ( .D(o[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][1] ) );
  DFF \min_val_reg_reg[2][2]  ( .D(o[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][2] ) );
  DFF \min_val_reg_reg[2][3]  ( .D(o[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][3] ) );
  DFF \min_val_reg_reg[2][4]  ( .D(o[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][4] ) );
  DFF \min_val_reg_reg[2][5]  ( .D(o[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][5] ) );
  DFF \min_val_reg_reg[2][6]  ( .D(o[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][6] ) );
  DFF \min_val_reg_reg[2][7]  ( .D(o[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][7] ) );
  DFF \min_val_reg_reg[2][8]  ( .D(o[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][8] ) );
  DFF \min_val_reg_reg[2][9]  ( .D(o[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][9] ) );
  DFF \min_val_reg_reg[2][10]  ( .D(o[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][10] ) );
  DFF \min_val_reg_reg[2][11]  ( .D(o[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][11] ) );
  DFF \min_val_reg_reg[2][12]  ( .D(o[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][12] ) );
  DFF \min_val_reg_reg[2][13]  ( .D(o[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][13] ) );
  DFF \min_val_reg_reg[2][14]  ( .D(o[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][14] ) );
  DFF \min_val_reg_reg[2][15]  ( .D(o[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][15] ) );
  DFF \min_val_reg_reg[2][16]  ( .D(o[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][16] ) );
  DFF \min_val_reg_reg[2][17]  ( .D(o[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][17] ) );
  DFF \min_val_reg_reg[2][18]  ( .D(o[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][18] ) );
  DFF \min_val_reg_reg[2][19]  ( .D(o[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][19] ) );
  DFF \min_val_reg_reg[2][20]  ( .D(o[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][20] ) );
  DFF \min_val_reg_reg[2][21]  ( .D(o[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][21] ) );
  DFF \min_val_reg_reg[2][22]  ( .D(o[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][22] ) );
  DFF \min_val_reg_reg[2][23]  ( .D(o[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][23] ) );
  DFF \min_val_reg_reg[2][24]  ( .D(o[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][24] ) );
  DFF \min_val_reg_reg[2][25]  ( .D(o[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][25] ) );
  DFF \min_val_reg_reg[2][26]  ( .D(o[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][26] ) );
  DFF \min_val_reg_reg[2][27]  ( .D(o[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][27] ) );
  DFF \min_val_reg_reg[2][28]  ( .D(o[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][28] ) );
  DFF \min_val_reg_reg[2][29]  ( .D(o[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][29] ) );
  DFF \min_val_reg_reg[2][30]  ( .D(o[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][30] ) );
  DFF \min_val_reg_reg[2][31]  ( .D(o[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][31] ) );
  DFF \min_val_reg_reg[2][32]  ( .D(o[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][32] ) );
  DFF \min_val_reg_reg[2][33]  ( .D(o[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][33] ) );
  DFF \min_val_reg_reg[2][34]  ( .D(o[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][34] ) );
  DFF \min_val_reg_reg[2][35]  ( .D(o[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][35] ) );
  DFF \min_val_reg_reg[2][36]  ( .D(o[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][36] ) );
  DFF \min_val_reg_reg[2][37]  ( .D(o[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][37] ) );
  DFF \min_val_reg_reg[2][38]  ( .D(o[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][38] ) );
  DFF \min_val_reg_reg[2][39]  ( .D(o[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][39] ) );
  DFF \min_val_reg_reg[2][40]  ( .D(o[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][40] ) );
  DFF \min_val_reg_reg[2][41]  ( .D(o[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][41] ) );
  DFF \min_val_reg_reg[2][42]  ( .D(o[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][42] ) );
  DFF \min_val_reg_reg[2][43]  ( .D(o[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][43] ) );
  DFF \min_val_reg_reg[2][44]  ( .D(o[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][44] ) );
  DFF \min_val_reg_reg[2][45]  ( .D(o[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][45] ) );
  DFF \min_val_reg_reg[2][46]  ( .D(o[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][46] ) );
  DFF \min_val_reg_reg[2][47]  ( .D(o[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][47] ) );
  DFF \min_val_reg_reg[2][48]  ( .D(o[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][48] ) );
  DFF \min_val_reg_reg[2][49]  ( .D(o[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][49] ) );
  DFF \min_val_reg_reg[2][50]  ( .D(o[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][50] ) );
  DFF \min_val_reg_reg[2][51]  ( .D(o[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][51] ) );
  DFF \min_val_reg_reg[2][52]  ( .D(o[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][52] ) );
  DFF \min_val_reg_reg[2][53]  ( .D(o[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][53] ) );
  DFF \min_val_reg_reg[2][54]  ( .D(o[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][54] ) );
  DFF \min_val_reg_reg[2][55]  ( .D(o[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][55] ) );
  DFF \min_val_reg_reg[2][56]  ( .D(o[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][56] ) );
  DFF \min_val_reg_reg[2][57]  ( .D(o[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][57] ) );
  DFF \min_val_reg_reg[2][58]  ( .D(o[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][58] ) );
  DFF \min_val_reg_reg[2][59]  ( .D(o[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][59] ) );
  DFF \min_val_reg_reg[2][60]  ( .D(o[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][60] ) );
  DFF \min_val_reg_reg[2][61]  ( .D(o[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][61] ) );
  DFF \min_val_reg_reg[2][62]  ( .D(o[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][62] ) );
  DFF \min_val_reg_reg[2][63]  ( .D(o[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][63] ) );
  DFF \min_val_reg_reg[3][0]  ( .D(o[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][0] ) );
  DFF \min_val_reg_reg[3][1]  ( .D(o[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][1] ) );
  DFF \min_val_reg_reg[3][2]  ( .D(o[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][2] ) );
  DFF \min_val_reg_reg[3][3]  ( .D(o[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][3] ) );
  DFF \min_val_reg_reg[3][4]  ( .D(o[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][4] ) );
  DFF \min_val_reg_reg[3][5]  ( .D(o[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][5] ) );
  DFF \min_val_reg_reg[3][6]  ( .D(o[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][6] ) );
  DFF \min_val_reg_reg[3][7]  ( .D(o[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][7] ) );
  DFF \min_val_reg_reg[3][8]  ( .D(o[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][8] ) );
  DFF \min_val_reg_reg[3][9]  ( .D(o[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][9] ) );
  DFF \min_val_reg_reg[3][10]  ( .D(o[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][10] ) );
  DFF \min_val_reg_reg[3][11]  ( .D(o[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][11] ) );
  DFF \min_val_reg_reg[3][12]  ( .D(o[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][12] ) );
  DFF \min_val_reg_reg[3][13]  ( .D(o[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][13] ) );
  DFF \min_val_reg_reg[3][14]  ( .D(o[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][14] ) );
  DFF \min_val_reg_reg[3][15]  ( .D(o[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][15] ) );
  DFF \min_val_reg_reg[3][16]  ( .D(o[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][16] ) );
  DFF \min_val_reg_reg[3][17]  ( .D(o[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][17] ) );
  DFF \min_val_reg_reg[3][18]  ( .D(o[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][18] ) );
  DFF \min_val_reg_reg[3][19]  ( .D(o[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][19] ) );
  DFF \min_val_reg_reg[3][20]  ( .D(o[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][20] ) );
  DFF \min_val_reg_reg[3][21]  ( .D(o[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][21] ) );
  DFF \min_val_reg_reg[3][22]  ( .D(o[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][22] ) );
  DFF \min_val_reg_reg[3][23]  ( .D(o[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][23] ) );
  DFF \min_val_reg_reg[3][24]  ( .D(o[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][24] ) );
  DFF \min_val_reg_reg[3][25]  ( .D(o[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][25] ) );
  DFF \min_val_reg_reg[3][26]  ( .D(o[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][26] ) );
  DFF \min_val_reg_reg[3][27]  ( .D(o[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][27] ) );
  DFF \min_val_reg_reg[3][28]  ( .D(o[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][28] ) );
  DFF \min_val_reg_reg[3][29]  ( .D(o[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][29] ) );
  DFF \min_val_reg_reg[3][30]  ( .D(o[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][30] ) );
  DFF \min_val_reg_reg[3][31]  ( .D(o[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][31] ) );
  DFF \min_val_reg_reg[3][32]  ( .D(o[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][32] ) );
  DFF \min_val_reg_reg[3][33]  ( .D(o[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][33] ) );
  DFF \min_val_reg_reg[3][34]  ( .D(o[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][34] ) );
  DFF \min_val_reg_reg[3][35]  ( .D(o[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][35] ) );
  DFF \min_val_reg_reg[3][36]  ( .D(o[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][36] ) );
  DFF \min_val_reg_reg[3][37]  ( .D(o[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][37] ) );
  DFF \min_val_reg_reg[3][38]  ( .D(o[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][38] ) );
  DFF \min_val_reg_reg[3][39]  ( .D(o[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][39] ) );
  DFF \min_val_reg_reg[3][40]  ( .D(o[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][40] ) );
  DFF \min_val_reg_reg[3][41]  ( .D(o[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][41] ) );
  DFF \min_val_reg_reg[3][42]  ( .D(o[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][42] ) );
  DFF \min_val_reg_reg[3][43]  ( .D(o[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][43] ) );
  DFF \min_val_reg_reg[3][44]  ( .D(o[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][44] ) );
  DFF \min_val_reg_reg[3][45]  ( .D(o[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][45] ) );
  DFF \min_val_reg_reg[3][46]  ( .D(o[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][46] ) );
  DFF \min_val_reg_reg[3][47]  ( .D(o[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][47] ) );
  DFF \min_val_reg_reg[3][48]  ( .D(o[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][48] ) );
  DFF \min_val_reg_reg[3][49]  ( .D(o[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][49] ) );
  DFF \min_val_reg_reg[3][50]  ( .D(o[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][50] ) );
  DFF \min_val_reg_reg[3][51]  ( .D(o[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][51] ) );
  DFF \min_val_reg_reg[3][52]  ( .D(o[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][52] ) );
  DFF \min_val_reg_reg[3][53]  ( .D(o[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][53] ) );
  DFF \min_val_reg_reg[3][54]  ( .D(o[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][54] ) );
  DFF \min_val_reg_reg[3][55]  ( .D(o[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][55] ) );
  DFF \min_val_reg_reg[3][56]  ( .D(o[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][56] ) );
  DFF \min_val_reg_reg[3][57]  ( .D(o[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][57] ) );
  DFF \min_val_reg_reg[3][58]  ( .D(o[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][58] ) );
  DFF \min_val_reg_reg[3][59]  ( .D(o[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][59] ) );
  DFF \min_val_reg_reg[3][60]  ( .D(o[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][60] ) );
  DFF \min_val_reg_reg[3][61]  ( .D(o[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][61] ) );
  DFF \min_val_reg_reg[3][62]  ( .D(o[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][62] ) );
  DFF \min_val_reg_reg[3][63]  ( .D(o[255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][63] ) );
  XNOR U395 ( .A(n1418), .B(n1419), .Z(n393) );
  XNOR U396 ( .A(n2762), .B(n2763), .Z(n394) );
  XNOR U397 ( .A(n2777), .B(n2778), .Z(n395) );
  XOR U398 ( .A(\min_val_reg[0][9] ), .B(n396), .Z(o[9]) );
  AND U399 ( .A(n397), .B(n398), .Z(n396) );
  XOR U400 ( .A(n399), .B(n400), .Z(o[99]) );
  AND U401 ( .A(n401), .B(n402), .Z(n399) );
  XOR U402 ( .A(n403), .B(n404), .Z(o[98]) );
  AND U403 ( .A(n401), .B(n405), .Z(n403) );
  XOR U404 ( .A(n406), .B(n407), .Z(o[97]) );
  AND U405 ( .A(n401), .B(n408), .Z(n406) );
  XOR U406 ( .A(n409), .B(n410), .Z(o[96]) );
  AND U407 ( .A(n401), .B(n411), .Z(n409) );
  XOR U408 ( .A(n412), .B(n413), .Z(o[95]) );
  AND U409 ( .A(n401), .B(n414), .Z(n412) );
  XOR U410 ( .A(n415), .B(n416), .Z(o[94]) );
  AND U411 ( .A(n401), .B(n417), .Z(n415) );
  XOR U412 ( .A(n418), .B(n419), .Z(o[93]) );
  AND U413 ( .A(n401), .B(n420), .Z(n418) );
  XOR U414 ( .A(n421), .B(n422), .Z(o[92]) );
  AND U415 ( .A(n401), .B(n423), .Z(n421) );
  XOR U416 ( .A(n424), .B(n425), .Z(o[91]) );
  AND U417 ( .A(n401), .B(n426), .Z(n424) );
  XOR U418 ( .A(n427), .B(n428), .Z(o[90]) );
  AND U419 ( .A(n401), .B(n429), .Z(n427) );
  XOR U420 ( .A(\min_val_reg[0][8] ), .B(n430), .Z(o[8]) );
  AND U421 ( .A(n397), .B(n431), .Z(n430) );
  XOR U422 ( .A(n432), .B(n433), .Z(o[89]) );
  AND U423 ( .A(n401), .B(n434), .Z(n432) );
  XOR U424 ( .A(n435), .B(n436), .Z(o[88]) );
  AND U425 ( .A(n401), .B(n437), .Z(n435) );
  XOR U426 ( .A(n438), .B(n439), .Z(o[87]) );
  AND U427 ( .A(n401), .B(n440), .Z(n438) );
  XOR U428 ( .A(n441), .B(n442), .Z(o[86]) );
  AND U429 ( .A(n401), .B(n443), .Z(n441) );
  XOR U430 ( .A(n444), .B(n445), .Z(o[85]) );
  AND U431 ( .A(n401), .B(n446), .Z(n444) );
  XOR U432 ( .A(n447), .B(n448), .Z(o[84]) );
  AND U433 ( .A(n401), .B(n449), .Z(n447) );
  XOR U434 ( .A(n450), .B(n451), .Z(o[83]) );
  AND U435 ( .A(n401), .B(n452), .Z(n450) );
  XOR U436 ( .A(n453), .B(n454), .Z(o[82]) );
  AND U437 ( .A(n401), .B(n455), .Z(n453) );
  XOR U438 ( .A(n456), .B(n457), .Z(o[81]) );
  AND U439 ( .A(n401), .B(n458), .Z(n456) );
  XOR U440 ( .A(n459), .B(n460), .Z(o[80]) );
  AND U441 ( .A(n401), .B(n461), .Z(n459) );
  XOR U442 ( .A(\min_val_reg[0][7] ), .B(n462), .Z(o[7]) );
  AND U443 ( .A(n397), .B(n463), .Z(n462) );
  XOR U444 ( .A(n464), .B(n465), .Z(o[79]) );
  AND U445 ( .A(n401), .B(n466), .Z(n464) );
  XOR U446 ( .A(n467), .B(n468), .Z(o[78]) );
  AND U447 ( .A(n401), .B(n469), .Z(n467) );
  XOR U448 ( .A(n470), .B(n471), .Z(o[77]) );
  AND U449 ( .A(n401), .B(n472), .Z(n470) );
  XOR U450 ( .A(n473), .B(n474), .Z(o[76]) );
  AND U451 ( .A(n401), .B(n475), .Z(n473) );
  XOR U452 ( .A(n476), .B(n477), .Z(o[75]) );
  AND U453 ( .A(n401), .B(n478), .Z(n476) );
  XOR U454 ( .A(n479), .B(n480), .Z(o[74]) );
  AND U455 ( .A(n401), .B(n481), .Z(n479) );
  XOR U456 ( .A(n482), .B(n483), .Z(o[73]) );
  AND U457 ( .A(n401), .B(n398), .Z(n482) );
  XOR U458 ( .A(\min_val_reg[0][9] ), .B(n483), .Z(n398) );
  XNOR U459 ( .A(n484), .B(\min_val_reg[1][9] ), .Z(n483) );
  NAND U460 ( .A(n485), .B(n486), .Z(n484) );
  XOR U461 ( .A(n487), .B(n488), .Z(o[72]) );
  AND U462 ( .A(n401), .B(n431), .Z(n487) );
  XOR U463 ( .A(\min_val_reg[0][8] ), .B(n488), .Z(n431) );
  XNOR U464 ( .A(n489), .B(\min_val_reg[1][8] ), .Z(n488) );
  NAND U465 ( .A(n490), .B(n486), .Z(n489) );
  XOR U466 ( .A(n491), .B(n492), .Z(o[71]) );
  AND U467 ( .A(n401), .B(n463), .Z(n491) );
  XOR U468 ( .A(\min_val_reg[0][7] ), .B(n492), .Z(n463) );
  XNOR U469 ( .A(n493), .B(\min_val_reg[1][7] ), .Z(n492) );
  NAND U470 ( .A(n494), .B(n486), .Z(n493) );
  XOR U471 ( .A(n495), .B(n496), .Z(o[70]) );
  AND U472 ( .A(n401), .B(n497), .Z(n495) );
  XOR U473 ( .A(\min_val_reg[0][6] ), .B(n498), .Z(o[6]) );
  AND U474 ( .A(n397), .B(n497), .Z(n498) );
  XOR U475 ( .A(\min_val_reg[0][6] ), .B(n496), .Z(n497) );
  XNOR U476 ( .A(n499), .B(\min_val_reg[1][6] ), .Z(n496) );
  NAND U477 ( .A(n500), .B(n486), .Z(n499) );
  XOR U478 ( .A(n501), .B(n502), .Z(o[69]) );
  AND U479 ( .A(n401), .B(n503), .Z(n501) );
  XOR U480 ( .A(n504), .B(n505), .Z(o[68]) );
  AND U481 ( .A(n401), .B(n506), .Z(n504) );
  XOR U482 ( .A(n507), .B(n508), .Z(o[67]) );
  AND U483 ( .A(n401), .B(n509), .Z(n507) );
  XOR U484 ( .A(n510), .B(n511), .Z(o[66]) );
  AND U485 ( .A(n401), .B(n512), .Z(n510) );
  XOR U486 ( .A(n513), .B(n514), .Z(o[65]) );
  AND U487 ( .A(n401), .B(n515), .Z(n513) );
  XOR U488 ( .A(n516), .B(n517), .Z(o[64]) );
  AND U489 ( .A(n401), .B(n518), .Z(n516) );
  XOR U490 ( .A(\min_val_reg[0][63] ), .B(n519), .Z(o[63]) );
  AND U491 ( .A(n397), .B(n520), .Z(n519) );
  XOR U492 ( .A(\min_val_reg[0][62] ), .B(n521), .Z(o[62]) );
  AND U493 ( .A(n397), .B(n522), .Z(n521) );
  XOR U494 ( .A(\min_val_reg[0][61] ), .B(n523), .Z(o[61]) );
  AND U495 ( .A(n397), .B(n524), .Z(n523) );
  XOR U496 ( .A(\min_val_reg[0][60] ), .B(n525), .Z(o[60]) );
  AND U497 ( .A(n397), .B(n526), .Z(n525) );
  XOR U498 ( .A(\min_val_reg[0][5] ), .B(n527), .Z(o[5]) );
  AND U499 ( .A(n397), .B(n503), .Z(n527) );
  XOR U500 ( .A(\min_val_reg[0][5] ), .B(n502), .Z(n503) );
  XNOR U501 ( .A(n528), .B(\min_val_reg[1][5] ), .Z(n502) );
  NAND U502 ( .A(n529), .B(n486), .Z(n528) );
  XOR U503 ( .A(\min_val_reg[0][59] ), .B(n530), .Z(o[59]) );
  AND U504 ( .A(n397), .B(n531), .Z(n530) );
  XOR U505 ( .A(\min_val_reg[0][58] ), .B(n532), .Z(o[58]) );
  AND U506 ( .A(n397), .B(n533), .Z(n532) );
  XOR U507 ( .A(\min_val_reg[0][57] ), .B(n534), .Z(o[57]) );
  AND U508 ( .A(n397), .B(n535), .Z(n534) );
  XOR U509 ( .A(\min_val_reg[0][56] ), .B(n536), .Z(o[56]) );
  AND U510 ( .A(n397), .B(n537), .Z(n536) );
  XOR U511 ( .A(\min_val_reg[0][55] ), .B(n538), .Z(o[55]) );
  AND U512 ( .A(n397), .B(n539), .Z(n538) );
  XOR U513 ( .A(\min_val_reg[0][54] ), .B(n540), .Z(o[54]) );
  AND U514 ( .A(n397), .B(n541), .Z(n540) );
  XOR U515 ( .A(\min_val_reg[0][53] ), .B(n542), .Z(o[53]) );
  AND U516 ( .A(n397), .B(n543), .Z(n542) );
  XOR U517 ( .A(\min_val_reg[0][52] ), .B(n544), .Z(o[52]) );
  AND U518 ( .A(n397), .B(n545), .Z(n544) );
  XOR U519 ( .A(\min_val_reg[0][51] ), .B(n546), .Z(o[51]) );
  AND U520 ( .A(n397), .B(n547), .Z(n546) );
  XOR U521 ( .A(\min_val_reg[0][50] ), .B(n548), .Z(o[50]) );
  AND U522 ( .A(n397), .B(n549), .Z(n548) );
  XOR U523 ( .A(\min_val_reg[0][4] ), .B(n550), .Z(o[4]) );
  AND U524 ( .A(n397), .B(n506), .Z(n550) );
  XOR U525 ( .A(\min_val_reg[0][4] ), .B(n505), .Z(n506) );
  XNOR U526 ( .A(n551), .B(\min_val_reg[1][4] ), .Z(n505) );
  NAND U527 ( .A(n552), .B(n486), .Z(n551) );
  XOR U528 ( .A(\min_val_reg[0][49] ), .B(n553), .Z(o[49]) );
  AND U529 ( .A(n397), .B(n554), .Z(n553) );
  XOR U530 ( .A(\min_val_reg[0][48] ), .B(n555), .Z(o[48]) );
  AND U531 ( .A(n397), .B(n556), .Z(n555) );
  XOR U532 ( .A(\min_val_reg[0][47] ), .B(n557), .Z(o[47]) );
  AND U533 ( .A(n397), .B(n558), .Z(n557) );
  XOR U534 ( .A(\min_val_reg[0][46] ), .B(n559), .Z(o[46]) );
  AND U535 ( .A(n397), .B(n560), .Z(n559) );
  XOR U536 ( .A(\min_val_reg[0][45] ), .B(n561), .Z(o[45]) );
  AND U537 ( .A(n397), .B(n562), .Z(n561) );
  XOR U538 ( .A(\min_val_reg[0][44] ), .B(n563), .Z(o[44]) );
  AND U539 ( .A(n397), .B(n564), .Z(n563) );
  XOR U540 ( .A(\min_val_reg[0][43] ), .B(n565), .Z(o[43]) );
  AND U541 ( .A(n397), .B(n566), .Z(n565) );
  XOR U542 ( .A(\min_val_reg[0][42] ), .B(n567), .Z(o[42]) );
  AND U543 ( .A(n397), .B(n568), .Z(n567) );
  XOR U544 ( .A(\min_val_reg[0][41] ), .B(n569), .Z(o[41]) );
  AND U545 ( .A(n397), .B(n570), .Z(n569) );
  XOR U546 ( .A(\min_val_reg[0][40] ), .B(n571), .Z(o[40]) );
  AND U547 ( .A(n397), .B(n572), .Z(n571) );
  XOR U548 ( .A(\min_val_reg[0][3] ), .B(n573), .Z(o[3]) );
  AND U549 ( .A(n397), .B(n509), .Z(n573) );
  XOR U550 ( .A(\min_val_reg[0][3] ), .B(n508), .Z(n509) );
  XNOR U551 ( .A(n574), .B(\min_val_reg[1][3] ), .Z(n508) );
  NAND U552 ( .A(n575), .B(n486), .Z(n574) );
  XOR U553 ( .A(\min_val_reg[0][39] ), .B(n576), .Z(o[39]) );
  AND U554 ( .A(n397), .B(n577), .Z(n576) );
  XOR U555 ( .A(\min_val_reg[0][38] ), .B(n578), .Z(o[38]) );
  AND U556 ( .A(n397), .B(n579), .Z(n578) );
  XOR U557 ( .A(\min_val_reg[0][37] ), .B(n580), .Z(o[37]) );
  AND U558 ( .A(n397), .B(n581), .Z(n580) );
  XOR U559 ( .A(\min_val_reg[0][36] ), .B(n582), .Z(o[36]) );
  AND U560 ( .A(n397), .B(n583), .Z(n582) );
  XOR U561 ( .A(\min_val_reg[0][35] ), .B(n584), .Z(o[35]) );
  AND U562 ( .A(n397), .B(n402), .Z(n584) );
  XOR U563 ( .A(\min_val_reg[0][35] ), .B(n400), .Z(n402) );
  XNOR U564 ( .A(n585), .B(\min_val_reg[1][35] ), .Z(n400) );
  NAND U565 ( .A(n586), .B(n486), .Z(n585) );
  XOR U566 ( .A(\min_val_reg[0][34] ), .B(n587), .Z(o[34]) );
  AND U567 ( .A(n397), .B(n405), .Z(n587) );
  XOR U568 ( .A(\min_val_reg[0][34] ), .B(n404), .Z(n405) );
  XNOR U569 ( .A(n588), .B(\min_val_reg[1][34] ), .Z(n404) );
  NAND U570 ( .A(n589), .B(n486), .Z(n588) );
  XOR U571 ( .A(\min_val_reg[0][33] ), .B(n590), .Z(o[33]) );
  AND U572 ( .A(n397), .B(n408), .Z(n590) );
  XOR U573 ( .A(\min_val_reg[0][33] ), .B(n407), .Z(n408) );
  XNOR U574 ( .A(n591), .B(\min_val_reg[1][33] ), .Z(n407) );
  NAND U575 ( .A(n592), .B(n486), .Z(n591) );
  XOR U576 ( .A(\min_val_reg[0][32] ), .B(n593), .Z(o[32]) );
  AND U577 ( .A(n397), .B(n411), .Z(n593) );
  XOR U578 ( .A(\min_val_reg[0][32] ), .B(n410), .Z(n411) );
  XNOR U579 ( .A(n594), .B(\min_val_reg[1][32] ), .Z(n410) );
  NAND U580 ( .A(n595), .B(n486), .Z(n594) );
  XOR U581 ( .A(\min_val_reg[0][31] ), .B(n596), .Z(o[31]) );
  AND U582 ( .A(n397), .B(n414), .Z(n596) );
  XOR U583 ( .A(\min_val_reg[0][31] ), .B(n413), .Z(n414) );
  XNOR U584 ( .A(n597), .B(\min_val_reg[1][31] ), .Z(n413) );
  NAND U585 ( .A(n598), .B(n486), .Z(n597) );
  XOR U586 ( .A(\min_val_reg[0][30] ), .B(n599), .Z(o[30]) );
  AND U587 ( .A(n397), .B(n417), .Z(n599) );
  XOR U588 ( .A(\min_val_reg[0][30] ), .B(n416), .Z(n417) );
  XNOR U589 ( .A(n600), .B(\min_val_reg[1][30] ), .Z(n416) );
  NAND U590 ( .A(n601), .B(n486), .Z(n600) );
  XOR U591 ( .A(\min_val_reg[0][2] ), .B(n602), .Z(o[2]) );
  AND U592 ( .A(n397), .B(n512), .Z(n602) );
  XOR U593 ( .A(\min_val_reg[0][2] ), .B(n511), .Z(n512) );
  XNOR U594 ( .A(n603), .B(\min_val_reg[1][2] ), .Z(n511) );
  NAND U595 ( .A(n604), .B(n486), .Z(n603) );
  XOR U596 ( .A(\min_val_reg[0][29] ), .B(n605), .Z(o[29]) );
  AND U597 ( .A(n397), .B(n420), .Z(n605) );
  XOR U598 ( .A(\min_val_reg[0][29] ), .B(n419), .Z(n420) );
  XNOR U599 ( .A(n606), .B(\min_val_reg[1][29] ), .Z(n419) );
  NAND U600 ( .A(n607), .B(n486), .Z(n606) );
  XOR U601 ( .A(\min_val_reg[0][28] ), .B(n608), .Z(o[28]) );
  AND U602 ( .A(n397), .B(n423), .Z(n608) );
  XOR U603 ( .A(\min_val_reg[0][28] ), .B(n422), .Z(n423) );
  XNOR U604 ( .A(n609), .B(\min_val_reg[1][28] ), .Z(n422) );
  NAND U605 ( .A(n610), .B(n486), .Z(n609) );
  XOR U606 ( .A(\min_val_reg[0][27] ), .B(n611), .Z(o[27]) );
  AND U607 ( .A(n397), .B(n426), .Z(n611) );
  XOR U608 ( .A(\min_val_reg[0][27] ), .B(n425), .Z(n426) );
  XNOR U609 ( .A(n612), .B(\min_val_reg[1][27] ), .Z(n425) );
  NAND U610 ( .A(n613), .B(n486), .Z(n612) );
  XOR U611 ( .A(\min_val_reg[0][26] ), .B(n614), .Z(o[26]) );
  AND U612 ( .A(n397), .B(n429), .Z(n614) );
  XOR U613 ( .A(\min_val_reg[0][26] ), .B(n428), .Z(n429) );
  XNOR U614 ( .A(n615), .B(\min_val_reg[1][26] ), .Z(n428) );
  NAND U615 ( .A(n616), .B(n486), .Z(n615) );
  XOR U616 ( .A(\min_val_reg[0][25] ), .B(n617), .Z(o[25]) );
  AND U617 ( .A(n397), .B(n434), .Z(n617) );
  XOR U618 ( .A(\min_val_reg[0][25] ), .B(n433), .Z(n434) );
  XNOR U619 ( .A(n618), .B(\min_val_reg[1][25] ), .Z(n433) );
  NAND U620 ( .A(n619), .B(n486), .Z(n618) );
  XNOR U621 ( .A(n620), .B(n621), .Z(o[255]) );
  AND U622 ( .A(n622), .B(n623), .Z(n620) );
  XNOR U623 ( .A(n624), .B(n625), .Z(o[254]) );
  AND U624 ( .A(n622), .B(n626), .Z(n624) );
  XNOR U625 ( .A(n627), .B(n628), .Z(o[253]) );
  AND U626 ( .A(n622), .B(n629), .Z(n627) );
  XNOR U627 ( .A(n630), .B(n631), .Z(o[252]) );
  AND U628 ( .A(n622), .B(n632), .Z(n630) );
  XNOR U629 ( .A(n633), .B(n634), .Z(o[251]) );
  AND U630 ( .A(n622), .B(n635), .Z(n633) );
  XNOR U631 ( .A(n636), .B(n637), .Z(o[250]) );
  AND U632 ( .A(n622), .B(n638), .Z(n636) );
  XOR U633 ( .A(\min_val_reg[0][24] ), .B(n639), .Z(o[24]) );
  AND U634 ( .A(n397), .B(n437), .Z(n639) );
  XOR U635 ( .A(\min_val_reg[0][24] ), .B(n436), .Z(n437) );
  XNOR U636 ( .A(n640), .B(\min_val_reg[1][24] ), .Z(n436) );
  NAND U637 ( .A(n641), .B(n486), .Z(n640) );
  XNOR U638 ( .A(n642), .B(n643), .Z(o[249]) );
  AND U639 ( .A(n622), .B(n644), .Z(n642) );
  XNOR U640 ( .A(n645), .B(n646), .Z(o[248]) );
  AND U641 ( .A(n622), .B(n647), .Z(n645) );
  XNOR U642 ( .A(n648), .B(n649), .Z(o[247]) );
  AND U643 ( .A(n622), .B(n650), .Z(n648) );
  XNOR U644 ( .A(n651), .B(n652), .Z(o[246]) );
  AND U645 ( .A(n622), .B(n653), .Z(n651) );
  XNOR U646 ( .A(n654), .B(n655), .Z(o[245]) );
  AND U647 ( .A(n622), .B(n656), .Z(n654) );
  XNOR U648 ( .A(n657), .B(n658), .Z(o[244]) );
  AND U649 ( .A(n622), .B(n659), .Z(n657) );
  XNOR U650 ( .A(n660), .B(n661), .Z(o[243]) );
  AND U651 ( .A(n622), .B(n662), .Z(n660) );
  XNOR U652 ( .A(n663), .B(n664), .Z(o[242]) );
  AND U653 ( .A(n622), .B(n665), .Z(n663) );
  XNOR U654 ( .A(n666), .B(n667), .Z(o[241]) );
  AND U655 ( .A(n622), .B(n668), .Z(n666) );
  XNOR U656 ( .A(n669), .B(n670), .Z(o[240]) );
  AND U657 ( .A(n622), .B(n671), .Z(n669) );
  XOR U658 ( .A(\min_val_reg[0][23] ), .B(n672), .Z(o[23]) );
  AND U659 ( .A(n397), .B(n440), .Z(n672) );
  XOR U660 ( .A(\min_val_reg[0][23] ), .B(n439), .Z(n440) );
  XNOR U661 ( .A(n673), .B(\min_val_reg[1][23] ), .Z(n439) );
  NAND U662 ( .A(n674), .B(n486), .Z(n673) );
  XNOR U663 ( .A(n675), .B(n676), .Z(o[239]) );
  AND U664 ( .A(n622), .B(n677), .Z(n675) );
  XNOR U665 ( .A(n678), .B(n679), .Z(o[238]) );
  AND U666 ( .A(n622), .B(n680), .Z(n678) );
  XNOR U667 ( .A(n681), .B(n682), .Z(o[237]) );
  AND U668 ( .A(n622), .B(n683), .Z(n681) );
  XNOR U669 ( .A(n684), .B(n685), .Z(o[236]) );
  AND U670 ( .A(n622), .B(n686), .Z(n684) );
  XNOR U671 ( .A(n687), .B(n688), .Z(o[235]) );
  AND U672 ( .A(n622), .B(n689), .Z(n687) );
  XNOR U673 ( .A(n690), .B(n691), .Z(o[234]) );
  AND U674 ( .A(n622), .B(n692), .Z(n690) );
  XNOR U675 ( .A(n693), .B(n694), .Z(o[233]) );
  AND U676 ( .A(n622), .B(n695), .Z(n693) );
  XNOR U677 ( .A(n696), .B(n697), .Z(o[232]) );
  AND U678 ( .A(n622), .B(n698), .Z(n696) );
  XNOR U679 ( .A(n699), .B(n700), .Z(o[231]) );
  AND U680 ( .A(n622), .B(n701), .Z(n699) );
  XNOR U681 ( .A(n702), .B(n703), .Z(o[230]) );
  AND U682 ( .A(n622), .B(n704), .Z(n702) );
  XOR U683 ( .A(\min_val_reg[0][22] ), .B(n705), .Z(o[22]) );
  AND U684 ( .A(n397), .B(n443), .Z(n705) );
  XOR U685 ( .A(\min_val_reg[0][22] ), .B(n442), .Z(n443) );
  XNOR U686 ( .A(n706), .B(\min_val_reg[1][22] ), .Z(n442) );
  NAND U687 ( .A(n707), .B(n486), .Z(n706) );
  XNOR U688 ( .A(n708), .B(n709), .Z(o[229]) );
  AND U689 ( .A(n622), .B(n710), .Z(n708) );
  XNOR U690 ( .A(n711), .B(n712), .Z(o[228]) );
  AND U691 ( .A(n622), .B(n713), .Z(n711) );
  XNOR U692 ( .A(n714), .B(n715), .Z(o[227]) );
  AND U693 ( .A(n622), .B(n716), .Z(n714) );
  XNOR U694 ( .A(n717), .B(n718), .Z(o[226]) );
  AND U695 ( .A(n622), .B(n719), .Z(n717) );
  XNOR U696 ( .A(n720), .B(n721), .Z(o[225]) );
  AND U697 ( .A(n622), .B(n722), .Z(n720) );
  XNOR U698 ( .A(n723), .B(n724), .Z(o[224]) );
  AND U699 ( .A(n622), .B(n725), .Z(n723) );
  XNOR U700 ( .A(n726), .B(n727), .Z(o[223]) );
  AND U701 ( .A(n622), .B(n728), .Z(n726) );
  XNOR U702 ( .A(n729), .B(n730), .Z(o[222]) );
  AND U703 ( .A(n622), .B(n731), .Z(n729) );
  XNOR U704 ( .A(n732), .B(n733), .Z(o[221]) );
  AND U705 ( .A(n622), .B(n734), .Z(n732) );
  XNOR U706 ( .A(n735), .B(n736), .Z(o[220]) );
  AND U707 ( .A(n622), .B(n737), .Z(n735) );
  XOR U708 ( .A(\min_val_reg[0][21] ), .B(n738), .Z(o[21]) );
  AND U709 ( .A(n397), .B(n446), .Z(n738) );
  XOR U710 ( .A(\min_val_reg[0][21] ), .B(n445), .Z(n446) );
  XNOR U711 ( .A(n739), .B(\min_val_reg[1][21] ), .Z(n445) );
  NAND U712 ( .A(n740), .B(n486), .Z(n739) );
  XNOR U713 ( .A(n741), .B(n742), .Z(o[219]) );
  AND U714 ( .A(n622), .B(n743), .Z(n741) );
  XNOR U715 ( .A(n744), .B(n745), .Z(o[218]) );
  AND U716 ( .A(n622), .B(n746), .Z(n744) );
  XNOR U717 ( .A(n747), .B(n748), .Z(o[217]) );
  AND U718 ( .A(n622), .B(n749), .Z(n747) );
  XNOR U719 ( .A(n750), .B(n751), .Z(o[216]) );
  AND U720 ( .A(n622), .B(n752), .Z(n750) );
  XNOR U721 ( .A(n753), .B(n754), .Z(o[215]) );
  AND U722 ( .A(n622), .B(n755), .Z(n753) );
  XNOR U723 ( .A(n756), .B(n757), .Z(o[214]) );
  AND U724 ( .A(n622), .B(n758), .Z(n756) );
  XNOR U725 ( .A(n759), .B(n760), .Z(o[213]) );
  AND U726 ( .A(n622), .B(n761), .Z(n759) );
  XNOR U727 ( .A(n762), .B(n763), .Z(o[212]) );
  AND U728 ( .A(n622), .B(n764), .Z(n762) );
  XNOR U729 ( .A(n765), .B(n766), .Z(o[211]) );
  AND U730 ( .A(n622), .B(n767), .Z(n765) );
  XNOR U731 ( .A(n768), .B(n769), .Z(o[210]) );
  AND U732 ( .A(n622), .B(n770), .Z(n768) );
  XOR U733 ( .A(\min_val_reg[0][20] ), .B(n771), .Z(o[20]) );
  AND U734 ( .A(n397), .B(n449), .Z(n771) );
  XOR U735 ( .A(\min_val_reg[0][20] ), .B(n448), .Z(n449) );
  XNOR U736 ( .A(n772), .B(\min_val_reg[1][20] ), .Z(n448) );
  NAND U737 ( .A(n773), .B(n486), .Z(n772) );
  XNOR U738 ( .A(n774), .B(n775), .Z(o[209]) );
  AND U739 ( .A(n622), .B(n776), .Z(n774) );
  XNOR U740 ( .A(n777), .B(n778), .Z(o[208]) );
  AND U741 ( .A(n622), .B(n779), .Z(n777) );
  XNOR U742 ( .A(n780), .B(n781), .Z(o[207]) );
  AND U743 ( .A(n622), .B(n782), .Z(n780) );
  XNOR U744 ( .A(n783), .B(n784), .Z(o[206]) );
  AND U745 ( .A(n622), .B(n785), .Z(n783) );
  XNOR U746 ( .A(n786), .B(n787), .Z(o[205]) );
  AND U747 ( .A(n622), .B(n788), .Z(n786) );
  XNOR U748 ( .A(n789), .B(n790), .Z(o[204]) );
  AND U749 ( .A(n622), .B(n791), .Z(n789) );
  XNOR U750 ( .A(n792), .B(n793), .Z(o[203]) );
  AND U751 ( .A(n622), .B(n794), .Z(n792) );
  XNOR U752 ( .A(n795), .B(n796), .Z(o[202]) );
  AND U753 ( .A(n622), .B(n797), .Z(n795) );
  XNOR U754 ( .A(n798), .B(n799), .Z(o[201]) );
  AND U755 ( .A(n622), .B(n800), .Z(n798) );
  XNOR U756 ( .A(n801), .B(n802), .Z(o[200]) );
  AND U757 ( .A(n622), .B(n803), .Z(n801) );
  XOR U758 ( .A(\min_val_reg[0][1] ), .B(n804), .Z(o[1]) );
  AND U759 ( .A(n397), .B(n515), .Z(n804) );
  XOR U760 ( .A(\min_val_reg[0][1] ), .B(n514), .Z(n515) );
  XNOR U761 ( .A(n805), .B(\min_val_reg[1][1] ), .Z(n514) );
  NAND U762 ( .A(n806), .B(n486), .Z(n805) );
  XOR U763 ( .A(\min_val_reg[0][19] ), .B(n807), .Z(o[19]) );
  AND U764 ( .A(n397), .B(n452), .Z(n807) );
  XOR U765 ( .A(\min_val_reg[0][19] ), .B(n451), .Z(n452) );
  XNOR U766 ( .A(n808), .B(\min_val_reg[1][19] ), .Z(n451) );
  NAND U767 ( .A(n809), .B(n486), .Z(n808) );
  XNOR U768 ( .A(n810), .B(n811), .Z(o[199]) );
  AND U769 ( .A(n622), .B(n812), .Z(n810) );
  XNOR U770 ( .A(n813), .B(n814), .Z(o[198]) );
  AND U771 ( .A(n622), .B(n815), .Z(n813) );
  XNOR U772 ( .A(n816), .B(n817), .Z(o[197]) );
  AND U773 ( .A(n622), .B(n818), .Z(n816) );
  XNOR U774 ( .A(n819), .B(n820), .Z(o[196]) );
  AND U775 ( .A(n622), .B(n821), .Z(n819) );
  XNOR U776 ( .A(n822), .B(n823), .Z(o[195]) );
  AND U777 ( .A(n622), .B(n824), .Z(n822) );
  XNOR U778 ( .A(n825), .B(n826), .Z(o[194]) );
  AND U779 ( .A(n622), .B(n827), .Z(n825) );
  XNOR U780 ( .A(n828), .B(n829), .Z(o[193]) );
  AND U781 ( .A(n622), .B(n830), .Z(n828) );
  XNOR U782 ( .A(n831), .B(n832), .Z(o[192]) );
  AND U783 ( .A(n622), .B(n833), .Z(n831) );
  XOR U784 ( .A(n834), .B(n835), .Z(o[191]) );
  AND U785 ( .A(n486), .B(n836), .Z(n834) );
  XOR U786 ( .A(n837), .B(n838), .Z(o[190]) );
  AND U787 ( .A(n486), .B(n839), .Z(n837) );
  XOR U788 ( .A(\min_val_reg[0][18] ), .B(n840), .Z(o[18]) );
  AND U789 ( .A(n397), .B(n455), .Z(n840) );
  XOR U790 ( .A(\min_val_reg[0][18] ), .B(n454), .Z(n455) );
  XNOR U791 ( .A(n841), .B(\min_val_reg[1][18] ), .Z(n454) );
  NAND U792 ( .A(n842), .B(n486), .Z(n841) );
  XOR U793 ( .A(n843), .B(n844), .Z(o[189]) );
  AND U794 ( .A(n486), .B(n845), .Z(n843) );
  XOR U795 ( .A(n846), .B(n847), .Z(o[188]) );
  AND U796 ( .A(n486), .B(n848), .Z(n846) );
  XOR U797 ( .A(n849), .B(n850), .Z(o[187]) );
  AND U798 ( .A(n486), .B(n851), .Z(n849) );
  XOR U799 ( .A(n852), .B(n853), .Z(o[186]) );
  AND U800 ( .A(n486), .B(n854), .Z(n852) );
  XOR U801 ( .A(n855), .B(n856), .Z(o[185]) );
  AND U802 ( .A(n486), .B(n857), .Z(n855) );
  XOR U803 ( .A(n858), .B(n859), .Z(o[184]) );
  AND U804 ( .A(n486), .B(n860), .Z(n858) );
  XOR U805 ( .A(n861), .B(n862), .Z(o[183]) );
  AND U806 ( .A(n486), .B(n863), .Z(n861) );
  XOR U807 ( .A(n864), .B(n865), .Z(o[182]) );
  AND U808 ( .A(n486), .B(n866), .Z(n864) );
  XOR U809 ( .A(n867), .B(n868), .Z(o[181]) );
  AND U810 ( .A(n486), .B(n869), .Z(n867) );
  XOR U811 ( .A(n870), .B(n871), .Z(o[180]) );
  AND U812 ( .A(n486), .B(n872), .Z(n870) );
  XOR U813 ( .A(\min_val_reg[0][17] ), .B(n873), .Z(o[17]) );
  AND U814 ( .A(n397), .B(n458), .Z(n873) );
  XOR U815 ( .A(\min_val_reg[0][17] ), .B(n457), .Z(n458) );
  XNOR U816 ( .A(n874), .B(\min_val_reg[1][17] ), .Z(n457) );
  NAND U817 ( .A(n875), .B(n486), .Z(n874) );
  XOR U818 ( .A(n876), .B(n877), .Z(o[179]) );
  AND U819 ( .A(n486), .B(n878), .Z(n876) );
  XOR U820 ( .A(n879), .B(n880), .Z(o[178]) );
  AND U821 ( .A(n486), .B(n881), .Z(n879) );
  XOR U822 ( .A(n882), .B(n883), .Z(o[177]) );
  AND U823 ( .A(n486), .B(n884), .Z(n882) );
  XOR U824 ( .A(n885), .B(n886), .Z(o[176]) );
  AND U825 ( .A(n486), .B(n887), .Z(n885) );
  XOR U826 ( .A(n888), .B(n889), .Z(o[175]) );
  AND U827 ( .A(n486), .B(n890), .Z(n888) );
  XOR U828 ( .A(n891), .B(n892), .Z(o[174]) );
  AND U829 ( .A(n486), .B(n893), .Z(n891) );
  XOR U830 ( .A(n894), .B(n895), .Z(o[173]) );
  AND U831 ( .A(n486), .B(n896), .Z(n894) );
  XOR U832 ( .A(n897), .B(n898), .Z(o[172]) );
  AND U833 ( .A(n486), .B(n899), .Z(n897) );
  XOR U834 ( .A(n900), .B(n901), .Z(o[171]) );
  AND U835 ( .A(n486), .B(n902), .Z(n900) );
  XOR U836 ( .A(n903), .B(n904), .Z(o[170]) );
  AND U837 ( .A(n486), .B(n905), .Z(n903) );
  XOR U838 ( .A(\min_val_reg[0][16] ), .B(n906), .Z(o[16]) );
  AND U839 ( .A(n397), .B(n461), .Z(n906) );
  XOR U840 ( .A(\min_val_reg[0][16] ), .B(n460), .Z(n461) );
  XNOR U841 ( .A(n907), .B(\min_val_reg[1][16] ), .Z(n460) );
  NAND U842 ( .A(n908), .B(n486), .Z(n907) );
  XOR U843 ( .A(n909), .B(n910), .Z(o[169]) );
  AND U844 ( .A(n486), .B(n911), .Z(n909) );
  XOR U845 ( .A(n912), .B(n913), .Z(o[168]) );
  AND U846 ( .A(n486), .B(n914), .Z(n912) );
  XOR U847 ( .A(n915), .B(n916), .Z(o[167]) );
  AND U848 ( .A(n486), .B(n917), .Z(n915) );
  XOR U849 ( .A(n918), .B(n919), .Z(o[166]) );
  AND U850 ( .A(n486), .B(n920), .Z(n918) );
  XOR U851 ( .A(n921), .B(n922), .Z(o[165]) );
  AND U852 ( .A(n486), .B(n923), .Z(n921) );
  XOR U853 ( .A(n924), .B(n925), .Z(o[164]) );
  AND U854 ( .A(n486), .B(n926), .Z(n924) );
  XOR U855 ( .A(n927), .B(n928), .Z(o[163]) );
  AND U856 ( .A(n486), .B(n586), .Z(n927) );
  XOR U857 ( .A(\min_val_reg[1][35] ), .B(n928), .Z(n586) );
  XNOR U858 ( .A(n929), .B(\min_val_reg[2][35] ), .Z(n928) );
  NAND U859 ( .A(n716), .B(n930), .Z(n929) );
  XNOR U860 ( .A(\min_val_reg[2][35] ), .B(n715), .Z(n716) );
  XOR U861 ( .A(n931), .B(\min_val_reg[3][35] ), .Z(n715) );
  NAND U862 ( .A(n932), .B(n933), .Z(n931) );
  XOR U863 ( .A(\min_val_reg[3][35] ), .B(g_input[35]), .Z(n932) );
  XOR U864 ( .A(n934), .B(n935), .Z(o[162]) );
  AND U865 ( .A(n486), .B(n589), .Z(n934) );
  XOR U866 ( .A(\min_val_reg[1][34] ), .B(n935), .Z(n589) );
  XNOR U867 ( .A(n936), .B(\min_val_reg[2][34] ), .Z(n935) );
  NAND U868 ( .A(n719), .B(n930), .Z(n936) );
  XNOR U869 ( .A(\min_val_reg[2][34] ), .B(n718), .Z(n719) );
  XOR U870 ( .A(n937), .B(\min_val_reg[3][34] ), .Z(n718) );
  NAND U871 ( .A(n938), .B(n933), .Z(n937) );
  XOR U872 ( .A(\min_val_reg[3][34] ), .B(g_input[34]), .Z(n938) );
  XOR U873 ( .A(n939), .B(n940), .Z(o[161]) );
  AND U874 ( .A(n486), .B(n592), .Z(n939) );
  XOR U875 ( .A(\min_val_reg[1][33] ), .B(n940), .Z(n592) );
  XNOR U876 ( .A(n941), .B(\min_val_reg[2][33] ), .Z(n940) );
  NAND U877 ( .A(n722), .B(n930), .Z(n941) );
  XNOR U878 ( .A(\min_val_reg[2][33] ), .B(n721), .Z(n722) );
  XOR U879 ( .A(n942), .B(\min_val_reg[3][33] ), .Z(n721) );
  NAND U880 ( .A(n943), .B(n933), .Z(n942) );
  XOR U881 ( .A(\min_val_reg[3][33] ), .B(g_input[33]), .Z(n943) );
  XOR U882 ( .A(n944), .B(n945), .Z(o[160]) );
  AND U883 ( .A(n486), .B(n595), .Z(n944) );
  XOR U884 ( .A(\min_val_reg[1][32] ), .B(n945), .Z(n595) );
  XNOR U885 ( .A(n946), .B(\min_val_reg[2][32] ), .Z(n945) );
  NAND U886 ( .A(n725), .B(n930), .Z(n946) );
  XNOR U887 ( .A(\min_val_reg[2][32] ), .B(n724), .Z(n725) );
  XOR U888 ( .A(n947), .B(\min_val_reg[3][32] ), .Z(n724) );
  NAND U889 ( .A(n948), .B(n933), .Z(n947) );
  XNOR U890 ( .A(\min_val_reg[3][32] ), .B(n949), .Z(n948) );
  XOR U891 ( .A(\min_val_reg[0][15] ), .B(n950), .Z(o[15]) );
  AND U892 ( .A(n397), .B(n466), .Z(n950) );
  XOR U893 ( .A(\min_val_reg[0][15] ), .B(n465), .Z(n466) );
  XNOR U894 ( .A(n951), .B(\min_val_reg[1][15] ), .Z(n465) );
  NAND U895 ( .A(n952), .B(n486), .Z(n951) );
  XOR U896 ( .A(n953), .B(n954), .Z(o[159]) );
  AND U897 ( .A(n486), .B(n598), .Z(n953) );
  XOR U898 ( .A(\min_val_reg[1][31] ), .B(n954), .Z(n598) );
  XNOR U899 ( .A(n955), .B(\min_val_reg[2][31] ), .Z(n954) );
  NAND U900 ( .A(n728), .B(n930), .Z(n955) );
  XNOR U901 ( .A(\min_val_reg[2][31] ), .B(n727), .Z(n728) );
  XOR U902 ( .A(n956), .B(\min_val_reg[3][31] ), .Z(n727) );
  NAND U903 ( .A(n957), .B(n933), .Z(n956) );
  XOR U904 ( .A(\min_val_reg[3][31] ), .B(g_input[31]), .Z(n957) );
  XOR U905 ( .A(n958), .B(n959), .Z(o[158]) );
  AND U906 ( .A(n486), .B(n601), .Z(n958) );
  XOR U907 ( .A(\min_val_reg[1][30] ), .B(n959), .Z(n601) );
  XNOR U908 ( .A(n960), .B(\min_val_reg[2][30] ), .Z(n959) );
  NAND U909 ( .A(n731), .B(n930), .Z(n960) );
  XNOR U910 ( .A(\min_val_reg[2][30] ), .B(n730), .Z(n731) );
  XOR U911 ( .A(n961), .B(\min_val_reg[3][30] ), .Z(n730) );
  NAND U912 ( .A(n962), .B(n933), .Z(n961) );
  XOR U913 ( .A(\min_val_reg[3][30] ), .B(g_input[30]), .Z(n962) );
  XOR U914 ( .A(n963), .B(n964), .Z(o[157]) );
  AND U915 ( .A(n486), .B(n607), .Z(n963) );
  XOR U916 ( .A(\min_val_reg[1][29] ), .B(n964), .Z(n607) );
  XNOR U917 ( .A(n965), .B(\min_val_reg[2][29] ), .Z(n964) );
  NAND U918 ( .A(n734), .B(n930), .Z(n965) );
  XNOR U919 ( .A(\min_val_reg[2][29] ), .B(n733), .Z(n734) );
  XOR U920 ( .A(n966), .B(\min_val_reg[3][29] ), .Z(n733) );
  NAND U921 ( .A(n967), .B(n933), .Z(n966) );
  XOR U922 ( .A(\min_val_reg[3][29] ), .B(g_input[29]), .Z(n967) );
  XOR U923 ( .A(n968), .B(n969), .Z(o[156]) );
  AND U924 ( .A(n486), .B(n610), .Z(n968) );
  XOR U925 ( .A(\min_val_reg[1][28] ), .B(n969), .Z(n610) );
  XNOR U926 ( .A(n970), .B(\min_val_reg[2][28] ), .Z(n969) );
  NAND U927 ( .A(n737), .B(n930), .Z(n970) );
  XNOR U928 ( .A(\min_val_reg[2][28] ), .B(n736), .Z(n737) );
  XOR U929 ( .A(n971), .B(\min_val_reg[3][28] ), .Z(n736) );
  NAND U930 ( .A(n972), .B(n933), .Z(n971) );
  XOR U931 ( .A(\min_val_reg[3][28] ), .B(g_input[28]), .Z(n972) );
  XOR U932 ( .A(n973), .B(n974), .Z(o[155]) );
  AND U933 ( .A(n486), .B(n613), .Z(n973) );
  XOR U934 ( .A(\min_val_reg[1][27] ), .B(n974), .Z(n613) );
  XNOR U935 ( .A(n975), .B(\min_val_reg[2][27] ), .Z(n974) );
  NAND U936 ( .A(n743), .B(n930), .Z(n975) );
  XNOR U937 ( .A(\min_val_reg[2][27] ), .B(n742), .Z(n743) );
  XOR U938 ( .A(n976), .B(\min_val_reg[3][27] ), .Z(n742) );
  NAND U939 ( .A(n977), .B(n933), .Z(n976) );
  XOR U940 ( .A(\min_val_reg[3][27] ), .B(g_input[27]), .Z(n977) );
  XOR U941 ( .A(n978), .B(n979), .Z(o[154]) );
  AND U942 ( .A(n486), .B(n616), .Z(n978) );
  XOR U943 ( .A(\min_val_reg[1][26] ), .B(n979), .Z(n616) );
  XNOR U944 ( .A(n980), .B(\min_val_reg[2][26] ), .Z(n979) );
  NAND U945 ( .A(n746), .B(n930), .Z(n980) );
  XNOR U946 ( .A(\min_val_reg[2][26] ), .B(n745), .Z(n746) );
  XOR U947 ( .A(n981), .B(\min_val_reg[3][26] ), .Z(n745) );
  NAND U948 ( .A(n982), .B(n933), .Z(n981) );
  XOR U949 ( .A(\min_val_reg[3][26] ), .B(g_input[26]), .Z(n982) );
  XOR U950 ( .A(n983), .B(n984), .Z(o[153]) );
  AND U951 ( .A(n486), .B(n619), .Z(n983) );
  XOR U952 ( .A(\min_val_reg[1][25] ), .B(n984), .Z(n619) );
  XNOR U953 ( .A(n985), .B(\min_val_reg[2][25] ), .Z(n984) );
  NAND U954 ( .A(n749), .B(n930), .Z(n985) );
  XNOR U955 ( .A(\min_val_reg[2][25] ), .B(n748), .Z(n749) );
  XOR U956 ( .A(n986), .B(\min_val_reg[3][25] ), .Z(n748) );
  NAND U957 ( .A(n987), .B(n933), .Z(n986) );
  XOR U958 ( .A(\min_val_reg[3][25] ), .B(g_input[25]), .Z(n987) );
  XOR U959 ( .A(n988), .B(n989), .Z(o[152]) );
  AND U960 ( .A(n486), .B(n641), .Z(n988) );
  XOR U961 ( .A(\min_val_reg[1][24] ), .B(n989), .Z(n641) );
  XNOR U962 ( .A(n990), .B(\min_val_reg[2][24] ), .Z(n989) );
  NAND U963 ( .A(n752), .B(n930), .Z(n990) );
  XNOR U964 ( .A(\min_val_reg[2][24] ), .B(n751), .Z(n752) );
  XOR U965 ( .A(n991), .B(\min_val_reg[3][24] ), .Z(n751) );
  NAND U966 ( .A(n992), .B(n933), .Z(n991) );
  XOR U967 ( .A(\min_val_reg[3][24] ), .B(g_input[24]), .Z(n992) );
  XOR U968 ( .A(n993), .B(n994), .Z(o[151]) );
  AND U969 ( .A(n486), .B(n674), .Z(n993) );
  XOR U970 ( .A(\min_val_reg[1][23] ), .B(n994), .Z(n674) );
  XNOR U971 ( .A(n995), .B(\min_val_reg[2][23] ), .Z(n994) );
  NAND U972 ( .A(n755), .B(n930), .Z(n995) );
  XNOR U973 ( .A(\min_val_reg[2][23] ), .B(n754), .Z(n755) );
  XOR U974 ( .A(n996), .B(\min_val_reg[3][23] ), .Z(n754) );
  NAND U975 ( .A(n997), .B(n933), .Z(n996) );
  XOR U976 ( .A(\min_val_reg[3][23] ), .B(g_input[23]), .Z(n997) );
  XOR U977 ( .A(n998), .B(n999), .Z(o[150]) );
  AND U978 ( .A(n486), .B(n707), .Z(n998) );
  XOR U979 ( .A(\min_val_reg[1][22] ), .B(n999), .Z(n707) );
  XNOR U980 ( .A(n1000), .B(\min_val_reg[2][22] ), .Z(n999) );
  NAND U981 ( .A(n758), .B(n930), .Z(n1000) );
  XNOR U982 ( .A(\min_val_reg[2][22] ), .B(n757), .Z(n758) );
  XOR U983 ( .A(n1001), .B(\min_val_reg[3][22] ), .Z(n757) );
  NAND U984 ( .A(n1002), .B(n933), .Z(n1001) );
  XOR U985 ( .A(\min_val_reg[3][22] ), .B(g_input[22]), .Z(n1002) );
  XOR U986 ( .A(\min_val_reg[0][14] ), .B(n1003), .Z(o[14]) );
  AND U987 ( .A(n397), .B(n469), .Z(n1003) );
  XOR U988 ( .A(\min_val_reg[0][14] ), .B(n468), .Z(n469) );
  XNOR U989 ( .A(n1004), .B(\min_val_reg[1][14] ), .Z(n468) );
  NAND U990 ( .A(n1005), .B(n486), .Z(n1004) );
  XOR U991 ( .A(n1006), .B(n1007), .Z(o[149]) );
  AND U992 ( .A(n486), .B(n740), .Z(n1006) );
  XOR U993 ( .A(\min_val_reg[1][21] ), .B(n1007), .Z(n740) );
  XNOR U994 ( .A(n1008), .B(\min_val_reg[2][21] ), .Z(n1007) );
  NAND U995 ( .A(n761), .B(n930), .Z(n1008) );
  XNOR U996 ( .A(\min_val_reg[2][21] ), .B(n760), .Z(n761) );
  XOR U997 ( .A(n1009), .B(\min_val_reg[3][21] ), .Z(n760) );
  NAND U998 ( .A(n1010), .B(n933), .Z(n1009) );
  XOR U999 ( .A(\min_val_reg[3][21] ), .B(g_input[21]), .Z(n1010) );
  XOR U1000 ( .A(n1011), .B(n1012), .Z(o[148]) );
  AND U1001 ( .A(n486), .B(n773), .Z(n1011) );
  XOR U1002 ( .A(\min_val_reg[1][20] ), .B(n1012), .Z(n773) );
  XNOR U1003 ( .A(n1013), .B(\min_val_reg[2][20] ), .Z(n1012) );
  NAND U1004 ( .A(n764), .B(n930), .Z(n1013) );
  XNOR U1005 ( .A(\min_val_reg[2][20] ), .B(n763), .Z(n764) );
  XOR U1006 ( .A(n1014), .B(\min_val_reg[3][20] ), .Z(n763) );
  NAND U1007 ( .A(n1015), .B(n933), .Z(n1014) );
  XOR U1008 ( .A(\min_val_reg[3][20] ), .B(g_input[20]), .Z(n1015) );
  XOR U1009 ( .A(n1016), .B(n1017), .Z(o[147]) );
  AND U1010 ( .A(n486), .B(n809), .Z(n1016) );
  XOR U1011 ( .A(\min_val_reg[1][19] ), .B(n1017), .Z(n809) );
  XNOR U1012 ( .A(n1018), .B(\min_val_reg[2][19] ), .Z(n1017) );
  NAND U1013 ( .A(n767), .B(n930), .Z(n1018) );
  XNOR U1014 ( .A(\min_val_reg[2][19] ), .B(n766), .Z(n767) );
  XOR U1015 ( .A(n1019), .B(\min_val_reg[3][19] ), .Z(n766) );
  NAND U1016 ( .A(n1020), .B(n933), .Z(n1019) );
  XOR U1017 ( .A(\min_val_reg[3][19] ), .B(g_input[19]), .Z(n1020) );
  XOR U1018 ( .A(n1021), .B(n1022), .Z(o[146]) );
  AND U1019 ( .A(n486), .B(n842), .Z(n1021) );
  XOR U1020 ( .A(\min_val_reg[1][18] ), .B(n1022), .Z(n842) );
  XNOR U1021 ( .A(n1023), .B(\min_val_reg[2][18] ), .Z(n1022) );
  NAND U1022 ( .A(n770), .B(n930), .Z(n1023) );
  XNOR U1023 ( .A(\min_val_reg[2][18] ), .B(n769), .Z(n770) );
  XOR U1024 ( .A(n1024), .B(\min_val_reg[3][18] ), .Z(n769) );
  NAND U1025 ( .A(n1025), .B(n933), .Z(n1024) );
  XOR U1026 ( .A(\min_val_reg[3][18] ), .B(g_input[18]), .Z(n1025) );
  XOR U1027 ( .A(n1026), .B(n1027), .Z(o[145]) );
  AND U1028 ( .A(n486), .B(n875), .Z(n1026) );
  XOR U1029 ( .A(\min_val_reg[1][17] ), .B(n1027), .Z(n875) );
  XNOR U1030 ( .A(n1028), .B(\min_val_reg[2][17] ), .Z(n1027) );
  NAND U1031 ( .A(n776), .B(n930), .Z(n1028) );
  XNOR U1032 ( .A(\min_val_reg[2][17] ), .B(n775), .Z(n776) );
  XOR U1033 ( .A(n1029), .B(\min_val_reg[3][17] ), .Z(n775) );
  NAND U1034 ( .A(n1030), .B(n933), .Z(n1029) );
  XOR U1035 ( .A(\min_val_reg[3][17] ), .B(g_input[17]), .Z(n1030) );
  XOR U1036 ( .A(n1031), .B(n1032), .Z(o[144]) );
  AND U1037 ( .A(n486), .B(n908), .Z(n1031) );
  XOR U1038 ( .A(\min_val_reg[1][16] ), .B(n1032), .Z(n908) );
  XNOR U1039 ( .A(n1033), .B(\min_val_reg[2][16] ), .Z(n1032) );
  NAND U1040 ( .A(n779), .B(n930), .Z(n1033) );
  XNOR U1041 ( .A(\min_val_reg[2][16] ), .B(n778), .Z(n779) );
  XOR U1042 ( .A(n1034), .B(\min_val_reg[3][16] ), .Z(n778) );
  NAND U1043 ( .A(n1035), .B(n933), .Z(n1034) );
  XOR U1044 ( .A(\min_val_reg[3][16] ), .B(g_input[16]), .Z(n1035) );
  XOR U1045 ( .A(n1036), .B(n1037), .Z(o[143]) );
  AND U1046 ( .A(n486), .B(n952), .Z(n1036) );
  XOR U1047 ( .A(\min_val_reg[1][15] ), .B(n1037), .Z(n952) );
  XNOR U1048 ( .A(n1038), .B(\min_val_reg[2][15] ), .Z(n1037) );
  NAND U1049 ( .A(n782), .B(n930), .Z(n1038) );
  XNOR U1050 ( .A(\min_val_reg[2][15] ), .B(n781), .Z(n782) );
  XOR U1051 ( .A(n1039), .B(\min_val_reg[3][15] ), .Z(n781) );
  NAND U1052 ( .A(n1040), .B(n933), .Z(n1039) );
  XOR U1053 ( .A(\min_val_reg[3][15] ), .B(g_input[15]), .Z(n1040) );
  XOR U1054 ( .A(n1041), .B(n1042), .Z(o[142]) );
  AND U1055 ( .A(n486), .B(n1005), .Z(n1041) );
  XOR U1056 ( .A(\min_val_reg[1][14] ), .B(n1042), .Z(n1005) );
  XNOR U1057 ( .A(n1043), .B(\min_val_reg[2][14] ), .Z(n1042) );
  NAND U1058 ( .A(n785), .B(n930), .Z(n1043) );
  XNOR U1059 ( .A(\min_val_reg[2][14] ), .B(n784), .Z(n785) );
  XOR U1060 ( .A(n1044), .B(\min_val_reg[3][14] ), .Z(n784) );
  NAND U1061 ( .A(n1045), .B(n933), .Z(n1044) );
  XOR U1062 ( .A(\min_val_reg[3][14] ), .B(g_input[14]), .Z(n1045) );
  XOR U1063 ( .A(n1046), .B(n1047), .Z(o[141]) );
  AND U1064 ( .A(n486), .B(n1048), .Z(n1046) );
  XOR U1065 ( .A(n1049), .B(n1050), .Z(o[140]) );
  AND U1066 ( .A(n486), .B(n1051), .Z(n1049) );
  XOR U1067 ( .A(\min_val_reg[0][13] ), .B(n1052), .Z(o[13]) );
  AND U1068 ( .A(n397), .B(n472), .Z(n1052) );
  XOR U1069 ( .A(\min_val_reg[0][13] ), .B(n471), .Z(n472) );
  XNOR U1070 ( .A(n1053), .B(\min_val_reg[1][13] ), .Z(n471) );
  NAND U1071 ( .A(n1048), .B(n486), .Z(n1053) );
  XOR U1072 ( .A(\min_val_reg[1][13] ), .B(n1047), .Z(n1048) );
  XNOR U1073 ( .A(n1054), .B(\min_val_reg[2][13] ), .Z(n1047) );
  NAND U1074 ( .A(n788), .B(n930), .Z(n1054) );
  XNOR U1075 ( .A(\min_val_reg[2][13] ), .B(n787), .Z(n788) );
  XOR U1076 ( .A(n1055), .B(\min_val_reg[3][13] ), .Z(n787) );
  NAND U1077 ( .A(n1056), .B(n933), .Z(n1055) );
  XOR U1078 ( .A(\min_val_reg[3][13] ), .B(g_input[13]), .Z(n1056) );
  XOR U1079 ( .A(n1057), .B(n1058), .Z(o[139]) );
  AND U1080 ( .A(n486), .B(n1059), .Z(n1057) );
  XOR U1081 ( .A(n1060), .B(n1061), .Z(o[138]) );
  AND U1082 ( .A(n486), .B(n1062), .Z(n1060) );
  XOR U1083 ( .A(n1063), .B(n1064), .Z(o[137]) );
  AND U1084 ( .A(n486), .B(n485), .Z(n1063) );
  XOR U1085 ( .A(\min_val_reg[1][9] ), .B(n1064), .Z(n485) );
  XNOR U1086 ( .A(n1065), .B(\min_val_reg[2][9] ), .Z(n1064) );
  NAND U1087 ( .A(n800), .B(n930), .Z(n1065) );
  XNOR U1088 ( .A(\min_val_reg[2][9] ), .B(n799), .Z(n800) );
  XOR U1089 ( .A(n1066), .B(\min_val_reg[3][9] ), .Z(n799) );
  NAND U1090 ( .A(n1067), .B(n933), .Z(n1066) );
  XOR U1091 ( .A(\min_val_reg[3][9] ), .B(g_input[9]), .Z(n1067) );
  XOR U1092 ( .A(n1068), .B(n1069), .Z(o[136]) );
  AND U1093 ( .A(n486), .B(n490), .Z(n1068) );
  XOR U1094 ( .A(\min_val_reg[1][8] ), .B(n1069), .Z(n490) );
  XNOR U1095 ( .A(n1070), .B(\min_val_reg[2][8] ), .Z(n1069) );
  NAND U1096 ( .A(n803), .B(n930), .Z(n1070) );
  XNOR U1097 ( .A(\min_val_reg[2][8] ), .B(n802), .Z(n803) );
  XOR U1098 ( .A(n1071), .B(\min_val_reg[3][8] ), .Z(n802) );
  NAND U1099 ( .A(n1072), .B(n933), .Z(n1071) );
  XOR U1100 ( .A(\min_val_reg[3][8] ), .B(g_input[8]), .Z(n1072) );
  XOR U1101 ( .A(n1073), .B(n1074), .Z(o[135]) );
  AND U1102 ( .A(n486), .B(n494), .Z(n1073) );
  XOR U1103 ( .A(\min_val_reg[1][7] ), .B(n1074), .Z(n494) );
  XNOR U1104 ( .A(n1075), .B(\min_val_reg[2][7] ), .Z(n1074) );
  NAND U1105 ( .A(n812), .B(n930), .Z(n1075) );
  XNOR U1106 ( .A(\min_val_reg[2][7] ), .B(n811), .Z(n812) );
  XOR U1107 ( .A(n1076), .B(\min_val_reg[3][7] ), .Z(n811) );
  NAND U1108 ( .A(n1077), .B(n933), .Z(n1076) );
  XOR U1109 ( .A(\min_val_reg[3][7] ), .B(g_input[7]), .Z(n1077) );
  XOR U1110 ( .A(n1078), .B(n1079), .Z(o[134]) );
  AND U1111 ( .A(n486), .B(n500), .Z(n1078) );
  XOR U1112 ( .A(\min_val_reg[1][6] ), .B(n1079), .Z(n500) );
  XNOR U1113 ( .A(n1080), .B(\min_val_reg[2][6] ), .Z(n1079) );
  NAND U1114 ( .A(n815), .B(n930), .Z(n1080) );
  XNOR U1115 ( .A(\min_val_reg[2][6] ), .B(n814), .Z(n815) );
  XOR U1116 ( .A(n1081), .B(\min_val_reg[3][6] ), .Z(n814) );
  NAND U1117 ( .A(n1082), .B(n933), .Z(n1081) );
  XOR U1118 ( .A(\min_val_reg[3][6] ), .B(g_input[6]), .Z(n1082) );
  XOR U1119 ( .A(n1083), .B(n1084), .Z(o[133]) );
  AND U1120 ( .A(n486), .B(n529), .Z(n1083) );
  XOR U1121 ( .A(\min_val_reg[1][5] ), .B(n1084), .Z(n529) );
  XNOR U1122 ( .A(n1085), .B(\min_val_reg[2][5] ), .Z(n1084) );
  NAND U1123 ( .A(n818), .B(n930), .Z(n1085) );
  XNOR U1124 ( .A(\min_val_reg[2][5] ), .B(n817), .Z(n818) );
  XOR U1125 ( .A(n1086), .B(\min_val_reg[3][5] ), .Z(n817) );
  NAND U1126 ( .A(n1087), .B(n933), .Z(n1086) );
  XOR U1127 ( .A(\min_val_reg[3][5] ), .B(g_input[5]), .Z(n1087) );
  XOR U1128 ( .A(n1088), .B(n1089), .Z(o[132]) );
  AND U1129 ( .A(n486), .B(n552), .Z(n1088) );
  XOR U1130 ( .A(\min_val_reg[1][4] ), .B(n1089), .Z(n552) );
  XNOR U1131 ( .A(n1090), .B(\min_val_reg[2][4] ), .Z(n1089) );
  NAND U1132 ( .A(n821), .B(n930), .Z(n1090) );
  XNOR U1133 ( .A(\min_val_reg[2][4] ), .B(n820), .Z(n821) );
  XOR U1134 ( .A(n1091), .B(\min_val_reg[3][4] ), .Z(n820) );
  NAND U1135 ( .A(n1092), .B(n933), .Z(n1091) );
  XOR U1136 ( .A(\min_val_reg[3][4] ), .B(g_input[4]), .Z(n1092) );
  XOR U1137 ( .A(n1093), .B(n1094), .Z(o[131]) );
  AND U1138 ( .A(n486), .B(n575), .Z(n1093) );
  XOR U1139 ( .A(\min_val_reg[1][3] ), .B(n1094), .Z(n575) );
  XNOR U1140 ( .A(n1095), .B(\min_val_reg[2][3] ), .Z(n1094) );
  NAND U1141 ( .A(n824), .B(n930), .Z(n1095) );
  XNOR U1142 ( .A(\min_val_reg[2][3] ), .B(n823), .Z(n824) );
  XOR U1143 ( .A(n1096), .B(\min_val_reg[3][3] ), .Z(n823) );
  NAND U1144 ( .A(n1097), .B(n933), .Z(n1096) );
  XOR U1145 ( .A(\min_val_reg[3][3] ), .B(g_input[3]), .Z(n1097) );
  XOR U1146 ( .A(n1098), .B(n1099), .Z(o[130]) );
  AND U1147 ( .A(n486), .B(n604), .Z(n1098) );
  XOR U1148 ( .A(\min_val_reg[1][2] ), .B(n1099), .Z(n604) );
  XNOR U1149 ( .A(n1100), .B(\min_val_reg[2][2] ), .Z(n1099) );
  NAND U1150 ( .A(n827), .B(n930), .Z(n1100) );
  XNOR U1151 ( .A(\min_val_reg[2][2] ), .B(n826), .Z(n827) );
  XOR U1152 ( .A(n1101), .B(\min_val_reg[3][2] ), .Z(n826) );
  NAND U1153 ( .A(n1102), .B(n933), .Z(n1101) );
  XOR U1154 ( .A(\min_val_reg[3][2] ), .B(g_input[2]), .Z(n1102) );
  XOR U1155 ( .A(\min_val_reg[0][12] ), .B(n1103), .Z(o[12]) );
  AND U1156 ( .A(n397), .B(n475), .Z(n1103) );
  XOR U1157 ( .A(\min_val_reg[0][12] ), .B(n474), .Z(n475) );
  XNOR U1158 ( .A(n1104), .B(\min_val_reg[1][12] ), .Z(n474) );
  NAND U1159 ( .A(n1051), .B(n486), .Z(n1104) );
  XOR U1160 ( .A(\min_val_reg[1][12] ), .B(n1050), .Z(n1051) );
  XNOR U1161 ( .A(n1105), .B(\min_val_reg[2][12] ), .Z(n1050) );
  NAND U1162 ( .A(n791), .B(n930), .Z(n1105) );
  XNOR U1163 ( .A(\min_val_reg[2][12] ), .B(n790), .Z(n791) );
  XOR U1164 ( .A(n1106), .B(\min_val_reg[3][12] ), .Z(n790) );
  NAND U1165 ( .A(n1107), .B(n933), .Z(n1106) );
  XOR U1166 ( .A(\min_val_reg[3][12] ), .B(g_input[12]), .Z(n1107) );
  XOR U1167 ( .A(n1108), .B(n1109), .Z(o[129]) );
  AND U1168 ( .A(n486), .B(n806), .Z(n1108) );
  XOR U1169 ( .A(\min_val_reg[1][1] ), .B(n1109), .Z(n806) );
  XNOR U1170 ( .A(n1110), .B(\min_val_reg[2][1] ), .Z(n1109) );
  NAND U1171 ( .A(n830), .B(n930), .Z(n1110) );
  XNOR U1172 ( .A(\min_val_reg[2][1] ), .B(n829), .Z(n830) );
  XOR U1173 ( .A(n1111), .B(\min_val_reg[3][1] ), .Z(n829) );
  NAND U1174 ( .A(n1112), .B(n933), .Z(n1111) );
  XOR U1175 ( .A(\min_val_reg[3][1] ), .B(g_input[1]), .Z(n1112) );
  XOR U1176 ( .A(n1113), .B(n1114), .Z(o[128]) );
  AND U1177 ( .A(n486), .B(n1115), .Z(n1113) );
  XOR U1178 ( .A(n1116), .B(n1117), .Z(o[127]) );
  AND U1179 ( .A(n401), .B(n520), .Z(n1116) );
  XOR U1180 ( .A(\min_val_reg[0][63] ), .B(n1117), .Z(n520) );
  XNOR U1181 ( .A(n1118), .B(\min_val_reg[1][63] ), .Z(n1117) );
  NAND U1182 ( .A(n836), .B(n486), .Z(n1118) );
  XOR U1183 ( .A(\min_val_reg[1][63] ), .B(n835), .Z(n836) );
  XNOR U1184 ( .A(n1119), .B(\min_val_reg[2][63] ), .Z(n835) );
  NAND U1185 ( .A(n623), .B(n930), .Z(n1119) );
  XNOR U1186 ( .A(\min_val_reg[2][63] ), .B(n621), .Z(n623) );
  XOR U1187 ( .A(n1120), .B(\min_val_reg[3][63] ), .Z(n621) );
  NAND U1188 ( .A(n1121), .B(n933), .Z(n1120) );
  XOR U1189 ( .A(\min_val_reg[3][63] ), .B(g_input[63]), .Z(n1121) );
  XOR U1190 ( .A(n1122), .B(n1123), .Z(o[126]) );
  AND U1191 ( .A(n401), .B(n522), .Z(n1122) );
  XOR U1192 ( .A(\min_val_reg[0][62] ), .B(n1123), .Z(n522) );
  XNOR U1193 ( .A(n1124), .B(\min_val_reg[1][62] ), .Z(n1123) );
  NAND U1194 ( .A(n839), .B(n486), .Z(n1124) );
  XOR U1195 ( .A(\min_val_reg[1][62] ), .B(n838), .Z(n839) );
  XNOR U1196 ( .A(n1125), .B(\min_val_reg[2][62] ), .Z(n838) );
  NAND U1197 ( .A(n626), .B(n930), .Z(n1125) );
  XNOR U1198 ( .A(\min_val_reg[2][62] ), .B(n625), .Z(n626) );
  XOR U1199 ( .A(n1126), .B(\min_val_reg[3][62] ), .Z(n625) );
  NAND U1200 ( .A(n1127), .B(n933), .Z(n1126) );
  XOR U1201 ( .A(\min_val_reg[3][62] ), .B(g_input[62]), .Z(n1127) );
  XOR U1202 ( .A(n1128), .B(n1129), .Z(o[125]) );
  AND U1203 ( .A(n401), .B(n524), .Z(n1128) );
  XOR U1204 ( .A(\min_val_reg[0][61] ), .B(n1129), .Z(n524) );
  XNOR U1205 ( .A(n1130), .B(\min_val_reg[1][61] ), .Z(n1129) );
  NAND U1206 ( .A(n845), .B(n486), .Z(n1130) );
  XOR U1207 ( .A(\min_val_reg[1][61] ), .B(n844), .Z(n845) );
  XNOR U1208 ( .A(n1131), .B(\min_val_reg[2][61] ), .Z(n844) );
  NAND U1209 ( .A(n629), .B(n930), .Z(n1131) );
  XNOR U1210 ( .A(\min_val_reg[2][61] ), .B(n628), .Z(n629) );
  XOR U1211 ( .A(n1132), .B(\min_val_reg[3][61] ), .Z(n628) );
  NAND U1212 ( .A(n1133), .B(n933), .Z(n1132) );
  XOR U1213 ( .A(\min_val_reg[3][61] ), .B(g_input[61]), .Z(n1133) );
  XOR U1214 ( .A(n1134), .B(n1135), .Z(o[124]) );
  AND U1215 ( .A(n401), .B(n526), .Z(n1134) );
  XOR U1216 ( .A(\min_val_reg[0][60] ), .B(n1135), .Z(n526) );
  XNOR U1217 ( .A(n1136), .B(\min_val_reg[1][60] ), .Z(n1135) );
  NAND U1218 ( .A(n848), .B(n486), .Z(n1136) );
  XOR U1219 ( .A(\min_val_reg[1][60] ), .B(n847), .Z(n848) );
  XNOR U1220 ( .A(n1137), .B(\min_val_reg[2][60] ), .Z(n847) );
  NAND U1221 ( .A(n632), .B(n930), .Z(n1137) );
  XNOR U1222 ( .A(\min_val_reg[2][60] ), .B(n631), .Z(n632) );
  XOR U1223 ( .A(n1138), .B(\min_val_reg[3][60] ), .Z(n631) );
  NAND U1224 ( .A(n1139), .B(n933), .Z(n1138) );
  XOR U1225 ( .A(\min_val_reg[3][60] ), .B(g_input[60]), .Z(n1139) );
  XOR U1226 ( .A(n1140), .B(n1141), .Z(o[123]) );
  AND U1227 ( .A(n401), .B(n531), .Z(n1140) );
  XOR U1228 ( .A(\min_val_reg[0][59] ), .B(n1141), .Z(n531) );
  XNOR U1229 ( .A(n1142), .B(\min_val_reg[1][59] ), .Z(n1141) );
  NAND U1230 ( .A(n851), .B(n486), .Z(n1142) );
  XOR U1231 ( .A(\min_val_reg[1][59] ), .B(n850), .Z(n851) );
  XNOR U1232 ( .A(n1143), .B(\min_val_reg[2][59] ), .Z(n850) );
  NAND U1233 ( .A(n635), .B(n930), .Z(n1143) );
  XNOR U1234 ( .A(\min_val_reg[2][59] ), .B(n634), .Z(n635) );
  XOR U1235 ( .A(n1144), .B(\min_val_reg[3][59] ), .Z(n634) );
  NAND U1236 ( .A(n1145), .B(n933), .Z(n1144) );
  XOR U1237 ( .A(\min_val_reg[3][59] ), .B(g_input[59]), .Z(n1145) );
  XOR U1238 ( .A(n1146), .B(n1147), .Z(o[122]) );
  AND U1239 ( .A(n401), .B(n533), .Z(n1146) );
  XOR U1240 ( .A(\min_val_reg[0][58] ), .B(n1147), .Z(n533) );
  XNOR U1241 ( .A(n1148), .B(\min_val_reg[1][58] ), .Z(n1147) );
  NAND U1242 ( .A(n854), .B(n486), .Z(n1148) );
  XOR U1243 ( .A(\min_val_reg[1][58] ), .B(n853), .Z(n854) );
  XNOR U1244 ( .A(n1149), .B(\min_val_reg[2][58] ), .Z(n853) );
  NAND U1245 ( .A(n638), .B(n930), .Z(n1149) );
  XNOR U1246 ( .A(\min_val_reg[2][58] ), .B(n637), .Z(n638) );
  XOR U1247 ( .A(n1150), .B(\min_val_reg[3][58] ), .Z(n637) );
  NAND U1248 ( .A(n1151), .B(n933), .Z(n1150) );
  XOR U1249 ( .A(\min_val_reg[3][58] ), .B(g_input[58]), .Z(n1151) );
  XOR U1250 ( .A(n1152), .B(n1153), .Z(o[121]) );
  AND U1251 ( .A(n401), .B(n535), .Z(n1152) );
  XOR U1252 ( .A(\min_val_reg[0][57] ), .B(n1153), .Z(n535) );
  XNOR U1253 ( .A(n1154), .B(\min_val_reg[1][57] ), .Z(n1153) );
  NAND U1254 ( .A(n857), .B(n486), .Z(n1154) );
  XOR U1255 ( .A(\min_val_reg[1][57] ), .B(n856), .Z(n857) );
  XNOR U1256 ( .A(n1155), .B(\min_val_reg[2][57] ), .Z(n856) );
  NAND U1257 ( .A(n644), .B(n930), .Z(n1155) );
  XNOR U1258 ( .A(\min_val_reg[2][57] ), .B(n643), .Z(n644) );
  XOR U1259 ( .A(n1156), .B(\min_val_reg[3][57] ), .Z(n643) );
  NAND U1260 ( .A(n1157), .B(n933), .Z(n1156) );
  XOR U1261 ( .A(\min_val_reg[3][57] ), .B(g_input[57]), .Z(n1157) );
  XOR U1262 ( .A(n1158), .B(n1159), .Z(o[120]) );
  AND U1263 ( .A(n401), .B(n537), .Z(n1158) );
  XOR U1264 ( .A(\min_val_reg[0][56] ), .B(n1159), .Z(n537) );
  XNOR U1265 ( .A(n1160), .B(\min_val_reg[1][56] ), .Z(n1159) );
  NAND U1266 ( .A(n860), .B(n486), .Z(n1160) );
  XOR U1267 ( .A(\min_val_reg[1][56] ), .B(n859), .Z(n860) );
  XNOR U1268 ( .A(n1161), .B(\min_val_reg[2][56] ), .Z(n859) );
  NAND U1269 ( .A(n647), .B(n930), .Z(n1161) );
  XNOR U1270 ( .A(\min_val_reg[2][56] ), .B(n646), .Z(n647) );
  XOR U1271 ( .A(n1162), .B(\min_val_reg[3][56] ), .Z(n646) );
  NAND U1272 ( .A(n1163), .B(n933), .Z(n1162) );
  XOR U1273 ( .A(\min_val_reg[3][56] ), .B(g_input[56]), .Z(n1163) );
  XOR U1274 ( .A(\min_val_reg[0][11] ), .B(n1164), .Z(o[11]) );
  AND U1275 ( .A(n397), .B(n478), .Z(n1164) );
  XOR U1276 ( .A(\min_val_reg[0][11] ), .B(n477), .Z(n478) );
  XNOR U1277 ( .A(n1165), .B(\min_val_reg[1][11] ), .Z(n477) );
  NAND U1278 ( .A(n1059), .B(n486), .Z(n1165) );
  XOR U1279 ( .A(\min_val_reg[1][11] ), .B(n1058), .Z(n1059) );
  XNOR U1280 ( .A(n1166), .B(\min_val_reg[2][11] ), .Z(n1058) );
  NAND U1281 ( .A(n794), .B(n930), .Z(n1166) );
  XNOR U1282 ( .A(\min_val_reg[2][11] ), .B(n793), .Z(n794) );
  XOR U1283 ( .A(n1167), .B(\min_val_reg[3][11] ), .Z(n793) );
  NAND U1284 ( .A(n1168), .B(n933), .Z(n1167) );
  XOR U1285 ( .A(\min_val_reg[3][11] ), .B(g_input[11]), .Z(n1168) );
  XOR U1286 ( .A(n1169), .B(n1170), .Z(o[119]) );
  AND U1287 ( .A(n401), .B(n539), .Z(n1169) );
  XOR U1288 ( .A(\min_val_reg[0][55] ), .B(n1170), .Z(n539) );
  XNOR U1289 ( .A(n1171), .B(\min_val_reg[1][55] ), .Z(n1170) );
  NAND U1290 ( .A(n863), .B(n486), .Z(n1171) );
  XOR U1291 ( .A(\min_val_reg[1][55] ), .B(n862), .Z(n863) );
  XNOR U1292 ( .A(n1172), .B(\min_val_reg[2][55] ), .Z(n862) );
  NAND U1293 ( .A(n650), .B(n930), .Z(n1172) );
  XNOR U1294 ( .A(\min_val_reg[2][55] ), .B(n649), .Z(n650) );
  XOR U1295 ( .A(n1173), .B(\min_val_reg[3][55] ), .Z(n649) );
  NAND U1296 ( .A(n1174), .B(n933), .Z(n1173) );
  XOR U1297 ( .A(\min_val_reg[3][55] ), .B(g_input[55]), .Z(n1174) );
  XOR U1298 ( .A(n1175), .B(n1176), .Z(o[118]) );
  AND U1299 ( .A(n401), .B(n541), .Z(n1175) );
  XOR U1300 ( .A(\min_val_reg[0][54] ), .B(n1176), .Z(n541) );
  XNOR U1301 ( .A(n1177), .B(\min_val_reg[1][54] ), .Z(n1176) );
  NAND U1302 ( .A(n866), .B(n486), .Z(n1177) );
  XOR U1303 ( .A(\min_val_reg[1][54] ), .B(n865), .Z(n866) );
  XNOR U1304 ( .A(n1178), .B(\min_val_reg[2][54] ), .Z(n865) );
  NAND U1305 ( .A(n653), .B(n930), .Z(n1178) );
  XNOR U1306 ( .A(\min_val_reg[2][54] ), .B(n652), .Z(n653) );
  XOR U1307 ( .A(n1179), .B(\min_val_reg[3][54] ), .Z(n652) );
  NAND U1308 ( .A(n1180), .B(n933), .Z(n1179) );
  XOR U1309 ( .A(\min_val_reg[3][54] ), .B(g_input[54]), .Z(n1180) );
  XOR U1310 ( .A(n1181), .B(n1182), .Z(o[117]) );
  AND U1311 ( .A(n401), .B(n543), .Z(n1181) );
  XOR U1312 ( .A(\min_val_reg[0][53] ), .B(n1182), .Z(n543) );
  XNOR U1313 ( .A(n1183), .B(\min_val_reg[1][53] ), .Z(n1182) );
  NAND U1314 ( .A(n869), .B(n486), .Z(n1183) );
  XOR U1315 ( .A(\min_val_reg[1][53] ), .B(n868), .Z(n869) );
  XNOR U1316 ( .A(n1184), .B(\min_val_reg[2][53] ), .Z(n868) );
  NAND U1317 ( .A(n656), .B(n930), .Z(n1184) );
  XNOR U1318 ( .A(\min_val_reg[2][53] ), .B(n655), .Z(n656) );
  XOR U1319 ( .A(n1185), .B(\min_val_reg[3][53] ), .Z(n655) );
  NAND U1320 ( .A(n1186), .B(n933), .Z(n1185) );
  XOR U1321 ( .A(\min_val_reg[3][53] ), .B(g_input[53]), .Z(n1186) );
  XOR U1322 ( .A(n1187), .B(n1188), .Z(o[116]) );
  AND U1323 ( .A(n401), .B(n545), .Z(n1187) );
  XOR U1324 ( .A(\min_val_reg[0][52] ), .B(n1188), .Z(n545) );
  XNOR U1325 ( .A(n1189), .B(\min_val_reg[1][52] ), .Z(n1188) );
  NAND U1326 ( .A(n872), .B(n486), .Z(n1189) );
  XOR U1327 ( .A(\min_val_reg[1][52] ), .B(n871), .Z(n872) );
  XNOR U1328 ( .A(n1190), .B(\min_val_reg[2][52] ), .Z(n871) );
  NAND U1329 ( .A(n659), .B(n930), .Z(n1190) );
  XNOR U1330 ( .A(\min_val_reg[2][52] ), .B(n658), .Z(n659) );
  XOR U1331 ( .A(n1191), .B(\min_val_reg[3][52] ), .Z(n658) );
  NAND U1332 ( .A(n1192), .B(n933), .Z(n1191) );
  XOR U1333 ( .A(\min_val_reg[3][52] ), .B(g_input[52]), .Z(n1192) );
  XOR U1334 ( .A(n1193), .B(n1194), .Z(o[115]) );
  AND U1335 ( .A(n401), .B(n547), .Z(n1193) );
  XOR U1336 ( .A(\min_val_reg[0][51] ), .B(n1194), .Z(n547) );
  XNOR U1337 ( .A(n1195), .B(\min_val_reg[1][51] ), .Z(n1194) );
  NAND U1338 ( .A(n878), .B(n486), .Z(n1195) );
  XOR U1339 ( .A(\min_val_reg[1][51] ), .B(n877), .Z(n878) );
  XNOR U1340 ( .A(n1196), .B(\min_val_reg[2][51] ), .Z(n877) );
  NAND U1341 ( .A(n662), .B(n930), .Z(n1196) );
  XNOR U1342 ( .A(\min_val_reg[2][51] ), .B(n661), .Z(n662) );
  XOR U1343 ( .A(n1197), .B(\min_val_reg[3][51] ), .Z(n661) );
  NAND U1344 ( .A(n1198), .B(n933), .Z(n1197) );
  XOR U1345 ( .A(\min_val_reg[3][51] ), .B(g_input[51]), .Z(n1198) );
  XOR U1346 ( .A(n1199), .B(n1200), .Z(o[114]) );
  AND U1347 ( .A(n401), .B(n549), .Z(n1199) );
  XOR U1348 ( .A(\min_val_reg[0][50] ), .B(n1200), .Z(n549) );
  XNOR U1349 ( .A(n1201), .B(\min_val_reg[1][50] ), .Z(n1200) );
  NAND U1350 ( .A(n881), .B(n486), .Z(n1201) );
  XOR U1351 ( .A(\min_val_reg[1][50] ), .B(n880), .Z(n881) );
  XNOR U1352 ( .A(n1202), .B(\min_val_reg[2][50] ), .Z(n880) );
  NAND U1353 ( .A(n665), .B(n930), .Z(n1202) );
  XNOR U1354 ( .A(\min_val_reg[2][50] ), .B(n664), .Z(n665) );
  XOR U1355 ( .A(n1203), .B(\min_val_reg[3][50] ), .Z(n664) );
  NAND U1356 ( .A(n1204), .B(n933), .Z(n1203) );
  XOR U1357 ( .A(\min_val_reg[3][50] ), .B(g_input[50]), .Z(n1204) );
  XOR U1358 ( .A(n1205), .B(n1206), .Z(o[113]) );
  AND U1359 ( .A(n401), .B(n554), .Z(n1205) );
  XOR U1360 ( .A(\min_val_reg[0][49] ), .B(n1206), .Z(n554) );
  XNOR U1361 ( .A(n1207), .B(\min_val_reg[1][49] ), .Z(n1206) );
  NAND U1362 ( .A(n884), .B(n486), .Z(n1207) );
  XOR U1363 ( .A(\min_val_reg[1][49] ), .B(n883), .Z(n884) );
  XNOR U1364 ( .A(n1208), .B(\min_val_reg[2][49] ), .Z(n883) );
  NAND U1365 ( .A(n668), .B(n930), .Z(n1208) );
  XNOR U1366 ( .A(\min_val_reg[2][49] ), .B(n667), .Z(n668) );
  XOR U1367 ( .A(n1209), .B(\min_val_reg[3][49] ), .Z(n667) );
  NAND U1368 ( .A(n1210), .B(n933), .Z(n1209) );
  XOR U1369 ( .A(\min_val_reg[3][49] ), .B(g_input[49]), .Z(n1210) );
  XOR U1370 ( .A(n1211), .B(n1212), .Z(o[112]) );
  AND U1371 ( .A(n401), .B(n556), .Z(n1211) );
  XOR U1372 ( .A(\min_val_reg[0][48] ), .B(n1212), .Z(n556) );
  XNOR U1373 ( .A(n1213), .B(\min_val_reg[1][48] ), .Z(n1212) );
  NAND U1374 ( .A(n887), .B(n486), .Z(n1213) );
  XOR U1375 ( .A(\min_val_reg[1][48] ), .B(n886), .Z(n887) );
  XNOR U1376 ( .A(n1214), .B(\min_val_reg[2][48] ), .Z(n886) );
  NAND U1377 ( .A(n671), .B(n930), .Z(n1214) );
  XNOR U1378 ( .A(\min_val_reg[2][48] ), .B(n670), .Z(n671) );
  XOR U1379 ( .A(n1215), .B(\min_val_reg[3][48] ), .Z(n670) );
  NAND U1380 ( .A(n1216), .B(n933), .Z(n1215) );
  XOR U1381 ( .A(\min_val_reg[3][48] ), .B(g_input[48]), .Z(n1216) );
  XOR U1382 ( .A(n1217), .B(n1218), .Z(o[111]) );
  AND U1383 ( .A(n401), .B(n558), .Z(n1217) );
  XOR U1384 ( .A(\min_val_reg[0][47] ), .B(n1218), .Z(n558) );
  XNOR U1385 ( .A(n1219), .B(\min_val_reg[1][47] ), .Z(n1218) );
  NAND U1386 ( .A(n890), .B(n486), .Z(n1219) );
  XOR U1387 ( .A(\min_val_reg[1][47] ), .B(n889), .Z(n890) );
  XNOR U1388 ( .A(n1220), .B(\min_val_reg[2][47] ), .Z(n889) );
  NAND U1389 ( .A(n677), .B(n930), .Z(n1220) );
  XNOR U1390 ( .A(\min_val_reg[2][47] ), .B(n676), .Z(n677) );
  XOR U1391 ( .A(n1221), .B(\min_val_reg[3][47] ), .Z(n676) );
  NAND U1392 ( .A(n1222), .B(n933), .Z(n1221) );
  XOR U1393 ( .A(\min_val_reg[3][47] ), .B(g_input[47]), .Z(n1222) );
  XOR U1394 ( .A(n1223), .B(n1224), .Z(o[110]) );
  AND U1395 ( .A(n401), .B(n560), .Z(n1223) );
  XOR U1396 ( .A(\min_val_reg[0][46] ), .B(n1224), .Z(n560) );
  XNOR U1397 ( .A(n1225), .B(\min_val_reg[1][46] ), .Z(n1224) );
  NAND U1398 ( .A(n893), .B(n486), .Z(n1225) );
  XOR U1399 ( .A(\min_val_reg[1][46] ), .B(n892), .Z(n893) );
  XNOR U1400 ( .A(n1226), .B(\min_val_reg[2][46] ), .Z(n892) );
  NAND U1401 ( .A(n680), .B(n930), .Z(n1226) );
  XNOR U1402 ( .A(\min_val_reg[2][46] ), .B(n679), .Z(n680) );
  XOR U1403 ( .A(n1227), .B(\min_val_reg[3][46] ), .Z(n679) );
  NAND U1404 ( .A(n1228), .B(n933), .Z(n1227) );
  XOR U1405 ( .A(\min_val_reg[3][46] ), .B(g_input[46]), .Z(n1228) );
  XOR U1406 ( .A(\min_val_reg[0][10] ), .B(n1229), .Z(o[10]) );
  AND U1407 ( .A(n397), .B(n481), .Z(n1229) );
  XOR U1408 ( .A(\min_val_reg[0][10] ), .B(n480), .Z(n481) );
  XNOR U1409 ( .A(n1230), .B(\min_val_reg[1][10] ), .Z(n480) );
  NAND U1410 ( .A(n1062), .B(n486), .Z(n1230) );
  XOR U1411 ( .A(\min_val_reg[1][10] ), .B(n1061), .Z(n1062) );
  XNOR U1412 ( .A(n1231), .B(\min_val_reg[2][10] ), .Z(n1061) );
  NAND U1413 ( .A(n797), .B(n930), .Z(n1231) );
  XNOR U1414 ( .A(\min_val_reg[2][10] ), .B(n796), .Z(n797) );
  XOR U1415 ( .A(n1232), .B(\min_val_reg[3][10] ), .Z(n796) );
  NAND U1416 ( .A(n1233), .B(n933), .Z(n1232) );
  XOR U1417 ( .A(\min_val_reg[3][10] ), .B(g_input[10]), .Z(n1233) );
  XOR U1418 ( .A(n1234), .B(n1235), .Z(o[109]) );
  AND U1419 ( .A(n401), .B(n562), .Z(n1234) );
  XOR U1420 ( .A(\min_val_reg[0][45] ), .B(n1235), .Z(n562) );
  XNOR U1421 ( .A(n1236), .B(\min_val_reg[1][45] ), .Z(n1235) );
  NAND U1422 ( .A(n896), .B(n486), .Z(n1236) );
  XOR U1423 ( .A(\min_val_reg[1][45] ), .B(n895), .Z(n896) );
  XNOR U1424 ( .A(n1237), .B(\min_val_reg[2][45] ), .Z(n895) );
  NAND U1425 ( .A(n683), .B(n930), .Z(n1237) );
  XNOR U1426 ( .A(\min_val_reg[2][45] ), .B(n682), .Z(n683) );
  XOR U1427 ( .A(n1238), .B(\min_val_reg[3][45] ), .Z(n682) );
  NAND U1428 ( .A(n1239), .B(n933), .Z(n1238) );
  XOR U1429 ( .A(\min_val_reg[3][45] ), .B(g_input[45]), .Z(n1239) );
  XOR U1430 ( .A(n1240), .B(n1241), .Z(o[108]) );
  AND U1431 ( .A(n401), .B(n564), .Z(n1240) );
  XOR U1432 ( .A(\min_val_reg[0][44] ), .B(n1241), .Z(n564) );
  XNOR U1433 ( .A(n1242), .B(\min_val_reg[1][44] ), .Z(n1241) );
  NAND U1434 ( .A(n899), .B(n486), .Z(n1242) );
  XOR U1435 ( .A(\min_val_reg[1][44] ), .B(n898), .Z(n899) );
  XNOR U1436 ( .A(n1243), .B(\min_val_reg[2][44] ), .Z(n898) );
  NAND U1437 ( .A(n686), .B(n930), .Z(n1243) );
  XNOR U1438 ( .A(\min_val_reg[2][44] ), .B(n685), .Z(n686) );
  XOR U1439 ( .A(n1244), .B(\min_val_reg[3][44] ), .Z(n685) );
  NAND U1440 ( .A(n1245), .B(n933), .Z(n1244) );
  XOR U1441 ( .A(\min_val_reg[3][44] ), .B(g_input[44]), .Z(n1245) );
  XOR U1442 ( .A(n1246), .B(n1247), .Z(o[107]) );
  AND U1443 ( .A(n401), .B(n566), .Z(n1246) );
  XOR U1444 ( .A(\min_val_reg[0][43] ), .B(n1247), .Z(n566) );
  XNOR U1445 ( .A(n1248), .B(\min_val_reg[1][43] ), .Z(n1247) );
  NAND U1446 ( .A(n902), .B(n486), .Z(n1248) );
  XOR U1447 ( .A(\min_val_reg[1][43] ), .B(n901), .Z(n902) );
  XNOR U1448 ( .A(n1249), .B(\min_val_reg[2][43] ), .Z(n901) );
  NAND U1449 ( .A(n689), .B(n930), .Z(n1249) );
  XNOR U1450 ( .A(\min_val_reg[2][43] ), .B(n688), .Z(n689) );
  XOR U1451 ( .A(n1250), .B(\min_val_reg[3][43] ), .Z(n688) );
  NAND U1452 ( .A(n1251), .B(n933), .Z(n1250) );
  XOR U1453 ( .A(\min_val_reg[3][43] ), .B(g_input[43]), .Z(n1251) );
  XOR U1454 ( .A(n1252), .B(n1253), .Z(o[106]) );
  AND U1455 ( .A(n401), .B(n568), .Z(n1252) );
  XOR U1456 ( .A(\min_val_reg[0][42] ), .B(n1253), .Z(n568) );
  XNOR U1457 ( .A(n1254), .B(\min_val_reg[1][42] ), .Z(n1253) );
  NAND U1458 ( .A(n905), .B(n486), .Z(n1254) );
  XOR U1459 ( .A(\min_val_reg[1][42] ), .B(n904), .Z(n905) );
  XNOR U1460 ( .A(n1255), .B(\min_val_reg[2][42] ), .Z(n904) );
  NAND U1461 ( .A(n692), .B(n930), .Z(n1255) );
  XNOR U1462 ( .A(\min_val_reg[2][42] ), .B(n691), .Z(n692) );
  XOR U1463 ( .A(n1256), .B(\min_val_reg[3][42] ), .Z(n691) );
  NAND U1464 ( .A(n1257), .B(n933), .Z(n1256) );
  XOR U1465 ( .A(\min_val_reg[3][42] ), .B(g_input[42]), .Z(n1257) );
  XOR U1466 ( .A(n1258), .B(n1259), .Z(o[105]) );
  AND U1467 ( .A(n401), .B(n570), .Z(n1258) );
  XOR U1468 ( .A(\min_val_reg[0][41] ), .B(n1259), .Z(n570) );
  XNOR U1469 ( .A(n1260), .B(\min_val_reg[1][41] ), .Z(n1259) );
  NAND U1470 ( .A(n911), .B(n486), .Z(n1260) );
  XOR U1471 ( .A(\min_val_reg[1][41] ), .B(n910), .Z(n911) );
  XNOR U1472 ( .A(n1261), .B(\min_val_reg[2][41] ), .Z(n910) );
  NAND U1473 ( .A(n695), .B(n930), .Z(n1261) );
  XNOR U1474 ( .A(\min_val_reg[2][41] ), .B(n694), .Z(n695) );
  XOR U1475 ( .A(n1262), .B(\min_val_reg[3][41] ), .Z(n694) );
  NAND U1476 ( .A(n1263), .B(n933), .Z(n1262) );
  XOR U1477 ( .A(\min_val_reg[3][41] ), .B(g_input[41]), .Z(n1263) );
  XOR U1478 ( .A(n1264), .B(n1265), .Z(o[104]) );
  AND U1479 ( .A(n401), .B(n572), .Z(n1264) );
  XOR U1480 ( .A(\min_val_reg[0][40] ), .B(n1265), .Z(n572) );
  XNOR U1481 ( .A(n1266), .B(\min_val_reg[1][40] ), .Z(n1265) );
  NAND U1482 ( .A(n914), .B(n486), .Z(n1266) );
  XOR U1483 ( .A(\min_val_reg[1][40] ), .B(n913), .Z(n914) );
  XNOR U1484 ( .A(n1267), .B(\min_val_reg[2][40] ), .Z(n913) );
  NAND U1485 ( .A(n698), .B(n930), .Z(n1267) );
  XNOR U1486 ( .A(\min_val_reg[2][40] ), .B(n697), .Z(n698) );
  XOR U1487 ( .A(n1268), .B(\min_val_reg[3][40] ), .Z(n697) );
  NAND U1488 ( .A(n1269), .B(n933), .Z(n1268) );
  XOR U1489 ( .A(\min_val_reg[3][40] ), .B(g_input[40]), .Z(n1269) );
  XOR U1490 ( .A(n1270), .B(n1271), .Z(o[103]) );
  AND U1491 ( .A(n401), .B(n577), .Z(n1270) );
  XOR U1492 ( .A(\min_val_reg[0][39] ), .B(n1271), .Z(n577) );
  XNOR U1493 ( .A(n1272), .B(\min_val_reg[1][39] ), .Z(n1271) );
  NAND U1494 ( .A(n917), .B(n486), .Z(n1272) );
  XOR U1495 ( .A(\min_val_reg[1][39] ), .B(n916), .Z(n917) );
  XNOR U1496 ( .A(n1273), .B(\min_val_reg[2][39] ), .Z(n916) );
  NAND U1497 ( .A(n701), .B(n930), .Z(n1273) );
  XNOR U1498 ( .A(\min_val_reg[2][39] ), .B(n700), .Z(n701) );
  XOR U1499 ( .A(n1274), .B(\min_val_reg[3][39] ), .Z(n700) );
  NAND U1500 ( .A(n1275), .B(n933), .Z(n1274) );
  XOR U1501 ( .A(\min_val_reg[3][39] ), .B(g_input[39]), .Z(n1275) );
  XOR U1502 ( .A(n1276), .B(n1277), .Z(o[102]) );
  AND U1503 ( .A(n401), .B(n579), .Z(n1276) );
  XOR U1504 ( .A(\min_val_reg[0][38] ), .B(n1277), .Z(n579) );
  XNOR U1505 ( .A(n1278), .B(\min_val_reg[1][38] ), .Z(n1277) );
  NAND U1506 ( .A(n920), .B(n486), .Z(n1278) );
  XOR U1507 ( .A(\min_val_reg[1][38] ), .B(n919), .Z(n920) );
  XNOR U1508 ( .A(n1279), .B(\min_val_reg[2][38] ), .Z(n919) );
  NAND U1509 ( .A(n704), .B(n930), .Z(n1279) );
  XNOR U1510 ( .A(\min_val_reg[2][38] ), .B(n703), .Z(n704) );
  XOR U1511 ( .A(n1280), .B(\min_val_reg[3][38] ), .Z(n703) );
  NAND U1512 ( .A(n1281), .B(n933), .Z(n1280) );
  XOR U1513 ( .A(\min_val_reg[3][38] ), .B(g_input[38]), .Z(n1281) );
  XOR U1514 ( .A(n1282), .B(n1283), .Z(o[101]) );
  AND U1515 ( .A(n401), .B(n581), .Z(n1282) );
  XOR U1516 ( .A(\min_val_reg[0][37] ), .B(n1283), .Z(n581) );
  XNOR U1517 ( .A(n1284), .B(\min_val_reg[1][37] ), .Z(n1283) );
  NAND U1518 ( .A(n923), .B(n486), .Z(n1284) );
  XOR U1519 ( .A(\min_val_reg[1][37] ), .B(n922), .Z(n923) );
  XNOR U1520 ( .A(n1285), .B(\min_val_reg[2][37] ), .Z(n922) );
  NAND U1521 ( .A(n710), .B(n930), .Z(n1285) );
  XNOR U1522 ( .A(\min_val_reg[2][37] ), .B(n709), .Z(n710) );
  XOR U1523 ( .A(n1286), .B(\min_val_reg[3][37] ), .Z(n709) );
  NAND U1524 ( .A(n1287), .B(n933), .Z(n1286) );
  XOR U1525 ( .A(\min_val_reg[3][37] ), .B(g_input[37]), .Z(n1287) );
  XOR U1526 ( .A(n1288), .B(n1289), .Z(o[100]) );
  AND U1527 ( .A(n401), .B(n583), .Z(n1288) );
  XOR U1528 ( .A(\min_val_reg[0][36] ), .B(n1289), .Z(n583) );
  XNOR U1529 ( .A(n1290), .B(\min_val_reg[1][36] ), .Z(n1289) );
  NAND U1530 ( .A(n926), .B(n486), .Z(n1290) );
  XOR U1531 ( .A(\min_val_reg[1][36] ), .B(n925), .Z(n926) );
  XNOR U1532 ( .A(n1291), .B(\min_val_reg[2][36] ), .Z(n925) );
  NAND U1533 ( .A(n713), .B(n930), .Z(n1291) );
  XNOR U1534 ( .A(\min_val_reg[2][36] ), .B(n712), .Z(n713) );
  XOR U1535 ( .A(n1292), .B(\min_val_reg[3][36] ), .Z(n712) );
  NAND U1536 ( .A(n1293), .B(n933), .Z(n1292) );
  XOR U1537 ( .A(\min_val_reg[3][36] ), .B(g_input[36]), .Z(n1293) );
  XOR U1538 ( .A(\min_val_reg[0][0] ), .B(n1294), .Z(o[0]) );
  AND U1539 ( .A(n397), .B(n518), .Z(n1294) );
  XOR U1540 ( .A(\min_val_reg[0][0] ), .B(n517), .Z(n518) );
  XNOR U1541 ( .A(n1295), .B(\min_val_reg[1][0] ), .Z(n517) );
  NAND U1542 ( .A(n1115), .B(n486), .Z(n1295) );
  XOR U1543 ( .A(\min_val_reg[1][0] ), .B(n1114), .Z(n1115) );
  XNOR U1544 ( .A(n1296), .B(\min_val_reg[2][0] ), .Z(n1114) );
  NAND U1545 ( .A(n833), .B(n930), .Z(n1296) );
  XNOR U1546 ( .A(\min_val_reg[2][0] ), .B(n832), .Z(n833) );
  XOR U1547 ( .A(n1297), .B(\min_val_reg[3][0] ), .Z(n832) );
  NAND U1548 ( .A(n1298), .B(n933), .Z(n1297) );
  XNOR U1549 ( .A(\min_val_reg[3][0] ), .B(n1299), .Z(n1298) );
  XOR U1550 ( .A(n1300), .B(n1301), .Z(\min_dist[3][9] ) );
  AND U1551 ( .A(n622), .B(n1302), .Z(n1300) );
  XOR U1552 ( .A(n1303), .B(n1304), .Z(\min_dist[3][8] ) );
  AND U1553 ( .A(n622), .B(n1305), .Z(n1303) );
  XOR U1554 ( .A(n1306), .B(n1307), .Z(\min_dist[3][7] ) );
  AND U1555 ( .A(n622), .B(n1308), .Z(n1306) );
  XOR U1556 ( .A(n1309), .B(n1310), .Z(\min_dist[3][6] ) );
  AND U1557 ( .A(n622), .B(n1311), .Z(n1309) );
  XOR U1558 ( .A(n1312), .B(n1313), .Z(\min_dist[3][5] ) );
  AND U1559 ( .A(n622), .B(n1314), .Z(n1312) );
  XOR U1560 ( .A(n1315), .B(n1316), .Z(\min_dist[3][4] ) );
  AND U1561 ( .A(n622), .B(n1317), .Z(n1315) );
  XOR U1562 ( .A(n1318), .B(n1319), .Z(\min_dist[3][3] ) );
  AND U1563 ( .A(n622), .B(n1320), .Z(n1318) );
  XOR U1564 ( .A(n1321), .B(n1322), .Z(\min_dist[3][33] ) );
  AND U1565 ( .A(n622), .B(n1323), .Z(n1321) );
  XOR U1566 ( .A(n1324), .B(n1325), .Z(\min_dist[3][32] ) );
  AND U1567 ( .A(n622), .B(n1326), .Z(n1324) );
  XOR U1568 ( .A(n1327), .B(n1328), .Z(\min_dist[3][31] ) );
  AND U1569 ( .A(n622), .B(n1329), .Z(n1327) );
  XOR U1570 ( .A(n1330), .B(n1331), .Z(\min_dist[3][30] ) );
  AND U1571 ( .A(n622), .B(n1332), .Z(n1330) );
  XOR U1572 ( .A(n1333), .B(n1334), .Z(\min_dist[3][2] ) );
  AND U1573 ( .A(n622), .B(n1335), .Z(n1333) );
  XNOR U1574 ( .A(\min_dist_reg[2][2] ), .B(n1336), .Z(n1335) );
  XOR U1575 ( .A(n1337), .B(n1338), .Z(\min_dist[3][29] ) );
  AND U1576 ( .A(n622), .B(n1339), .Z(n1337) );
  XOR U1577 ( .A(n1340), .B(n1341), .Z(\min_dist[3][28] ) );
  AND U1578 ( .A(n622), .B(n1342), .Z(n1340) );
  XOR U1579 ( .A(n1343), .B(n1344), .Z(\min_dist[3][27] ) );
  AND U1580 ( .A(n622), .B(n1345), .Z(n1343) );
  XOR U1581 ( .A(n1346), .B(n1347), .Z(\min_dist[3][26] ) );
  AND U1582 ( .A(n622), .B(n1348), .Z(n1346) );
  XOR U1583 ( .A(n1349), .B(n1350), .Z(\min_dist[3][25] ) );
  AND U1584 ( .A(n622), .B(n1351), .Z(n1349) );
  XOR U1585 ( .A(n1352), .B(n1353), .Z(\min_dist[3][24] ) );
  AND U1586 ( .A(n622), .B(n1354), .Z(n1352) );
  XOR U1587 ( .A(n1355), .B(n1356), .Z(\min_dist[3][23] ) );
  AND U1588 ( .A(n622), .B(n1357), .Z(n1355) );
  XOR U1589 ( .A(n1358), .B(n1359), .Z(\min_dist[3][22] ) );
  AND U1590 ( .A(n622), .B(n1360), .Z(n1358) );
  XOR U1591 ( .A(n1361), .B(n1362), .Z(\min_dist[3][21] ) );
  AND U1592 ( .A(n622), .B(n1363), .Z(n1361) );
  XOR U1593 ( .A(n1364), .B(n1365), .Z(\min_dist[3][20] ) );
  AND U1594 ( .A(n622), .B(n1366), .Z(n1364) );
  XOR U1595 ( .A(n1367), .B(n1368), .Z(\min_dist[3][1] ) );
  AND U1596 ( .A(n622), .B(n1369), .Z(n1367) );
  XNOR U1597 ( .A(\min_dist_reg[2][1] ), .B(n1370), .Z(n1369) );
  XOR U1598 ( .A(n1371), .B(n1372), .Z(\min_dist[3][19] ) );
  AND U1599 ( .A(n622), .B(n1373), .Z(n1371) );
  XOR U1600 ( .A(n1374), .B(n1375), .Z(\min_dist[3][18] ) );
  AND U1601 ( .A(n622), .B(n1376), .Z(n1374) );
  XOR U1602 ( .A(n1377), .B(n1378), .Z(\min_dist[3][17] ) );
  AND U1603 ( .A(n622), .B(n1379), .Z(n1377) );
  XOR U1604 ( .A(n1380), .B(n1381), .Z(\min_dist[3][16] ) );
  AND U1605 ( .A(n622), .B(n1382), .Z(n1380) );
  XOR U1606 ( .A(n1383), .B(n1384), .Z(\min_dist[3][15] ) );
  AND U1607 ( .A(n622), .B(n1385), .Z(n1383) );
  XOR U1608 ( .A(n1386), .B(n1387), .Z(\min_dist[3][14] ) );
  AND U1609 ( .A(n622), .B(n1388), .Z(n1386) );
  XOR U1610 ( .A(n1389), .B(n1390), .Z(\min_dist[3][13] ) );
  AND U1611 ( .A(n622), .B(n1391), .Z(n1389) );
  XOR U1612 ( .A(n1392), .B(n1393), .Z(\min_dist[3][12] ) );
  AND U1613 ( .A(n622), .B(n1394), .Z(n1392) );
  XOR U1614 ( .A(n1395), .B(n1396), .Z(\min_dist[3][11] ) );
  AND U1615 ( .A(n622), .B(n1397), .Z(n1395) );
  XOR U1616 ( .A(n1398), .B(n1399), .Z(\min_dist[3][10] ) );
  AND U1617 ( .A(n622), .B(n1400), .Z(n1398) );
  XOR U1618 ( .A(n1401), .B(n1402), .Z(\min_dist[3][0] ) );
  AND U1619 ( .A(n622), .B(n1403), .Z(n1401) );
  XNOR U1620 ( .A(n1404), .B(n1405), .Z(n622) );
  AND U1621 ( .A(n1406), .B(n1407), .Z(n1405) );
  XNOR U1622 ( .A(n1408), .B(n1404), .Z(n1407) );
  XNOR U1623 ( .A(n1404), .B(\min_dist_reg[2][33] ), .Z(n1406) );
  XOR U1624 ( .A(n1409), .B(n1410), .Z(n1404) );
  AND U1625 ( .A(n1411), .B(n1412), .Z(n1410) );
  XNOR U1626 ( .A(n1413), .B(n1409), .Z(n1412) );
  XNOR U1627 ( .A(n1409), .B(\min_dist_reg[2][32] ), .Z(n1411) );
  XOR U1628 ( .A(n393), .B(n1414), .Z(n1409) );
  AND U1629 ( .A(n1415), .B(n1416), .Z(n1414) );
  XNOR U1630 ( .A(n1417), .B(n393), .Z(n1416) );
  XNOR U1631 ( .A(n393), .B(\min_dist_reg[2][31] ), .Z(n1415) );
  AND U1632 ( .A(n1420), .B(n1421), .Z(n1419) );
  XNOR U1633 ( .A(n1422), .B(n1423), .Z(n1421) );
  XNOR U1634 ( .A(n1423), .B(\min_dist_reg[2][30] ), .Z(n1420) );
  IV U1635 ( .A(n1418), .Z(n1423) );
  XOR U1636 ( .A(n1424), .B(n1425), .Z(n1418) );
  AND U1637 ( .A(n1426), .B(n1427), .Z(n1425) );
  XNOR U1638 ( .A(n1428), .B(n1429), .Z(n1427) );
  XNOR U1639 ( .A(n1429), .B(\min_dist_reg[2][29] ), .Z(n1426) );
  IV U1640 ( .A(n1424), .Z(n1429) );
  XOR U1641 ( .A(n1430), .B(n1431), .Z(n1424) );
  AND U1642 ( .A(n1432), .B(n1433), .Z(n1431) );
  XNOR U1643 ( .A(n1434), .B(n1435), .Z(n1433) );
  XNOR U1644 ( .A(n1435), .B(\min_dist_reg[2][28] ), .Z(n1432) );
  IV U1645 ( .A(n1430), .Z(n1435) );
  XOR U1646 ( .A(n1436), .B(n1437), .Z(n1430) );
  AND U1647 ( .A(n1438), .B(n1439), .Z(n1437) );
  XNOR U1648 ( .A(n1440), .B(n1441), .Z(n1439) );
  XNOR U1649 ( .A(n1441), .B(\min_dist_reg[2][27] ), .Z(n1438) );
  IV U1650 ( .A(n1436), .Z(n1441) );
  XOR U1651 ( .A(n1442), .B(n1443), .Z(n1436) );
  AND U1652 ( .A(n1444), .B(n1445), .Z(n1443) );
  XNOR U1653 ( .A(n1446), .B(n1447), .Z(n1445) );
  XNOR U1654 ( .A(n1447), .B(\min_dist_reg[2][26] ), .Z(n1444) );
  IV U1655 ( .A(n1442), .Z(n1447) );
  XOR U1656 ( .A(n1448), .B(n1449), .Z(n1442) );
  AND U1657 ( .A(n1450), .B(n1451), .Z(n1449) );
  XNOR U1658 ( .A(n1452), .B(n1453), .Z(n1451) );
  XNOR U1659 ( .A(n1453), .B(\min_dist_reg[2][25] ), .Z(n1450) );
  IV U1660 ( .A(n1448), .Z(n1453) );
  XOR U1661 ( .A(n1454), .B(n1455), .Z(n1448) );
  AND U1662 ( .A(n1456), .B(n1457), .Z(n1455) );
  XNOR U1663 ( .A(n1458), .B(n1459), .Z(n1457) );
  XNOR U1664 ( .A(n1459), .B(\min_dist_reg[2][24] ), .Z(n1456) );
  IV U1665 ( .A(n1454), .Z(n1459) );
  XOR U1666 ( .A(n1460), .B(n1461), .Z(n1454) );
  AND U1667 ( .A(n1462), .B(n1463), .Z(n1461) );
  XNOR U1668 ( .A(n1464), .B(n1465), .Z(n1463) );
  XNOR U1669 ( .A(n1465), .B(\min_dist_reg[2][23] ), .Z(n1462) );
  IV U1670 ( .A(n1460), .Z(n1465) );
  XOR U1671 ( .A(n1466), .B(n1467), .Z(n1460) );
  AND U1672 ( .A(n1468), .B(n1469), .Z(n1467) );
  XNOR U1673 ( .A(n1470), .B(n1471), .Z(n1469) );
  XNOR U1674 ( .A(n1471), .B(\min_dist_reg[2][22] ), .Z(n1468) );
  IV U1675 ( .A(n1466), .Z(n1471) );
  XOR U1676 ( .A(n1472), .B(n1473), .Z(n1466) );
  AND U1677 ( .A(n1474), .B(n1475), .Z(n1473) );
  XNOR U1678 ( .A(n1476), .B(n1477), .Z(n1475) );
  XNOR U1679 ( .A(n1477), .B(\min_dist_reg[2][21] ), .Z(n1474) );
  IV U1680 ( .A(n1472), .Z(n1477) );
  XOR U1681 ( .A(n1478), .B(n1479), .Z(n1472) );
  AND U1682 ( .A(n1480), .B(n1481), .Z(n1479) );
  XNOR U1683 ( .A(n1482), .B(n1483), .Z(n1481) );
  XNOR U1684 ( .A(n1483), .B(\min_dist_reg[2][20] ), .Z(n1480) );
  IV U1685 ( .A(n1478), .Z(n1483) );
  XOR U1686 ( .A(n1484), .B(n1485), .Z(n1478) );
  AND U1687 ( .A(n1486), .B(n1487), .Z(n1485) );
  XNOR U1688 ( .A(n1488), .B(n1489), .Z(n1487) );
  XNOR U1689 ( .A(n1489), .B(\min_dist_reg[2][19] ), .Z(n1486) );
  IV U1690 ( .A(n1484), .Z(n1489) );
  XOR U1691 ( .A(n1490), .B(n1491), .Z(n1484) );
  AND U1692 ( .A(n1492), .B(n1493), .Z(n1491) );
  XNOR U1693 ( .A(n1494), .B(n1495), .Z(n1493) );
  XNOR U1694 ( .A(n1495), .B(\min_dist_reg[2][18] ), .Z(n1492) );
  IV U1695 ( .A(n1490), .Z(n1495) );
  XOR U1696 ( .A(n1496), .B(n1497), .Z(n1490) );
  AND U1697 ( .A(n1498), .B(n1499), .Z(n1497) );
  XNOR U1698 ( .A(n1500), .B(n1501), .Z(n1499) );
  XNOR U1699 ( .A(n1501), .B(\min_dist_reg[2][17] ), .Z(n1498) );
  IV U1700 ( .A(n1496), .Z(n1501) );
  XOR U1701 ( .A(n1502), .B(n1503), .Z(n1496) );
  AND U1702 ( .A(n1504), .B(n1505), .Z(n1503) );
  XNOR U1703 ( .A(n1506), .B(n1507), .Z(n1505) );
  XNOR U1704 ( .A(n1507), .B(\min_dist_reg[2][16] ), .Z(n1504) );
  IV U1705 ( .A(n1502), .Z(n1507) );
  XOR U1706 ( .A(n1508), .B(n1509), .Z(n1502) );
  AND U1707 ( .A(n1510), .B(n1511), .Z(n1509) );
  XNOR U1708 ( .A(n1512), .B(n1513), .Z(n1511) );
  XNOR U1709 ( .A(n1513), .B(\min_dist_reg[2][15] ), .Z(n1510) );
  IV U1710 ( .A(n1508), .Z(n1513) );
  XOR U1711 ( .A(n1514), .B(n1515), .Z(n1508) );
  AND U1712 ( .A(n1516), .B(n1517), .Z(n1515) );
  XNOR U1713 ( .A(n1518), .B(n1519), .Z(n1517) );
  XNOR U1714 ( .A(n1519), .B(\min_dist_reg[2][14] ), .Z(n1516) );
  IV U1715 ( .A(n1514), .Z(n1519) );
  XOR U1716 ( .A(n1520), .B(n1521), .Z(n1514) );
  AND U1717 ( .A(n1522), .B(n1523), .Z(n1521) );
  XNOR U1718 ( .A(n1524), .B(n1525), .Z(n1523) );
  XNOR U1719 ( .A(n1525), .B(\min_dist_reg[2][13] ), .Z(n1522) );
  IV U1720 ( .A(n1520), .Z(n1525) );
  XOR U1721 ( .A(n1526), .B(n1527), .Z(n1520) );
  AND U1722 ( .A(n1528), .B(n1529), .Z(n1527) );
  XNOR U1723 ( .A(n1530), .B(n1531), .Z(n1529) );
  XNOR U1724 ( .A(n1531), .B(\min_dist_reg[2][12] ), .Z(n1528) );
  IV U1725 ( .A(n1526), .Z(n1531) );
  XOR U1726 ( .A(n1532), .B(n1533), .Z(n1526) );
  AND U1727 ( .A(n1534), .B(n1535), .Z(n1533) );
  XNOR U1728 ( .A(n1536), .B(n1537), .Z(n1535) );
  XNOR U1729 ( .A(n1537), .B(\min_dist_reg[2][11] ), .Z(n1534) );
  IV U1730 ( .A(n1532), .Z(n1537) );
  XOR U1731 ( .A(n1538), .B(n1539), .Z(n1532) );
  AND U1732 ( .A(n1540), .B(n1541), .Z(n1539) );
  XNOR U1733 ( .A(n1542), .B(n1543), .Z(n1541) );
  XNOR U1734 ( .A(n1543), .B(\min_dist_reg[2][10] ), .Z(n1540) );
  IV U1735 ( .A(n1538), .Z(n1543) );
  XOR U1736 ( .A(n1544), .B(n1545), .Z(n1538) );
  AND U1737 ( .A(n1546), .B(n1547), .Z(n1545) );
  XNOR U1738 ( .A(n1548), .B(n1549), .Z(n1547) );
  XNOR U1739 ( .A(n1549), .B(\min_dist_reg[2][9] ), .Z(n1546) );
  IV U1740 ( .A(n1544), .Z(n1549) );
  XOR U1741 ( .A(n1550), .B(n1551), .Z(n1544) );
  AND U1742 ( .A(n1552), .B(n1553), .Z(n1551) );
  XNOR U1743 ( .A(n1554), .B(n1555), .Z(n1553) );
  XNOR U1744 ( .A(n1555), .B(\min_dist_reg[2][8] ), .Z(n1552) );
  IV U1745 ( .A(n1550), .Z(n1555) );
  XOR U1746 ( .A(n1556), .B(n1557), .Z(n1550) );
  AND U1747 ( .A(n1558), .B(n1559), .Z(n1557) );
  XNOR U1748 ( .A(n1560), .B(n1561), .Z(n1559) );
  XNOR U1749 ( .A(n1561), .B(\min_dist_reg[2][7] ), .Z(n1558) );
  IV U1750 ( .A(n1556), .Z(n1561) );
  XOR U1751 ( .A(n1562), .B(n1563), .Z(n1556) );
  AND U1752 ( .A(n1564), .B(n1565), .Z(n1563) );
  XNOR U1753 ( .A(n1566), .B(n1567), .Z(n1565) );
  XNOR U1754 ( .A(n1567), .B(\min_dist_reg[2][6] ), .Z(n1564) );
  IV U1755 ( .A(n1562), .Z(n1567) );
  XOR U1756 ( .A(n1568), .B(n1569), .Z(n1562) );
  AND U1757 ( .A(n1570), .B(n1571), .Z(n1569) );
  XNOR U1758 ( .A(n1572), .B(n1573), .Z(n1571) );
  XNOR U1759 ( .A(n1573), .B(\min_dist_reg[2][5] ), .Z(n1570) );
  IV U1760 ( .A(n1568), .Z(n1573) );
  XOR U1761 ( .A(n1574), .B(n1575), .Z(n1568) );
  AND U1762 ( .A(n1576), .B(n1577), .Z(n1575) );
  XNOR U1763 ( .A(n1578), .B(n1579), .Z(n1577) );
  XNOR U1764 ( .A(n1579), .B(\min_dist_reg[2][4] ), .Z(n1576) );
  IV U1765 ( .A(n1574), .Z(n1579) );
  XOR U1766 ( .A(n1580), .B(n1581), .Z(n1574) );
  AND U1767 ( .A(n1582), .B(n1583), .Z(n1581) );
  XNOR U1768 ( .A(n1584), .B(n1585), .Z(n1583) );
  XOR U1769 ( .A(n1586), .B(n1587), .Z(\min_dist[2][9] ) );
  AND U1770 ( .A(n486), .B(n1588), .Z(n1586) );
  XOR U1771 ( .A(n1589), .B(n1590), .Z(\min_dist[2][8] ) );
  AND U1772 ( .A(n486), .B(n1591), .Z(n1589) );
  XOR U1773 ( .A(n1592), .B(n1593), .Z(\min_dist[2][7] ) );
  AND U1774 ( .A(n486), .B(n1594), .Z(n1592) );
  XOR U1775 ( .A(n1595), .B(n1596), .Z(\min_dist[2][6] ) );
  AND U1776 ( .A(n486), .B(n1597), .Z(n1595) );
  XOR U1777 ( .A(n1598), .B(n1599), .Z(\min_dist[2][5] ) );
  AND U1778 ( .A(n486), .B(n1600), .Z(n1598) );
  XOR U1779 ( .A(n1601), .B(n1602), .Z(\min_dist[2][4] ) );
  AND U1780 ( .A(n486), .B(n1603), .Z(n1601) );
  XOR U1781 ( .A(n1604), .B(n1605), .Z(\min_dist[2][3] ) );
  AND U1782 ( .A(n486), .B(n1606), .Z(n1604) );
  XOR U1783 ( .A(n1607), .B(n1608), .Z(\min_dist[2][33] ) );
  AND U1784 ( .A(n486), .B(n1609), .Z(n1607) );
  XOR U1785 ( .A(n1610), .B(n1611), .Z(\min_dist[2][32] ) );
  AND U1786 ( .A(n486), .B(n1612), .Z(n1610) );
  XOR U1787 ( .A(n1613), .B(n1614), .Z(\min_dist[2][31] ) );
  AND U1788 ( .A(n486), .B(n1615), .Z(n1613) );
  XOR U1789 ( .A(n1616), .B(n1617), .Z(\min_dist[2][30] ) );
  AND U1790 ( .A(n486), .B(n1618), .Z(n1616) );
  XOR U1791 ( .A(n1619), .B(n1620), .Z(\min_dist[2][2] ) );
  AND U1792 ( .A(n486), .B(n1621), .Z(n1619) );
  XOR U1793 ( .A(\min_dist_reg[1][2] ), .B(n1620), .Z(n1621) );
  XOR U1794 ( .A(n1622), .B(n1623), .Z(\min_dist[2][29] ) );
  AND U1795 ( .A(n486), .B(n1624), .Z(n1622) );
  XOR U1796 ( .A(n1625), .B(n1626), .Z(\min_dist[2][28] ) );
  AND U1797 ( .A(n486), .B(n1627), .Z(n1625) );
  XOR U1798 ( .A(n1628), .B(n1629), .Z(\min_dist[2][27] ) );
  AND U1799 ( .A(n486), .B(n1630), .Z(n1628) );
  XOR U1800 ( .A(n1631), .B(n1632), .Z(\min_dist[2][26] ) );
  AND U1801 ( .A(n486), .B(n1633), .Z(n1631) );
  XOR U1802 ( .A(n1634), .B(n1635), .Z(\min_dist[2][25] ) );
  AND U1803 ( .A(n486), .B(n1636), .Z(n1634) );
  XOR U1804 ( .A(n1637), .B(n1638), .Z(\min_dist[2][24] ) );
  AND U1805 ( .A(n486), .B(n1639), .Z(n1637) );
  XOR U1806 ( .A(n1640), .B(n1641), .Z(\min_dist[2][23] ) );
  AND U1807 ( .A(n486), .B(n1642), .Z(n1640) );
  XOR U1808 ( .A(n1643), .B(n1644), .Z(\min_dist[2][22] ) );
  AND U1809 ( .A(n486), .B(n1645), .Z(n1643) );
  XOR U1810 ( .A(n1646), .B(n1647), .Z(\min_dist[2][21] ) );
  AND U1811 ( .A(n486), .B(n1648), .Z(n1646) );
  XOR U1812 ( .A(n1649), .B(n1650), .Z(\min_dist[2][20] ) );
  AND U1813 ( .A(n486), .B(n1651), .Z(n1649) );
  XOR U1814 ( .A(n1652), .B(n1653), .Z(\min_dist[2][1] ) );
  AND U1815 ( .A(n486), .B(n1654), .Z(n1652) );
  XOR U1816 ( .A(\min_dist_reg[1][1] ), .B(n1653), .Z(n1654) );
  XOR U1817 ( .A(n1655), .B(n1656), .Z(\min_dist[2][19] ) );
  AND U1818 ( .A(n486), .B(n1657), .Z(n1655) );
  XOR U1819 ( .A(n1658), .B(n1659), .Z(\min_dist[2][18] ) );
  AND U1820 ( .A(n486), .B(n1660), .Z(n1658) );
  XOR U1821 ( .A(n1661), .B(n1662), .Z(\min_dist[2][17] ) );
  AND U1822 ( .A(n486), .B(n1663), .Z(n1661) );
  XOR U1823 ( .A(n1664), .B(n1665), .Z(\min_dist[2][16] ) );
  AND U1824 ( .A(n486), .B(n1666), .Z(n1664) );
  XOR U1825 ( .A(n1667), .B(n1668), .Z(\min_dist[2][15] ) );
  AND U1826 ( .A(n486), .B(n1669), .Z(n1667) );
  XOR U1827 ( .A(n1670), .B(n1671), .Z(\min_dist[2][14] ) );
  AND U1828 ( .A(n486), .B(n1672), .Z(n1670) );
  XOR U1829 ( .A(n1673), .B(n1674), .Z(\min_dist[2][13] ) );
  AND U1830 ( .A(n486), .B(n1675), .Z(n1673) );
  XOR U1831 ( .A(n1676), .B(n1677), .Z(\min_dist[2][12] ) );
  AND U1832 ( .A(n486), .B(n1678), .Z(n1676) );
  XOR U1833 ( .A(n1679), .B(n1680), .Z(\min_dist[2][11] ) );
  AND U1834 ( .A(n486), .B(n1681), .Z(n1679) );
  XOR U1835 ( .A(n1682), .B(n1683), .Z(\min_dist[2][10] ) );
  AND U1836 ( .A(n486), .B(n1684), .Z(n1682) );
  XOR U1837 ( .A(n1685), .B(n1686), .Z(\min_dist[2][0] ) );
  AND U1838 ( .A(n486), .B(n1687), .Z(n1685) );
  XOR U1839 ( .A(n1688), .B(n1689), .Z(\min_dist[1][9] ) );
  AND U1840 ( .A(n401), .B(n1690), .Z(n1688) );
  XOR U1841 ( .A(n1691), .B(n1692), .Z(\min_dist[1][8] ) );
  AND U1842 ( .A(n401), .B(n1693), .Z(n1691) );
  XOR U1843 ( .A(n1694), .B(n1695), .Z(\min_dist[1][7] ) );
  AND U1844 ( .A(n401), .B(n1696), .Z(n1694) );
  XOR U1845 ( .A(n1697), .B(n1698), .Z(\min_dist[1][6] ) );
  AND U1846 ( .A(n401), .B(n1699), .Z(n1697) );
  XOR U1847 ( .A(n1700), .B(n1701), .Z(\min_dist[1][5] ) );
  AND U1848 ( .A(n401), .B(n1702), .Z(n1700) );
  XOR U1849 ( .A(n1703), .B(n1704), .Z(\min_dist[1][4] ) );
  AND U1850 ( .A(n401), .B(n1705), .Z(n1703) );
  XOR U1851 ( .A(n1706), .B(n1707), .Z(\min_dist[1][3] ) );
  AND U1852 ( .A(n401), .B(n1708), .Z(n1706) );
  XOR U1853 ( .A(n1709), .B(n1710), .Z(\min_dist[1][33] ) );
  AND U1854 ( .A(n401), .B(n1711), .Z(n1709) );
  XOR U1855 ( .A(n1712), .B(n1713), .Z(\min_dist[1][32] ) );
  AND U1856 ( .A(n401), .B(n1714), .Z(n1712) );
  XOR U1857 ( .A(n1715), .B(n1716), .Z(\min_dist[1][31] ) );
  AND U1858 ( .A(n401), .B(n1717), .Z(n1715) );
  XOR U1859 ( .A(n1718), .B(n1719), .Z(\min_dist[1][30] ) );
  AND U1860 ( .A(n401), .B(n1720), .Z(n1718) );
  XOR U1861 ( .A(n1721), .B(n1722), .Z(\min_dist[1][2] ) );
  AND U1862 ( .A(n401), .B(n1723), .Z(n1721) );
  XOR U1863 ( .A(n1724), .B(n1725), .Z(\min_dist[1][29] ) );
  AND U1864 ( .A(n401), .B(n1726), .Z(n1724) );
  XOR U1865 ( .A(n1727), .B(n1728), .Z(\min_dist[1][28] ) );
  AND U1866 ( .A(n401), .B(n1729), .Z(n1727) );
  XOR U1867 ( .A(n1730), .B(n1731), .Z(\min_dist[1][27] ) );
  AND U1868 ( .A(n401), .B(n1732), .Z(n1730) );
  XOR U1869 ( .A(n1733), .B(n1734), .Z(\min_dist[1][26] ) );
  AND U1870 ( .A(n401), .B(n1735), .Z(n1733) );
  XOR U1871 ( .A(n1736), .B(n1737), .Z(\min_dist[1][25] ) );
  AND U1872 ( .A(n401), .B(n1738), .Z(n1736) );
  XOR U1873 ( .A(n1739), .B(n1740), .Z(\min_dist[1][24] ) );
  AND U1874 ( .A(n401), .B(n1741), .Z(n1739) );
  XOR U1875 ( .A(n1742), .B(n1743), .Z(\min_dist[1][23] ) );
  AND U1876 ( .A(n401), .B(n1744), .Z(n1742) );
  XOR U1877 ( .A(n1745), .B(n1746), .Z(\min_dist[1][22] ) );
  AND U1878 ( .A(n401), .B(n1747), .Z(n1745) );
  XOR U1879 ( .A(n1748), .B(n1749), .Z(\min_dist[1][21] ) );
  AND U1880 ( .A(n401), .B(n1750), .Z(n1748) );
  XOR U1881 ( .A(n1751), .B(n1752), .Z(\min_dist[1][20] ) );
  AND U1882 ( .A(n401), .B(n1753), .Z(n1751) );
  XOR U1883 ( .A(n1754), .B(n1755), .Z(\min_dist[1][1] ) );
  AND U1884 ( .A(n401), .B(n1756), .Z(n1754) );
  XOR U1885 ( .A(n1757), .B(n1758), .Z(\min_dist[1][19] ) );
  AND U1886 ( .A(n401), .B(n1759), .Z(n1757) );
  XOR U1887 ( .A(n1760), .B(n1761), .Z(\min_dist[1][18] ) );
  AND U1888 ( .A(n401), .B(n1762), .Z(n1760) );
  XOR U1889 ( .A(n1763), .B(n1764), .Z(\min_dist[1][17] ) );
  AND U1890 ( .A(n401), .B(n1765), .Z(n1763) );
  XOR U1891 ( .A(n1766), .B(n1767), .Z(\min_dist[1][16] ) );
  AND U1892 ( .A(n401), .B(n1768), .Z(n1766) );
  XOR U1893 ( .A(n1769), .B(n1770), .Z(\min_dist[1][15] ) );
  AND U1894 ( .A(n401), .B(n1771), .Z(n1769) );
  XOR U1895 ( .A(n1772), .B(n1773), .Z(\min_dist[1][14] ) );
  AND U1896 ( .A(n401), .B(n1774), .Z(n1772) );
  XOR U1897 ( .A(n1775), .B(n1776), .Z(\min_dist[1][13] ) );
  AND U1898 ( .A(n401), .B(n1777), .Z(n1775) );
  XOR U1899 ( .A(n1778), .B(n1779), .Z(\min_dist[1][12] ) );
  AND U1900 ( .A(n401), .B(n1780), .Z(n1778) );
  XOR U1901 ( .A(n1781), .B(n1782), .Z(\min_dist[1][11] ) );
  AND U1902 ( .A(n401), .B(n1783), .Z(n1781) );
  XOR U1903 ( .A(n1784), .B(n1785), .Z(\min_dist[1][10] ) );
  AND U1904 ( .A(n401), .B(n1786), .Z(n1784) );
  XNOR U1905 ( .A(n1787), .B(n1788), .Z(\min_dist[1][0] ) );
  AND U1906 ( .A(n401), .B(n1789), .Z(n1787) );
  XNOR U1907 ( .A(\min_dist_reg[0][0] ), .B(n1788), .Z(n1789) );
  XNOR U1908 ( .A(n1790), .B(n1791), .Z(n401) );
  AND U1909 ( .A(n1792), .B(n1793), .Z(n1791) );
  XNOR U1910 ( .A(n1710), .B(n1794), .Z(n1793) );
  XNOR U1911 ( .A(n1790), .B(\min_dist_reg[0][33] ), .Z(n1792) );
  IV U1912 ( .A(n1794), .Z(n1790) );
  XOR U1913 ( .A(n1795), .B(n1796), .Z(n1794) );
  AND U1914 ( .A(n1797), .B(n1798), .Z(n1796) );
  XNOR U1915 ( .A(n1713), .B(n1795), .Z(n1798) );
  XNOR U1916 ( .A(n1799), .B(\min_dist_reg[0][32] ), .Z(n1797) );
  IV U1917 ( .A(n1795), .Z(n1799) );
  XOR U1918 ( .A(n1800), .B(n1801), .Z(n1795) );
  AND U1919 ( .A(n1802), .B(n1803), .Z(n1801) );
  XNOR U1920 ( .A(n1716), .B(n1800), .Z(n1803) );
  XNOR U1921 ( .A(n1804), .B(\min_dist_reg[0][31] ), .Z(n1802) );
  IV U1922 ( .A(n1800), .Z(n1804) );
  XOR U1923 ( .A(n1805), .B(n1806), .Z(n1800) );
  AND U1924 ( .A(n1807), .B(n1808), .Z(n1806) );
  XNOR U1925 ( .A(n1719), .B(n1805), .Z(n1808) );
  XNOR U1926 ( .A(n1809), .B(\min_dist_reg[0][30] ), .Z(n1807) );
  IV U1927 ( .A(n1805), .Z(n1809) );
  XOR U1928 ( .A(n1810), .B(n1811), .Z(n1805) );
  AND U1929 ( .A(n1812), .B(n1813), .Z(n1811) );
  XNOR U1930 ( .A(n1725), .B(n1810), .Z(n1813) );
  XNOR U1931 ( .A(n1814), .B(\min_dist_reg[0][29] ), .Z(n1812) );
  IV U1932 ( .A(n1810), .Z(n1814) );
  XOR U1933 ( .A(n1815), .B(n1816), .Z(n1810) );
  AND U1934 ( .A(n1817), .B(n1818), .Z(n1816) );
  XNOR U1935 ( .A(n1728), .B(n1815), .Z(n1818) );
  XNOR U1936 ( .A(n1819), .B(\min_dist_reg[0][28] ), .Z(n1817) );
  IV U1937 ( .A(n1815), .Z(n1819) );
  XOR U1938 ( .A(n1820), .B(n1821), .Z(n1815) );
  AND U1939 ( .A(n1822), .B(n1823), .Z(n1821) );
  XNOR U1940 ( .A(n1731), .B(n1820), .Z(n1823) );
  XNOR U1941 ( .A(n1824), .B(\min_dist_reg[0][27] ), .Z(n1822) );
  IV U1942 ( .A(n1820), .Z(n1824) );
  XOR U1943 ( .A(n1825), .B(n1826), .Z(n1820) );
  AND U1944 ( .A(n1827), .B(n1828), .Z(n1826) );
  XNOR U1945 ( .A(n1734), .B(n1825), .Z(n1828) );
  XNOR U1946 ( .A(n1829), .B(\min_dist_reg[0][26] ), .Z(n1827) );
  IV U1947 ( .A(n1825), .Z(n1829) );
  XOR U1948 ( .A(n1830), .B(n1831), .Z(n1825) );
  AND U1949 ( .A(n1832), .B(n1833), .Z(n1831) );
  XNOR U1950 ( .A(n1737), .B(n1830), .Z(n1833) );
  XNOR U1951 ( .A(n1834), .B(\min_dist_reg[0][25] ), .Z(n1832) );
  IV U1952 ( .A(n1830), .Z(n1834) );
  XOR U1953 ( .A(n1835), .B(n1836), .Z(n1830) );
  AND U1954 ( .A(n1837), .B(n1838), .Z(n1836) );
  XNOR U1955 ( .A(n1740), .B(n1835), .Z(n1838) );
  XNOR U1956 ( .A(n1839), .B(\min_dist_reg[0][24] ), .Z(n1837) );
  IV U1957 ( .A(n1835), .Z(n1839) );
  XOR U1958 ( .A(n1840), .B(n1841), .Z(n1835) );
  AND U1959 ( .A(n1842), .B(n1843), .Z(n1841) );
  XNOR U1960 ( .A(n1743), .B(n1840), .Z(n1843) );
  XNOR U1961 ( .A(n1844), .B(\min_dist_reg[0][23] ), .Z(n1842) );
  IV U1962 ( .A(n1840), .Z(n1844) );
  XOR U1963 ( .A(n1845), .B(n1846), .Z(n1840) );
  AND U1964 ( .A(n1847), .B(n1848), .Z(n1846) );
  XNOR U1965 ( .A(n1746), .B(n1845), .Z(n1848) );
  XNOR U1966 ( .A(n1849), .B(\min_dist_reg[0][22] ), .Z(n1847) );
  IV U1967 ( .A(n1845), .Z(n1849) );
  XOR U1968 ( .A(n1850), .B(n1851), .Z(n1845) );
  AND U1969 ( .A(n1852), .B(n1853), .Z(n1851) );
  XNOR U1970 ( .A(n1749), .B(n1850), .Z(n1853) );
  XNOR U1971 ( .A(n1854), .B(\min_dist_reg[0][21] ), .Z(n1852) );
  IV U1972 ( .A(n1850), .Z(n1854) );
  XOR U1973 ( .A(n1855), .B(n1856), .Z(n1850) );
  AND U1974 ( .A(n1857), .B(n1858), .Z(n1856) );
  XNOR U1975 ( .A(n1752), .B(n1855), .Z(n1858) );
  XNOR U1976 ( .A(n1859), .B(\min_dist_reg[0][20] ), .Z(n1857) );
  IV U1977 ( .A(n1855), .Z(n1859) );
  XOR U1978 ( .A(n1860), .B(n1861), .Z(n1855) );
  AND U1979 ( .A(n1862), .B(n1863), .Z(n1861) );
  XNOR U1980 ( .A(n1758), .B(n1860), .Z(n1863) );
  XNOR U1981 ( .A(n1864), .B(\min_dist_reg[0][19] ), .Z(n1862) );
  IV U1982 ( .A(n1860), .Z(n1864) );
  XOR U1983 ( .A(n1865), .B(n1866), .Z(n1860) );
  AND U1984 ( .A(n1867), .B(n1868), .Z(n1866) );
  XNOR U1985 ( .A(n1761), .B(n1865), .Z(n1868) );
  XNOR U1986 ( .A(n1869), .B(\min_dist_reg[0][18] ), .Z(n1867) );
  IV U1987 ( .A(n1865), .Z(n1869) );
  XOR U1988 ( .A(n1870), .B(n1871), .Z(n1865) );
  AND U1989 ( .A(n1872), .B(n1873), .Z(n1871) );
  XNOR U1990 ( .A(n1764), .B(n1870), .Z(n1873) );
  XNOR U1991 ( .A(n1874), .B(\min_dist_reg[0][17] ), .Z(n1872) );
  IV U1992 ( .A(n1870), .Z(n1874) );
  XOR U1993 ( .A(n1875), .B(n1876), .Z(n1870) );
  AND U1994 ( .A(n1877), .B(n1878), .Z(n1876) );
  XNOR U1995 ( .A(n1767), .B(n1875), .Z(n1878) );
  XNOR U1996 ( .A(n1879), .B(\min_dist_reg[0][16] ), .Z(n1877) );
  IV U1997 ( .A(n1875), .Z(n1879) );
  XOR U1998 ( .A(n1880), .B(n1881), .Z(n1875) );
  AND U1999 ( .A(n1882), .B(n1883), .Z(n1881) );
  XNOR U2000 ( .A(n1770), .B(n1880), .Z(n1883) );
  XNOR U2001 ( .A(n1884), .B(\min_dist_reg[0][15] ), .Z(n1882) );
  IV U2002 ( .A(n1880), .Z(n1884) );
  XOR U2003 ( .A(n1885), .B(n1886), .Z(n1880) );
  AND U2004 ( .A(n1887), .B(n1888), .Z(n1886) );
  XNOR U2005 ( .A(n1773), .B(n1885), .Z(n1888) );
  XNOR U2006 ( .A(n1889), .B(\min_dist_reg[0][14] ), .Z(n1887) );
  IV U2007 ( .A(n1885), .Z(n1889) );
  XOR U2008 ( .A(n1890), .B(n1891), .Z(n1885) );
  AND U2009 ( .A(n1892), .B(n1893), .Z(n1891) );
  XNOR U2010 ( .A(n1776), .B(n1890), .Z(n1893) );
  XNOR U2011 ( .A(n1894), .B(\min_dist_reg[0][13] ), .Z(n1892) );
  IV U2012 ( .A(n1890), .Z(n1894) );
  XOR U2013 ( .A(n1895), .B(n1896), .Z(n1890) );
  AND U2014 ( .A(n1897), .B(n1898), .Z(n1896) );
  XNOR U2015 ( .A(n1779), .B(n1895), .Z(n1898) );
  XNOR U2016 ( .A(n1899), .B(\min_dist_reg[0][12] ), .Z(n1897) );
  IV U2017 ( .A(n1895), .Z(n1899) );
  XOR U2018 ( .A(n1900), .B(n1901), .Z(n1895) );
  AND U2019 ( .A(n1902), .B(n1903), .Z(n1901) );
  XNOR U2020 ( .A(n1782), .B(n1900), .Z(n1903) );
  XNOR U2021 ( .A(n1904), .B(\min_dist_reg[0][11] ), .Z(n1902) );
  IV U2022 ( .A(n1900), .Z(n1904) );
  XOR U2023 ( .A(n1905), .B(n1906), .Z(n1900) );
  AND U2024 ( .A(n1907), .B(n1908), .Z(n1906) );
  XNOR U2025 ( .A(n1785), .B(n1905), .Z(n1908) );
  XNOR U2026 ( .A(n1909), .B(\min_dist_reg[0][10] ), .Z(n1907) );
  IV U2027 ( .A(n1905), .Z(n1909) );
  XOR U2028 ( .A(n1910), .B(n1911), .Z(n1905) );
  AND U2029 ( .A(n1912), .B(n1913), .Z(n1911) );
  XNOR U2030 ( .A(n1689), .B(n1910), .Z(n1913) );
  XNOR U2031 ( .A(n1914), .B(\min_dist_reg[0][9] ), .Z(n1912) );
  IV U2032 ( .A(n1910), .Z(n1914) );
  XOR U2033 ( .A(n1915), .B(n1916), .Z(n1910) );
  AND U2034 ( .A(n1917), .B(n1918), .Z(n1916) );
  XNOR U2035 ( .A(n1692), .B(n1915), .Z(n1918) );
  XNOR U2036 ( .A(n1919), .B(\min_dist_reg[0][8] ), .Z(n1917) );
  IV U2037 ( .A(n1915), .Z(n1919) );
  XOR U2038 ( .A(n1920), .B(n1921), .Z(n1915) );
  AND U2039 ( .A(n1922), .B(n1923), .Z(n1921) );
  XNOR U2040 ( .A(n1695), .B(n1920), .Z(n1923) );
  XNOR U2041 ( .A(n1924), .B(\min_dist_reg[0][7] ), .Z(n1922) );
  IV U2042 ( .A(n1920), .Z(n1924) );
  XOR U2043 ( .A(n1925), .B(n1926), .Z(n1920) );
  AND U2044 ( .A(n1927), .B(n1928), .Z(n1926) );
  XNOR U2045 ( .A(n1698), .B(n1925), .Z(n1928) );
  XNOR U2046 ( .A(n1929), .B(\min_dist_reg[0][6] ), .Z(n1927) );
  IV U2047 ( .A(n1925), .Z(n1929) );
  XOR U2048 ( .A(n1930), .B(n1931), .Z(n1925) );
  AND U2049 ( .A(n1932), .B(n1933), .Z(n1931) );
  XNOR U2050 ( .A(n1701), .B(n1930), .Z(n1933) );
  XNOR U2051 ( .A(n1934), .B(\min_dist_reg[0][5] ), .Z(n1932) );
  IV U2052 ( .A(n1930), .Z(n1934) );
  XOR U2053 ( .A(n1935), .B(n1936), .Z(n1930) );
  AND U2054 ( .A(n1937), .B(n1938), .Z(n1936) );
  XNOR U2055 ( .A(n1704), .B(n1935), .Z(n1938) );
  XNOR U2056 ( .A(n1939), .B(\min_dist_reg[0][4] ), .Z(n1937) );
  IV U2057 ( .A(n1935), .Z(n1939) );
  XOR U2058 ( .A(n1940), .B(n1941), .Z(n1935) );
  AND U2059 ( .A(n1942), .B(n1943), .Z(n1941) );
  XNOR U2060 ( .A(n1707), .B(n1940), .Z(n1943) );
  XNOR U2061 ( .A(n1944), .B(\min_dist_reg[0][3] ), .Z(n1942) );
  IV U2062 ( .A(n1940), .Z(n1944) );
  XOR U2063 ( .A(n1945), .B(n1946), .Z(n1940) );
  AND U2064 ( .A(n1947), .B(n1948), .Z(n1946) );
  XNOR U2065 ( .A(n1722), .B(n1945), .Z(n1948) );
  XOR U2066 ( .A(n1945), .B(\min_dist_reg[0][2] ), .Z(n1947) );
  XOR U2067 ( .A(n1949), .B(n1950), .Z(n1945) );
  NAND U2068 ( .A(n1951), .B(n1952), .Z(n1949) );
  XOR U2069 ( .A(n1950), .B(n1755), .Z(n1952) );
  XNOR U2070 ( .A(n1950), .B(\min_dist_reg[0][1] ), .Z(n1951) );
  NOR U2071 ( .A(n1788), .B(\min_dist_reg[0][0] ), .Z(n1950) );
  XOR U2072 ( .A(\min_dist_reg[0][9] ), .B(n1953), .Z(\local_min_dist[0][9] )
         );
  AND U2073 ( .A(n397), .B(n1690), .Z(n1953) );
  XOR U2074 ( .A(\min_dist_reg[0][9] ), .B(n1689), .Z(n1690) );
  XOR U2075 ( .A(\min_dist_reg[0][8] ), .B(n1954), .Z(\local_min_dist[0][8] )
         );
  AND U2076 ( .A(n397), .B(n1693), .Z(n1954) );
  XOR U2077 ( .A(\min_dist_reg[0][8] ), .B(n1692), .Z(n1693) );
  XOR U2078 ( .A(\min_dist_reg[0][7] ), .B(n1955), .Z(\local_min_dist[0][7] )
         );
  AND U2079 ( .A(n397), .B(n1696), .Z(n1955) );
  XOR U2080 ( .A(\min_dist_reg[0][7] ), .B(n1695), .Z(n1696) );
  XOR U2081 ( .A(\min_dist_reg[0][6] ), .B(n1956), .Z(\local_min_dist[0][6] )
         );
  AND U2082 ( .A(n397), .B(n1699), .Z(n1956) );
  XOR U2083 ( .A(\min_dist_reg[0][6] ), .B(n1698), .Z(n1699) );
  XOR U2084 ( .A(\min_dist_reg[0][5] ), .B(n1957), .Z(\local_min_dist[0][5] )
         );
  AND U2085 ( .A(n397), .B(n1702), .Z(n1957) );
  XOR U2086 ( .A(\min_dist_reg[0][5] ), .B(n1701), .Z(n1702) );
  XOR U2087 ( .A(\min_dist_reg[0][4] ), .B(n1958), .Z(\local_min_dist[0][4] )
         );
  AND U2088 ( .A(n397), .B(n1705), .Z(n1958) );
  XOR U2089 ( .A(\min_dist_reg[0][4] ), .B(n1704), .Z(n1705) );
  XOR U2090 ( .A(\min_dist_reg[0][3] ), .B(n1959), .Z(\local_min_dist[0][3] )
         );
  AND U2091 ( .A(n397), .B(n1708), .Z(n1959) );
  XOR U2092 ( .A(\min_dist_reg[0][3] ), .B(n1707), .Z(n1708) );
  XOR U2093 ( .A(\min_dist_reg[0][33] ), .B(n1960), .Z(\local_min_dist[0][33] ) );
  AND U2094 ( .A(n397), .B(n1711), .Z(n1960) );
  XOR U2095 ( .A(\min_dist_reg[0][33] ), .B(n1710), .Z(n1711) );
  XOR U2096 ( .A(\min_dist_reg[0][32] ), .B(n1961), .Z(\local_min_dist[0][32] ) );
  AND U2097 ( .A(n397), .B(n1714), .Z(n1961) );
  XOR U2098 ( .A(\min_dist_reg[0][32] ), .B(n1713), .Z(n1714) );
  XOR U2099 ( .A(\min_dist_reg[0][31] ), .B(n1962), .Z(\local_min_dist[0][31] ) );
  AND U2100 ( .A(n397), .B(n1717), .Z(n1962) );
  XOR U2101 ( .A(\min_dist_reg[0][31] ), .B(n1716), .Z(n1717) );
  XOR U2102 ( .A(\min_dist_reg[0][30] ), .B(n1963), .Z(\local_min_dist[0][30] ) );
  AND U2103 ( .A(n397), .B(n1720), .Z(n1963) );
  XOR U2104 ( .A(\min_dist_reg[0][30] ), .B(n1719), .Z(n1720) );
  XOR U2105 ( .A(\min_dist_reg[0][2] ), .B(n1964), .Z(\local_min_dist[0][2] )
         );
  AND U2106 ( .A(n397), .B(n1723), .Z(n1964) );
  XOR U2107 ( .A(\min_dist_reg[0][2] ), .B(n1722), .Z(n1723) );
  XOR U2108 ( .A(\min_dist_reg[0][29] ), .B(n1965), .Z(\local_min_dist[0][29] ) );
  AND U2109 ( .A(n397), .B(n1726), .Z(n1965) );
  XOR U2110 ( .A(\min_dist_reg[0][29] ), .B(n1725), .Z(n1726) );
  XOR U2111 ( .A(\min_dist_reg[0][28] ), .B(n1966), .Z(\local_min_dist[0][28] ) );
  AND U2112 ( .A(n397), .B(n1729), .Z(n1966) );
  XOR U2113 ( .A(\min_dist_reg[0][28] ), .B(n1728), .Z(n1729) );
  XOR U2114 ( .A(\min_dist_reg[0][27] ), .B(n1967), .Z(\local_min_dist[0][27] ) );
  AND U2115 ( .A(n397), .B(n1732), .Z(n1967) );
  XOR U2116 ( .A(\min_dist_reg[0][27] ), .B(n1731), .Z(n1732) );
  XOR U2117 ( .A(\min_dist_reg[0][26] ), .B(n1968), .Z(\local_min_dist[0][26] ) );
  AND U2118 ( .A(n397), .B(n1735), .Z(n1968) );
  XOR U2119 ( .A(\min_dist_reg[0][26] ), .B(n1734), .Z(n1735) );
  XOR U2120 ( .A(\min_dist_reg[0][25] ), .B(n1969), .Z(\local_min_dist[0][25] ) );
  AND U2121 ( .A(n397), .B(n1738), .Z(n1969) );
  XOR U2122 ( .A(\min_dist_reg[0][25] ), .B(n1737), .Z(n1738) );
  XOR U2123 ( .A(\min_dist_reg[0][24] ), .B(n1970), .Z(\local_min_dist[0][24] ) );
  AND U2124 ( .A(n397), .B(n1741), .Z(n1970) );
  XOR U2125 ( .A(\min_dist_reg[0][24] ), .B(n1740), .Z(n1741) );
  XOR U2126 ( .A(\min_dist_reg[0][23] ), .B(n1971), .Z(\local_min_dist[0][23] ) );
  AND U2127 ( .A(n397), .B(n1744), .Z(n1971) );
  XOR U2128 ( .A(\min_dist_reg[0][23] ), .B(n1743), .Z(n1744) );
  XOR U2129 ( .A(\min_dist_reg[0][22] ), .B(n1972), .Z(\local_min_dist[0][22] ) );
  AND U2130 ( .A(n397), .B(n1747), .Z(n1972) );
  XOR U2131 ( .A(\min_dist_reg[0][22] ), .B(n1746), .Z(n1747) );
  XOR U2132 ( .A(\min_dist_reg[0][21] ), .B(n1973), .Z(\local_min_dist[0][21] ) );
  AND U2133 ( .A(n397), .B(n1750), .Z(n1973) );
  XOR U2134 ( .A(\min_dist_reg[0][21] ), .B(n1749), .Z(n1750) );
  XOR U2135 ( .A(\min_dist_reg[0][20] ), .B(n1974), .Z(\local_min_dist[0][20] ) );
  AND U2136 ( .A(n397), .B(n1753), .Z(n1974) );
  XOR U2137 ( .A(\min_dist_reg[0][20] ), .B(n1752), .Z(n1753) );
  XOR U2138 ( .A(\min_dist_reg[0][1] ), .B(n1975), .Z(\local_min_dist[0][1] )
         );
  AND U2139 ( .A(n397), .B(n1756), .Z(n1975) );
  XOR U2140 ( .A(\min_dist_reg[0][1] ), .B(n1755), .Z(n1756) );
  XOR U2141 ( .A(\min_dist_reg[0][19] ), .B(n1976), .Z(\local_min_dist[0][19] ) );
  AND U2142 ( .A(n397), .B(n1759), .Z(n1976) );
  XOR U2143 ( .A(\min_dist_reg[0][19] ), .B(n1758), .Z(n1759) );
  XOR U2144 ( .A(\min_dist_reg[0][18] ), .B(n1977), .Z(\local_min_dist[0][18] ) );
  AND U2145 ( .A(n397), .B(n1762), .Z(n1977) );
  XOR U2146 ( .A(\min_dist_reg[0][18] ), .B(n1761), .Z(n1762) );
  XOR U2147 ( .A(\min_dist_reg[0][17] ), .B(n1978), .Z(\local_min_dist[0][17] ) );
  AND U2148 ( .A(n397), .B(n1765), .Z(n1978) );
  XOR U2149 ( .A(\min_dist_reg[0][17] ), .B(n1764), .Z(n1765) );
  XOR U2150 ( .A(\min_dist_reg[0][16] ), .B(n1979), .Z(\local_min_dist[0][16] ) );
  AND U2151 ( .A(n397), .B(n1768), .Z(n1979) );
  XOR U2152 ( .A(\min_dist_reg[0][16] ), .B(n1767), .Z(n1768) );
  XOR U2153 ( .A(\min_dist_reg[0][15] ), .B(n1980), .Z(\local_min_dist[0][15] ) );
  AND U2154 ( .A(n397), .B(n1771), .Z(n1980) );
  XOR U2155 ( .A(\min_dist_reg[0][15] ), .B(n1770), .Z(n1771) );
  XOR U2156 ( .A(\min_dist_reg[0][14] ), .B(n1981), .Z(\local_min_dist[0][14] ) );
  AND U2157 ( .A(n397), .B(n1774), .Z(n1981) );
  XOR U2158 ( .A(\min_dist_reg[0][14] ), .B(n1773), .Z(n1774) );
  XOR U2159 ( .A(\min_dist_reg[0][13] ), .B(n1982), .Z(\local_min_dist[0][13] ) );
  AND U2160 ( .A(n397), .B(n1777), .Z(n1982) );
  XOR U2161 ( .A(\min_dist_reg[0][13] ), .B(n1776), .Z(n1777) );
  XOR U2162 ( .A(\min_dist_reg[0][12] ), .B(n1983), .Z(\local_min_dist[0][12] ) );
  AND U2163 ( .A(n397), .B(n1780), .Z(n1983) );
  XOR U2164 ( .A(\min_dist_reg[0][12] ), .B(n1779), .Z(n1780) );
  XOR U2165 ( .A(\min_dist_reg[0][11] ), .B(n1984), .Z(\local_min_dist[0][11] ) );
  AND U2166 ( .A(n397), .B(n1783), .Z(n1984) );
  XOR U2167 ( .A(\min_dist_reg[0][11] ), .B(n1782), .Z(n1783) );
  XOR U2168 ( .A(\min_dist_reg[0][10] ), .B(n1985), .Z(\local_min_dist[0][10] ) );
  AND U2169 ( .A(n397), .B(n1786), .Z(n1985) );
  XOR U2170 ( .A(\min_dist_reg[0][10] ), .B(n1785), .Z(n1786) );
  XOR U2171 ( .A(\min_dist_reg[0][0] ), .B(n1986), .Z(\local_min_dist[0][0] )
         );
  AND U2172 ( .A(n397), .B(n1987), .Z(n1986) );
  XOR U2173 ( .A(\min_dist_reg[0][0] ), .B(n1988), .Z(n1987) );
  XNOR U2174 ( .A(n1989), .B(n1990), .Z(n397) );
  AND U2175 ( .A(n1991), .B(n1992), .Z(n1990) );
  XNOR U2176 ( .A(n1993), .B(n1710), .Z(n1992) );
  XNOR U2177 ( .A(n1994), .B(\min_dist_reg[1][33] ), .Z(n1710) );
  NAND U2178 ( .A(n1609), .B(n486), .Z(n1994) );
  XOR U2179 ( .A(\min_dist_reg[1][33] ), .B(n1608), .Z(n1609) );
  XNOR U2180 ( .A(n1989), .B(\min_dist_reg[0][33] ), .Z(n1991) );
  IV U2181 ( .A(n1993), .Z(n1989) );
  XOR U2182 ( .A(n1995), .B(n1996), .Z(n1993) );
  AND U2183 ( .A(n1997), .B(n1998), .Z(n1996) );
  XNOR U2184 ( .A(n1995), .B(n1713), .Z(n1998) );
  XNOR U2185 ( .A(n1999), .B(\min_dist_reg[1][32] ), .Z(n1713) );
  NAND U2186 ( .A(n1612), .B(n486), .Z(n1999) );
  XOR U2187 ( .A(\min_dist_reg[1][32] ), .B(n1611), .Z(n1612) );
  XNOR U2188 ( .A(n2000), .B(\min_dist_reg[0][32] ), .Z(n1997) );
  IV U2189 ( .A(n1995), .Z(n2000) );
  XOR U2190 ( .A(n2001), .B(n2002), .Z(n1995) );
  AND U2191 ( .A(n2003), .B(n2004), .Z(n2002) );
  XNOR U2192 ( .A(n2001), .B(n1716), .Z(n2004) );
  XNOR U2193 ( .A(n2005), .B(\min_dist_reg[1][31] ), .Z(n1716) );
  NAND U2194 ( .A(n1615), .B(n486), .Z(n2005) );
  XOR U2195 ( .A(\min_dist_reg[1][31] ), .B(n1614), .Z(n1615) );
  XNOR U2196 ( .A(n2006), .B(\min_dist_reg[0][31] ), .Z(n2003) );
  IV U2197 ( .A(n2001), .Z(n2006) );
  XOR U2198 ( .A(n2007), .B(n2008), .Z(n2001) );
  AND U2199 ( .A(n2009), .B(n2010), .Z(n2008) );
  XNOR U2200 ( .A(n2007), .B(n1719), .Z(n2010) );
  XNOR U2201 ( .A(n2011), .B(\min_dist_reg[1][30] ), .Z(n1719) );
  NAND U2202 ( .A(n1618), .B(n486), .Z(n2011) );
  XOR U2203 ( .A(\min_dist_reg[1][30] ), .B(n1617), .Z(n1618) );
  XNOR U2204 ( .A(n2012), .B(\min_dist_reg[0][30] ), .Z(n2009) );
  IV U2205 ( .A(n2007), .Z(n2012) );
  XOR U2206 ( .A(n2013), .B(n2014), .Z(n2007) );
  AND U2207 ( .A(n2015), .B(n2016), .Z(n2014) );
  XNOR U2208 ( .A(n2013), .B(n1725), .Z(n2016) );
  XNOR U2209 ( .A(n2017), .B(\min_dist_reg[1][29] ), .Z(n1725) );
  NAND U2210 ( .A(n1624), .B(n486), .Z(n2017) );
  XOR U2211 ( .A(\min_dist_reg[1][29] ), .B(n1623), .Z(n1624) );
  XNOR U2212 ( .A(n2018), .B(\min_dist_reg[0][29] ), .Z(n2015) );
  IV U2213 ( .A(n2013), .Z(n2018) );
  XOR U2214 ( .A(n2019), .B(n2020), .Z(n2013) );
  AND U2215 ( .A(n2021), .B(n2022), .Z(n2020) );
  XNOR U2216 ( .A(n2019), .B(n1728), .Z(n2022) );
  XNOR U2217 ( .A(n2023), .B(\min_dist_reg[1][28] ), .Z(n1728) );
  NAND U2218 ( .A(n1627), .B(n486), .Z(n2023) );
  XOR U2219 ( .A(\min_dist_reg[1][28] ), .B(n1626), .Z(n1627) );
  XNOR U2220 ( .A(n2024), .B(\min_dist_reg[0][28] ), .Z(n2021) );
  IV U2221 ( .A(n2019), .Z(n2024) );
  XOR U2222 ( .A(n2025), .B(n2026), .Z(n2019) );
  AND U2223 ( .A(n2027), .B(n2028), .Z(n2026) );
  XNOR U2224 ( .A(n2025), .B(n1731), .Z(n2028) );
  XNOR U2225 ( .A(n2029), .B(\min_dist_reg[1][27] ), .Z(n1731) );
  NAND U2226 ( .A(n1630), .B(n486), .Z(n2029) );
  XOR U2227 ( .A(\min_dist_reg[1][27] ), .B(n1629), .Z(n1630) );
  XNOR U2228 ( .A(n2030), .B(\min_dist_reg[0][27] ), .Z(n2027) );
  IV U2229 ( .A(n2025), .Z(n2030) );
  XOR U2230 ( .A(n2031), .B(n2032), .Z(n2025) );
  AND U2231 ( .A(n2033), .B(n2034), .Z(n2032) );
  XNOR U2232 ( .A(n2031), .B(n1734), .Z(n2034) );
  XNOR U2233 ( .A(n2035), .B(\min_dist_reg[1][26] ), .Z(n1734) );
  NAND U2234 ( .A(n1633), .B(n486), .Z(n2035) );
  XOR U2235 ( .A(\min_dist_reg[1][26] ), .B(n1632), .Z(n1633) );
  XNOR U2236 ( .A(n2036), .B(\min_dist_reg[0][26] ), .Z(n2033) );
  IV U2237 ( .A(n2031), .Z(n2036) );
  XOR U2238 ( .A(n2037), .B(n2038), .Z(n2031) );
  AND U2239 ( .A(n2039), .B(n2040), .Z(n2038) );
  XNOR U2240 ( .A(n2037), .B(n1737), .Z(n2040) );
  XNOR U2241 ( .A(n2041), .B(\min_dist_reg[1][25] ), .Z(n1737) );
  NAND U2242 ( .A(n1636), .B(n486), .Z(n2041) );
  XOR U2243 ( .A(\min_dist_reg[1][25] ), .B(n1635), .Z(n1636) );
  XNOR U2244 ( .A(n2042), .B(\min_dist_reg[0][25] ), .Z(n2039) );
  IV U2245 ( .A(n2037), .Z(n2042) );
  XOR U2246 ( .A(n2043), .B(n2044), .Z(n2037) );
  AND U2247 ( .A(n2045), .B(n2046), .Z(n2044) );
  XNOR U2248 ( .A(n2043), .B(n1740), .Z(n2046) );
  XNOR U2249 ( .A(n2047), .B(\min_dist_reg[1][24] ), .Z(n1740) );
  NAND U2250 ( .A(n1639), .B(n486), .Z(n2047) );
  XOR U2251 ( .A(\min_dist_reg[1][24] ), .B(n1638), .Z(n1639) );
  XNOR U2252 ( .A(n2048), .B(\min_dist_reg[0][24] ), .Z(n2045) );
  IV U2253 ( .A(n2043), .Z(n2048) );
  XOR U2254 ( .A(n2049), .B(n2050), .Z(n2043) );
  AND U2255 ( .A(n2051), .B(n2052), .Z(n2050) );
  XNOR U2256 ( .A(n2049), .B(n1743), .Z(n2052) );
  XNOR U2257 ( .A(n2053), .B(\min_dist_reg[1][23] ), .Z(n1743) );
  NAND U2258 ( .A(n1642), .B(n486), .Z(n2053) );
  XOR U2259 ( .A(\min_dist_reg[1][23] ), .B(n1641), .Z(n1642) );
  XNOR U2260 ( .A(n2054), .B(\min_dist_reg[0][23] ), .Z(n2051) );
  IV U2261 ( .A(n2049), .Z(n2054) );
  XOR U2262 ( .A(n2055), .B(n2056), .Z(n2049) );
  AND U2263 ( .A(n2057), .B(n2058), .Z(n2056) );
  XNOR U2264 ( .A(n2055), .B(n1746), .Z(n2058) );
  XNOR U2265 ( .A(n2059), .B(\min_dist_reg[1][22] ), .Z(n1746) );
  NAND U2266 ( .A(n1645), .B(n486), .Z(n2059) );
  XOR U2267 ( .A(\min_dist_reg[1][22] ), .B(n1644), .Z(n1645) );
  XNOR U2268 ( .A(n2060), .B(\min_dist_reg[0][22] ), .Z(n2057) );
  IV U2269 ( .A(n2055), .Z(n2060) );
  XOR U2270 ( .A(n2061), .B(n2062), .Z(n2055) );
  AND U2271 ( .A(n2063), .B(n2064), .Z(n2062) );
  XNOR U2272 ( .A(n2061), .B(n1749), .Z(n2064) );
  XNOR U2273 ( .A(n2065), .B(\min_dist_reg[1][21] ), .Z(n1749) );
  NAND U2274 ( .A(n1648), .B(n486), .Z(n2065) );
  XOR U2275 ( .A(\min_dist_reg[1][21] ), .B(n1647), .Z(n1648) );
  XNOR U2276 ( .A(n2066), .B(\min_dist_reg[0][21] ), .Z(n2063) );
  IV U2277 ( .A(n2061), .Z(n2066) );
  XOR U2278 ( .A(n2067), .B(n2068), .Z(n2061) );
  AND U2279 ( .A(n2069), .B(n2070), .Z(n2068) );
  XNOR U2280 ( .A(n2067), .B(n1752), .Z(n2070) );
  XNOR U2281 ( .A(n2071), .B(\min_dist_reg[1][20] ), .Z(n1752) );
  NAND U2282 ( .A(n1651), .B(n486), .Z(n2071) );
  XOR U2283 ( .A(\min_dist_reg[1][20] ), .B(n1650), .Z(n1651) );
  XNOR U2284 ( .A(n2072), .B(\min_dist_reg[0][20] ), .Z(n2069) );
  IV U2285 ( .A(n2067), .Z(n2072) );
  XOR U2286 ( .A(n2073), .B(n2074), .Z(n2067) );
  AND U2287 ( .A(n2075), .B(n2076), .Z(n2074) );
  XNOR U2288 ( .A(n2073), .B(n1758), .Z(n2076) );
  XNOR U2289 ( .A(n2077), .B(\min_dist_reg[1][19] ), .Z(n1758) );
  NAND U2290 ( .A(n1657), .B(n486), .Z(n2077) );
  XOR U2291 ( .A(\min_dist_reg[1][19] ), .B(n1656), .Z(n1657) );
  XNOR U2292 ( .A(n2078), .B(\min_dist_reg[0][19] ), .Z(n2075) );
  IV U2293 ( .A(n2073), .Z(n2078) );
  XOR U2294 ( .A(n2079), .B(n2080), .Z(n2073) );
  AND U2295 ( .A(n2081), .B(n2082), .Z(n2080) );
  XNOR U2296 ( .A(n2079), .B(n1761), .Z(n2082) );
  XNOR U2297 ( .A(n2083), .B(\min_dist_reg[1][18] ), .Z(n1761) );
  NAND U2298 ( .A(n1660), .B(n486), .Z(n2083) );
  XOR U2299 ( .A(\min_dist_reg[1][18] ), .B(n1659), .Z(n1660) );
  XNOR U2300 ( .A(n2084), .B(\min_dist_reg[0][18] ), .Z(n2081) );
  IV U2301 ( .A(n2079), .Z(n2084) );
  XOR U2302 ( .A(n2085), .B(n2086), .Z(n2079) );
  AND U2303 ( .A(n2087), .B(n2088), .Z(n2086) );
  XNOR U2304 ( .A(n2085), .B(n1764), .Z(n2088) );
  XNOR U2305 ( .A(n2089), .B(\min_dist_reg[1][17] ), .Z(n1764) );
  NAND U2306 ( .A(n1663), .B(n486), .Z(n2089) );
  XOR U2307 ( .A(\min_dist_reg[1][17] ), .B(n1662), .Z(n1663) );
  XNOR U2308 ( .A(n2090), .B(\min_dist_reg[0][17] ), .Z(n2087) );
  IV U2309 ( .A(n2085), .Z(n2090) );
  XOR U2310 ( .A(n2091), .B(n2092), .Z(n2085) );
  AND U2311 ( .A(n2093), .B(n2094), .Z(n2092) );
  XNOR U2312 ( .A(n2091), .B(n1767), .Z(n2094) );
  XNOR U2313 ( .A(n2095), .B(\min_dist_reg[1][16] ), .Z(n1767) );
  NAND U2314 ( .A(n1666), .B(n486), .Z(n2095) );
  XOR U2315 ( .A(\min_dist_reg[1][16] ), .B(n1665), .Z(n1666) );
  XNOR U2316 ( .A(n2096), .B(\min_dist_reg[0][16] ), .Z(n2093) );
  IV U2317 ( .A(n2091), .Z(n2096) );
  XOR U2318 ( .A(n2097), .B(n2098), .Z(n2091) );
  AND U2319 ( .A(n2099), .B(n2100), .Z(n2098) );
  XNOR U2320 ( .A(n2097), .B(n1770), .Z(n2100) );
  XNOR U2321 ( .A(n2101), .B(\min_dist_reg[1][15] ), .Z(n1770) );
  NAND U2322 ( .A(n1669), .B(n486), .Z(n2101) );
  XOR U2323 ( .A(\min_dist_reg[1][15] ), .B(n1668), .Z(n1669) );
  XNOR U2324 ( .A(n2102), .B(\min_dist_reg[0][15] ), .Z(n2099) );
  IV U2325 ( .A(n2097), .Z(n2102) );
  XOR U2326 ( .A(n2103), .B(n2104), .Z(n2097) );
  AND U2327 ( .A(n2105), .B(n2106), .Z(n2104) );
  XNOR U2328 ( .A(n2103), .B(n1773), .Z(n2106) );
  XNOR U2329 ( .A(n2107), .B(\min_dist_reg[1][14] ), .Z(n1773) );
  NAND U2330 ( .A(n1672), .B(n486), .Z(n2107) );
  XOR U2331 ( .A(\min_dist_reg[1][14] ), .B(n1671), .Z(n1672) );
  XNOR U2332 ( .A(n2108), .B(\min_dist_reg[0][14] ), .Z(n2105) );
  IV U2333 ( .A(n2103), .Z(n2108) );
  XOR U2334 ( .A(n2109), .B(n2110), .Z(n2103) );
  AND U2335 ( .A(n2111), .B(n2112), .Z(n2110) );
  XNOR U2336 ( .A(n2109), .B(n1776), .Z(n2112) );
  XNOR U2337 ( .A(n2113), .B(\min_dist_reg[1][13] ), .Z(n1776) );
  NAND U2338 ( .A(n1675), .B(n486), .Z(n2113) );
  XOR U2339 ( .A(\min_dist_reg[1][13] ), .B(n1674), .Z(n1675) );
  XNOR U2340 ( .A(n2114), .B(\min_dist_reg[0][13] ), .Z(n2111) );
  IV U2341 ( .A(n2109), .Z(n2114) );
  XOR U2342 ( .A(n2115), .B(n2116), .Z(n2109) );
  AND U2343 ( .A(n2117), .B(n2118), .Z(n2116) );
  XNOR U2344 ( .A(n2115), .B(n1779), .Z(n2118) );
  XNOR U2345 ( .A(n2119), .B(\min_dist_reg[1][12] ), .Z(n1779) );
  NAND U2346 ( .A(n1678), .B(n486), .Z(n2119) );
  XOR U2347 ( .A(\min_dist_reg[1][12] ), .B(n1677), .Z(n1678) );
  XNOR U2348 ( .A(n2120), .B(\min_dist_reg[0][12] ), .Z(n2117) );
  IV U2349 ( .A(n2115), .Z(n2120) );
  XOR U2350 ( .A(n2121), .B(n2122), .Z(n2115) );
  AND U2351 ( .A(n2123), .B(n2124), .Z(n2122) );
  XNOR U2352 ( .A(n2121), .B(n1782), .Z(n2124) );
  XNOR U2353 ( .A(n2125), .B(\min_dist_reg[1][11] ), .Z(n1782) );
  NAND U2354 ( .A(n1681), .B(n486), .Z(n2125) );
  XOR U2355 ( .A(\min_dist_reg[1][11] ), .B(n1680), .Z(n1681) );
  XNOR U2356 ( .A(n2126), .B(\min_dist_reg[0][11] ), .Z(n2123) );
  IV U2357 ( .A(n2121), .Z(n2126) );
  XOR U2358 ( .A(n2127), .B(n2128), .Z(n2121) );
  AND U2359 ( .A(n2129), .B(n2130), .Z(n2128) );
  XNOR U2360 ( .A(n2127), .B(n1785), .Z(n2130) );
  XNOR U2361 ( .A(n2131), .B(\min_dist_reg[1][10] ), .Z(n1785) );
  NAND U2362 ( .A(n1684), .B(n486), .Z(n2131) );
  XOR U2363 ( .A(\min_dist_reg[1][10] ), .B(n1683), .Z(n1684) );
  XNOR U2364 ( .A(n2132), .B(\min_dist_reg[0][10] ), .Z(n2129) );
  IV U2365 ( .A(n2127), .Z(n2132) );
  XOR U2366 ( .A(n2133), .B(n2134), .Z(n2127) );
  AND U2367 ( .A(n2135), .B(n2136), .Z(n2134) );
  XNOR U2368 ( .A(n2133), .B(n1689), .Z(n2136) );
  XNOR U2369 ( .A(n2137), .B(\min_dist_reg[1][9] ), .Z(n1689) );
  NAND U2370 ( .A(n1588), .B(n486), .Z(n2137) );
  XOR U2371 ( .A(\min_dist_reg[1][9] ), .B(n1587), .Z(n1588) );
  XNOR U2372 ( .A(n2138), .B(\min_dist_reg[0][9] ), .Z(n2135) );
  IV U2373 ( .A(n2133), .Z(n2138) );
  XOR U2374 ( .A(n2139), .B(n2140), .Z(n2133) );
  AND U2375 ( .A(n2141), .B(n2142), .Z(n2140) );
  XNOR U2376 ( .A(n2139), .B(n1692), .Z(n2142) );
  XNOR U2377 ( .A(n2143), .B(\min_dist_reg[1][8] ), .Z(n1692) );
  NAND U2378 ( .A(n1591), .B(n486), .Z(n2143) );
  XOR U2379 ( .A(\min_dist_reg[1][8] ), .B(n1590), .Z(n1591) );
  XNOR U2380 ( .A(n2144), .B(\min_dist_reg[0][8] ), .Z(n2141) );
  IV U2381 ( .A(n2139), .Z(n2144) );
  XOR U2382 ( .A(n2145), .B(n2146), .Z(n2139) );
  AND U2383 ( .A(n2147), .B(n2148), .Z(n2146) );
  XNOR U2384 ( .A(n2145), .B(n1695), .Z(n2148) );
  XNOR U2385 ( .A(n2149), .B(\min_dist_reg[1][7] ), .Z(n1695) );
  NAND U2386 ( .A(n1594), .B(n486), .Z(n2149) );
  XOR U2387 ( .A(\min_dist_reg[1][7] ), .B(n1593), .Z(n1594) );
  XNOR U2388 ( .A(n2150), .B(\min_dist_reg[0][7] ), .Z(n2147) );
  IV U2389 ( .A(n2145), .Z(n2150) );
  XOR U2390 ( .A(n2151), .B(n2152), .Z(n2145) );
  AND U2391 ( .A(n2153), .B(n2154), .Z(n2152) );
  XNOR U2392 ( .A(n2151), .B(n1698), .Z(n2154) );
  XNOR U2393 ( .A(n2155), .B(\min_dist_reg[1][6] ), .Z(n1698) );
  NAND U2394 ( .A(n1597), .B(n486), .Z(n2155) );
  XOR U2395 ( .A(\min_dist_reg[1][6] ), .B(n1596), .Z(n1597) );
  XNOR U2396 ( .A(n2156), .B(\min_dist_reg[0][6] ), .Z(n2153) );
  IV U2397 ( .A(n2151), .Z(n2156) );
  XOR U2398 ( .A(n2157), .B(n2158), .Z(n2151) );
  AND U2399 ( .A(n2159), .B(n2160), .Z(n2158) );
  XNOR U2400 ( .A(n2157), .B(n1701), .Z(n2160) );
  XNOR U2401 ( .A(n2161), .B(\min_dist_reg[1][5] ), .Z(n1701) );
  NAND U2402 ( .A(n1600), .B(n486), .Z(n2161) );
  XOR U2403 ( .A(\min_dist_reg[1][5] ), .B(n1599), .Z(n1600) );
  XNOR U2404 ( .A(n2162), .B(\min_dist_reg[0][5] ), .Z(n2159) );
  IV U2405 ( .A(n2157), .Z(n2162) );
  XOR U2406 ( .A(n2163), .B(n2164), .Z(n2157) );
  AND U2407 ( .A(n2165), .B(n2166), .Z(n2164) );
  XNOR U2408 ( .A(n2163), .B(n1704), .Z(n2166) );
  XNOR U2409 ( .A(n2167), .B(\min_dist_reg[1][4] ), .Z(n1704) );
  NAND U2410 ( .A(n1603), .B(n486), .Z(n2167) );
  XOR U2411 ( .A(\min_dist_reg[1][4] ), .B(n1602), .Z(n1603) );
  XNOR U2412 ( .A(n2168), .B(\min_dist_reg[0][4] ), .Z(n2165) );
  IV U2413 ( .A(n2163), .Z(n2168) );
  XOR U2414 ( .A(n2169), .B(n2170), .Z(n2163) );
  AND U2415 ( .A(n2171), .B(n2172), .Z(n2170) );
  XNOR U2416 ( .A(n2169), .B(n1707), .Z(n2172) );
  XNOR U2417 ( .A(n2173), .B(\min_dist_reg[1][3] ), .Z(n1707) );
  NAND U2418 ( .A(n1606), .B(n486), .Z(n2173) );
  XOR U2419 ( .A(\min_dist_reg[1][3] ), .B(n1605), .Z(n1606) );
  XNOR U2420 ( .A(n2174), .B(\min_dist_reg[0][3] ), .Z(n2171) );
  IV U2421 ( .A(n2169), .Z(n2174) );
  XOR U2422 ( .A(n2175), .B(n2176), .Z(n2169) );
  AND U2423 ( .A(n2177), .B(n2178), .Z(n2176) );
  XNOR U2424 ( .A(n2175), .B(n1722), .Z(n2178) );
  XNOR U2425 ( .A(n2179), .B(\min_dist_reg[1][2] ), .Z(n1722) );
  NAND U2426 ( .A(n2180), .B(n486), .Z(n2179) );
  XNOR U2427 ( .A(n2181), .B(n1620), .Z(n2180) );
  XOR U2428 ( .A(n2175), .B(\min_dist_reg[0][2] ), .Z(n2177) );
  XOR U2429 ( .A(n2182), .B(n2183), .Z(n2175) );
  NAND U2430 ( .A(n2184), .B(n2185), .Z(n2182) );
  XOR U2431 ( .A(n2183), .B(n1755), .Z(n2185) );
  XNOR U2432 ( .A(n2186), .B(\min_dist_reg[1][1] ), .Z(n1755) );
  NAND U2433 ( .A(n2187), .B(n486), .Z(n2186) );
  XNOR U2434 ( .A(n2188), .B(n1653), .Z(n2187) );
  XNOR U2435 ( .A(n2183), .B(\min_dist_reg[0][1] ), .Z(n2184) );
  ANDN U2436 ( .A(n1988), .B(\min_dist_reg[0][0] ), .Z(n2183) );
  IV U2437 ( .A(n1788), .Z(n1988) );
  XOR U2438 ( .A(n2189), .B(\min_dist_reg[1][0] ), .Z(n1788) );
  NAND U2439 ( .A(n1687), .B(n486), .Z(n2189) );
  XNOR U2440 ( .A(n2190), .B(n2191), .Z(n486) );
  AND U2441 ( .A(n2192), .B(n2193), .Z(n2191) );
  XNOR U2442 ( .A(n1608), .B(n2194), .Z(n2193) );
  XNOR U2443 ( .A(n2195), .B(\min_dist_reg[2][33] ), .Z(n1608) );
  NAND U2444 ( .A(n1323), .B(n930), .Z(n2195) );
  XNOR U2445 ( .A(\min_dist_reg[2][33] ), .B(n1408), .Z(n1323) );
  IV U2446 ( .A(n1322), .Z(n1408) );
  XNOR U2447 ( .A(n2190), .B(\min_dist_reg[1][33] ), .Z(n2192) );
  IV U2448 ( .A(n2194), .Z(n2190) );
  XOR U2449 ( .A(n2196), .B(n2197), .Z(n2194) );
  AND U2450 ( .A(n2198), .B(n2199), .Z(n2197) );
  XNOR U2451 ( .A(n1611), .B(n2196), .Z(n2199) );
  XNOR U2452 ( .A(n2200), .B(\min_dist_reg[2][32] ), .Z(n1611) );
  NAND U2453 ( .A(n1326), .B(n930), .Z(n2200) );
  XNOR U2454 ( .A(\min_dist_reg[2][32] ), .B(n1413), .Z(n1326) );
  IV U2455 ( .A(n1325), .Z(n1413) );
  XNOR U2456 ( .A(n2201), .B(\min_dist_reg[1][32] ), .Z(n2198) );
  IV U2457 ( .A(n2196), .Z(n2201) );
  XOR U2458 ( .A(n2202), .B(n2203), .Z(n2196) );
  AND U2459 ( .A(n2204), .B(n2205), .Z(n2203) );
  XNOR U2460 ( .A(n1614), .B(n2202), .Z(n2205) );
  XNOR U2461 ( .A(n2206), .B(\min_dist_reg[2][31] ), .Z(n1614) );
  NAND U2462 ( .A(n1329), .B(n930), .Z(n2206) );
  XNOR U2463 ( .A(\min_dist_reg[2][31] ), .B(n1417), .Z(n1329) );
  IV U2464 ( .A(n1328), .Z(n1417) );
  XNOR U2465 ( .A(n2207), .B(\min_dist_reg[1][31] ), .Z(n2204) );
  IV U2466 ( .A(n2202), .Z(n2207) );
  XOR U2467 ( .A(n2208), .B(n2209), .Z(n2202) );
  AND U2468 ( .A(n2210), .B(n2211), .Z(n2209) );
  XNOR U2469 ( .A(n1617), .B(n2208), .Z(n2211) );
  XNOR U2470 ( .A(n2212), .B(\min_dist_reg[2][30] ), .Z(n1617) );
  NAND U2471 ( .A(n1332), .B(n930), .Z(n2212) );
  XNOR U2472 ( .A(\min_dist_reg[2][30] ), .B(n1422), .Z(n1332) );
  IV U2473 ( .A(n1331), .Z(n1422) );
  XNOR U2474 ( .A(n2213), .B(\min_dist_reg[1][30] ), .Z(n2210) );
  IV U2475 ( .A(n2208), .Z(n2213) );
  XOR U2476 ( .A(n2214), .B(n2215), .Z(n2208) );
  AND U2477 ( .A(n2216), .B(n2217), .Z(n2215) );
  XNOR U2478 ( .A(n1623), .B(n2214), .Z(n2217) );
  XNOR U2479 ( .A(n2218), .B(\min_dist_reg[2][29] ), .Z(n1623) );
  NAND U2480 ( .A(n1339), .B(n930), .Z(n2218) );
  XNOR U2481 ( .A(\min_dist_reg[2][29] ), .B(n1428), .Z(n1339) );
  IV U2482 ( .A(n1338), .Z(n1428) );
  XNOR U2483 ( .A(n2219), .B(\min_dist_reg[1][29] ), .Z(n2216) );
  IV U2484 ( .A(n2214), .Z(n2219) );
  XOR U2485 ( .A(n2220), .B(n2221), .Z(n2214) );
  AND U2486 ( .A(n2222), .B(n2223), .Z(n2221) );
  XNOR U2487 ( .A(n1626), .B(n2220), .Z(n2223) );
  XNOR U2488 ( .A(n2224), .B(\min_dist_reg[2][28] ), .Z(n1626) );
  NAND U2489 ( .A(n1342), .B(n930), .Z(n2224) );
  XNOR U2490 ( .A(\min_dist_reg[2][28] ), .B(n1434), .Z(n1342) );
  IV U2491 ( .A(n1341), .Z(n1434) );
  XNOR U2492 ( .A(n2225), .B(\min_dist_reg[1][28] ), .Z(n2222) );
  IV U2493 ( .A(n2220), .Z(n2225) );
  XOR U2494 ( .A(n2226), .B(n2227), .Z(n2220) );
  AND U2495 ( .A(n2228), .B(n2229), .Z(n2227) );
  XNOR U2496 ( .A(n1629), .B(n2226), .Z(n2229) );
  XNOR U2497 ( .A(n2230), .B(\min_dist_reg[2][27] ), .Z(n1629) );
  NAND U2498 ( .A(n1345), .B(n930), .Z(n2230) );
  XNOR U2499 ( .A(\min_dist_reg[2][27] ), .B(n1440), .Z(n1345) );
  IV U2500 ( .A(n1344), .Z(n1440) );
  XNOR U2501 ( .A(n2231), .B(\min_dist_reg[1][27] ), .Z(n2228) );
  IV U2502 ( .A(n2226), .Z(n2231) );
  XOR U2503 ( .A(n2232), .B(n2233), .Z(n2226) );
  AND U2504 ( .A(n2234), .B(n2235), .Z(n2233) );
  XNOR U2505 ( .A(n1632), .B(n2232), .Z(n2235) );
  XNOR U2506 ( .A(n2236), .B(\min_dist_reg[2][26] ), .Z(n1632) );
  NAND U2507 ( .A(n1348), .B(n930), .Z(n2236) );
  XNOR U2508 ( .A(\min_dist_reg[2][26] ), .B(n1446), .Z(n1348) );
  IV U2509 ( .A(n1347), .Z(n1446) );
  XNOR U2510 ( .A(n2237), .B(\min_dist_reg[1][26] ), .Z(n2234) );
  IV U2511 ( .A(n2232), .Z(n2237) );
  XOR U2512 ( .A(n2238), .B(n2239), .Z(n2232) );
  AND U2513 ( .A(n2240), .B(n2241), .Z(n2239) );
  XNOR U2514 ( .A(n1635), .B(n2238), .Z(n2241) );
  XNOR U2515 ( .A(n2242), .B(\min_dist_reg[2][25] ), .Z(n1635) );
  NAND U2516 ( .A(n1351), .B(n930), .Z(n2242) );
  XNOR U2517 ( .A(\min_dist_reg[2][25] ), .B(n1452), .Z(n1351) );
  IV U2518 ( .A(n1350), .Z(n1452) );
  XNOR U2519 ( .A(n2243), .B(\min_dist_reg[1][25] ), .Z(n2240) );
  IV U2520 ( .A(n2238), .Z(n2243) );
  XOR U2521 ( .A(n2244), .B(n2245), .Z(n2238) );
  AND U2522 ( .A(n2246), .B(n2247), .Z(n2245) );
  XNOR U2523 ( .A(n1638), .B(n2244), .Z(n2247) );
  XNOR U2524 ( .A(n2248), .B(\min_dist_reg[2][24] ), .Z(n1638) );
  NAND U2525 ( .A(n1354), .B(n930), .Z(n2248) );
  XNOR U2526 ( .A(\min_dist_reg[2][24] ), .B(n1458), .Z(n1354) );
  IV U2527 ( .A(n1353), .Z(n1458) );
  XNOR U2528 ( .A(n2249), .B(\min_dist_reg[1][24] ), .Z(n2246) );
  IV U2529 ( .A(n2244), .Z(n2249) );
  XOR U2530 ( .A(n2250), .B(n2251), .Z(n2244) );
  AND U2531 ( .A(n2252), .B(n2253), .Z(n2251) );
  XNOR U2532 ( .A(n1641), .B(n2250), .Z(n2253) );
  XNOR U2533 ( .A(n2254), .B(\min_dist_reg[2][23] ), .Z(n1641) );
  NAND U2534 ( .A(n1357), .B(n930), .Z(n2254) );
  XNOR U2535 ( .A(\min_dist_reg[2][23] ), .B(n1464), .Z(n1357) );
  IV U2536 ( .A(n1356), .Z(n1464) );
  XNOR U2537 ( .A(n2255), .B(\min_dist_reg[1][23] ), .Z(n2252) );
  IV U2538 ( .A(n2250), .Z(n2255) );
  XOR U2539 ( .A(n2256), .B(n2257), .Z(n2250) );
  AND U2540 ( .A(n2258), .B(n2259), .Z(n2257) );
  XNOR U2541 ( .A(n1644), .B(n2256), .Z(n2259) );
  XNOR U2542 ( .A(n2260), .B(\min_dist_reg[2][22] ), .Z(n1644) );
  NAND U2543 ( .A(n1360), .B(n930), .Z(n2260) );
  XNOR U2544 ( .A(\min_dist_reg[2][22] ), .B(n1470), .Z(n1360) );
  IV U2545 ( .A(n1359), .Z(n1470) );
  XNOR U2546 ( .A(n2261), .B(\min_dist_reg[1][22] ), .Z(n2258) );
  IV U2547 ( .A(n2256), .Z(n2261) );
  XOR U2548 ( .A(n2262), .B(n2263), .Z(n2256) );
  AND U2549 ( .A(n2264), .B(n2265), .Z(n2263) );
  XNOR U2550 ( .A(n1647), .B(n2262), .Z(n2265) );
  XNOR U2551 ( .A(n2266), .B(\min_dist_reg[2][21] ), .Z(n1647) );
  NAND U2552 ( .A(n1363), .B(n930), .Z(n2266) );
  XNOR U2553 ( .A(\min_dist_reg[2][21] ), .B(n1476), .Z(n1363) );
  IV U2554 ( .A(n1362), .Z(n1476) );
  XNOR U2555 ( .A(n2267), .B(\min_dist_reg[1][21] ), .Z(n2264) );
  IV U2556 ( .A(n2262), .Z(n2267) );
  XOR U2557 ( .A(n2268), .B(n2269), .Z(n2262) );
  AND U2558 ( .A(n2270), .B(n2271), .Z(n2269) );
  XNOR U2559 ( .A(n1650), .B(n2268), .Z(n2271) );
  XNOR U2560 ( .A(n2272), .B(\min_dist_reg[2][20] ), .Z(n1650) );
  NAND U2561 ( .A(n1366), .B(n930), .Z(n2272) );
  XNOR U2562 ( .A(\min_dist_reg[2][20] ), .B(n1482), .Z(n1366) );
  IV U2563 ( .A(n1365), .Z(n1482) );
  XNOR U2564 ( .A(n2273), .B(\min_dist_reg[1][20] ), .Z(n2270) );
  IV U2565 ( .A(n2268), .Z(n2273) );
  XOR U2566 ( .A(n2274), .B(n2275), .Z(n2268) );
  AND U2567 ( .A(n2276), .B(n2277), .Z(n2275) );
  XNOR U2568 ( .A(n1656), .B(n2274), .Z(n2277) );
  XNOR U2569 ( .A(n2278), .B(\min_dist_reg[2][19] ), .Z(n1656) );
  NAND U2570 ( .A(n1373), .B(n930), .Z(n2278) );
  XNOR U2571 ( .A(\min_dist_reg[2][19] ), .B(n1488), .Z(n1373) );
  IV U2572 ( .A(n1372), .Z(n1488) );
  XNOR U2573 ( .A(n2279), .B(\min_dist_reg[1][19] ), .Z(n2276) );
  IV U2574 ( .A(n2274), .Z(n2279) );
  XOR U2575 ( .A(n2280), .B(n2281), .Z(n2274) );
  AND U2576 ( .A(n2282), .B(n2283), .Z(n2281) );
  XNOR U2577 ( .A(n1659), .B(n2280), .Z(n2283) );
  XNOR U2578 ( .A(n2284), .B(\min_dist_reg[2][18] ), .Z(n1659) );
  NAND U2579 ( .A(n1376), .B(n930), .Z(n2284) );
  XNOR U2580 ( .A(\min_dist_reg[2][18] ), .B(n1494), .Z(n1376) );
  IV U2581 ( .A(n1375), .Z(n1494) );
  XNOR U2582 ( .A(n2285), .B(\min_dist_reg[1][18] ), .Z(n2282) );
  IV U2583 ( .A(n2280), .Z(n2285) );
  XOR U2584 ( .A(n2286), .B(n2287), .Z(n2280) );
  AND U2585 ( .A(n2288), .B(n2289), .Z(n2287) );
  XNOR U2586 ( .A(n1662), .B(n2286), .Z(n2289) );
  XNOR U2587 ( .A(n2290), .B(\min_dist_reg[2][17] ), .Z(n1662) );
  NAND U2588 ( .A(n1379), .B(n930), .Z(n2290) );
  XNOR U2589 ( .A(\min_dist_reg[2][17] ), .B(n1500), .Z(n1379) );
  IV U2590 ( .A(n1378), .Z(n1500) );
  XNOR U2591 ( .A(n2291), .B(\min_dist_reg[1][17] ), .Z(n2288) );
  IV U2592 ( .A(n2286), .Z(n2291) );
  XOR U2593 ( .A(n2292), .B(n2293), .Z(n2286) );
  AND U2594 ( .A(n2294), .B(n2295), .Z(n2293) );
  XNOR U2595 ( .A(n1665), .B(n2292), .Z(n2295) );
  XNOR U2596 ( .A(n2296), .B(\min_dist_reg[2][16] ), .Z(n1665) );
  NAND U2597 ( .A(n1382), .B(n930), .Z(n2296) );
  XNOR U2598 ( .A(\min_dist_reg[2][16] ), .B(n1506), .Z(n1382) );
  IV U2599 ( .A(n1381), .Z(n1506) );
  XNOR U2600 ( .A(n2297), .B(\min_dist_reg[1][16] ), .Z(n2294) );
  IV U2601 ( .A(n2292), .Z(n2297) );
  XOR U2602 ( .A(n2298), .B(n2299), .Z(n2292) );
  AND U2603 ( .A(n2300), .B(n2301), .Z(n2299) );
  XNOR U2604 ( .A(n1668), .B(n2298), .Z(n2301) );
  XNOR U2605 ( .A(n2302), .B(\min_dist_reg[2][15] ), .Z(n1668) );
  NAND U2606 ( .A(n1385), .B(n930), .Z(n2302) );
  XNOR U2607 ( .A(\min_dist_reg[2][15] ), .B(n1512), .Z(n1385) );
  IV U2608 ( .A(n1384), .Z(n1512) );
  XNOR U2609 ( .A(n2303), .B(\min_dist_reg[1][15] ), .Z(n2300) );
  IV U2610 ( .A(n2298), .Z(n2303) );
  XOR U2611 ( .A(n2304), .B(n2305), .Z(n2298) );
  AND U2612 ( .A(n2306), .B(n2307), .Z(n2305) );
  XNOR U2613 ( .A(n1671), .B(n2304), .Z(n2307) );
  XNOR U2614 ( .A(n2308), .B(\min_dist_reg[2][14] ), .Z(n1671) );
  NAND U2615 ( .A(n1388), .B(n930), .Z(n2308) );
  XNOR U2616 ( .A(\min_dist_reg[2][14] ), .B(n1518), .Z(n1388) );
  IV U2617 ( .A(n1387), .Z(n1518) );
  XNOR U2618 ( .A(n2309), .B(\min_dist_reg[1][14] ), .Z(n2306) );
  IV U2619 ( .A(n2304), .Z(n2309) );
  XOR U2620 ( .A(n2310), .B(n2311), .Z(n2304) );
  AND U2621 ( .A(n2312), .B(n2313), .Z(n2311) );
  XNOR U2622 ( .A(n1674), .B(n2310), .Z(n2313) );
  XNOR U2623 ( .A(n2314), .B(\min_dist_reg[2][13] ), .Z(n1674) );
  NAND U2624 ( .A(n1391), .B(n930), .Z(n2314) );
  XNOR U2625 ( .A(\min_dist_reg[2][13] ), .B(n1524), .Z(n1391) );
  IV U2626 ( .A(n1390), .Z(n1524) );
  XNOR U2627 ( .A(n2315), .B(\min_dist_reg[1][13] ), .Z(n2312) );
  IV U2628 ( .A(n2310), .Z(n2315) );
  XOR U2629 ( .A(n2316), .B(n2317), .Z(n2310) );
  AND U2630 ( .A(n2318), .B(n2319), .Z(n2317) );
  XNOR U2631 ( .A(n1677), .B(n2316), .Z(n2319) );
  XNOR U2632 ( .A(n2320), .B(\min_dist_reg[2][12] ), .Z(n1677) );
  NAND U2633 ( .A(n1394), .B(n930), .Z(n2320) );
  XNOR U2634 ( .A(\min_dist_reg[2][12] ), .B(n1530), .Z(n1394) );
  IV U2635 ( .A(n1393), .Z(n1530) );
  XNOR U2636 ( .A(n2321), .B(\min_dist_reg[1][12] ), .Z(n2318) );
  IV U2637 ( .A(n2316), .Z(n2321) );
  XOR U2638 ( .A(n2322), .B(n2323), .Z(n2316) );
  AND U2639 ( .A(n2324), .B(n2325), .Z(n2323) );
  XNOR U2640 ( .A(n1680), .B(n2322), .Z(n2325) );
  XNOR U2641 ( .A(n2326), .B(\min_dist_reg[2][11] ), .Z(n1680) );
  NAND U2642 ( .A(n1397), .B(n930), .Z(n2326) );
  XNOR U2643 ( .A(\min_dist_reg[2][11] ), .B(n1536), .Z(n1397) );
  IV U2644 ( .A(n1396), .Z(n1536) );
  XNOR U2645 ( .A(n2327), .B(\min_dist_reg[1][11] ), .Z(n2324) );
  IV U2646 ( .A(n2322), .Z(n2327) );
  XOR U2647 ( .A(n2328), .B(n2329), .Z(n2322) );
  AND U2648 ( .A(n2330), .B(n2331), .Z(n2329) );
  XNOR U2649 ( .A(n1683), .B(n2328), .Z(n2331) );
  XNOR U2650 ( .A(n2332), .B(\min_dist_reg[2][10] ), .Z(n1683) );
  NAND U2651 ( .A(n1400), .B(n930), .Z(n2332) );
  XNOR U2652 ( .A(\min_dist_reg[2][10] ), .B(n1542), .Z(n1400) );
  IV U2653 ( .A(n1399), .Z(n1542) );
  XNOR U2654 ( .A(n2333), .B(\min_dist_reg[1][10] ), .Z(n2330) );
  IV U2655 ( .A(n2328), .Z(n2333) );
  XOR U2656 ( .A(n2334), .B(n2335), .Z(n2328) );
  AND U2657 ( .A(n2336), .B(n2337), .Z(n2335) );
  XNOR U2658 ( .A(n1587), .B(n2334), .Z(n2337) );
  XNOR U2659 ( .A(n2338), .B(\min_dist_reg[2][9] ), .Z(n1587) );
  NAND U2660 ( .A(n1302), .B(n930), .Z(n2338) );
  XNOR U2661 ( .A(\min_dist_reg[2][9] ), .B(n1548), .Z(n1302) );
  IV U2662 ( .A(n1301), .Z(n1548) );
  XNOR U2663 ( .A(n2339), .B(\min_dist_reg[1][9] ), .Z(n2336) );
  IV U2664 ( .A(n2334), .Z(n2339) );
  XOR U2665 ( .A(n2340), .B(n2341), .Z(n2334) );
  AND U2666 ( .A(n2342), .B(n2343), .Z(n2341) );
  XNOR U2667 ( .A(n1590), .B(n2340), .Z(n2343) );
  XNOR U2668 ( .A(n2344), .B(\min_dist_reg[2][8] ), .Z(n1590) );
  NAND U2669 ( .A(n1305), .B(n930), .Z(n2344) );
  XNOR U2670 ( .A(\min_dist_reg[2][8] ), .B(n1554), .Z(n1305) );
  IV U2671 ( .A(n1304), .Z(n1554) );
  XNOR U2672 ( .A(n2345), .B(\min_dist_reg[1][8] ), .Z(n2342) );
  IV U2673 ( .A(n2340), .Z(n2345) );
  XOR U2674 ( .A(n2346), .B(n2347), .Z(n2340) );
  AND U2675 ( .A(n2348), .B(n2349), .Z(n2347) );
  XNOR U2676 ( .A(n1593), .B(n2346), .Z(n2349) );
  XNOR U2677 ( .A(n2350), .B(\min_dist_reg[2][7] ), .Z(n1593) );
  NAND U2678 ( .A(n1308), .B(n930), .Z(n2350) );
  XNOR U2679 ( .A(\min_dist_reg[2][7] ), .B(n1560), .Z(n1308) );
  IV U2680 ( .A(n1307), .Z(n1560) );
  XNOR U2681 ( .A(n2351), .B(\min_dist_reg[1][7] ), .Z(n2348) );
  IV U2682 ( .A(n2346), .Z(n2351) );
  XOR U2683 ( .A(n2352), .B(n2353), .Z(n2346) );
  AND U2684 ( .A(n2354), .B(n2355), .Z(n2353) );
  XNOR U2685 ( .A(n1596), .B(n2352), .Z(n2355) );
  XNOR U2686 ( .A(n2356), .B(\min_dist_reg[2][6] ), .Z(n1596) );
  NAND U2687 ( .A(n1311), .B(n930), .Z(n2356) );
  XNOR U2688 ( .A(\min_dist_reg[2][6] ), .B(n1566), .Z(n1311) );
  IV U2689 ( .A(n1310), .Z(n1566) );
  XNOR U2690 ( .A(n2357), .B(\min_dist_reg[1][6] ), .Z(n2354) );
  IV U2691 ( .A(n2352), .Z(n2357) );
  XOR U2692 ( .A(n2358), .B(n2359), .Z(n2352) );
  AND U2693 ( .A(n2360), .B(n2361), .Z(n2359) );
  XNOR U2694 ( .A(n1599), .B(n2358), .Z(n2361) );
  XNOR U2695 ( .A(n2362), .B(\min_dist_reg[2][5] ), .Z(n1599) );
  NAND U2696 ( .A(n1314), .B(n930), .Z(n2362) );
  XNOR U2697 ( .A(\min_dist_reg[2][5] ), .B(n1572), .Z(n1314) );
  IV U2698 ( .A(n1313), .Z(n1572) );
  XNOR U2699 ( .A(n2363), .B(\min_dist_reg[1][5] ), .Z(n2360) );
  IV U2700 ( .A(n2358), .Z(n2363) );
  XOR U2701 ( .A(n2364), .B(n2365), .Z(n2358) );
  AND U2702 ( .A(n2366), .B(n2367), .Z(n2365) );
  XNOR U2703 ( .A(n1602), .B(n2364), .Z(n2367) );
  XNOR U2704 ( .A(n2368), .B(\min_dist_reg[2][4] ), .Z(n1602) );
  NAND U2705 ( .A(n1317), .B(n930), .Z(n2368) );
  XNOR U2706 ( .A(\min_dist_reg[2][4] ), .B(n1578), .Z(n1317) );
  IV U2707 ( .A(n1316), .Z(n1578) );
  XNOR U2708 ( .A(n2369), .B(\min_dist_reg[1][4] ), .Z(n2366) );
  IV U2709 ( .A(n2364), .Z(n2369) );
  XOR U2710 ( .A(n2370), .B(n2371), .Z(n2364) );
  AND U2711 ( .A(n2372), .B(n2373), .Z(n2371) );
  XNOR U2712 ( .A(n1605), .B(n2370), .Z(n2373) );
  XNOR U2713 ( .A(n2374), .B(\min_dist_reg[2][3] ), .Z(n1605) );
  NAND U2714 ( .A(n1320), .B(n930), .Z(n2374) );
  XNOR U2715 ( .A(\min_dist_reg[2][3] ), .B(n1584), .Z(n1320) );
  IV U2716 ( .A(n1319), .Z(n1584) );
  XNOR U2717 ( .A(n2375), .B(\min_dist_reg[1][3] ), .Z(n2372) );
  IV U2718 ( .A(n2370), .Z(n2375) );
  XOR U2719 ( .A(n2376), .B(n2377), .Z(n2370) );
  AND U2720 ( .A(n2378), .B(n2379), .Z(n2377) );
  XNOR U2721 ( .A(n1620), .B(n2376), .Z(n2379) );
  XNOR U2722 ( .A(n2380), .B(\min_dist_reg[2][2] ), .Z(n1620) );
  NAND U2723 ( .A(n2381), .B(n930), .Z(n2380) );
  XNOR U2724 ( .A(n2382), .B(n1334), .Z(n2381) );
  XNOR U2725 ( .A(n2376), .B(n2181), .Z(n2378) );
  IV U2726 ( .A(\min_dist_reg[1][2] ), .Z(n2181) );
  XOR U2727 ( .A(n2383), .B(n2384), .Z(n2376) );
  NAND U2728 ( .A(n2385), .B(n2386), .Z(n2383) );
  XOR U2729 ( .A(n2384), .B(n1653), .Z(n2386) );
  XNOR U2730 ( .A(n2387), .B(\min_dist_reg[2][1] ), .Z(n1653) );
  NAND U2731 ( .A(n2388), .B(n930), .Z(n2387) );
  XNOR U2732 ( .A(n2389), .B(n1368), .Z(n2388) );
  XOR U2733 ( .A(n2384), .B(n2188), .Z(n2385) );
  IV U2734 ( .A(\min_dist_reg[1][1] ), .Z(n2188) );
  AND U2735 ( .A(n1686), .B(n2390), .Z(n2384) );
  XNOR U2736 ( .A(n2390), .B(n1686), .Z(n1687) );
  XNOR U2737 ( .A(n2391), .B(\min_dist_reg[2][0] ), .Z(n1686) );
  NAND U2738 ( .A(n1403), .B(n930), .Z(n2391) );
  XNOR U2739 ( .A(n2392), .B(n2393), .Z(n930) );
  AND U2740 ( .A(n2394), .B(n2395), .Z(n2393) );
  XNOR U2741 ( .A(n2396), .B(n1322), .Z(n2395) );
  XNOR U2742 ( .A(n2397), .B(\min_dist_reg[3][33] ), .Z(n1322) );
  NAND U2743 ( .A(n2398), .B(n933), .Z(n2397) );
  XOR U2744 ( .A(\min_dist_reg[3][33] ), .B(n2399), .Z(n2398) );
  XNOR U2745 ( .A(n2392), .B(\min_dist_reg[2][33] ), .Z(n2394) );
  IV U2746 ( .A(n2396), .Z(n2392) );
  XOR U2747 ( .A(n2400), .B(n2401), .Z(n2396) );
  AND U2748 ( .A(n2402), .B(n2403), .Z(n2401) );
  XNOR U2749 ( .A(n2400), .B(n1325), .Z(n2403) );
  XNOR U2750 ( .A(n2404), .B(\min_dist_reg[3][32] ), .Z(n1325) );
  NAND U2751 ( .A(n2405), .B(n933), .Z(n2404) );
  XOR U2752 ( .A(\min_dist_reg[3][32] ), .B(n2406), .Z(n2405) );
  XNOR U2753 ( .A(n2407), .B(\min_dist_reg[2][32] ), .Z(n2402) );
  IV U2754 ( .A(n2400), .Z(n2407) );
  XOR U2755 ( .A(n2408), .B(n2409), .Z(n2400) );
  AND U2756 ( .A(n2410), .B(n2411), .Z(n2409) );
  XNOR U2757 ( .A(n2408), .B(n1328), .Z(n2411) );
  XNOR U2758 ( .A(n2412), .B(\min_dist_reg[3][31] ), .Z(n1328) );
  NAND U2759 ( .A(n2413), .B(n933), .Z(n2412) );
  XOR U2760 ( .A(\min_dist_reg[3][31] ), .B(n2414), .Z(n2413) );
  XNOR U2761 ( .A(n2415), .B(\min_dist_reg[2][31] ), .Z(n2410) );
  IV U2762 ( .A(n2408), .Z(n2415) );
  XOR U2763 ( .A(n2416), .B(n2417), .Z(n2408) );
  AND U2764 ( .A(n2418), .B(n2419), .Z(n2417) );
  XNOR U2765 ( .A(n2416), .B(n1331), .Z(n2419) );
  XNOR U2766 ( .A(n2420), .B(\min_dist_reg[3][30] ), .Z(n1331) );
  NAND U2767 ( .A(n2421), .B(n933), .Z(n2420) );
  XOR U2768 ( .A(\min_dist_reg[3][30] ), .B(n2422), .Z(n2421) );
  XNOR U2769 ( .A(n2423), .B(\min_dist_reg[2][30] ), .Z(n2418) );
  IV U2770 ( .A(n2416), .Z(n2423) );
  XOR U2771 ( .A(n2424), .B(n2425), .Z(n2416) );
  AND U2772 ( .A(n2426), .B(n2427), .Z(n2425) );
  XNOR U2773 ( .A(n2424), .B(n1338), .Z(n2427) );
  XNOR U2774 ( .A(n2428), .B(\min_dist_reg[3][29] ), .Z(n1338) );
  NAND U2775 ( .A(n2429), .B(n933), .Z(n2428) );
  XOR U2776 ( .A(\min_dist_reg[3][29] ), .B(n2430), .Z(n2429) );
  XNOR U2777 ( .A(n2431), .B(\min_dist_reg[2][29] ), .Z(n2426) );
  IV U2778 ( .A(n2424), .Z(n2431) );
  XOR U2779 ( .A(n2432), .B(n2433), .Z(n2424) );
  AND U2780 ( .A(n2434), .B(n2435), .Z(n2433) );
  XNOR U2781 ( .A(n2432), .B(n1341), .Z(n2435) );
  XNOR U2782 ( .A(n2436), .B(\min_dist_reg[3][28] ), .Z(n1341) );
  NAND U2783 ( .A(n2437), .B(n933), .Z(n2436) );
  XOR U2784 ( .A(\min_dist_reg[3][28] ), .B(n2438), .Z(n2437) );
  XNOR U2785 ( .A(n2439), .B(\min_dist_reg[2][28] ), .Z(n2434) );
  IV U2786 ( .A(n2432), .Z(n2439) );
  XOR U2787 ( .A(n2440), .B(n2441), .Z(n2432) );
  AND U2788 ( .A(n2442), .B(n2443), .Z(n2441) );
  XNOR U2789 ( .A(n2440), .B(n1344), .Z(n2443) );
  XNOR U2790 ( .A(n2444), .B(\min_dist_reg[3][27] ), .Z(n1344) );
  NAND U2791 ( .A(n2445), .B(n933), .Z(n2444) );
  XOR U2792 ( .A(\min_dist_reg[3][27] ), .B(n2446), .Z(n2445) );
  XNOR U2793 ( .A(n2447), .B(\min_dist_reg[2][27] ), .Z(n2442) );
  IV U2794 ( .A(n2440), .Z(n2447) );
  XOR U2795 ( .A(n2448), .B(n2449), .Z(n2440) );
  AND U2796 ( .A(n2450), .B(n2451), .Z(n2449) );
  XNOR U2797 ( .A(n2448), .B(n1347), .Z(n2451) );
  XNOR U2798 ( .A(n2452), .B(\min_dist_reg[3][26] ), .Z(n1347) );
  NAND U2799 ( .A(n2453), .B(n933), .Z(n2452) );
  XOR U2800 ( .A(\min_dist_reg[3][26] ), .B(n2454), .Z(n2453) );
  XNOR U2801 ( .A(n2455), .B(\min_dist_reg[2][26] ), .Z(n2450) );
  IV U2802 ( .A(n2448), .Z(n2455) );
  XOR U2803 ( .A(n2456), .B(n2457), .Z(n2448) );
  AND U2804 ( .A(n2458), .B(n2459), .Z(n2457) );
  XNOR U2805 ( .A(n2456), .B(n1350), .Z(n2459) );
  XNOR U2806 ( .A(n2460), .B(\min_dist_reg[3][25] ), .Z(n1350) );
  NAND U2807 ( .A(n2461), .B(n933), .Z(n2460) );
  XOR U2808 ( .A(\min_dist_reg[3][25] ), .B(n2462), .Z(n2461) );
  XNOR U2809 ( .A(n2463), .B(\min_dist_reg[2][25] ), .Z(n2458) );
  IV U2810 ( .A(n2456), .Z(n2463) );
  XOR U2811 ( .A(n2464), .B(n2465), .Z(n2456) );
  AND U2812 ( .A(n2466), .B(n2467), .Z(n2465) );
  XNOR U2813 ( .A(n2464), .B(n1353), .Z(n2467) );
  XNOR U2814 ( .A(n2468), .B(\min_dist_reg[3][24] ), .Z(n1353) );
  NAND U2815 ( .A(n2469), .B(n933), .Z(n2468) );
  XOR U2816 ( .A(\min_dist_reg[3][24] ), .B(n2470), .Z(n2469) );
  XNOR U2817 ( .A(n2471), .B(\min_dist_reg[2][24] ), .Z(n2466) );
  IV U2818 ( .A(n2464), .Z(n2471) );
  XOR U2819 ( .A(n2472), .B(n2473), .Z(n2464) );
  AND U2820 ( .A(n2474), .B(n2475), .Z(n2473) );
  XNOR U2821 ( .A(n2472), .B(n1356), .Z(n2475) );
  XNOR U2822 ( .A(n2476), .B(\min_dist_reg[3][23] ), .Z(n1356) );
  NAND U2823 ( .A(n2477), .B(n933), .Z(n2476) );
  XOR U2824 ( .A(\min_dist_reg[3][23] ), .B(n2478), .Z(n2477) );
  XNOR U2825 ( .A(n2479), .B(\min_dist_reg[2][23] ), .Z(n2474) );
  IV U2826 ( .A(n2472), .Z(n2479) );
  XOR U2827 ( .A(n2480), .B(n2481), .Z(n2472) );
  AND U2828 ( .A(n2482), .B(n2483), .Z(n2481) );
  XNOR U2829 ( .A(n2480), .B(n1359), .Z(n2483) );
  XNOR U2830 ( .A(n2484), .B(\min_dist_reg[3][22] ), .Z(n1359) );
  NAND U2831 ( .A(n2485), .B(n933), .Z(n2484) );
  XOR U2832 ( .A(\min_dist_reg[3][22] ), .B(n2486), .Z(n2485) );
  XNOR U2833 ( .A(n2487), .B(\min_dist_reg[2][22] ), .Z(n2482) );
  IV U2834 ( .A(n2480), .Z(n2487) );
  XOR U2835 ( .A(n2488), .B(n2489), .Z(n2480) );
  AND U2836 ( .A(n2490), .B(n2491), .Z(n2489) );
  XNOR U2837 ( .A(n2488), .B(n1362), .Z(n2491) );
  XNOR U2838 ( .A(n2492), .B(\min_dist_reg[3][21] ), .Z(n1362) );
  NAND U2839 ( .A(n2493), .B(n933), .Z(n2492) );
  XOR U2840 ( .A(\min_dist_reg[3][21] ), .B(n2494), .Z(n2493) );
  XNOR U2841 ( .A(n2495), .B(\min_dist_reg[2][21] ), .Z(n2490) );
  IV U2842 ( .A(n2488), .Z(n2495) );
  XOR U2843 ( .A(n2496), .B(n2497), .Z(n2488) );
  AND U2844 ( .A(n2498), .B(n2499), .Z(n2497) );
  XNOR U2845 ( .A(n2496), .B(n1365), .Z(n2499) );
  XNOR U2846 ( .A(n2500), .B(\min_dist_reg[3][20] ), .Z(n1365) );
  NAND U2847 ( .A(n2501), .B(n933), .Z(n2500) );
  XOR U2848 ( .A(\min_dist_reg[3][20] ), .B(n2502), .Z(n2501) );
  XNOR U2849 ( .A(n2503), .B(\min_dist_reg[2][20] ), .Z(n2498) );
  IV U2850 ( .A(n2496), .Z(n2503) );
  XOR U2851 ( .A(n2504), .B(n2505), .Z(n2496) );
  AND U2852 ( .A(n2506), .B(n2507), .Z(n2505) );
  XNOR U2853 ( .A(n2504), .B(n1372), .Z(n2507) );
  XNOR U2854 ( .A(n2508), .B(\min_dist_reg[3][19] ), .Z(n1372) );
  NAND U2855 ( .A(n2509), .B(n933), .Z(n2508) );
  XOR U2856 ( .A(\min_dist_reg[3][19] ), .B(n2510), .Z(n2509) );
  XNOR U2857 ( .A(n2511), .B(\min_dist_reg[2][19] ), .Z(n2506) );
  IV U2858 ( .A(n2504), .Z(n2511) );
  XOR U2859 ( .A(n2512), .B(n2513), .Z(n2504) );
  AND U2860 ( .A(n2514), .B(n2515), .Z(n2513) );
  XNOR U2861 ( .A(n2512), .B(n1375), .Z(n2515) );
  XNOR U2862 ( .A(n2516), .B(\min_dist_reg[3][18] ), .Z(n1375) );
  NAND U2863 ( .A(n2517), .B(n933), .Z(n2516) );
  XOR U2864 ( .A(\min_dist_reg[3][18] ), .B(n2518), .Z(n2517) );
  XNOR U2865 ( .A(n2519), .B(\min_dist_reg[2][18] ), .Z(n2514) );
  IV U2866 ( .A(n2512), .Z(n2519) );
  XOR U2867 ( .A(n2520), .B(n2521), .Z(n2512) );
  AND U2868 ( .A(n2522), .B(n2523), .Z(n2521) );
  XNOR U2869 ( .A(n2520), .B(n1378), .Z(n2523) );
  XNOR U2870 ( .A(n2524), .B(\min_dist_reg[3][17] ), .Z(n1378) );
  NAND U2871 ( .A(n2525), .B(n933), .Z(n2524) );
  XOR U2872 ( .A(\min_dist_reg[3][17] ), .B(n2526), .Z(n2525) );
  XNOR U2873 ( .A(n2527), .B(\min_dist_reg[2][17] ), .Z(n2522) );
  IV U2874 ( .A(n2520), .Z(n2527) );
  XOR U2875 ( .A(n2528), .B(n2529), .Z(n2520) );
  AND U2876 ( .A(n2530), .B(n2531), .Z(n2529) );
  XNOR U2877 ( .A(n2528), .B(n1381), .Z(n2531) );
  XNOR U2878 ( .A(n2532), .B(\min_dist_reg[3][16] ), .Z(n1381) );
  NAND U2879 ( .A(n2533), .B(n933), .Z(n2532) );
  XOR U2880 ( .A(\min_dist_reg[3][16] ), .B(n2534), .Z(n2533) );
  XNOR U2881 ( .A(n2535), .B(\min_dist_reg[2][16] ), .Z(n2530) );
  IV U2882 ( .A(n2528), .Z(n2535) );
  XOR U2883 ( .A(n2536), .B(n2537), .Z(n2528) );
  AND U2884 ( .A(n2538), .B(n2539), .Z(n2537) );
  XNOR U2885 ( .A(n2536), .B(n1384), .Z(n2539) );
  XNOR U2886 ( .A(n2540), .B(\min_dist_reg[3][15] ), .Z(n1384) );
  NAND U2887 ( .A(n2541), .B(n933), .Z(n2540) );
  XOR U2888 ( .A(\min_dist_reg[3][15] ), .B(n2542), .Z(n2541) );
  XNOR U2889 ( .A(n2543), .B(\min_dist_reg[2][15] ), .Z(n2538) );
  IV U2890 ( .A(n2536), .Z(n2543) );
  XOR U2891 ( .A(n2544), .B(n2545), .Z(n2536) );
  AND U2892 ( .A(n2546), .B(n2547), .Z(n2545) );
  XNOR U2893 ( .A(n2544), .B(n1387), .Z(n2547) );
  XNOR U2894 ( .A(n2548), .B(\min_dist_reg[3][14] ), .Z(n1387) );
  NAND U2895 ( .A(n2549), .B(n933), .Z(n2548) );
  XOR U2896 ( .A(\min_dist_reg[3][14] ), .B(n2550), .Z(n2549) );
  XNOR U2897 ( .A(n2551), .B(\min_dist_reg[2][14] ), .Z(n2546) );
  IV U2898 ( .A(n2544), .Z(n2551) );
  XOR U2899 ( .A(n2552), .B(n2553), .Z(n2544) );
  AND U2900 ( .A(n2554), .B(n2555), .Z(n2553) );
  XNOR U2901 ( .A(n2552), .B(n1390), .Z(n2555) );
  XNOR U2902 ( .A(n2556), .B(\min_dist_reg[3][13] ), .Z(n1390) );
  NAND U2903 ( .A(n2557), .B(n933), .Z(n2556) );
  XOR U2904 ( .A(\min_dist_reg[3][13] ), .B(n2558), .Z(n2557) );
  XNOR U2905 ( .A(n2559), .B(\min_dist_reg[2][13] ), .Z(n2554) );
  IV U2906 ( .A(n2552), .Z(n2559) );
  XOR U2907 ( .A(n2560), .B(n2561), .Z(n2552) );
  AND U2908 ( .A(n2562), .B(n2563), .Z(n2561) );
  XNOR U2909 ( .A(n2560), .B(n1393), .Z(n2563) );
  XNOR U2910 ( .A(n2564), .B(\min_dist_reg[3][12] ), .Z(n1393) );
  NAND U2911 ( .A(n2565), .B(n933), .Z(n2564) );
  XOR U2912 ( .A(\min_dist_reg[3][12] ), .B(n2566), .Z(n2565) );
  XNOR U2913 ( .A(n2567), .B(\min_dist_reg[2][12] ), .Z(n2562) );
  IV U2914 ( .A(n2560), .Z(n2567) );
  XOR U2915 ( .A(n2568), .B(n2569), .Z(n2560) );
  AND U2916 ( .A(n2570), .B(n2571), .Z(n2569) );
  XNOR U2917 ( .A(n2568), .B(n1396), .Z(n2571) );
  XNOR U2918 ( .A(n2572), .B(\min_dist_reg[3][11] ), .Z(n1396) );
  NAND U2919 ( .A(n2573), .B(n933), .Z(n2572) );
  XOR U2920 ( .A(\min_dist_reg[3][11] ), .B(n2574), .Z(n2573) );
  XNOR U2921 ( .A(n2575), .B(\min_dist_reg[2][11] ), .Z(n2570) );
  IV U2922 ( .A(n2568), .Z(n2575) );
  XOR U2923 ( .A(n2576), .B(n2577), .Z(n2568) );
  AND U2924 ( .A(n2578), .B(n2579), .Z(n2577) );
  XNOR U2925 ( .A(n2576), .B(n1399), .Z(n2579) );
  XNOR U2926 ( .A(n2580), .B(\min_dist_reg[3][10] ), .Z(n1399) );
  NAND U2927 ( .A(n2581), .B(n933), .Z(n2580) );
  XOR U2928 ( .A(\min_dist_reg[3][10] ), .B(n2582), .Z(n2581) );
  XNOR U2929 ( .A(n2583), .B(\min_dist_reg[2][10] ), .Z(n2578) );
  IV U2930 ( .A(n2576), .Z(n2583) );
  XOR U2931 ( .A(n2584), .B(n2585), .Z(n2576) );
  AND U2932 ( .A(n2586), .B(n2587), .Z(n2585) );
  XNOR U2933 ( .A(n2584), .B(n1301), .Z(n2587) );
  XNOR U2934 ( .A(n2588), .B(\min_dist_reg[3][9] ), .Z(n1301) );
  NAND U2935 ( .A(n2589), .B(n933), .Z(n2588) );
  XOR U2936 ( .A(\min_dist_reg[3][9] ), .B(n2590), .Z(n2589) );
  XNOR U2937 ( .A(n2591), .B(\min_dist_reg[2][9] ), .Z(n2586) );
  IV U2938 ( .A(n2584), .Z(n2591) );
  XOR U2939 ( .A(n2592), .B(n2593), .Z(n2584) );
  AND U2940 ( .A(n2594), .B(n2595), .Z(n2593) );
  XNOR U2941 ( .A(n2592), .B(n1304), .Z(n2595) );
  XNOR U2942 ( .A(n2596), .B(\min_dist_reg[3][8] ), .Z(n1304) );
  NAND U2943 ( .A(n2597), .B(n933), .Z(n2596) );
  XOR U2944 ( .A(\min_dist_reg[3][8] ), .B(n2598), .Z(n2597) );
  XNOR U2945 ( .A(n2599), .B(\min_dist_reg[2][8] ), .Z(n2594) );
  IV U2946 ( .A(n2592), .Z(n2599) );
  XOR U2947 ( .A(n2600), .B(n2601), .Z(n2592) );
  AND U2948 ( .A(n2602), .B(n2603), .Z(n2601) );
  XNOR U2949 ( .A(n2600), .B(n1307), .Z(n2603) );
  XNOR U2950 ( .A(n2604), .B(\min_dist_reg[3][7] ), .Z(n1307) );
  NAND U2951 ( .A(n2605), .B(n933), .Z(n2604) );
  XOR U2952 ( .A(\min_dist_reg[3][7] ), .B(n2606), .Z(n2605) );
  XNOR U2953 ( .A(n2607), .B(\min_dist_reg[2][7] ), .Z(n2602) );
  IV U2954 ( .A(n2600), .Z(n2607) );
  XOR U2955 ( .A(n2608), .B(n2609), .Z(n2600) );
  AND U2956 ( .A(n2610), .B(n2611), .Z(n2609) );
  XNOR U2957 ( .A(n2608), .B(n1310), .Z(n2611) );
  XNOR U2958 ( .A(n2612), .B(\min_dist_reg[3][6] ), .Z(n1310) );
  NAND U2959 ( .A(n2613), .B(n933), .Z(n2612) );
  XOR U2960 ( .A(\min_dist_reg[3][6] ), .B(n2614), .Z(n2613) );
  XNOR U2961 ( .A(n2615), .B(\min_dist_reg[2][6] ), .Z(n2610) );
  IV U2962 ( .A(n2608), .Z(n2615) );
  XOR U2963 ( .A(n2616), .B(n2617), .Z(n2608) );
  AND U2964 ( .A(n2618), .B(n2619), .Z(n2617) );
  XNOR U2965 ( .A(n2616), .B(n1313), .Z(n2619) );
  XNOR U2966 ( .A(n2620), .B(\min_dist_reg[3][5] ), .Z(n1313) );
  NAND U2967 ( .A(n2621), .B(n933), .Z(n2620) );
  XOR U2968 ( .A(\min_dist_reg[3][5] ), .B(n2622), .Z(n2621) );
  XNOR U2969 ( .A(n2623), .B(\min_dist_reg[2][5] ), .Z(n2618) );
  IV U2970 ( .A(n2616), .Z(n2623) );
  XOR U2971 ( .A(n2624), .B(n2625), .Z(n2616) );
  AND U2972 ( .A(n2626), .B(n2627), .Z(n2625) );
  XNOR U2973 ( .A(n2624), .B(n1316), .Z(n2627) );
  XNOR U2974 ( .A(n2628), .B(\min_dist_reg[3][4] ), .Z(n1316) );
  NAND U2975 ( .A(n2629), .B(n933), .Z(n2628) );
  XOR U2976 ( .A(\min_dist_reg[3][4] ), .B(n2630), .Z(n2629) );
  XNOR U2977 ( .A(n2631), .B(\min_dist_reg[2][4] ), .Z(n2626) );
  IV U2978 ( .A(n2624), .Z(n2631) );
  XOR U2979 ( .A(n1580), .B(n2632), .Z(n2624) );
  AND U2980 ( .A(n1582), .B(n2633), .Z(n2632) );
  XNOR U2981 ( .A(n1580), .B(n1319), .Z(n2633) );
  XNOR U2982 ( .A(n2634), .B(\min_dist_reg[3][3] ), .Z(n1319) );
  NAND U2983 ( .A(n2635), .B(n933), .Z(n2634) );
  XOR U2984 ( .A(\min_dist_reg[3][3] ), .B(n2636), .Z(n2635) );
  XNOR U2985 ( .A(n1585), .B(\min_dist_reg[2][3] ), .Z(n1582) );
  IV U2986 ( .A(n1580), .Z(n1585) );
  XOR U2987 ( .A(n2637), .B(n2638), .Z(n1580) );
  AND U2988 ( .A(n2639), .B(n2640), .Z(n2638) );
  XOR U2989 ( .A(n1336), .B(n2637), .Z(n2640) );
  IV U2990 ( .A(n1334), .Z(n1336) );
  XNOR U2991 ( .A(n2641), .B(\min_dist_reg[3][2] ), .Z(n1334) );
  NAND U2992 ( .A(n2642), .B(n933), .Z(n2641) );
  XOR U2993 ( .A(\min_dist_reg[3][2] ), .B(n2643), .Z(n2642) );
  XNOR U2994 ( .A(n2637), .B(n2382), .Z(n2639) );
  IV U2995 ( .A(\min_dist_reg[2][2] ), .Z(n2382) );
  XOR U2996 ( .A(n2644), .B(n2645), .Z(n2637) );
  NAND U2997 ( .A(n2646), .B(n2647), .Z(n2644) );
  XNOR U2998 ( .A(n2645), .B(n1370), .Z(n2647) );
  IV U2999 ( .A(n1368), .Z(n1370) );
  XNOR U3000 ( .A(n2648), .B(\min_dist_reg[3][1] ), .Z(n1368) );
  NAND U3001 ( .A(n2649), .B(n933), .Z(n2648) );
  XOR U3002 ( .A(\min_dist_reg[3][1] ), .B(n2650), .Z(n2649) );
  XOR U3003 ( .A(n2645), .B(n2389), .Z(n2646) );
  IV U3004 ( .A(\min_dist_reg[2][1] ), .Z(n2389) );
  ANDN U3005 ( .A(n1402), .B(\min_dist_reg[2][0] ), .Z(n2645) );
  XOR U3006 ( .A(\min_dist_reg[2][0] ), .B(n1402), .Z(n1403) );
  XOR U3007 ( .A(n2651), .B(n2652), .Z(n1402) );
  NAND U3008 ( .A(n2653), .B(n933), .Z(n2651) );
  XNOR U3009 ( .A(n2654), .B(n2655), .Z(n933) );
  AND U3010 ( .A(n2656), .B(n2657), .Z(n2655) );
  XNOR U3011 ( .A(n2658), .B(n2399), .Z(n2657) );
  XOR U3012 ( .A(n2659), .B(n2660), .Z(n2399) );
  ANDN U3013 ( .A(n2661), .B(n2662), .Z(n2660) );
  XNOR U3014 ( .A(n2663), .B(n2659), .Z(n2661) );
  XNOR U3015 ( .A(n2654), .B(\min_dist_reg[3][33] ), .Z(n2656) );
  IV U3016 ( .A(n2658), .Z(n2654) );
  XOR U3017 ( .A(n2664), .B(n2665), .Z(n2658) );
  AND U3018 ( .A(n2666), .B(n2667), .Z(n2665) );
  XNOR U3019 ( .A(n2664), .B(n2406), .Z(n2667) );
  XNOR U3020 ( .A(n2668), .B(n2663), .Z(n2406) );
  NAND U3021 ( .A(n2669), .B(n2670), .Z(n2663) );
  XOR U3022 ( .A(n2671), .B(n2672), .Z(n2669) );
  AND U3023 ( .A(n2673), .B(n2674), .Z(n2671) );
  XOR U3024 ( .A(e_input[31]), .B(n2672), .Z(n2674) );
  IV U3025 ( .A(n2662), .Z(n2668) );
  XNOR U3026 ( .A(n2659), .B(n2675), .Z(n2662) );
  AND U3027 ( .A(n2676), .B(n2677), .Z(n2675) );
  XOR U3028 ( .A(n2678), .B(n2679), .Z(n2677) );
  AND U3029 ( .A(n2680), .B(n2681), .Z(n2678) );
  XOR U3030 ( .A(e_input[63]), .B(n2679), .Z(n2681) );
  XNOR U3031 ( .A(n2682), .B(n2683), .Z(n2659) );
  ANDN U3032 ( .A(n2684), .B(n2685), .Z(n2683) );
  XOR U3033 ( .A(n2682), .B(n2686), .Z(n2684) );
  XNOR U3034 ( .A(n2687), .B(\min_dist_reg[3][32] ), .Z(n2666) );
  IV U3035 ( .A(n2664), .Z(n2687) );
  XOR U3036 ( .A(n2688), .B(n2689), .Z(n2664) );
  AND U3037 ( .A(n2690), .B(n2691), .Z(n2689) );
  XNOR U3038 ( .A(n2688), .B(n2414), .Z(n2691) );
  XOR U3039 ( .A(n2686), .B(n2685), .Z(n2414) );
  XNOR U3040 ( .A(n2692), .B(n2693), .Z(n2685) );
  XNOR U3041 ( .A(n2694), .B(n2695), .Z(n2692) );
  AND U3042 ( .A(n2676), .B(n2696), .Z(n2695) );
  XNOR U3043 ( .A(n2697), .B(n2680), .Z(n2696) );
  XOR U3044 ( .A(n2679), .B(n2698), .Z(n2680) );
  XOR U3045 ( .A(n2699), .B(n2700), .Z(n2679) );
  AND U3046 ( .A(n2701), .B(n2702), .Z(n2700) );
  XOR U3047 ( .A(e_input[62]), .B(n2699), .Z(n2702) );
  NOR U3048 ( .A(e_input[63]), .B(n2693), .Z(n2697) );
  XNOR U3049 ( .A(n2703), .B(g_input[63]), .Z(n2693) );
  IV U3050 ( .A(n2682), .Z(n2694) );
  XOR U3051 ( .A(n2704), .B(n2705), .Z(n2682) );
  ANDN U3052 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U3053 ( .A(n2704), .B(n2708), .Z(n2706) );
  XOR U3054 ( .A(n2709), .B(n2710), .Z(n2686) );
  AND U3055 ( .A(n2670), .B(n2711), .Z(n2710) );
  XNOR U3056 ( .A(n2712), .B(n2673), .Z(n2711) );
  XOR U3057 ( .A(n2672), .B(n2713), .Z(n2673) );
  XOR U3058 ( .A(n2714), .B(n2715), .Z(n2672) );
  AND U3059 ( .A(n2716), .B(n2717), .Z(n2715) );
  XOR U3060 ( .A(e_input[30]), .B(n2714), .Z(n2717) );
  NOR U3061 ( .A(e_input[31]), .B(n2709), .Z(n2712) );
  XNOR U3062 ( .A(n2718), .B(g_input[31]), .Z(n2709) );
  XNOR U3063 ( .A(n2719), .B(\min_dist_reg[3][31] ), .Z(n2690) );
  IV U3064 ( .A(n2688), .Z(n2719) );
  XOR U3065 ( .A(n2720), .B(n2721), .Z(n2688) );
  AND U3066 ( .A(n2722), .B(n2723), .Z(n2721) );
  XNOR U3067 ( .A(n2720), .B(n2422), .Z(n2723) );
  XOR U3068 ( .A(n2708), .B(n2707), .Z(n2422) );
  XNOR U3069 ( .A(n2724), .B(n2725), .Z(n2707) );
  XNOR U3070 ( .A(n2726), .B(n2727), .Z(n2724) );
  AND U3071 ( .A(n2676), .B(n2728), .Z(n2727) );
  XNOR U3072 ( .A(n2701), .B(n2729), .Z(n2728) );
  XOR U3073 ( .A(n2730), .B(n2725), .Z(n2729) );
  XNOR U3074 ( .A(n2731), .B(g_input[62]), .Z(n2725) );
  IV U3075 ( .A(e_input[62]), .Z(n2730) );
  XNOR U3076 ( .A(n2699), .B(g_input[62]), .Z(n2701) );
  XOR U3077 ( .A(n394), .B(n2732), .Z(n2699) );
  AND U3078 ( .A(n2733), .B(n2734), .Z(n2732) );
  XOR U3079 ( .A(e_input[61]), .B(n394), .Z(n2734) );
  IV U3080 ( .A(n2704), .Z(n2726) );
  XOR U3081 ( .A(n2735), .B(n2736), .Z(n2704) );
  ANDN U3082 ( .A(n2737), .B(n2738), .Z(n2736) );
  XOR U3083 ( .A(n2735), .B(n2739), .Z(n2737) );
  XOR U3084 ( .A(n2740), .B(n2741), .Z(n2708) );
  AND U3085 ( .A(n2670), .B(n2742), .Z(n2741) );
  XNOR U3086 ( .A(n2716), .B(n2743), .Z(n2742) );
  XOR U3087 ( .A(n2744), .B(n2740), .Z(n2743) );
  IV U3088 ( .A(e_input[30]), .Z(n2744) );
  XNOR U3089 ( .A(n2714), .B(g_input[30]), .Z(n2716) );
  XOR U3090 ( .A(n395), .B(n2745), .Z(n2714) );
  AND U3091 ( .A(n2746), .B(n2747), .Z(n2745) );
  XOR U3092 ( .A(e_input[29]), .B(n395), .Z(n2747) );
  XNOR U3093 ( .A(n2748), .B(g_input[30]), .Z(n2740) );
  XNOR U3094 ( .A(n2749), .B(\min_dist_reg[3][30] ), .Z(n2722) );
  IV U3095 ( .A(n2720), .Z(n2749) );
  XOR U3096 ( .A(n2750), .B(n2751), .Z(n2720) );
  AND U3097 ( .A(n2752), .B(n2753), .Z(n2751) );
  XNOR U3098 ( .A(n2750), .B(n2430), .Z(n2753) );
  XOR U3099 ( .A(n2739), .B(n2738), .Z(n2430) );
  XNOR U3100 ( .A(n2754), .B(n2755), .Z(n2738) );
  XNOR U3101 ( .A(n2756), .B(n2757), .Z(n2754) );
  AND U3102 ( .A(n2676), .B(n2758), .Z(n2757) );
  XNOR U3103 ( .A(n2733), .B(n2759), .Z(n2758) );
  XOR U3104 ( .A(n2760), .B(n2755), .Z(n2759) );
  XNOR U3105 ( .A(n2761), .B(g_input[61]), .Z(n2755) );
  IV U3106 ( .A(e_input[61]), .Z(n2760) );
  XNOR U3107 ( .A(n394), .B(g_input[61]), .Z(n2733) );
  AND U3108 ( .A(n2764), .B(n2765), .Z(n2763) );
  XOR U3109 ( .A(e_input[60]), .B(n2766), .Z(n2765) );
  IV U3110 ( .A(n2735), .Z(n2756) );
  XOR U3111 ( .A(n2767), .B(n2768), .Z(n2735) );
  ANDN U3112 ( .A(n2769), .B(n2770), .Z(n2768) );
  XOR U3113 ( .A(n2767), .B(n2771), .Z(n2769) );
  XOR U3114 ( .A(n2772), .B(n2773), .Z(n2739) );
  AND U3115 ( .A(n2670), .B(n2774), .Z(n2773) );
  XNOR U3116 ( .A(n2746), .B(n2775), .Z(n2774) );
  XOR U3117 ( .A(n2776), .B(n2772), .Z(n2775) );
  IV U3118 ( .A(e_input[29]), .Z(n2776) );
  XNOR U3119 ( .A(n395), .B(g_input[29]), .Z(n2746) );
  AND U3120 ( .A(n2779), .B(n2780), .Z(n2778) );
  XOR U3121 ( .A(e_input[28]), .B(n2781), .Z(n2780) );
  XNOR U3122 ( .A(n2782), .B(g_input[29]), .Z(n2772) );
  XNOR U3123 ( .A(n2783), .B(\min_dist_reg[3][29] ), .Z(n2752) );
  IV U3124 ( .A(n2750), .Z(n2783) );
  XOR U3125 ( .A(n2784), .B(n2785), .Z(n2750) );
  AND U3126 ( .A(n2786), .B(n2787), .Z(n2785) );
  XNOR U3127 ( .A(n2784), .B(n2438), .Z(n2787) );
  XOR U3128 ( .A(n2771), .B(n2770), .Z(n2438) );
  XNOR U3129 ( .A(n2788), .B(n2789), .Z(n2770) );
  XNOR U3130 ( .A(n2790), .B(n2791), .Z(n2788) );
  AND U3131 ( .A(n2676), .B(n2792), .Z(n2791) );
  XNOR U3132 ( .A(n2764), .B(n2793), .Z(n2792) );
  XOR U3133 ( .A(n2794), .B(n2789), .Z(n2793) );
  XNOR U3134 ( .A(n2795), .B(g_input[60]), .Z(n2789) );
  IV U3135 ( .A(e_input[60]), .Z(n2794) );
  XNOR U3136 ( .A(n2766), .B(g_input[60]), .Z(n2764) );
  IV U3137 ( .A(n2762), .Z(n2766) );
  XOR U3138 ( .A(n2796), .B(n2797), .Z(n2762) );
  AND U3139 ( .A(n2798), .B(n2799), .Z(n2797) );
  XOR U3140 ( .A(e_input[59]), .B(n2800), .Z(n2799) );
  IV U3141 ( .A(n2767), .Z(n2790) );
  XOR U3142 ( .A(n2801), .B(n2802), .Z(n2767) );
  ANDN U3143 ( .A(n2803), .B(n2804), .Z(n2802) );
  XOR U3144 ( .A(n2801), .B(n2805), .Z(n2803) );
  XOR U3145 ( .A(n2806), .B(n2807), .Z(n2771) );
  AND U3146 ( .A(n2670), .B(n2808), .Z(n2807) );
  XNOR U3147 ( .A(n2779), .B(n2809), .Z(n2808) );
  XOR U3148 ( .A(n2810), .B(n2806), .Z(n2809) );
  IV U3149 ( .A(e_input[28]), .Z(n2810) );
  XNOR U3150 ( .A(n2781), .B(g_input[28]), .Z(n2779) );
  IV U3151 ( .A(n2777), .Z(n2781) );
  XOR U3152 ( .A(n2811), .B(n2812), .Z(n2777) );
  AND U3153 ( .A(n2813), .B(n2814), .Z(n2812) );
  XOR U3154 ( .A(e_input[27]), .B(n2815), .Z(n2814) );
  XNOR U3155 ( .A(n2816), .B(g_input[28]), .Z(n2806) );
  XNOR U3156 ( .A(n2817), .B(\min_dist_reg[3][28] ), .Z(n2786) );
  IV U3157 ( .A(n2784), .Z(n2817) );
  XOR U3158 ( .A(n2818), .B(n2819), .Z(n2784) );
  AND U3159 ( .A(n2820), .B(n2821), .Z(n2819) );
  XNOR U3160 ( .A(n2818), .B(n2446), .Z(n2821) );
  XOR U3161 ( .A(n2805), .B(n2804), .Z(n2446) );
  XNOR U3162 ( .A(n2822), .B(n2823), .Z(n2804) );
  XNOR U3163 ( .A(n2824), .B(n2825), .Z(n2822) );
  AND U3164 ( .A(n2676), .B(n2826), .Z(n2825) );
  XNOR U3165 ( .A(n2798), .B(n2827), .Z(n2826) );
  XOR U3166 ( .A(n2828), .B(n2823), .Z(n2827) );
  XNOR U3167 ( .A(n2829), .B(g_input[59]), .Z(n2823) );
  IV U3168 ( .A(e_input[59]), .Z(n2828) );
  XNOR U3169 ( .A(n2800), .B(g_input[59]), .Z(n2798) );
  IV U3170 ( .A(n2796), .Z(n2800) );
  XOR U3171 ( .A(n2830), .B(n2831), .Z(n2796) );
  AND U3172 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U3173 ( .A(e_input[58]), .B(n2834), .Z(n2833) );
  IV U3174 ( .A(n2801), .Z(n2824) );
  XOR U3175 ( .A(n2835), .B(n2836), .Z(n2801) );
  ANDN U3176 ( .A(n2837), .B(n2838), .Z(n2836) );
  XOR U3177 ( .A(n2835), .B(n2839), .Z(n2837) );
  XOR U3178 ( .A(n2840), .B(n2841), .Z(n2805) );
  AND U3179 ( .A(n2670), .B(n2842), .Z(n2841) );
  XNOR U3180 ( .A(n2813), .B(n2843), .Z(n2842) );
  XOR U3181 ( .A(n2844), .B(n2840), .Z(n2843) );
  IV U3182 ( .A(e_input[27]), .Z(n2844) );
  XNOR U3183 ( .A(n2815), .B(g_input[27]), .Z(n2813) );
  IV U3184 ( .A(n2811), .Z(n2815) );
  XOR U3185 ( .A(n2845), .B(n2846), .Z(n2811) );
  AND U3186 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U3187 ( .A(e_input[26]), .B(n2849), .Z(n2848) );
  XNOR U3188 ( .A(n2850), .B(g_input[27]), .Z(n2840) );
  XNOR U3189 ( .A(n2851), .B(\min_dist_reg[3][27] ), .Z(n2820) );
  IV U3190 ( .A(n2818), .Z(n2851) );
  XOR U3191 ( .A(n2852), .B(n2853), .Z(n2818) );
  AND U3192 ( .A(n2854), .B(n2855), .Z(n2853) );
  XNOR U3193 ( .A(n2852), .B(n2454), .Z(n2855) );
  XOR U3194 ( .A(n2839), .B(n2838), .Z(n2454) );
  XNOR U3195 ( .A(n2856), .B(n2857), .Z(n2838) );
  XNOR U3196 ( .A(n2858), .B(n2859), .Z(n2856) );
  AND U3197 ( .A(n2676), .B(n2860), .Z(n2859) );
  XNOR U3198 ( .A(n2832), .B(n2861), .Z(n2860) );
  XOR U3199 ( .A(n2862), .B(n2857), .Z(n2861) );
  XNOR U3200 ( .A(n2863), .B(g_input[58]), .Z(n2857) );
  IV U3201 ( .A(e_input[58]), .Z(n2862) );
  XNOR U3202 ( .A(n2834), .B(g_input[58]), .Z(n2832) );
  IV U3203 ( .A(n2830), .Z(n2834) );
  XOR U3204 ( .A(n2864), .B(n2865), .Z(n2830) );
  AND U3205 ( .A(n2866), .B(n2867), .Z(n2865) );
  XOR U3206 ( .A(e_input[57]), .B(n2868), .Z(n2867) );
  IV U3207 ( .A(n2835), .Z(n2858) );
  XOR U3208 ( .A(n2869), .B(n2870), .Z(n2835) );
  ANDN U3209 ( .A(n2871), .B(n2872), .Z(n2870) );
  XOR U3210 ( .A(n2869), .B(n2873), .Z(n2871) );
  XOR U3211 ( .A(n2874), .B(n2875), .Z(n2839) );
  AND U3212 ( .A(n2670), .B(n2876), .Z(n2875) );
  XNOR U3213 ( .A(n2847), .B(n2877), .Z(n2876) );
  XOR U3214 ( .A(n2878), .B(n2874), .Z(n2877) );
  IV U3215 ( .A(e_input[26]), .Z(n2878) );
  XNOR U3216 ( .A(n2849), .B(g_input[26]), .Z(n2847) );
  IV U3217 ( .A(n2845), .Z(n2849) );
  XOR U3218 ( .A(n2879), .B(n2880), .Z(n2845) );
  AND U3219 ( .A(n2881), .B(n2882), .Z(n2880) );
  XOR U3220 ( .A(e_input[25]), .B(n2883), .Z(n2882) );
  XNOR U3221 ( .A(n2884), .B(g_input[26]), .Z(n2874) );
  XNOR U3222 ( .A(n2885), .B(\min_dist_reg[3][26] ), .Z(n2854) );
  IV U3223 ( .A(n2852), .Z(n2885) );
  XOR U3224 ( .A(n2886), .B(n2887), .Z(n2852) );
  AND U3225 ( .A(n2888), .B(n2889), .Z(n2887) );
  XNOR U3226 ( .A(n2886), .B(n2462), .Z(n2889) );
  XOR U3227 ( .A(n2873), .B(n2872), .Z(n2462) );
  XNOR U3228 ( .A(n2890), .B(n2891), .Z(n2872) );
  XNOR U3229 ( .A(n2892), .B(n2893), .Z(n2890) );
  AND U3230 ( .A(n2676), .B(n2894), .Z(n2893) );
  XNOR U3231 ( .A(n2866), .B(n2895), .Z(n2894) );
  XOR U3232 ( .A(n2896), .B(n2891), .Z(n2895) );
  XNOR U3233 ( .A(n2897), .B(g_input[57]), .Z(n2891) );
  IV U3234 ( .A(e_input[57]), .Z(n2896) );
  XNOR U3235 ( .A(n2868), .B(g_input[57]), .Z(n2866) );
  IV U3236 ( .A(n2864), .Z(n2868) );
  XOR U3237 ( .A(n2898), .B(n2899), .Z(n2864) );
  AND U3238 ( .A(n2900), .B(n2901), .Z(n2899) );
  XOR U3239 ( .A(e_input[56]), .B(n2902), .Z(n2901) );
  IV U3240 ( .A(n2869), .Z(n2892) );
  XOR U3241 ( .A(n2903), .B(n2904), .Z(n2869) );
  ANDN U3242 ( .A(n2905), .B(n2906), .Z(n2904) );
  XOR U3243 ( .A(n2903), .B(n2907), .Z(n2905) );
  XOR U3244 ( .A(n2908), .B(n2909), .Z(n2873) );
  AND U3245 ( .A(n2670), .B(n2910), .Z(n2909) );
  XNOR U3246 ( .A(n2881), .B(n2911), .Z(n2910) );
  XOR U3247 ( .A(n2912), .B(n2908), .Z(n2911) );
  IV U3248 ( .A(e_input[25]), .Z(n2912) );
  XNOR U3249 ( .A(n2883), .B(g_input[25]), .Z(n2881) );
  IV U3250 ( .A(n2879), .Z(n2883) );
  XOR U3251 ( .A(n2913), .B(n2914), .Z(n2879) );
  AND U3252 ( .A(n2915), .B(n2916), .Z(n2914) );
  XOR U3253 ( .A(e_input[24]), .B(n2917), .Z(n2916) );
  XNOR U3254 ( .A(n2918), .B(g_input[25]), .Z(n2908) );
  XNOR U3255 ( .A(n2919), .B(\min_dist_reg[3][25] ), .Z(n2888) );
  IV U3256 ( .A(n2886), .Z(n2919) );
  XOR U3257 ( .A(n2920), .B(n2921), .Z(n2886) );
  AND U3258 ( .A(n2922), .B(n2923), .Z(n2921) );
  XNOR U3259 ( .A(n2920), .B(n2470), .Z(n2923) );
  XOR U3260 ( .A(n2907), .B(n2906), .Z(n2470) );
  XNOR U3261 ( .A(n2924), .B(n2925), .Z(n2906) );
  XNOR U3262 ( .A(n2926), .B(n2927), .Z(n2924) );
  AND U3263 ( .A(n2676), .B(n2928), .Z(n2927) );
  XNOR U3264 ( .A(n2900), .B(n2929), .Z(n2928) );
  XOR U3265 ( .A(n2930), .B(n2925), .Z(n2929) );
  XNOR U3266 ( .A(n2931), .B(g_input[56]), .Z(n2925) );
  IV U3267 ( .A(e_input[56]), .Z(n2930) );
  XNOR U3268 ( .A(n2902), .B(g_input[56]), .Z(n2900) );
  IV U3269 ( .A(n2898), .Z(n2902) );
  XOR U3270 ( .A(n2932), .B(n2933), .Z(n2898) );
  AND U3271 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR U3272 ( .A(e_input[55]), .B(n2936), .Z(n2935) );
  IV U3273 ( .A(n2903), .Z(n2926) );
  XOR U3274 ( .A(n2937), .B(n2938), .Z(n2903) );
  ANDN U3275 ( .A(n2939), .B(n2940), .Z(n2938) );
  XOR U3276 ( .A(n2937), .B(n2941), .Z(n2939) );
  XOR U3277 ( .A(n2942), .B(n2943), .Z(n2907) );
  AND U3278 ( .A(n2670), .B(n2944), .Z(n2943) );
  XNOR U3279 ( .A(n2915), .B(n2945), .Z(n2944) );
  XOR U3280 ( .A(n2946), .B(n2942), .Z(n2945) );
  IV U3281 ( .A(e_input[24]), .Z(n2946) );
  XNOR U3282 ( .A(n2917), .B(g_input[24]), .Z(n2915) );
  IV U3283 ( .A(n2913), .Z(n2917) );
  XOR U3284 ( .A(n2947), .B(n2948), .Z(n2913) );
  AND U3285 ( .A(n2949), .B(n2950), .Z(n2948) );
  XOR U3286 ( .A(e_input[23]), .B(n2951), .Z(n2950) );
  XNOR U3287 ( .A(n2952), .B(g_input[24]), .Z(n2942) );
  XNOR U3288 ( .A(n2953), .B(\min_dist_reg[3][24] ), .Z(n2922) );
  IV U3289 ( .A(n2920), .Z(n2953) );
  XOR U3290 ( .A(n2954), .B(n2955), .Z(n2920) );
  AND U3291 ( .A(n2956), .B(n2957), .Z(n2955) );
  XNOR U3292 ( .A(n2954), .B(n2478), .Z(n2957) );
  XOR U3293 ( .A(n2941), .B(n2940), .Z(n2478) );
  XNOR U3294 ( .A(n2958), .B(n2959), .Z(n2940) );
  XNOR U3295 ( .A(n2960), .B(n2961), .Z(n2958) );
  AND U3296 ( .A(n2676), .B(n2962), .Z(n2961) );
  XNOR U3297 ( .A(n2934), .B(n2963), .Z(n2962) );
  XOR U3298 ( .A(n2964), .B(n2959), .Z(n2963) );
  XNOR U3299 ( .A(n2965), .B(g_input[55]), .Z(n2959) );
  IV U3300 ( .A(e_input[55]), .Z(n2964) );
  XNOR U3301 ( .A(n2936), .B(g_input[55]), .Z(n2934) );
  IV U3302 ( .A(n2932), .Z(n2936) );
  XOR U3303 ( .A(n2966), .B(n2967), .Z(n2932) );
  AND U3304 ( .A(n2968), .B(n2969), .Z(n2967) );
  XOR U3305 ( .A(e_input[54]), .B(n2970), .Z(n2969) );
  IV U3306 ( .A(n2937), .Z(n2960) );
  XOR U3307 ( .A(n2971), .B(n2972), .Z(n2937) );
  ANDN U3308 ( .A(n2973), .B(n2974), .Z(n2972) );
  XOR U3309 ( .A(n2971), .B(n2975), .Z(n2973) );
  XOR U3310 ( .A(n2976), .B(n2977), .Z(n2941) );
  AND U3311 ( .A(n2670), .B(n2978), .Z(n2977) );
  XNOR U3312 ( .A(n2949), .B(n2979), .Z(n2978) );
  XOR U3313 ( .A(n2980), .B(n2976), .Z(n2979) );
  IV U3314 ( .A(e_input[23]), .Z(n2980) );
  XNOR U3315 ( .A(n2951), .B(g_input[23]), .Z(n2949) );
  IV U3316 ( .A(n2947), .Z(n2951) );
  XOR U3317 ( .A(n2981), .B(n2982), .Z(n2947) );
  AND U3318 ( .A(n2983), .B(n2984), .Z(n2982) );
  XOR U3319 ( .A(e_input[22]), .B(n2985), .Z(n2984) );
  XNOR U3320 ( .A(n2986), .B(g_input[23]), .Z(n2976) );
  XNOR U3321 ( .A(n2987), .B(\min_dist_reg[3][23] ), .Z(n2956) );
  IV U3322 ( .A(n2954), .Z(n2987) );
  XOR U3323 ( .A(n2988), .B(n2989), .Z(n2954) );
  AND U3324 ( .A(n2990), .B(n2991), .Z(n2989) );
  XNOR U3325 ( .A(n2988), .B(n2486), .Z(n2991) );
  XOR U3326 ( .A(n2975), .B(n2974), .Z(n2486) );
  XNOR U3327 ( .A(n2992), .B(n2993), .Z(n2974) );
  XNOR U3328 ( .A(n2994), .B(n2995), .Z(n2992) );
  AND U3329 ( .A(n2676), .B(n2996), .Z(n2995) );
  XNOR U3330 ( .A(n2968), .B(n2997), .Z(n2996) );
  XOR U3331 ( .A(n2998), .B(n2993), .Z(n2997) );
  XNOR U3332 ( .A(n2999), .B(g_input[54]), .Z(n2993) );
  IV U3333 ( .A(e_input[54]), .Z(n2998) );
  XNOR U3334 ( .A(n2970), .B(g_input[54]), .Z(n2968) );
  IV U3335 ( .A(n2966), .Z(n2970) );
  XOR U3336 ( .A(n3000), .B(n3001), .Z(n2966) );
  AND U3337 ( .A(n3002), .B(n3003), .Z(n3001) );
  XOR U3338 ( .A(e_input[53]), .B(n3004), .Z(n3003) );
  IV U3339 ( .A(n2971), .Z(n2994) );
  XOR U3340 ( .A(n3005), .B(n3006), .Z(n2971) );
  ANDN U3341 ( .A(n3007), .B(n3008), .Z(n3006) );
  XOR U3342 ( .A(n3005), .B(n3009), .Z(n3007) );
  XOR U3343 ( .A(n3010), .B(n3011), .Z(n2975) );
  AND U3344 ( .A(n2670), .B(n3012), .Z(n3011) );
  XNOR U3345 ( .A(n2983), .B(n3013), .Z(n3012) );
  XOR U3346 ( .A(n3014), .B(n3010), .Z(n3013) );
  IV U3347 ( .A(e_input[22]), .Z(n3014) );
  XNOR U3348 ( .A(n2985), .B(g_input[22]), .Z(n2983) );
  IV U3349 ( .A(n2981), .Z(n2985) );
  XOR U3350 ( .A(n3015), .B(n3016), .Z(n2981) );
  AND U3351 ( .A(n3017), .B(n3018), .Z(n3016) );
  XOR U3352 ( .A(e_input[21]), .B(n3019), .Z(n3018) );
  XNOR U3353 ( .A(n3020), .B(g_input[22]), .Z(n3010) );
  XNOR U3354 ( .A(n3021), .B(\min_dist_reg[3][22] ), .Z(n2990) );
  IV U3355 ( .A(n2988), .Z(n3021) );
  XOR U3356 ( .A(n3022), .B(n3023), .Z(n2988) );
  AND U3357 ( .A(n3024), .B(n3025), .Z(n3023) );
  XNOR U3358 ( .A(n3022), .B(n2494), .Z(n3025) );
  XOR U3359 ( .A(n3009), .B(n3008), .Z(n2494) );
  XNOR U3360 ( .A(n3026), .B(n3027), .Z(n3008) );
  XNOR U3361 ( .A(n3028), .B(n3029), .Z(n3026) );
  AND U3362 ( .A(n2676), .B(n3030), .Z(n3029) );
  XNOR U3363 ( .A(n3002), .B(n3031), .Z(n3030) );
  XOR U3364 ( .A(n3032), .B(n3027), .Z(n3031) );
  XNOR U3365 ( .A(n3033), .B(g_input[53]), .Z(n3027) );
  IV U3366 ( .A(e_input[53]), .Z(n3032) );
  XNOR U3367 ( .A(n3004), .B(g_input[53]), .Z(n3002) );
  IV U3368 ( .A(n3000), .Z(n3004) );
  XOR U3369 ( .A(n3034), .B(n3035), .Z(n3000) );
  AND U3370 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U3371 ( .A(e_input[52]), .B(n3038), .Z(n3037) );
  IV U3372 ( .A(n3005), .Z(n3028) );
  XOR U3373 ( .A(n3039), .B(n3040), .Z(n3005) );
  ANDN U3374 ( .A(n3041), .B(n3042), .Z(n3040) );
  XOR U3375 ( .A(n3039), .B(n3043), .Z(n3041) );
  XOR U3376 ( .A(n3044), .B(n3045), .Z(n3009) );
  AND U3377 ( .A(n2670), .B(n3046), .Z(n3045) );
  XNOR U3378 ( .A(n3017), .B(n3047), .Z(n3046) );
  XOR U3379 ( .A(n3048), .B(n3044), .Z(n3047) );
  IV U3380 ( .A(e_input[21]), .Z(n3048) );
  XNOR U3381 ( .A(n3019), .B(g_input[21]), .Z(n3017) );
  IV U3382 ( .A(n3015), .Z(n3019) );
  XOR U3383 ( .A(n3049), .B(n3050), .Z(n3015) );
  AND U3384 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U3385 ( .A(e_input[20]), .B(n3053), .Z(n3052) );
  XNOR U3386 ( .A(n3054), .B(g_input[21]), .Z(n3044) );
  XNOR U3387 ( .A(n3055), .B(\min_dist_reg[3][21] ), .Z(n3024) );
  IV U3388 ( .A(n3022), .Z(n3055) );
  XOR U3389 ( .A(n3056), .B(n3057), .Z(n3022) );
  AND U3390 ( .A(n3058), .B(n3059), .Z(n3057) );
  XNOR U3391 ( .A(n3056), .B(n2502), .Z(n3059) );
  XOR U3392 ( .A(n3043), .B(n3042), .Z(n2502) );
  XNOR U3393 ( .A(n3060), .B(n3061), .Z(n3042) );
  XNOR U3394 ( .A(n3062), .B(n3063), .Z(n3060) );
  AND U3395 ( .A(n2676), .B(n3064), .Z(n3063) );
  XNOR U3396 ( .A(n3036), .B(n3065), .Z(n3064) );
  XOR U3397 ( .A(n3066), .B(n3061), .Z(n3065) );
  XNOR U3398 ( .A(n3067), .B(g_input[52]), .Z(n3061) );
  IV U3399 ( .A(e_input[52]), .Z(n3066) );
  XNOR U3400 ( .A(n3038), .B(g_input[52]), .Z(n3036) );
  IV U3401 ( .A(n3034), .Z(n3038) );
  XOR U3402 ( .A(n3068), .B(n3069), .Z(n3034) );
  AND U3403 ( .A(n3070), .B(n3071), .Z(n3069) );
  XOR U3404 ( .A(e_input[51]), .B(n3072), .Z(n3071) );
  IV U3405 ( .A(n3039), .Z(n3062) );
  XOR U3406 ( .A(n3073), .B(n3074), .Z(n3039) );
  ANDN U3407 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR U3408 ( .A(n3073), .B(n3077), .Z(n3075) );
  XOR U3409 ( .A(n3078), .B(n3079), .Z(n3043) );
  AND U3410 ( .A(n2670), .B(n3080), .Z(n3079) );
  XNOR U3411 ( .A(n3051), .B(n3081), .Z(n3080) );
  XOR U3412 ( .A(n3082), .B(n3078), .Z(n3081) );
  IV U3413 ( .A(e_input[20]), .Z(n3082) );
  XNOR U3414 ( .A(n3053), .B(g_input[20]), .Z(n3051) );
  IV U3415 ( .A(n3049), .Z(n3053) );
  XOR U3416 ( .A(n3083), .B(n3084), .Z(n3049) );
  AND U3417 ( .A(n3085), .B(n3086), .Z(n3084) );
  XOR U3418 ( .A(e_input[19]), .B(n3087), .Z(n3086) );
  XNOR U3419 ( .A(n3088), .B(g_input[20]), .Z(n3078) );
  XNOR U3420 ( .A(n3089), .B(\min_dist_reg[3][20] ), .Z(n3058) );
  IV U3421 ( .A(n3056), .Z(n3089) );
  XOR U3422 ( .A(n3090), .B(n3091), .Z(n3056) );
  AND U3423 ( .A(n3092), .B(n3093), .Z(n3091) );
  XNOR U3424 ( .A(n3090), .B(n2510), .Z(n3093) );
  XOR U3425 ( .A(n3077), .B(n3076), .Z(n2510) );
  XNOR U3426 ( .A(n3094), .B(n3095), .Z(n3076) );
  XNOR U3427 ( .A(n3096), .B(n3097), .Z(n3094) );
  AND U3428 ( .A(n2676), .B(n3098), .Z(n3097) );
  XNOR U3429 ( .A(n3070), .B(n3099), .Z(n3098) );
  XOR U3430 ( .A(n3100), .B(n3095), .Z(n3099) );
  XNOR U3431 ( .A(n3101), .B(g_input[51]), .Z(n3095) );
  IV U3432 ( .A(e_input[51]), .Z(n3100) );
  XNOR U3433 ( .A(n3072), .B(g_input[51]), .Z(n3070) );
  IV U3434 ( .A(n3068), .Z(n3072) );
  XOR U3435 ( .A(n3102), .B(n3103), .Z(n3068) );
  AND U3436 ( .A(n3104), .B(n3105), .Z(n3103) );
  XOR U3437 ( .A(e_input[50]), .B(n3106), .Z(n3105) );
  IV U3438 ( .A(n3073), .Z(n3096) );
  XOR U3439 ( .A(n3107), .B(n3108), .Z(n3073) );
  ANDN U3440 ( .A(n3109), .B(n3110), .Z(n3108) );
  XOR U3441 ( .A(n3107), .B(n3111), .Z(n3109) );
  XOR U3442 ( .A(n3112), .B(n3113), .Z(n3077) );
  AND U3443 ( .A(n2670), .B(n3114), .Z(n3113) );
  XNOR U3444 ( .A(n3085), .B(n3115), .Z(n3114) );
  XOR U3445 ( .A(n3116), .B(n3112), .Z(n3115) );
  IV U3446 ( .A(e_input[19]), .Z(n3116) );
  XNOR U3447 ( .A(n3087), .B(g_input[19]), .Z(n3085) );
  IV U3448 ( .A(n3083), .Z(n3087) );
  XOR U3449 ( .A(n3117), .B(n3118), .Z(n3083) );
  AND U3450 ( .A(n3119), .B(n3120), .Z(n3118) );
  XOR U3451 ( .A(e_input[18]), .B(n3121), .Z(n3120) );
  XNOR U3452 ( .A(n3122), .B(g_input[19]), .Z(n3112) );
  XNOR U3453 ( .A(n3123), .B(\min_dist_reg[3][19] ), .Z(n3092) );
  IV U3454 ( .A(n3090), .Z(n3123) );
  XOR U3455 ( .A(n3124), .B(n3125), .Z(n3090) );
  AND U3456 ( .A(n3126), .B(n3127), .Z(n3125) );
  XNOR U3457 ( .A(n3124), .B(n2518), .Z(n3127) );
  XOR U3458 ( .A(n3111), .B(n3110), .Z(n2518) );
  XNOR U3459 ( .A(n3128), .B(n3129), .Z(n3110) );
  XNOR U3460 ( .A(n3130), .B(n3131), .Z(n3128) );
  AND U3461 ( .A(n2676), .B(n3132), .Z(n3131) );
  XNOR U3462 ( .A(n3104), .B(n3133), .Z(n3132) );
  XOR U3463 ( .A(n3134), .B(n3129), .Z(n3133) );
  XNOR U3464 ( .A(n3135), .B(g_input[50]), .Z(n3129) );
  IV U3465 ( .A(e_input[50]), .Z(n3134) );
  XNOR U3466 ( .A(n3106), .B(g_input[50]), .Z(n3104) );
  IV U3467 ( .A(n3102), .Z(n3106) );
  XOR U3468 ( .A(n3136), .B(n3137), .Z(n3102) );
  AND U3469 ( .A(n3138), .B(n3139), .Z(n3137) );
  XOR U3470 ( .A(e_input[49]), .B(n3140), .Z(n3139) );
  IV U3471 ( .A(n3107), .Z(n3130) );
  XOR U3472 ( .A(n3141), .B(n3142), .Z(n3107) );
  ANDN U3473 ( .A(n3143), .B(n3144), .Z(n3142) );
  XOR U3474 ( .A(n3141), .B(n3145), .Z(n3143) );
  XOR U3475 ( .A(n3146), .B(n3147), .Z(n3111) );
  AND U3476 ( .A(n2670), .B(n3148), .Z(n3147) );
  XNOR U3477 ( .A(n3119), .B(n3149), .Z(n3148) );
  XOR U3478 ( .A(n3150), .B(n3146), .Z(n3149) );
  IV U3479 ( .A(e_input[18]), .Z(n3150) );
  XNOR U3480 ( .A(n3121), .B(g_input[18]), .Z(n3119) );
  IV U3481 ( .A(n3117), .Z(n3121) );
  XOR U3482 ( .A(n3151), .B(n3152), .Z(n3117) );
  AND U3483 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U3484 ( .A(e_input[17]), .B(n3155), .Z(n3154) );
  XNOR U3485 ( .A(n3156), .B(g_input[18]), .Z(n3146) );
  XNOR U3486 ( .A(n3157), .B(\min_dist_reg[3][18] ), .Z(n3126) );
  IV U3487 ( .A(n3124), .Z(n3157) );
  XOR U3488 ( .A(n3158), .B(n3159), .Z(n3124) );
  AND U3489 ( .A(n3160), .B(n3161), .Z(n3159) );
  XNOR U3490 ( .A(n3158), .B(n2526), .Z(n3161) );
  XOR U3491 ( .A(n3145), .B(n3144), .Z(n2526) );
  XNOR U3492 ( .A(n3162), .B(n3163), .Z(n3144) );
  XNOR U3493 ( .A(n3164), .B(n3165), .Z(n3162) );
  AND U3494 ( .A(n2676), .B(n3166), .Z(n3165) );
  XNOR U3495 ( .A(n3138), .B(n3167), .Z(n3166) );
  XOR U3496 ( .A(n3168), .B(n3163), .Z(n3167) );
  XNOR U3497 ( .A(n3169), .B(g_input[49]), .Z(n3163) );
  IV U3498 ( .A(e_input[49]), .Z(n3168) );
  XNOR U3499 ( .A(n3140), .B(g_input[49]), .Z(n3138) );
  IV U3500 ( .A(n3136), .Z(n3140) );
  XOR U3501 ( .A(n3170), .B(n3171), .Z(n3136) );
  AND U3502 ( .A(n3172), .B(n3173), .Z(n3171) );
  XOR U3503 ( .A(e_input[48]), .B(n3174), .Z(n3173) );
  IV U3504 ( .A(n3141), .Z(n3164) );
  XOR U3505 ( .A(n3175), .B(n3176), .Z(n3141) );
  ANDN U3506 ( .A(n3177), .B(n3178), .Z(n3176) );
  XOR U3507 ( .A(n3175), .B(n3179), .Z(n3177) );
  XOR U3508 ( .A(n3180), .B(n3181), .Z(n3145) );
  AND U3509 ( .A(n2670), .B(n3182), .Z(n3181) );
  XNOR U3510 ( .A(n3153), .B(n3183), .Z(n3182) );
  XOR U3511 ( .A(n3184), .B(n3180), .Z(n3183) );
  IV U3512 ( .A(e_input[17]), .Z(n3184) );
  XNOR U3513 ( .A(n3155), .B(g_input[17]), .Z(n3153) );
  IV U3514 ( .A(n3151), .Z(n3155) );
  XOR U3515 ( .A(n3185), .B(n3186), .Z(n3151) );
  AND U3516 ( .A(n3187), .B(n3188), .Z(n3186) );
  XOR U3517 ( .A(e_input[16]), .B(n3189), .Z(n3188) );
  XNOR U3518 ( .A(n3190), .B(g_input[17]), .Z(n3180) );
  XNOR U3519 ( .A(n3191), .B(\min_dist_reg[3][17] ), .Z(n3160) );
  IV U3520 ( .A(n3158), .Z(n3191) );
  XOR U3521 ( .A(n3192), .B(n3193), .Z(n3158) );
  AND U3522 ( .A(n3194), .B(n3195), .Z(n3193) );
  XNOR U3523 ( .A(n3192), .B(n2534), .Z(n3195) );
  XOR U3524 ( .A(n3179), .B(n3178), .Z(n2534) );
  XNOR U3525 ( .A(n3196), .B(n3197), .Z(n3178) );
  XNOR U3526 ( .A(n3198), .B(n3199), .Z(n3196) );
  AND U3527 ( .A(n2676), .B(n3200), .Z(n3199) );
  XNOR U3528 ( .A(n3172), .B(n3201), .Z(n3200) );
  XOR U3529 ( .A(n3202), .B(n3197), .Z(n3201) );
  XNOR U3530 ( .A(n3203), .B(g_input[48]), .Z(n3197) );
  IV U3531 ( .A(e_input[48]), .Z(n3202) );
  XNOR U3532 ( .A(n3174), .B(g_input[48]), .Z(n3172) );
  IV U3533 ( .A(n3170), .Z(n3174) );
  XOR U3534 ( .A(n3204), .B(n3205), .Z(n3170) );
  AND U3535 ( .A(n3206), .B(n3207), .Z(n3205) );
  XOR U3536 ( .A(e_input[47]), .B(n3208), .Z(n3207) );
  IV U3537 ( .A(n3175), .Z(n3198) );
  XOR U3538 ( .A(n3209), .B(n3210), .Z(n3175) );
  ANDN U3539 ( .A(n3211), .B(n3212), .Z(n3210) );
  XOR U3540 ( .A(n3209), .B(n3213), .Z(n3211) );
  XOR U3541 ( .A(n3214), .B(n3215), .Z(n3179) );
  AND U3542 ( .A(n2670), .B(n3216), .Z(n3215) );
  XNOR U3543 ( .A(n3187), .B(n3217), .Z(n3216) );
  XOR U3544 ( .A(n3218), .B(n3214), .Z(n3217) );
  IV U3545 ( .A(e_input[16]), .Z(n3218) );
  XNOR U3546 ( .A(n3189), .B(g_input[16]), .Z(n3187) );
  IV U3547 ( .A(n3185), .Z(n3189) );
  XOR U3548 ( .A(n3219), .B(n3220), .Z(n3185) );
  AND U3549 ( .A(n3221), .B(n3222), .Z(n3220) );
  XOR U3550 ( .A(e_input[15]), .B(n3223), .Z(n3222) );
  XNOR U3551 ( .A(n3224), .B(g_input[16]), .Z(n3214) );
  XNOR U3552 ( .A(n3225), .B(\min_dist_reg[3][16] ), .Z(n3194) );
  IV U3553 ( .A(n3192), .Z(n3225) );
  XOR U3554 ( .A(n3226), .B(n3227), .Z(n3192) );
  AND U3555 ( .A(n3228), .B(n3229), .Z(n3227) );
  XNOR U3556 ( .A(n3226), .B(n2542), .Z(n3229) );
  XOR U3557 ( .A(n3213), .B(n3212), .Z(n2542) );
  XNOR U3558 ( .A(n3230), .B(n3231), .Z(n3212) );
  XNOR U3559 ( .A(n3232), .B(n3233), .Z(n3230) );
  AND U3560 ( .A(n2676), .B(n3234), .Z(n3233) );
  XNOR U3561 ( .A(n3206), .B(n3235), .Z(n3234) );
  XOR U3562 ( .A(n3236), .B(n3231), .Z(n3235) );
  XNOR U3563 ( .A(n3237), .B(g_input[47]), .Z(n3231) );
  IV U3564 ( .A(e_input[47]), .Z(n3236) );
  XNOR U3565 ( .A(n3208), .B(g_input[47]), .Z(n3206) );
  IV U3566 ( .A(n3204), .Z(n3208) );
  XOR U3567 ( .A(n3238), .B(n3239), .Z(n3204) );
  AND U3568 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U3569 ( .A(e_input[46]), .B(n3242), .Z(n3241) );
  IV U3570 ( .A(n3209), .Z(n3232) );
  XOR U3571 ( .A(n3243), .B(n3244), .Z(n3209) );
  ANDN U3572 ( .A(n3245), .B(n3246), .Z(n3244) );
  XOR U3573 ( .A(n3243), .B(n3247), .Z(n3245) );
  XOR U3574 ( .A(n3248), .B(n3249), .Z(n3213) );
  AND U3575 ( .A(n2670), .B(n3250), .Z(n3249) );
  XNOR U3576 ( .A(n3221), .B(n3251), .Z(n3250) );
  XOR U3577 ( .A(n3252), .B(n3248), .Z(n3251) );
  IV U3578 ( .A(e_input[15]), .Z(n3252) );
  XNOR U3579 ( .A(n3223), .B(g_input[15]), .Z(n3221) );
  IV U3580 ( .A(n3219), .Z(n3223) );
  XOR U3581 ( .A(n3253), .B(n3254), .Z(n3219) );
  AND U3582 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U3583 ( .A(e_input[14]), .B(n3257), .Z(n3256) );
  XNOR U3584 ( .A(n3258), .B(g_input[15]), .Z(n3248) );
  XNOR U3585 ( .A(n3259), .B(\min_dist_reg[3][15] ), .Z(n3228) );
  IV U3586 ( .A(n3226), .Z(n3259) );
  XOR U3587 ( .A(n3260), .B(n3261), .Z(n3226) );
  AND U3588 ( .A(n3262), .B(n3263), .Z(n3261) );
  XNOR U3589 ( .A(n3260), .B(n2550), .Z(n3263) );
  XOR U3590 ( .A(n3247), .B(n3246), .Z(n2550) );
  XNOR U3591 ( .A(n3264), .B(n3265), .Z(n3246) );
  XNOR U3592 ( .A(n3266), .B(n3267), .Z(n3264) );
  AND U3593 ( .A(n2676), .B(n3268), .Z(n3267) );
  XNOR U3594 ( .A(n3240), .B(n3269), .Z(n3268) );
  XOR U3595 ( .A(n3270), .B(n3265), .Z(n3269) );
  XNOR U3596 ( .A(n3271), .B(g_input[46]), .Z(n3265) );
  IV U3597 ( .A(e_input[46]), .Z(n3270) );
  XNOR U3598 ( .A(n3242), .B(g_input[46]), .Z(n3240) );
  IV U3599 ( .A(n3238), .Z(n3242) );
  XOR U3600 ( .A(n3272), .B(n3273), .Z(n3238) );
  AND U3601 ( .A(n3274), .B(n3275), .Z(n3273) );
  XOR U3602 ( .A(e_input[45]), .B(n3276), .Z(n3275) );
  IV U3603 ( .A(n3243), .Z(n3266) );
  XOR U3604 ( .A(n3277), .B(n3278), .Z(n3243) );
  ANDN U3605 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR U3606 ( .A(n3277), .B(n3281), .Z(n3279) );
  XOR U3607 ( .A(n3282), .B(n3283), .Z(n3247) );
  AND U3608 ( .A(n2670), .B(n3284), .Z(n3283) );
  XNOR U3609 ( .A(n3255), .B(n3285), .Z(n3284) );
  XOR U3610 ( .A(n3286), .B(n3282), .Z(n3285) );
  IV U3611 ( .A(e_input[14]), .Z(n3286) );
  XNOR U3612 ( .A(n3257), .B(g_input[14]), .Z(n3255) );
  IV U3613 ( .A(n3253), .Z(n3257) );
  XOR U3614 ( .A(n3287), .B(n3288), .Z(n3253) );
  AND U3615 ( .A(n3289), .B(n3290), .Z(n3288) );
  XOR U3616 ( .A(e_input[13]), .B(n3291), .Z(n3290) );
  XNOR U3617 ( .A(n3292), .B(g_input[14]), .Z(n3282) );
  XNOR U3618 ( .A(n3293), .B(\min_dist_reg[3][14] ), .Z(n3262) );
  IV U3619 ( .A(n3260), .Z(n3293) );
  XOR U3620 ( .A(n3294), .B(n3295), .Z(n3260) );
  AND U3621 ( .A(n3296), .B(n3297), .Z(n3295) );
  XNOR U3622 ( .A(n3294), .B(n2558), .Z(n3297) );
  XOR U3623 ( .A(n3281), .B(n3280), .Z(n2558) );
  XNOR U3624 ( .A(n3298), .B(n3299), .Z(n3280) );
  XNOR U3625 ( .A(n3300), .B(n3301), .Z(n3298) );
  AND U3626 ( .A(n2676), .B(n3302), .Z(n3301) );
  XNOR U3627 ( .A(n3274), .B(n3303), .Z(n3302) );
  XOR U3628 ( .A(n3304), .B(n3299), .Z(n3303) );
  XNOR U3629 ( .A(n3305), .B(g_input[45]), .Z(n3299) );
  IV U3630 ( .A(e_input[45]), .Z(n3304) );
  XNOR U3631 ( .A(n3276), .B(g_input[45]), .Z(n3274) );
  IV U3632 ( .A(n3272), .Z(n3276) );
  XOR U3633 ( .A(n3306), .B(n3307), .Z(n3272) );
  AND U3634 ( .A(n3308), .B(n3309), .Z(n3307) );
  XOR U3635 ( .A(e_input[44]), .B(n3310), .Z(n3309) );
  IV U3636 ( .A(n3277), .Z(n3300) );
  XOR U3637 ( .A(n3311), .B(n3312), .Z(n3277) );
  ANDN U3638 ( .A(n3313), .B(n3314), .Z(n3312) );
  XOR U3639 ( .A(n3311), .B(n3315), .Z(n3313) );
  XOR U3640 ( .A(n3316), .B(n3317), .Z(n3281) );
  AND U3641 ( .A(n2670), .B(n3318), .Z(n3317) );
  XNOR U3642 ( .A(n3289), .B(n3319), .Z(n3318) );
  XOR U3643 ( .A(n3320), .B(n3316), .Z(n3319) );
  IV U3644 ( .A(e_input[13]), .Z(n3320) );
  XNOR U3645 ( .A(n3291), .B(g_input[13]), .Z(n3289) );
  IV U3646 ( .A(n3287), .Z(n3291) );
  XOR U3647 ( .A(n3321), .B(n3322), .Z(n3287) );
  AND U3648 ( .A(n3323), .B(n3324), .Z(n3322) );
  XOR U3649 ( .A(e_input[12]), .B(n3325), .Z(n3324) );
  XNOR U3650 ( .A(n3326), .B(g_input[13]), .Z(n3316) );
  XNOR U3651 ( .A(n3327), .B(\min_dist_reg[3][13] ), .Z(n3296) );
  IV U3652 ( .A(n3294), .Z(n3327) );
  XOR U3653 ( .A(n3328), .B(n3329), .Z(n3294) );
  AND U3654 ( .A(n3330), .B(n3331), .Z(n3329) );
  XNOR U3655 ( .A(n3328), .B(n2566), .Z(n3331) );
  XOR U3656 ( .A(n3315), .B(n3314), .Z(n2566) );
  XNOR U3657 ( .A(n3332), .B(n3333), .Z(n3314) );
  XNOR U3658 ( .A(n3334), .B(n3335), .Z(n3332) );
  AND U3659 ( .A(n2676), .B(n3336), .Z(n3335) );
  XNOR U3660 ( .A(n3308), .B(n3337), .Z(n3336) );
  XOR U3661 ( .A(n3338), .B(n3333), .Z(n3337) );
  XNOR U3662 ( .A(n3339), .B(g_input[44]), .Z(n3333) );
  IV U3663 ( .A(e_input[44]), .Z(n3338) );
  XNOR U3664 ( .A(n3310), .B(g_input[44]), .Z(n3308) );
  IV U3665 ( .A(n3306), .Z(n3310) );
  XOR U3666 ( .A(n3340), .B(n3341), .Z(n3306) );
  AND U3667 ( .A(n3342), .B(n3343), .Z(n3341) );
  XOR U3668 ( .A(e_input[43]), .B(n3344), .Z(n3343) );
  IV U3669 ( .A(n3311), .Z(n3334) );
  XOR U3670 ( .A(n3345), .B(n3346), .Z(n3311) );
  ANDN U3671 ( .A(n3347), .B(n3348), .Z(n3346) );
  XOR U3672 ( .A(n3345), .B(n3349), .Z(n3347) );
  XOR U3673 ( .A(n3350), .B(n3351), .Z(n3315) );
  AND U3674 ( .A(n2670), .B(n3352), .Z(n3351) );
  XNOR U3675 ( .A(n3323), .B(n3353), .Z(n3352) );
  XOR U3676 ( .A(n3354), .B(n3350), .Z(n3353) );
  IV U3677 ( .A(e_input[12]), .Z(n3354) );
  XNOR U3678 ( .A(n3325), .B(g_input[12]), .Z(n3323) );
  IV U3679 ( .A(n3321), .Z(n3325) );
  XOR U3680 ( .A(n3355), .B(n3356), .Z(n3321) );
  AND U3681 ( .A(n3357), .B(n3358), .Z(n3356) );
  XOR U3682 ( .A(e_input[11]), .B(n3359), .Z(n3358) );
  XNOR U3683 ( .A(n3360), .B(g_input[12]), .Z(n3350) );
  XNOR U3684 ( .A(n3361), .B(\min_dist_reg[3][12] ), .Z(n3330) );
  IV U3685 ( .A(n3328), .Z(n3361) );
  XOR U3686 ( .A(n3362), .B(n3363), .Z(n3328) );
  AND U3687 ( .A(n3364), .B(n3365), .Z(n3363) );
  XNOR U3688 ( .A(n3362), .B(n2574), .Z(n3365) );
  XOR U3689 ( .A(n3349), .B(n3348), .Z(n2574) );
  XNOR U3690 ( .A(n3366), .B(n3367), .Z(n3348) );
  XNOR U3691 ( .A(n3368), .B(n3369), .Z(n3366) );
  AND U3692 ( .A(n2676), .B(n3370), .Z(n3369) );
  XNOR U3693 ( .A(n3342), .B(n3371), .Z(n3370) );
  XOR U3694 ( .A(n3372), .B(n3367), .Z(n3371) );
  XNOR U3695 ( .A(n3373), .B(g_input[43]), .Z(n3367) );
  IV U3696 ( .A(e_input[43]), .Z(n3372) );
  XNOR U3697 ( .A(n3344), .B(g_input[43]), .Z(n3342) );
  IV U3698 ( .A(n3340), .Z(n3344) );
  XOR U3699 ( .A(n3374), .B(n3375), .Z(n3340) );
  AND U3700 ( .A(n3376), .B(n3377), .Z(n3375) );
  XOR U3701 ( .A(e_input[42]), .B(n3378), .Z(n3377) );
  IV U3702 ( .A(n3345), .Z(n3368) );
  XOR U3703 ( .A(n3379), .B(n3380), .Z(n3345) );
  ANDN U3704 ( .A(n3381), .B(n3382), .Z(n3380) );
  XOR U3705 ( .A(n3379), .B(n3383), .Z(n3381) );
  XOR U3706 ( .A(n3384), .B(n3385), .Z(n3349) );
  AND U3707 ( .A(n2670), .B(n3386), .Z(n3385) );
  XNOR U3708 ( .A(n3357), .B(n3387), .Z(n3386) );
  XOR U3709 ( .A(n3388), .B(n3384), .Z(n3387) );
  IV U3710 ( .A(e_input[11]), .Z(n3388) );
  XNOR U3711 ( .A(n3359), .B(g_input[11]), .Z(n3357) );
  IV U3712 ( .A(n3355), .Z(n3359) );
  XOR U3713 ( .A(n3389), .B(n3390), .Z(n3355) );
  AND U3714 ( .A(n3391), .B(n3392), .Z(n3390) );
  XOR U3715 ( .A(e_input[10]), .B(n3393), .Z(n3392) );
  XNOR U3716 ( .A(n3394), .B(g_input[11]), .Z(n3384) );
  XNOR U3717 ( .A(n3395), .B(\min_dist_reg[3][11] ), .Z(n3364) );
  IV U3718 ( .A(n3362), .Z(n3395) );
  XOR U3719 ( .A(n3396), .B(n3397), .Z(n3362) );
  AND U3720 ( .A(n3398), .B(n3399), .Z(n3397) );
  XNOR U3721 ( .A(n3396), .B(n2582), .Z(n3399) );
  XOR U3722 ( .A(n3383), .B(n3382), .Z(n2582) );
  XNOR U3723 ( .A(n3400), .B(n3401), .Z(n3382) );
  XNOR U3724 ( .A(n3402), .B(n3403), .Z(n3400) );
  AND U3725 ( .A(n2676), .B(n3404), .Z(n3403) );
  XNOR U3726 ( .A(n3376), .B(n3405), .Z(n3404) );
  XOR U3727 ( .A(n3406), .B(n3401), .Z(n3405) );
  XNOR U3728 ( .A(n3407), .B(g_input[42]), .Z(n3401) );
  IV U3729 ( .A(e_input[42]), .Z(n3406) );
  XNOR U3730 ( .A(n3378), .B(g_input[42]), .Z(n3376) );
  IV U3731 ( .A(n3374), .Z(n3378) );
  XOR U3732 ( .A(n3408), .B(n3409), .Z(n3374) );
  AND U3733 ( .A(n3410), .B(n3411), .Z(n3409) );
  XOR U3734 ( .A(e_input[41]), .B(n3412), .Z(n3411) );
  IV U3735 ( .A(n3379), .Z(n3402) );
  XOR U3736 ( .A(n3413), .B(n3414), .Z(n3379) );
  ANDN U3737 ( .A(n3415), .B(n3416), .Z(n3414) );
  XOR U3738 ( .A(n3413), .B(n3417), .Z(n3415) );
  XOR U3739 ( .A(n3418), .B(n3419), .Z(n3383) );
  AND U3740 ( .A(n2670), .B(n3420), .Z(n3419) );
  XNOR U3741 ( .A(n3391), .B(n3421), .Z(n3420) );
  XOR U3742 ( .A(n3422), .B(n3418), .Z(n3421) );
  IV U3743 ( .A(e_input[10]), .Z(n3422) );
  XNOR U3744 ( .A(n3393), .B(g_input[10]), .Z(n3391) );
  IV U3745 ( .A(n3389), .Z(n3393) );
  XOR U3746 ( .A(n3423), .B(n3424), .Z(n3389) );
  AND U3747 ( .A(n3425), .B(n3426), .Z(n3424) );
  XOR U3748 ( .A(e_input[9]), .B(n3427), .Z(n3426) );
  XNOR U3749 ( .A(n3428), .B(g_input[10]), .Z(n3418) );
  XNOR U3750 ( .A(n3429), .B(\min_dist_reg[3][10] ), .Z(n3398) );
  IV U3751 ( .A(n3396), .Z(n3429) );
  XOR U3752 ( .A(n3430), .B(n3431), .Z(n3396) );
  AND U3753 ( .A(n3432), .B(n3433), .Z(n3431) );
  XNOR U3754 ( .A(n3430), .B(n2590), .Z(n3433) );
  XOR U3755 ( .A(n3417), .B(n3416), .Z(n2590) );
  XNOR U3756 ( .A(n3434), .B(n3435), .Z(n3416) );
  XNOR U3757 ( .A(n3436), .B(n3437), .Z(n3434) );
  AND U3758 ( .A(n2676), .B(n3438), .Z(n3437) );
  XNOR U3759 ( .A(n3410), .B(n3439), .Z(n3438) );
  XOR U3760 ( .A(n3440), .B(n3435), .Z(n3439) );
  XNOR U3761 ( .A(n3441), .B(g_input[41]), .Z(n3435) );
  IV U3762 ( .A(e_input[41]), .Z(n3440) );
  XNOR U3763 ( .A(n3412), .B(g_input[41]), .Z(n3410) );
  IV U3764 ( .A(n3408), .Z(n3412) );
  XOR U3765 ( .A(n3442), .B(n3443), .Z(n3408) );
  AND U3766 ( .A(n3444), .B(n3445), .Z(n3443) );
  XOR U3767 ( .A(e_input[40]), .B(n3446), .Z(n3445) );
  IV U3768 ( .A(n3413), .Z(n3436) );
  XOR U3769 ( .A(n3447), .B(n3448), .Z(n3413) );
  ANDN U3770 ( .A(n3449), .B(n3450), .Z(n3448) );
  XOR U3771 ( .A(n3447), .B(n3451), .Z(n3449) );
  XOR U3772 ( .A(n3452), .B(n3453), .Z(n3417) );
  AND U3773 ( .A(n2670), .B(n3454), .Z(n3453) );
  XNOR U3774 ( .A(n3425), .B(n3455), .Z(n3454) );
  XOR U3775 ( .A(n3456), .B(n3452), .Z(n3455) );
  IV U3776 ( .A(e_input[9]), .Z(n3456) );
  XNOR U3777 ( .A(n3427), .B(g_input[9]), .Z(n3425) );
  IV U3778 ( .A(n3423), .Z(n3427) );
  XOR U3779 ( .A(n3457), .B(n3458), .Z(n3423) );
  AND U3780 ( .A(n3459), .B(n3460), .Z(n3458) );
  XOR U3781 ( .A(e_input[8]), .B(n3461), .Z(n3460) );
  XNOR U3782 ( .A(n3462), .B(g_input[9]), .Z(n3452) );
  XNOR U3783 ( .A(n3463), .B(\min_dist_reg[3][9] ), .Z(n3432) );
  IV U3784 ( .A(n3430), .Z(n3463) );
  XOR U3785 ( .A(n3464), .B(n3465), .Z(n3430) );
  AND U3786 ( .A(n3466), .B(n3467), .Z(n3465) );
  XNOR U3787 ( .A(n3464), .B(n2598), .Z(n3467) );
  XOR U3788 ( .A(n3451), .B(n3450), .Z(n2598) );
  XNOR U3789 ( .A(n3468), .B(n3469), .Z(n3450) );
  XNOR U3790 ( .A(n3470), .B(n3471), .Z(n3468) );
  AND U3791 ( .A(n2676), .B(n3472), .Z(n3471) );
  XNOR U3792 ( .A(n3444), .B(n3473), .Z(n3472) );
  XOR U3793 ( .A(n3474), .B(n3469), .Z(n3473) );
  XNOR U3794 ( .A(n3475), .B(g_input[40]), .Z(n3469) );
  IV U3795 ( .A(e_input[40]), .Z(n3474) );
  XNOR U3796 ( .A(n3446), .B(g_input[40]), .Z(n3444) );
  IV U3797 ( .A(n3442), .Z(n3446) );
  XOR U3798 ( .A(n3476), .B(n3477), .Z(n3442) );
  AND U3799 ( .A(n3478), .B(n3479), .Z(n3477) );
  XOR U3800 ( .A(e_input[39]), .B(n3480), .Z(n3479) );
  IV U3801 ( .A(n3447), .Z(n3470) );
  XOR U3802 ( .A(n3481), .B(n3482), .Z(n3447) );
  ANDN U3803 ( .A(n3483), .B(n3484), .Z(n3482) );
  XOR U3804 ( .A(n3481), .B(n3485), .Z(n3483) );
  XOR U3805 ( .A(n3486), .B(n3487), .Z(n3451) );
  AND U3806 ( .A(n2670), .B(n3488), .Z(n3487) );
  XNOR U3807 ( .A(n3459), .B(n3489), .Z(n3488) );
  XOR U3808 ( .A(n3490), .B(n3486), .Z(n3489) );
  IV U3809 ( .A(e_input[8]), .Z(n3490) );
  XNOR U3810 ( .A(n3461), .B(g_input[8]), .Z(n3459) );
  IV U3811 ( .A(n3457), .Z(n3461) );
  XOR U3812 ( .A(n3491), .B(n3492), .Z(n3457) );
  AND U3813 ( .A(n3493), .B(n3494), .Z(n3492) );
  XOR U3814 ( .A(e_input[7]), .B(n3495), .Z(n3494) );
  XNOR U3815 ( .A(n3496), .B(g_input[8]), .Z(n3486) );
  XNOR U3816 ( .A(n3497), .B(\min_dist_reg[3][8] ), .Z(n3466) );
  IV U3817 ( .A(n3464), .Z(n3497) );
  XOR U3818 ( .A(n3498), .B(n3499), .Z(n3464) );
  AND U3819 ( .A(n3500), .B(n3501), .Z(n3499) );
  XNOR U3820 ( .A(n3498), .B(n2606), .Z(n3501) );
  XOR U3821 ( .A(n3485), .B(n3484), .Z(n2606) );
  XNOR U3822 ( .A(n3502), .B(n3503), .Z(n3484) );
  XNOR U3823 ( .A(n3504), .B(n3505), .Z(n3502) );
  AND U3824 ( .A(n2676), .B(n3506), .Z(n3505) );
  XNOR U3825 ( .A(n3478), .B(n3507), .Z(n3506) );
  XOR U3826 ( .A(n3508), .B(n3503), .Z(n3507) );
  XNOR U3827 ( .A(n3509), .B(g_input[39]), .Z(n3503) );
  IV U3828 ( .A(e_input[39]), .Z(n3508) );
  XNOR U3829 ( .A(n3480), .B(g_input[39]), .Z(n3478) );
  IV U3830 ( .A(n3476), .Z(n3480) );
  XOR U3831 ( .A(n3510), .B(n3511), .Z(n3476) );
  AND U3832 ( .A(n3512), .B(n3513), .Z(n3511) );
  XOR U3833 ( .A(e_input[38]), .B(n3514), .Z(n3513) );
  IV U3834 ( .A(n3481), .Z(n3504) );
  XOR U3835 ( .A(n3515), .B(n3516), .Z(n3481) );
  ANDN U3836 ( .A(n3517), .B(n3518), .Z(n3516) );
  XOR U3837 ( .A(n3515), .B(n3519), .Z(n3517) );
  XOR U3838 ( .A(n3520), .B(n3521), .Z(n3485) );
  AND U3839 ( .A(n2670), .B(n3522), .Z(n3521) );
  XNOR U3840 ( .A(n3493), .B(n3523), .Z(n3522) );
  XOR U3841 ( .A(n3524), .B(n3520), .Z(n3523) );
  IV U3842 ( .A(e_input[7]), .Z(n3524) );
  XNOR U3843 ( .A(n3495), .B(g_input[7]), .Z(n3493) );
  IV U3844 ( .A(n3491), .Z(n3495) );
  XOR U3845 ( .A(n3525), .B(n3526), .Z(n3491) );
  AND U3846 ( .A(n3527), .B(n3528), .Z(n3526) );
  XOR U3847 ( .A(e_input[6]), .B(n3529), .Z(n3528) );
  XNOR U3848 ( .A(n3530), .B(g_input[7]), .Z(n3520) );
  XNOR U3849 ( .A(n3531), .B(\min_dist_reg[3][7] ), .Z(n3500) );
  IV U3850 ( .A(n3498), .Z(n3531) );
  XOR U3851 ( .A(n3532), .B(n3533), .Z(n3498) );
  AND U3852 ( .A(n3534), .B(n3535), .Z(n3533) );
  XNOR U3853 ( .A(n3532), .B(n2614), .Z(n3535) );
  XOR U3854 ( .A(n3519), .B(n3518), .Z(n2614) );
  XNOR U3855 ( .A(n3536), .B(n3537), .Z(n3518) );
  XNOR U3856 ( .A(n3538), .B(n3539), .Z(n3536) );
  AND U3857 ( .A(n2676), .B(n3540), .Z(n3539) );
  XNOR U3858 ( .A(n3512), .B(n3541), .Z(n3540) );
  XOR U3859 ( .A(n3542), .B(n3537), .Z(n3541) );
  XNOR U3860 ( .A(n3543), .B(g_input[38]), .Z(n3537) );
  IV U3861 ( .A(e_input[38]), .Z(n3542) );
  XNOR U3862 ( .A(n3514), .B(g_input[38]), .Z(n3512) );
  IV U3863 ( .A(n3510), .Z(n3514) );
  XOR U3864 ( .A(n3544), .B(n3545), .Z(n3510) );
  AND U3865 ( .A(n3546), .B(n3547), .Z(n3545) );
  XOR U3866 ( .A(e_input[37]), .B(n3548), .Z(n3547) );
  IV U3867 ( .A(n3515), .Z(n3538) );
  XOR U3868 ( .A(n3549), .B(n3550), .Z(n3515) );
  ANDN U3869 ( .A(n3551), .B(n3552), .Z(n3550) );
  XOR U3870 ( .A(n3549), .B(n3553), .Z(n3551) );
  XOR U3871 ( .A(n3554), .B(n3555), .Z(n3519) );
  AND U3872 ( .A(n2670), .B(n3556), .Z(n3555) );
  XNOR U3873 ( .A(n3527), .B(n3557), .Z(n3556) );
  XOR U3874 ( .A(n3558), .B(n3554), .Z(n3557) );
  IV U3875 ( .A(e_input[6]), .Z(n3558) );
  XNOR U3876 ( .A(n3529), .B(g_input[6]), .Z(n3527) );
  IV U3877 ( .A(n3525), .Z(n3529) );
  XOR U3878 ( .A(n3559), .B(n3560), .Z(n3525) );
  AND U3879 ( .A(n3561), .B(n3562), .Z(n3560) );
  XOR U3880 ( .A(e_input[5]), .B(n3563), .Z(n3562) );
  XNOR U3881 ( .A(n3564), .B(g_input[6]), .Z(n3554) );
  XNOR U3882 ( .A(n3565), .B(\min_dist_reg[3][6] ), .Z(n3534) );
  IV U3883 ( .A(n3532), .Z(n3565) );
  XOR U3884 ( .A(n3566), .B(n3567), .Z(n3532) );
  AND U3885 ( .A(n3568), .B(n3569), .Z(n3567) );
  XNOR U3886 ( .A(n3566), .B(n2622), .Z(n3569) );
  XOR U3887 ( .A(n3553), .B(n3552), .Z(n2622) );
  XNOR U3888 ( .A(n3570), .B(n3571), .Z(n3552) );
  XNOR U3889 ( .A(n3572), .B(n3573), .Z(n3570) );
  AND U3890 ( .A(n2676), .B(n3574), .Z(n3573) );
  XNOR U3891 ( .A(n3546), .B(n3575), .Z(n3574) );
  XOR U3892 ( .A(n3576), .B(n3571), .Z(n3575) );
  XNOR U3893 ( .A(n3577), .B(g_input[37]), .Z(n3571) );
  IV U3894 ( .A(e_input[37]), .Z(n3576) );
  XNOR U3895 ( .A(n3548), .B(g_input[37]), .Z(n3546) );
  IV U3896 ( .A(n3544), .Z(n3548) );
  XOR U3897 ( .A(n3578), .B(n3579), .Z(n3544) );
  AND U3898 ( .A(n3580), .B(n3581), .Z(n3579) );
  XOR U3899 ( .A(e_input[36]), .B(n3582), .Z(n3581) );
  IV U3900 ( .A(n3549), .Z(n3572) );
  XOR U3901 ( .A(n3583), .B(n3584), .Z(n3549) );
  ANDN U3902 ( .A(n3585), .B(n3586), .Z(n3584) );
  XOR U3903 ( .A(n3583), .B(n3587), .Z(n3585) );
  XOR U3904 ( .A(n3588), .B(n3589), .Z(n3553) );
  AND U3905 ( .A(n2670), .B(n3590), .Z(n3589) );
  XNOR U3906 ( .A(n3561), .B(n3591), .Z(n3590) );
  XOR U3907 ( .A(n3592), .B(n3588), .Z(n3591) );
  IV U3908 ( .A(e_input[5]), .Z(n3592) );
  XNOR U3909 ( .A(n3563), .B(g_input[5]), .Z(n3561) );
  IV U3910 ( .A(n3559), .Z(n3563) );
  XOR U3911 ( .A(n3593), .B(n3594), .Z(n3559) );
  AND U3912 ( .A(n3595), .B(n3596), .Z(n3594) );
  XOR U3913 ( .A(e_input[4]), .B(n3597), .Z(n3596) );
  XNOR U3914 ( .A(n3598), .B(g_input[5]), .Z(n3588) );
  XNOR U3915 ( .A(n3599), .B(\min_dist_reg[3][5] ), .Z(n3568) );
  IV U3916 ( .A(n3566), .Z(n3599) );
  XOR U3917 ( .A(n3600), .B(n3601), .Z(n3566) );
  AND U3918 ( .A(n3602), .B(n3603), .Z(n3601) );
  XNOR U3919 ( .A(n3600), .B(n2630), .Z(n3603) );
  XOR U3920 ( .A(n3587), .B(n3586), .Z(n2630) );
  XNOR U3921 ( .A(n3604), .B(n3605), .Z(n3586) );
  XNOR U3922 ( .A(n3606), .B(n3607), .Z(n3604) );
  AND U3923 ( .A(n2676), .B(n3608), .Z(n3607) );
  XNOR U3924 ( .A(n3580), .B(n3609), .Z(n3608) );
  XOR U3925 ( .A(n3610), .B(n3605), .Z(n3609) );
  XNOR U3926 ( .A(n3611), .B(g_input[36]), .Z(n3605) );
  IV U3927 ( .A(e_input[36]), .Z(n3610) );
  XNOR U3928 ( .A(n3582), .B(g_input[36]), .Z(n3580) );
  IV U3929 ( .A(n3578), .Z(n3582) );
  XOR U3930 ( .A(n3612), .B(n3613), .Z(n3578) );
  AND U3931 ( .A(n3614), .B(n3615), .Z(n3613) );
  XOR U3932 ( .A(e_input[35]), .B(n3616), .Z(n3615) );
  IV U3933 ( .A(n3583), .Z(n3606) );
  XOR U3934 ( .A(n3617), .B(n3618), .Z(n3583) );
  ANDN U3935 ( .A(n3619), .B(n3620), .Z(n3618) );
  XOR U3936 ( .A(n3617), .B(n3621), .Z(n3619) );
  XOR U3937 ( .A(n3622), .B(n3623), .Z(n3587) );
  AND U3938 ( .A(n2670), .B(n3624), .Z(n3623) );
  XNOR U3939 ( .A(n3595), .B(n3625), .Z(n3624) );
  XOR U3940 ( .A(n3626), .B(n3622), .Z(n3625) );
  IV U3941 ( .A(e_input[4]), .Z(n3626) );
  XNOR U3942 ( .A(n3597), .B(g_input[4]), .Z(n3595) );
  IV U3943 ( .A(n3593), .Z(n3597) );
  XOR U3944 ( .A(n3627), .B(n3628), .Z(n3593) );
  AND U3945 ( .A(n3629), .B(n3630), .Z(n3628) );
  XOR U3946 ( .A(e_input[3]), .B(n3631), .Z(n3630) );
  XNOR U3947 ( .A(n3632), .B(g_input[4]), .Z(n3622) );
  XNOR U3948 ( .A(n3633), .B(\min_dist_reg[3][4] ), .Z(n3602) );
  IV U3949 ( .A(n3600), .Z(n3633) );
  XOR U3950 ( .A(n3634), .B(n3635), .Z(n3600) );
  AND U3951 ( .A(n3636), .B(n3637), .Z(n3635) );
  XNOR U3952 ( .A(n3634), .B(n2636), .Z(n3637) );
  XOR U3953 ( .A(n3621), .B(n3620), .Z(n2636) );
  XNOR U3954 ( .A(n3638), .B(n3639), .Z(n3620) );
  XNOR U3955 ( .A(n3640), .B(n3641), .Z(n3638) );
  AND U3956 ( .A(n2676), .B(n3642), .Z(n3641) );
  XNOR U3957 ( .A(n3614), .B(n3643), .Z(n3642) );
  XOR U3958 ( .A(n3644), .B(n3639), .Z(n3643) );
  XNOR U3959 ( .A(n3645), .B(g_input[35]), .Z(n3639) );
  IV U3960 ( .A(e_input[35]), .Z(n3644) );
  XNOR U3961 ( .A(n3616), .B(g_input[35]), .Z(n3614) );
  IV U3962 ( .A(n3612), .Z(n3616) );
  XOR U3963 ( .A(n3646), .B(n3647), .Z(n3612) );
  AND U3964 ( .A(n3648), .B(n3649), .Z(n3647) );
  XNOR U3965 ( .A(e_input[34]), .B(n3646), .Z(n3649) );
  IV U3966 ( .A(n3617), .Z(n3640) );
  XOR U3967 ( .A(n3650), .B(n3651), .Z(n3617) );
  ANDN U3968 ( .A(n3652), .B(n3653), .Z(n3651) );
  XOR U3969 ( .A(n3650), .B(n3654), .Z(n3652) );
  XOR U3970 ( .A(n3655), .B(n3656), .Z(n3621) );
  AND U3971 ( .A(n2670), .B(n3657), .Z(n3656) );
  XNOR U3972 ( .A(n3629), .B(n3658), .Z(n3657) );
  XOR U3973 ( .A(n3659), .B(n3655), .Z(n3658) );
  IV U3974 ( .A(e_input[3]), .Z(n3659) );
  XNOR U3975 ( .A(n3631), .B(g_input[3]), .Z(n3629) );
  IV U3976 ( .A(n3627), .Z(n3631) );
  XOR U3977 ( .A(n3660), .B(n3661), .Z(n3627) );
  AND U3978 ( .A(n3662), .B(n3663), .Z(n3661) );
  XNOR U3979 ( .A(e_input[2]), .B(n3660), .Z(n3663) );
  XNOR U3980 ( .A(n3664), .B(g_input[3]), .Z(n3655) );
  XNOR U3981 ( .A(n3665), .B(\min_dist_reg[3][3] ), .Z(n3636) );
  IV U3982 ( .A(n3634), .Z(n3665) );
  XOR U3983 ( .A(n3666), .B(n3667), .Z(n3634) );
  AND U3984 ( .A(n3668), .B(n3669), .Z(n3667) );
  XNOR U3985 ( .A(n3666), .B(n2643), .Z(n3669) );
  XOR U3986 ( .A(n3654), .B(n3653), .Z(n2643) );
  XNOR U3987 ( .A(n3670), .B(n3671), .Z(n3653) );
  XOR U3988 ( .A(n3650), .B(n3672), .Z(n3670) );
  AND U3989 ( .A(n2676), .B(n3673), .Z(n3672) );
  XNOR U3990 ( .A(n3648), .B(n3674), .Z(n3673) );
  XOR U3991 ( .A(n3675), .B(n3671), .Z(n3674) );
  XNOR U3992 ( .A(n3676), .B(g_input[34]), .Z(n3671) );
  IV U3993 ( .A(e_input[34]), .Z(n3675) );
  XOR U3994 ( .A(n3646), .B(g_input[34]), .Z(n3648) );
  XOR U3995 ( .A(n3677), .B(n3678), .Z(n3646) );
  NAND U3996 ( .A(n3679), .B(n3680), .Z(n3677) );
  XOR U3997 ( .A(e_input[33]), .B(n3678), .Z(n3679) );
  XNOR U3998 ( .A(n3681), .B(n3682), .Z(n3650) );
  NANDN U3999 ( .B(n3683), .A(n3684), .Z(n3681) );
  XOR U4000 ( .A(n3682), .B(n3685), .Z(n3684) );
  XOR U4001 ( .A(n3686), .B(n3687), .Z(n3654) );
  AND U4002 ( .A(n2670), .B(n3688), .Z(n3687) );
  XNOR U4003 ( .A(n3662), .B(n3689), .Z(n3688) );
  XOR U4004 ( .A(n3690), .B(n3686), .Z(n3689) );
  IV U4005 ( .A(e_input[2]), .Z(n3690) );
  XNOR U4006 ( .A(n3660), .B(n3691), .Z(n3662) );
  XOR U4007 ( .A(n3692), .B(n3693), .Z(n3660) );
  NAND U4008 ( .A(n3694), .B(n3695), .Z(n3692) );
  XOR U4009 ( .A(e_input[1]), .B(n3693), .Z(n3694) );
  XNOR U4010 ( .A(n3696), .B(g_input[2]), .Z(n3686) );
  XOR U4011 ( .A(n3666), .B(\min_dist_reg[3][2] ), .Z(n3668) );
  XOR U4012 ( .A(n3697), .B(n3698), .Z(n3666) );
  NAND U4013 ( .A(n3699), .B(n3700), .Z(n3697) );
  XOR U4014 ( .A(n3698), .B(n2650), .Z(n3700) );
  XOR U4015 ( .A(n3685), .B(n3683), .Z(n2650) );
  XNOR U4016 ( .A(n3701), .B(n3702), .Z(n3683) );
  XNOR U4017 ( .A(n3703), .B(n3682), .Z(n3701) );
  OR U4018 ( .A(n3704), .B(n3705), .Z(n3682) );
  NAND U4019 ( .A(n3706), .B(n2676), .Z(n3703) );
  XOR U4020 ( .A(n3707), .B(n3708), .Z(n2676) );
  ANDN U4021 ( .A(n3709), .B(n2703), .Z(n3708) );
  XOR U4022 ( .A(n3707), .B(e_input[63]), .Z(n2703) );
  XNOR U4023 ( .A(n2698), .B(n3707), .Z(n3709) );
  IV U4024 ( .A(g_input[63]), .Z(n2698) );
  XOR U4025 ( .A(n3710), .B(n3711), .Z(n3707) );
  ANDN U4026 ( .A(n3712), .B(n2731), .Z(n3711) );
  XOR U4027 ( .A(n3710), .B(e_input[62]), .Z(n2731) );
  XOR U4028 ( .A(g_input[62]), .B(n3710), .Z(n3712) );
  XOR U4029 ( .A(n3713), .B(n3714), .Z(n3710) );
  ANDN U4030 ( .A(n3715), .B(n2761), .Z(n3714) );
  XOR U4031 ( .A(n3713), .B(e_input[61]), .Z(n2761) );
  XOR U4032 ( .A(g_input[61]), .B(n3713), .Z(n3715) );
  XOR U4033 ( .A(n3716), .B(n3717), .Z(n3713) );
  ANDN U4034 ( .A(n3718), .B(n2795), .Z(n3717) );
  XOR U4035 ( .A(n3716), .B(e_input[60]), .Z(n2795) );
  XOR U4036 ( .A(g_input[60]), .B(n3716), .Z(n3718) );
  XOR U4037 ( .A(n3719), .B(n3720), .Z(n3716) );
  ANDN U4038 ( .A(n3721), .B(n2829), .Z(n3720) );
  XOR U4039 ( .A(n3719), .B(e_input[59]), .Z(n2829) );
  XOR U4040 ( .A(g_input[59]), .B(n3719), .Z(n3721) );
  XOR U4041 ( .A(n3722), .B(n3723), .Z(n3719) );
  ANDN U4042 ( .A(n3724), .B(n2863), .Z(n3723) );
  XOR U4043 ( .A(n3722), .B(e_input[58]), .Z(n2863) );
  XOR U4044 ( .A(g_input[58]), .B(n3722), .Z(n3724) );
  XOR U4045 ( .A(n3725), .B(n3726), .Z(n3722) );
  ANDN U4046 ( .A(n3727), .B(n2897), .Z(n3726) );
  XOR U4047 ( .A(n3725), .B(e_input[57]), .Z(n2897) );
  XOR U4048 ( .A(g_input[57]), .B(n3725), .Z(n3727) );
  XOR U4049 ( .A(n3728), .B(n3729), .Z(n3725) );
  ANDN U4050 ( .A(n3730), .B(n2931), .Z(n3729) );
  XOR U4051 ( .A(n3728), .B(e_input[56]), .Z(n2931) );
  XOR U4052 ( .A(g_input[56]), .B(n3728), .Z(n3730) );
  XOR U4053 ( .A(n3731), .B(n3732), .Z(n3728) );
  ANDN U4054 ( .A(n3733), .B(n2965), .Z(n3732) );
  XOR U4055 ( .A(n3731), .B(e_input[55]), .Z(n2965) );
  XOR U4056 ( .A(g_input[55]), .B(n3731), .Z(n3733) );
  XOR U4057 ( .A(n3734), .B(n3735), .Z(n3731) );
  ANDN U4058 ( .A(n3736), .B(n2999), .Z(n3735) );
  XOR U4059 ( .A(n3734), .B(e_input[54]), .Z(n2999) );
  XOR U4060 ( .A(g_input[54]), .B(n3734), .Z(n3736) );
  XOR U4061 ( .A(n3737), .B(n3738), .Z(n3734) );
  ANDN U4062 ( .A(n3739), .B(n3033), .Z(n3738) );
  XOR U4063 ( .A(n3737), .B(e_input[53]), .Z(n3033) );
  XOR U4064 ( .A(g_input[53]), .B(n3737), .Z(n3739) );
  XOR U4065 ( .A(n3740), .B(n3741), .Z(n3737) );
  ANDN U4066 ( .A(n3742), .B(n3067), .Z(n3741) );
  XOR U4067 ( .A(n3740), .B(e_input[52]), .Z(n3067) );
  XOR U4068 ( .A(g_input[52]), .B(n3740), .Z(n3742) );
  XOR U4069 ( .A(n3743), .B(n3744), .Z(n3740) );
  ANDN U4070 ( .A(n3745), .B(n3101), .Z(n3744) );
  XOR U4071 ( .A(n3743), .B(e_input[51]), .Z(n3101) );
  XOR U4072 ( .A(g_input[51]), .B(n3743), .Z(n3745) );
  XOR U4073 ( .A(n3746), .B(n3747), .Z(n3743) );
  ANDN U4074 ( .A(n3748), .B(n3135), .Z(n3747) );
  XOR U4075 ( .A(n3746), .B(e_input[50]), .Z(n3135) );
  XOR U4076 ( .A(g_input[50]), .B(n3746), .Z(n3748) );
  XOR U4077 ( .A(n3749), .B(n3750), .Z(n3746) );
  ANDN U4078 ( .A(n3751), .B(n3169), .Z(n3750) );
  XOR U4079 ( .A(n3749), .B(e_input[49]), .Z(n3169) );
  XOR U4080 ( .A(g_input[49]), .B(n3749), .Z(n3751) );
  XOR U4081 ( .A(n3752), .B(n3753), .Z(n3749) );
  ANDN U4082 ( .A(n3754), .B(n3203), .Z(n3753) );
  XOR U4083 ( .A(n3752), .B(e_input[48]), .Z(n3203) );
  XOR U4084 ( .A(g_input[48]), .B(n3752), .Z(n3754) );
  XOR U4085 ( .A(n3755), .B(n3756), .Z(n3752) );
  ANDN U4086 ( .A(n3757), .B(n3237), .Z(n3756) );
  XOR U4087 ( .A(n3755), .B(e_input[47]), .Z(n3237) );
  XOR U4088 ( .A(g_input[47]), .B(n3755), .Z(n3757) );
  XOR U4089 ( .A(n3758), .B(n3759), .Z(n3755) );
  ANDN U4090 ( .A(n3760), .B(n3271), .Z(n3759) );
  XOR U4091 ( .A(n3758), .B(e_input[46]), .Z(n3271) );
  XOR U4092 ( .A(g_input[46]), .B(n3758), .Z(n3760) );
  XOR U4093 ( .A(n3761), .B(n3762), .Z(n3758) );
  ANDN U4094 ( .A(n3763), .B(n3305), .Z(n3762) );
  XOR U4095 ( .A(n3761), .B(e_input[45]), .Z(n3305) );
  XOR U4096 ( .A(g_input[45]), .B(n3761), .Z(n3763) );
  XOR U4097 ( .A(n3764), .B(n3765), .Z(n3761) );
  ANDN U4098 ( .A(n3766), .B(n3339), .Z(n3765) );
  XOR U4099 ( .A(n3764), .B(e_input[44]), .Z(n3339) );
  XOR U4100 ( .A(g_input[44]), .B(n3764), .Z(n3766) );
  XOR U4101 ( .A(n3767), .B(n3768), .Z(n3764) );
  ANDN U4102 ( .A(n3769), .B(n3373), .Z(n3768) );
  XOR U4103 ( .A(n3767), .B(e_input[43]), .Z(n3373) );
  XOR U4104 ( .A(g_input[43]), .B(n3767), .Z(n3769) );
  XOR U4105 ( .A(n3770), .B(n3771), .Z(n3767) );
  ANDN U4106 ( .A(n3772), .B(n3407), .Z(n3771) );
  XOR U4107 ( .A(n3770), .B(e_input[42]), .Z(n3407) );
  XOR U4108 ( .A(g_input[42]), .B(n3770), .Z(n3772) );
  XOR U4109 ( .A(n3773), .B(n3774), .Z(n3770) );
  ANDN U4110 ( .A(n3775), .B(n3441), .Z(n3774) );
  XOR U4111 ( .A(n3773), .B(e_input[41]), .Z(n3441) );
  XOR U4112 ( .A(g_input[41]), .B(n3773), .Z(n3775) );
  XOR U4113 ( .A(n3776), .B(n3777), .Z(n3773) );
  ANDN U4114 ( .A(n3778), .B(n3475), .Z(n3777) );
  XOR U4115 ( .A(n3776), .B(e_input[40]), .Z(n3475) );
  XOR U4116 ( .A(g_input[40]), .B(n3776), .Z(n3778) );
  XOR U4117 ( .A(n3779), .B(n3780), .Z(n3776) );
  ANDN U4118 ( .A(n3781), .B(n3509), .Z(n3780) );
  XOR U4119 ( .A(n3779), .B(e_input[39]), .Z(n3509) );
  XOR U4120 ( .A(g_input[39]), .B(n3779), .Z(n3781) );
  XOR U4121 ( .A(n3782), .B(n3783), .Z(n3779) );
  ANDN U4122 ( .A(n3784), .B(n3543), .Z(n3783) );
  XOR U4123 ( .A(n3782), .B(e_input[38]), .Z(n3543) );
  XOR U4124 ( .A(g_input[38]), .B(n3782), .Z(n3784) );
  XOR U4125 ( .A(n3785), .B(n3786), .Z(n3782) );
  ANDN U4126 ( .A(n3787), .B(n3577), .Z(n3786) );
  XOR U4127 ( .A(n3785), .B(e_input[37]), .Z(n3577) );
  XOR U4128 ( .A(g_input[37]), .B(n3785), .Z(n3787) );
  XOR U4129 ( .A(n3788), .B(n3789), .Z(n3785) );
  ANDN U4130 ( .A(n3790), .B(n3611), .Z(n3789) );
  XOR U4131 ( .A(n3788), .B(e_input[36]), .Z(n3611) );
  XOR U4132 ( .A(g_input[36]), .B(n3788), .Z(n3790) );
  XOR U4133 ( .A(n3791), .B(n3792), .Z(n3788) );
  ANDN U4134 ( .A(n3793), .B(n3645), .Z(n3792) );
  XOR U4135 ( .A(n3791), .B(e_input[35]), .Z(n3645) );
  XOR U4136 ( .A(g_input[35]), .B(n3791), .Z(n3793) );
  XOR U4137 ( .A(n3794), .B(n3795), .Z(n3791) );
  ANDN U4138 ( .A(n3796), .B(n3676), .Z(n3795) );
  XOR U4139 ( .A(n3794), .B(e_input[34]), .Z(n3676) );
  XOR U4140 ( .A(g_input[34]), .B(n3794), .Z(n3796) );
  XNOR U4141 ( .A(n3797), .B(n3798), .Z(n3794) );
  NANDN U4142 ( .B(n3799), .A(n3800), .Z(n3797) );
  XOR U4143 ( .A(g_input[33]), .B(n3798), .Z(n3800) );
  XNOR U4144 ( .A(n3680), .B(n3801), .Z(n3706) );
  XNOR U4145 ( .A(e_input[33]), .B(n3702), .Z(n3801) );
  XNOR U4146 ( .A(n3799), .B(g_input[33]), .Z(n3702) );
  XOR U4147 ( .A(n3798), .B(e_input[33]), .Z(n3799) );
  ANDN U4148 ( .A(g_input[32]), .B(e_input[32]), .Z(n3798) );
  XNOR U4149 ( .A(n3678), .B(g_input[33]), .Z(n3680) );
  ANDN U4150 ( .A(e_input[32]), .B(g_input[32]), .Z(n3678) );
  XOR U4151 ( .A(n3802), .B(n3803), .Z(n3685) );
  AND U4152 ( .A(n2670), .B(n3804), .Z(n3803) );
  XNOR U4153 ( .A(n3695), .B(n3805), .Z(n3804) );
  XNOR U4154 ( .A(e_input[1]), .B(n3802), .Z(n3805) );
  XNOR U4155 ( .A(n3693), .B(g_input[1]), .Z(n3695) );
  ANDN U4156 ( .A(e_input[0]), .B(g_input[0]), .Z(n3693) );
  XOR U4157 ( .A(n3806), .B(n3807), .Z(n2670) );
  ANDN U4158 ( .A(n3808), .B(n2718), .Z(n3807) );
  XOR U4159 ( .A(n3806), .B(e_input[31]), .Z(n2718) );
  XNOR U4160 ( .A(n2713), .B(n3806), .Z(n3808) );
  IV U4161 ( .A(g_input[31]), .Z(n2713) );
  XOR U4162 ( .A(n3809), .B(n3810), .Z(n3806) );
  ANDN U4163 ( .A(n3811), .B(n2748), .Z(n3810) );
  XOR U4164 ( .A(n3809), .B(e_input[30]), .Z(n2748) );
  XOR U4165 ( .A(g_input[30]), .B(n3809), .Z(n3811) );
  XOR U4166 ( .A(n3812), .B(n3813), .Z(n3809) );
  ANDN U4167 ( .A(n3814), .B(n2782), .Z(n3813) );
  XOR U4168 ( .A(n3812), .B(e_input[29]), .Z(n2782) );
  XOR U4169 ( .A(g_input[29]), .B(n3812), .Z(n3814) );
  XOR U4170 ( .A(n3815), .B(n3816), .Z(n3812) );
  ANDN U4171 ( .A(n3817), .B(n2816), .Z(n3816) );
  XOR U4172 ( .A(n3815), .B(e_input[28]), .Z(n2816) );
  XOR U4173 ( .A(g_input[28]), .B(n3815), .Z(n3817) );
  XOR U4174 ( .A(n3818), .B(n3819), .Z(n3815) );
  ANDN U4175 ( .A(n3820), .B(n2850), .Z(n3819) );
  XOR U4176 ( .A(n3818), .B(e_input[27]), .Z(n2850) );
  XOR U4177 ( .A(g_input[27]), .B(n3818), .Z(n3820) );
  XOR U4178 ( .A(n3821), .B(n3822), .Z(n3818) );
  ANDN U4179 ( .A(n3823), .B(n2884), .Z(n3822) );
  XOR U4180 ( .A(n3821), .B(e_input[26]), .Z(n2884) );
  XOR U4181 ( .A(g_input[26]), .B(n3821), .Z(n3823) );
  XOR U4182 ( .A(n3824), .B(n3825), .Z(n3821) );
  ANDN U4183 ( .A(n3826), .B(n2918), .Z(n3825) );
  XOR U4184 ( .A(n3824), .B(e_input[25]), .Z(n2918) );
  XOR U4185 ( .A(g_input[25]), .B(n3824), .Z(n3826) );
  XOR U4186 ( .A(n3827), .B(n3828), .Z(n3824) );
  ANDN U4187 ( .A(n3829), .B(n2952), .Z(n3828) );
  XOR U4188 ( .A(n3827), .B(e_input[24]), .Z(n2952) );
  XOR U4189 ( .A(g_input[24]), .B(n3827), .Z(n3829) );
  XOR U4190 ( .A(n3830), .B(n3831), .Z(n3827) );
  ANDN U4191 ( .A(n3832), .B(n2986), .Z(n3831) );
  XOR U4192 ( .A(n3830), .B(e_input[23]), .Z(n2986) );
  XOR U4193 ( .A(g_input[23]), .B(n3830), .Z(n3832) );
  XOR U4194 ( .A(n3833), .B(n3834), .Z(n3830) );
  ANDN U4195 ( .A(n3835), .B(n3020), .Z(n3834) );
  XOR U4196 ( .A(n3833), .B(e_input[22]), .Z(n3020) );
  XOR U4197 ( .A(g_input[22]), .B(n3833), .Z(n3835) );
  XOR U4198 ( .A(n3836), .B(n3837), .Z(n3833) );
  ANDN U4199 ( .A(n3838), .B(n3054), .Z(n3837) );
  XOR U4200 ( .A(n3836), .B(e_input[21]), .Z(n3054) );
  XOR U4201 ( .A(g_input[21]), .B(n3836), .Z(n3838) );
  XOR U4202 ( .A(n3839), .B(n3840), .Z(n3836) );
  ANDN U4203 ( .A(n3841), .B(n3088), .Z(n3840) );
  XOR U4204 ( .A(n3839), .B(e_input[20]), .Z(n3088) );
  XOR U4205 ( .A(g_input[20]), .B(n3839), .Z(n3841) );
  XOR U4206 ( .A(n3842), .B(n3843), .Z(n3839) );
  ANDN U4207 ( .A(n3844), .B(n3122), .Z(n3843) );
  XOR U4208 ( .A(n3842), .B(e_input[19]), .Z(n3122) );
  XOR U4209 ( .A(g_input[19]), .B(n3842), .Z(n3844) );
  XOR U4210 ( .A(n3845), .B(n3846), .Z(n3842) );
  ANDN U4211 ( .A(n3847), .B(n3156), .Z(n3846) );
  XOR U4212 ( .A(n3845), .B(e_input[18]), .Z(n3156) );
  XOR U4213 ( .A(g_input[18]), .B(n3845), .Z(n3847) );
  XOR U4214 ( .A(n3848), .B(n3849), .Z(n3845) );
  ANDN U4215 ( .A(n3850), .B(n3190), .Z(n3849) );
  XOR U4216 ( .A(n3848), .B(e_input[17]), .Z(n3190) );
  XOR U4217 ( .A(g_input[17]), .B(n3848), .Z(n3850) );
  XOR U4218 ( .A(n3851), .B(n3852), .Z(n3848) );
  ANDN U4219 ( .A(n3853), .B(n3224), .Z(n3852) );
  XOR U4220 ( .A(n3851), .B(e_input[16]), .Z(n3224) );
  XOR U4221 ( .A(g_input[16]), .B(n3851), .Z(n3853) );
  XOR U4222 ( .A(n3854), .B(n3855), .Z(n3851) );
  ANDN U4223 ( .A(n3856), .B(n3258), .Z(n3855) );
  XOR U4224 ( .A(n3854), .B(e_input[15]), .Z(n3258) );
  XOR U4225 ( .A(g_input[15]), .B(n3854), .Z(n3856) );
  XOR U4226 ( .A(n3857), .B(n3858), .Z(n3854) );
  ANDN U4227 ( .A(n3859), .B(n3292), .Z(n3858) );
  XOR U4228 ( .A(n3857), .B(e_input[14]), .Z(n3292) );
  XOR U4229 ( .A(g_input[14]), .B(n3857), .Z(n3859) );
  XOR U4230 ( .A(n3860), .B(n3861), .Z(n3857) );
  ANDN U4231 ( .A(n3862), .B(n3326), .Z(n3861) );
  XOR U4232 ( .A(n3860), .B(e_input[13]), .Z(n3326) );
  XOR U4233 ( .A(g_input[13]), .B(n3860), .Z(n3862) );
  XOR U4234 ( .A(n3863), .B(n3864), .Z(n3860) );
  ANDN U4235 ( .A(n3865), .B(n3360), .Z(n3864) );
  XOR U4236 ( .A(n3863), .B(e_input[12]), .Z(n3360) );
  XOR U4237 ( .A(g_input[12]), .B(n3863), .Z(n3865) );
  XOR U4238 ( .A(n3866), .B(n3867), .Z(n3863) );
  ANDN U4239 ( .A(n3868), .B(n3394), .Z(n3867) );
  XOR U4240 ( .A(n3866), .B(e_input[11]), .Z(n3394) );
  XOR U4241 ( .A(g_input[11]), .B(n3866), .Z(n3868) );
  XOR U4242 ( .A(n3869), .B(n3870), .Z(n3866) );
  ANDN U4243 ( .A(n3871), .B(n3428), .Z(n3870) );
  XOR U4244 ( .A(n3869), .B(e_input[10]), .Z(n3428) );
  XOR U4245 ( .A(g_input[10]), .B(n3869), .Z(n3871) );
  XOR U4246 ( .A(n3872), .B(n3873), .Z(n3869) );
  ANDN U4247 ( .A(n3874), .B(n3462), .Z(n3873) );
  XOR U4248 ( .A(n3872), .B(e_input[9]), .Z(n3462) );
  XOR U4249 ( .A(g_input[9]), .B(n3872), .Z(n3874) );
  XOR U4250 ( .A(n3875), .B(n3876), .Z(n3872) );
  ANDN U4251 ( .A(n3877), .B(n3496), .Z(n3876) );
  XOR U4252 ( .A(n3875), .B(e_input[8]), .Z(n3496) );
  XOR U4253 ( .A(g_input[8]), .B(n3875), .Z(n3877) );
  XOR U4254 ( .A(n3878), .B(n3879), .Z(n3875) );
  ANDN U4255 ( .A(n3880), .B(n3530), .Z(n3879) );
  XOR U4256 ( .A(n3878), .B(e_input[7]), .Z(n3530) );
  XOR U4257 ( .A(g_input[7]), .B(n3878), .Z(n3880) );
  XOR U4258 ( .A(n3881), .B(n3882), .Z(n3878) );
  ANDN U4259 ( .A(n3883), .B(n3564), .Z(n3882) );
  XOR U4260 ( .A(n3881), .B(e_input[6]), .Z(n3564) );
  XOR U4261 ( .A(g_input[6]), .B(n3881), .Z(n3883) );
  XOR U4262 ( .A(n3884), .B(n3885), .Z(n3881) );
  ANDN U4263 ( .A(n3886), .B(n3598), .Z(n3885) );
  XOR U4264 ( .A(n3884), .B(e_input[5]), .Z(n3598) );
  XOR U4265 ( .A(g_input[5]), .B(n3884), .Z(n3886) );
  XOR U4266 ( .A(n3887), .B(n3888), .Z(n3884) );
  ANDN U4267 ( .A(n3889), .B(n3632), .Z(n3888) );
  XOR U4268 ( .A(n3887), .B(e_input[4]), .Z(n3632) );
  XOR U4269 ( .A(g_input[4]), .B(n3887), .Z(n3889) );
  XOR U4270 ( .A(n3890), .B(n3891), .Z(n3887) );
  ANDN U4271 ( .A(n3892), .B(n3664), .Z(n3891) );
  XOR U4272 ( .A(n3890), .B(e_input[3]), .Z(n3664) );
  XOR U4273 ( .A(g_input[3]), .B(n3890), .Z(n3892) );
  XOR U4274 ( .A(n3893), .B(n3894), .Z(n3890) );
  ANDN U4275 ( .A(n3895), .B(n3696), .Z(n3894) );
  XOR U4276 ( .A(n3893), .B(e_input[2]), .Z(n3696) );
  XNOR U4277 ( .A(n3691), .B(n3893), .Z(n3895) );
  IV U4278 ( .A(g_input[2]), .Z(n3691) );
  XNOR U4279 ( .A(n3896), .B(n3897), .Z(n3893) );
  NANDN U4280 ( .B(n3898), .A(n3899), .Z(n3896) );
  XOR U4281 ( .A(g_input[1]), .B(n3897), .Z(n3899) );
  XNOR U4282 ( .A(n3898), .B(g_input[1]), .Z(n3802) );
  XOR U4283 ( .A(n3897), .B(e_input[1]), .Z(n3898) );
  NOR U4284 ( .A(n1299), .B(e_input[0]), .Z(n3897) );
  XNOR U4285 ( .A(n3698), .B(\min_dist_reg[3][1] ), .Z(n3699) );
  NOR U4286 ( .A(\min_dist_reg[3][0] ), .B(n3900), .Z(n3698) );
  XOR U4287 ( .A(n2652), .B(n3900), .Z(n2653) );
  XNOR U4288 ( .A(n3704), .B(n3705), .Z(n3900) );
  XOR U4289 ( .A(e_input[32]), .B(n949), .Z(n3705) );
  IV U4290 ( .A(g_input[32]), .Z(n949) );
  XOR U4291 ( .A(e_input[0]), .B(n1299), .Z(n3704) );
  IV U4292 ( .A(g_input[0]), .Z(n1299) );
  IV U4293 ( .A(\min_dist_reg[3][0] ), .Z(n2652) );
  IV U4294 ( .A(\min_dist_reg[1][0] ), .Z(n2390) );
endmodule

